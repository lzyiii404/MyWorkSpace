//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_229(
  input  [1:0]  _EVAL,
  input         _EVAL_0,
  input  [29:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [1:0]  _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input  [29:0] _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  input  [1:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [31:0] _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input  [29:0] _EVAL_21,
  input         _EVAL_22,
  input  [29:0] _EVAL_23,
  input         _EVAL_24,
  input  [1:0]  _EVAL_25,
  input         _EVAL_26,
  input  [29:0] _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input  [31:0] _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  output [31:0] _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  input  [1:0]  _EVAL_40,
  input  [29:0] _EVAL_41,
  input         _EVAL_42,
  input  [29:0] _EVAL_43,
  input  [31:0] _EVAL_44,
  input         _EVAL_45,
  input  [1:0]  _EVAL_46,
  input  [31:0] _EVAL_47,
  input  [31:0] _EVAL_48,
  input  [1:0]  _EVAL_49,
  input  [29:0] _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  input  [31:0] _EVAL_57,
  input         _EVAL_58,
  input  [31:0] _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  input         _EVAL_62
);
  wire  pmp__EVAL;
  wire  pmp__EVAL_0;
  wire [29:0] pmp__EVAL_1;
  wire  pmp__EVAL_2;
  wire [1:0] pmp__EVAL_3;
  wire  pmp__EVAL_4;
  wire  pmp__EVAL_5;
  wire  pmp__EVAL_6;
  wire [31:0] pmp__EVAL_7;
  wire [1:0] pmp__EVAL_8;
  wire  pmp__EVAL_9;
  wire [31:0] pmp__EVAL_10;
  wire  pmp__EVAL_11;
  wire  pmp__EVAL_12;
  wire  pmp__EVAL_13;
  wire  pmp__EVAL_14;
  wire  pmp__EVAL_15;
  wire  pmp__EVAL_16;
  wire [1:0] pmp__EVAL_17;
  wire [29:0] pmp__EVAL_18;
  wire [1:0] pmp__EVAL_19;
  wire [31:0] pmp__EVAL_20;
  wire  pmp__EVAL_21;
  wire  pmp__EVAL_22;
  wire  pmp__EVAL_23;
  wire  pmp__EVAL_24;
  wire [1:0] pmp__EVAL_25;
  wire  pmp__EVAL_26;
  wire [31:0] pmp__EVAL_27;
  wire  pmp__EVAL_28;
  wire  pmp__EVAL_29;
  wire  pmp__EVAL_30;
  wire  pmp__EVAL_31;
  wire  pmp__EVAL_32;
  wire  pmp__EVAL_33;
  wire  pmp__EVAL_34;
  wire [1:0] pmp__EVAL_35;
  wire  pmp__EVAL_36;
  wire [31:0] pmp__EVAL_37;
  wire [1:0] pmp__EVAL_38;
  wire [31:0] pmp__EVAL_39;
  wire  pmp__EVAL_40;
  wire  pmp__EVAL_41;
  wire [29:0] pmp__EVAL_42;
  wire [29:0] pmp__EVAL_43;
  wire  pmp__EVAL_44;
  wire [29:0] pmp__EVAL_45;
  wire  pmp__EVAL_46;
  wire [29:0] pmp__EVAL_47;
  wire  pmp__EVAL_48;
  wire [31:0] pmp__EVAL_49;
  wire  pmp__EVAL_50;
  wire [1:0] pmp__EVAL_51;
  wire  pmp__EVAL_52;
  wire [29:0] pmp__EVAL_53;
  wire [31:0] pmp__EVAL_54;
  wire  pmp__EVAL_55;
  wire [1:0] pmp__EVAL_56;
  wire [29:0] pmp__EVAL_57;
  wire  pmp__EVAL_58;
  wire [31:0] pmp__EVAL_59;
  wire [19:0] _EVAL_110;
  wire [11:0] _EVAL_66;
  wire [31:0] _EVAL_159;
  wire [31:0] _EVAL_131;
  wire [31:0] _EVAL_141;
  wire [32:0] _EVAL_65;
  wire [32:0] _EVAL_112;
  wire [32:0] _EVAL_75;
  wire [31:0] _EVAL_149;
  wire [32:0] _EVAL_90;
  wire [32:0] _EVAL_146;
  wire [32:0] _EVAL_147;
  wire [32:0] _EVAL_132;
  wire [32:0] _EVAL_162;
  wire  _EVAL_88;
  wire [31:0] _EVAL_161;
  wire [32:0] _EVAL_117;
  wire [32:0] _EVAL_127;
  wire [32:0] _EVAL_64;
  wire  _EVAL_68;
  wire [32:0] _EVAL_98;
  wire  _EVAL_120;
  wire  _EVAL_126;
  wire [31:0] _EVAL_85;
  wire [32:0] _EVAL_70;
  wire [32:0] _EVAL_73;
  wire [32:0] _EVAL_152;
  wire  _EVAL_115;
  wire  _EVAL_139;
  wire [31:0] _EVAL_77;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_153;
  wire [32:0] _EVAL_107;
  wire  _EVAL_114;
  wire  _EVAL_136;
  wire [31:0] _EVAL_113;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_86;
  wire [32:0] _EVAL_74;
  wire  _EVAL_100;
  wire  _EVAL_142;
  wire [32:0] _EVAL_95;
  wire [32:0] _EVAL_69;
  wire  _EVAL_87;
  wire  _EVAL_76;
  wire [31:0] _EVAL_89;
  wire [32:0] _EVAL_101;
  wire [32:0] _EVAL_67;
  wire [32:0] _EVAL_83;
  wire  _EVAL_96;
  wire  _EVAL_154;
  wire [32:0] _EVAL_133;
  wire [32:0] _EVAL_63;
  wire [32:0] _EVAL_140;
  wire  _EVAL_105;
  wire  _EVAL_103;
  wire [31:0] _EVAL_155;
  wire [32:0] _EVAL_81;
  wire [32:0] _EVAL_125;
  wire [32:0] _EVAL_144;
  wire  _EVAL_123;
  wire  _EVAL_79;
  wire [31:0] _EVAL_157;
  wire [32:0] _EVAL_109;
  wire [32:0] _EVAL_91;
  wire [32:0] _EVAL_108;
  wire  _EVAL_137;
  wire  _EVAL_84;
  wire [32:0] _EVAL_72;
  wire [32:0] _EVAL_92;
  wire  _EVAL_78;
  wire  _EVAL_80;
  wire [1:0] _EVAL_82;
  wire [2:0] _EVAL_106;
  wire  _EVAL_121;
  wire [32:0] _EVAL_143;
  wire [32:0] _EVAL_71;
  wire  _EVAL_94;
  wire  _EVAL_160;
  wire  _EVAL_138;
  wire  _EVAL_128;
  wire [32:0] _EVAL_119;
  wire [32:0] _EVAL_145;
  wire  _EVAL_116;
  wire  _EVAL_122;
  wire [32:0] _EVAL_93;
  wire [32:0] _EVAL_111;
  wire  _EVAL_104;
  wire  _EVAL_148;
  wire  _EVAL_99;
  wire  _EVAL_124;
  wire  _EVAL_150;
  wire  _EVAL_135;
  wire [15:0] _EVAL_97;
  wire [15:0] _EVAL_156;
  wire  _EVAL_129;
  wire [1:0] _EVAL_158;
  wire [15:0] _EVAL_134;
  wire [15:0] _EVAL_151;
  wire [15:0] _EVAL_102;
  wire [19:0] _EVAL_118;
  SiFive__EVAL_228 pmp (
    ._EVAL(pmp__EVAL),
    ._EVAL_0(pmp__EVAL_0),
    ._EVAL_1(pmp__EVAL_1),
    ._EVAL_2(pmp__EVAL_2),
    ._EVAL_3(pmp__EVAL_3),
    ._EVAL_4(pmp__EVAL_4),
    ._EVAL_5(pmp__EVAL_5),
    ._EVAL_6(pmp__EVAL_6),
    ._EVAL_7(pmp__EVAL_7),
    ._EVAL_8(pmp__EVAL_8),
    ._EVAL_9(pmp__EVAL_9),
    ._EVAL_10(pmp__EVAL_10),
    ._EVAL_11(pmp__EVAL_11),
    ._EVAL_12(pmp__EVAL_12),
    ._EVAL_13(pmp__EVAL_13),
    ._EVAL_14(pmp__EVAL_14),
    ._EVAL_15(pmp__EVAL_15),
    ._EVAL_16(pmp__EVAL_16),
    ._EVAL_17(pmp__EVAL_17),
    ._EVAL_18(pmp__EVAL_18),
    ._EVAL_19(pmp__EVAL_19),
    ._EVAL_20(pmp__EVAL_20),
    ._EVAL_21(pmp__EVAL_21),
    ._EVAL_22(pmp__EVAL_22),
    ._EVAL_23(pmp__EVAL_23),
    ._EVAL_24(pmp__EVAL_24),
    ._EVAL_25(pmp__EVAL_25),
    ._EVAL_26(pmp__EVAL_26),
    ._EVAL_27(pmp__EVAL_27),
    ._EVAL_28(pmp__EVAL_28),
    ._EVAL_29(pmp__EVAL_29),
    ._EVAL_30(pmp__EVAL_30),
    ._EVAL_31(pmp__EVAL_31),
    ._EVAL_32(pmp__EVAL_32),
    ._EVAL_33(pmp__EVAL_33),
    ._EVAL_34(pmp__EVAL_34),
    ._EVAL_35(pmp__EVAL_35),
    ._EVAL_36(pmp__EVAL_36),
    ._EVAL_37(pmp__EVAL_37),
    ._EVAL_38(pmp__EVAL_38),
    ._EVAL_39(pmp__EVAL_39),
    ._EVAL_40(pmp__EVAL_40),
    ._EVAL_41(pmp__EVAL_41),
    ._EVAL_42(pmp__EVAL_42),
    ._EVAL_43(pmp__EVAL_43),
    ._EVAL_44(pmp__EVAL_44),
    ._EVAL_45(pmp__EVAL_45),
    ._EVAL_46(pmp__EVAL_46),
    ._EVAL_47(pmp__EVAL_47),
    ._EVAL_48(pmp__EVAL_48),
    ._EVAL_49(pmp__EVAL_49),
    ._EVAL_50(pmp__EVAL_50),
    ._EVAL_51(pmp__EVAL_51),
    ._EVAL_52(pmp__EVAL_52),
    ._EVAL_53(pmp__EVAL_53),
    ._EVAL_54(pmp__EVAL_54),
    ._EVAL_55(pmp__EVAL_55),
    ._EVAL_56(pmp__EVAL_56),
    ._EVAL_57(pmp__EVAL_57),
    ._EVAL_58(pmp__EVAL_58),
    ._EVAL_59(pmp__EVAL_59)
  );
  assign _EVAL_110 = _EVAL_57[31:12];
  assign _EVAL_66 = _EVAL_57[11:0];
  assign _EVAL_159 = {_EVAL_110,_EVAL_66};
  assign _EVAL_131 = _EVAL_159 ^ 32'h1900000;
  assign _EVAL_141 = _EVAL_159 ^ 32'h1000000;
  assign _EVAL_65 = {1'b0,$signed(_EVAL_141)};
  assign _EVAL_112 = $signed(_EVAL_65) & $signed(33'sheb000000);
  assign _EVAL_75 = $signed(_EVAL_112);
  assign _EVAL_149 = _EVAL_159 ^ 32'h80000000;
  assign _EVAL_90 = {1'b0,$signed(_EVAL_149)};
  assign _EVAL_146 = $signed(_EVAL_90) & $signed(-33'sh20000);
  assign _EVAL_147 = {1'b0,$signed(_EVAL_159)};
  assign _EVAL_132 = $signed(_EVAL_147) & $signed(33'shab004000);
  assign _EVAL_162 = $signed(_EVAL_132);
  assign _EVAL_88 = $signed(_EVAL_162) == $signed(33'sh0);
  assign _EVAL_161 = _EVAL_159 ^ 32'h40000000;
  assign _EVAL_117 = {1'b0,$signed(_EVAL_161)};
  assign _EVAL_127 = $signed(_EVAL_117) & $signed(-33'sh2000);
  assign _EVAL_64 = $signed(_EVAL_127);
  assign _EVAL_68 = $signed(_EVAL_64) == $signed(33'sh0);
  assign _EVAL_98 = $signed(_EVAL_146);
  assign _EVAL_120 = $signed(_EVAL_98) == $signed(33'sh0);
  assign _EVAL_126 = _EVAL_68 | _EVAL_120;
  assign _EVAL_85 = _EVAL_159 ^ 32'h3000;
  assign _EVAL_70 = {1'b0,$signed(_EVAL_85)};
  assign _EVAL_73 = $signed(_EVAL_70) & $signed(-33'sh1000);
  assign _EVAL_152 = $signed(_EVAL_73);
  assign _EVAL_115 = $signed(_EVAL_152) == $signed(33'sh0);
  assign _EVAL_139 = _EVAL_126 | _EVAL_115;
  assign _EVAL_77 = _EVAL_159 ^ 32'hc000000;
  assign _EVAL_163 = {1'b0,$signed(_EVAL_77)};
  assign _EVAL_153 = $signed(_EVAL_163) & $signed(-33'sh4000000);
  assign _EVAL_107 = $signed(_EVAL_153);
  assign _EVAL_114 = $signed(_EVAL_107) == $signed(33'sh0);
  assign _EVAL_136 = _EVAL_139 | _EVAL_114;
  assign _EVAL_113 = _EVAL_159 ^ 32'h2000000;
  assign _EVAL_130 = {1'b0,$signed(_EVAL_113)};
  assign _EVAL_86 = $signed(_EVAL_130) & $signed(-33'sh10000);
  assign _EVAL_74 = $signed(_EVAL_86);
  assign _EVAL_100 = $signed(_EVAL_74) == $signed(33'sh0);
  assign _EVAL_142 = _EVAL_136 | _EVAL_100;
  assign _EVAL_95 = $signed(_EVAL_147) & $signed(-33'sh1000);
  assign _EVAL_69 = $signed(_EVAL_95);
  assign _EVAL_87 = $signed(_EVAL_69) == $signed(33'sh0);
  assign _EVAL_76 = _EVAL_142 | _EVAL_87;
  assign _EVAL_89 = _EVAL_159 ^ 32'h1800000;
  assign _EVAL_101 = {1'b0,$signed(_EVAL_89)};
  assign _EVAL_67 = $signed(_EVAL_101) & $signed(-33'sh8000);
  assign _EVAL_83 = $signed(_EVAL_67);
  assign _EVAL_96 = $signed(_EVAL_83) == $signed(33'sh0);
  assign _EVAL_154 = _EVAL_76 | _EVAL_96;
  assign _EVAL_133 = {1'b0,$signed(_EVAL_131)};
  assign _EVAL_63 = $signed(_EVAL_133) & $signed(-33'sh2000);
  assign _EVAL_140 = $signed(_EVAL_63);
  assign _EVAL_105 = $signed(_EVAL_140) == $signed(33'sh0);
  assign _EVAL_103 = _EVAL_154 | _EVAL_105;
  assign _EVAL_155 = _EVAL_159 ^ 32'h4000;
  assign _EVAL_81 = {1'b0,$signed(_EVAL_155)};
  assign _EVAL_125 = $signed(_EVAL_81) & $signed(-33'sh1000);
  assign _EVAL_144 = $signed(_EVAL_125);
  assign _EVAL_123 = $signed(_EVAL_144) == $signed(33'sh0);
  assign _EVAL_79 = _EVAL_103 | _EVAL_123;
  assign _EVAL_157 = _EVAL_159 ^ 32'h20000000;
  assign _EVAL_109 = {1'b0,$signed(_EVAL_157)};
  assign _EVAL_91 = $signed(_EVAL_109) & $signed(-33'sh2000);
  assign _EVAL_108 = $signed(_EVAL_91);
  assign _EVAL_137 = $signed(_EVAL_108) == $signed(33'sh0);
  assign _EVAL_84 = _EVAL_79 | _EVAL_137;
  assign _EVAL_72 = $signed(_EVAL_90) & $signed(33'sh80000000);
  assign _EVAL_92 = $signed(_EVAL_72);
  assign _EVAL_78 = $signed(_EVAL_92) == $signed(33'sh0);
  assign _EVAL_80 = _EVAL_84 & _EVAL_78;
  assign _EVAL_82 = _EVAL_80 ? 2'h3 : 2'h0;
  assign _EVAL_106 = {_EVAL_2,_EVAL_16};
  assign _EVAL_121 = _EVAL_106 <= 3'h3;
  assign _EVAL_143 = $signed(_EVAL_90) & $signed(33'sheb000000);
  assign _EVAL_71 = $signed(_EVAL_143);
  assign _EVAL_94 = $signed(_EVAL_71) == $signed(33'sh0);
  assign _EVAL_160 = _EVAL_88 | _EVAL_94;
  assign _EVAL_138 = $signed(_EVAL_75) == $signed(33'sh0);
  assign _EVAL_128 = _EVAL_160 | _EVAL_138;
  assign _EVAL_119 = $signed(_EVAL_65) & $signed(33'sheb004000);
  assign _EVAL_145 = $signed(_EVAL_119);
  assign _EVAL_116 = $signed(_EVAL_145) == $signed(33'sh0);
  assign _EVAL_122 = _EVAL_128 | _EVAL_116;
  assign _EVAL_93 = $signed(_EVAL_109) & $signed(33'sheb004000);
  assign _EVAL_111 = $signed(_EVAL_93);
  assign _EVAL_104 = $signed(_EVAL_111) == $signed(33'sh0);
  assign _EVAL_148 = _EVAL_122 | _EVAL_104;
  assign _EVAL_99 = _EVAL_84 & _EVAL_148;
  assign _EVAL_124 = _EVAL_121 & _EVAL_87;
  assign _EVAL_150 = _EVAL_124 == 1'h0;
  assign _EVAL_135 = _EVAL_99 & _EVAL_150;
  assign _EVAL_97 = {_EVAL_82,14'h0};
  assign _EVAL_156 = _EVAL_97 & 16'h8000;
  assign _EVAL_129 = _EVAL_135 & pmp__EVAL_26;
  assign _EVAL_158 = _EVAL_129 ? 2'h3 : 2'h0;
  assign _EVAL_134 = {_EVAL_158,14'h0};
  assign _EVAL_151 = ~ _EVAL_134;
  assign _EVAL_102 = _EVAL_151 & 16'h8000;
  assign _EVAL_118 = _EVAL_57[31:12];
  assign pmp__EVAL_4 = _EVAL_62;
  assign pmp__EVAL_35 = _EVAL;
  assign pmp__EVAL_18 = _EVAL_50;
  assign pmp__EVAL_45 = _EVAL_23;
  assign pmp__EVAL_36 = _EVAL_26;
  assign pmp__EVAL_58 = _EVAL_53;
  assign _EVAL_10 = _EVAL_156 != 16'h0;
  assign pmp__EVAL_50 = _EVAL_11;
  assign pmp__EVAL_44 = _EVAL_3;
  assign pmp__EVAL_30 = _EVAL_12;
  assign pmp__EVAL_32 = _EVAL_28;
  assign pmp__EVAL_1 = _EVAL_43;
  assign pmp__EVAL_57 = _EVAL_27;
  assign pmp__EVAL_42 = _EVAL_1;
  assign pmp__EVAL_28 = _EVAL_29;
  assign pmp__EVAL_40 = _EVAL_32;
  assign pmp__EVAL_53 = _EVAL_9;
  assign pmp__EVAL_39 = _EVAL_44;
  assign pmp__EVAL_12 = _EVAL_33;
  assign pmp__EVAL_6 = _EVAL_58;
  assign pmp__EVAL_38 = _EVAL_106[1:0];
  assign pmp__EVAL_49 = _EVAL_8;
  assign pmp__EVAL_59 = _EVAL_48;
  assign pmp__EVAL_8 = _EVAL_15;
  assign pmp__EVAL_29 = _EVAL_35;
  assign pmp__EVAL_24 = _EVAL_54;
  assign pmp__EVAL_16 = _EVAL_42;
  assign pmp__EVAL_34 = _EVAL_13;
  assign pmp__EVAL_10 = {_EVAL_110,_EVAL_66};
  assign pmp__EVAL_47 = _EVAL_41;
  assign pmp__EVAL_22 = _EVAL_30;
  assign pmp__EVAL_43 = _EVAL_21;
  assign pmp__EVAL_48 = _EVAL_31;
  assign _EVAL_39 = _EVAL_102 != 16'h0;
  assign pmp__EVAL_9 = _EVAL_0;
  assign pmp__EVAL_51 = _EVAL_46;
  assign pmp__EVAL_5 = _EVAL_52;
  assign pmp__EVAL_20 = _EVAL_18;
  assign pmp__EVAL_37 = _EVAL_59;
  assign _EVAL_37 = {_EVAL_118,_EVAL_66};
  assign pmp__EVAL_2 = _EVAL_14;
  assign pmp__EVAL_41 = _EVAL_51;
  assign pmp__EVAL_19 = _EVAL_25;
  assign pmp__EVAL_46 = _EVAL_60;
  assign pmp__EVAL_0 = _EVAL_19;
  assign pmp__EVAL_52 = _EVAL_61;
  assign pmp__EVAL = _EVAL_4;
  assign pmp__EVAL_21 = _EVAL_56;
  assign pmp__EVAL_15 = _EVAL_55;
  assign pmp__EVAL_17 = _EVAL_49;
  assign pmp__EVAL_56 = _EVAL_7;
  assign pmp__EVAL_3 = _EVAL_40;
  assign pmp__EVAL_13 = _EVAL_22;
  assign pmp__EVAL_31 = _EVAL_24;
  assign pmp__EVAL_23 = _EVAL_36;
  assign pmp__EVAL_7 = _EVAL_34;
  assign pmp__EVAL_14 = _EVAL_38;
  assign pmp__EVAL_33 = _EVAL_6;
  assign pmp__EVAL_55 = _EVAL_45;
  assign pmp__EVAL_25 = _EVAL_5;
  assign pmp__EVAL_11 = _EVAL_20;
  assign pmp__EVAL_54 = _EVAL_47;
  assign pmp__EVAL_27 = _EVAL_17;
endmodule
