//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_273(
  output [63:0] _EVAL,
  output [31:0] _EVAL_0,
  output        _EVAL_1,
  output [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output [3:0]  _EVAL_5,
  output [63:0] _EVAL_6,
  input         _EVAL_7,
  output [3:0]  _EVAL_8,
  output [1:0]  _EVAL_9,
  output        _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  output [63:0] _EVAL_14,
  input  [63:0] _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  output [1:0]  _EVAL_18,
  output [31:0] _EVAL_19,
  output [3:0]  _EVAL_20,
  input  [3:0]  _EVAL_21,
  input  [3:0]  _EVAL_22,
  input         _EVAL_23,
  input  [1:0]  _EVAL_24,
  output [3:0]  _EVAL_25,
  input  [3:0]  _EVAL_26,
  input         _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  output [63:0] _EVAL_30,
  output [7:0]  _EVAL_31,
  output        _EVAL_32,
  input  [31:0] _EVAL_33,
  input  [3:0]  _EVAL_34,
  input  [63:0] _EVAL_35,
  output [2:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  output        _EVAL_38,
  output        _EVAL_39,
  output [7:0]  _EVAL_40,
  input  [1:0]  _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  input         _EVAL_44,
  output [1:0]  _EVAL_45,
  output [2:0]  _EVAL_46,
  output        _EVAL_47,
  output [3:0]  _EVAL_48,
  output [31:0] _EVAL_49,
  input  [1:0]  _EVAL_50,
  output [1:0]  _EVAL_51,
  input  [1:0]  _EVAL_52,
  output        _EVAL_53,
  input  [2:0]  _EVAL_54,
  output        _EVAL_55,
  input  [2:0]  _EVAL_56,
  output [1:0]  _EVAL_57,
  output        _EVAL_58,
  output        _EVAL_59,
  input  [63:0] _EVAL_60,
  input         _EVAL_61,
  input  [31:0] _EVAL_62,
  output [3:0]  _EVAL_63,
  output [3:0]  _EVAL_64,
  output [1:0]  _EVAL_65,
  input  [1:0]  _EVAL_66,
  input         _EVAL_67,
  input  [31:0] _EVAL_68,
  input  [2:0]  _EVAL_69,
  input  [1:0]  _EVAL_70,
  input  [31:0] _EVAL_71,
  output        _EVAL_72,
  output        _EVAL_73,
  input  [2:0]  _EVAL_74,
  input         _EVAL_75,
  output [63:0] _EVAL_76,
  input         _EVAL_77,
  input         _EVAL_78,
  output [31:0] _EVAL_79,
  output        _EVAL_80,
  output [2:0]  _EVAL_81,
  input  [2:0]  _EVAL_82,
  output        _EVAL_83,
  input  [2:0]  _EVAL_84,
  output [3:0]  _EVAL_85,
  input  [1:0]  _EVAL_86,
  output        _EVAL_87,
  input  [3:0]  _EVAL_88,
  input  [63:0] _EVAL_89,
  output [3:0]  _EVAL_90,
  output [2:0]  _EVAL_91,
  output [3:0]  _EVAL_92,
  input  [1:0]  _EVAL_93,
  output        _EVAL_94,
  output [31:0] _EVAL_95,
  input         _EVAL_96,
  output [2:0]  _EVAL_97,
  output [2:0]  _EVAL_98,
  output [1:0]  _EVAL_99,
  input  [7:0]  _EVAL_100,
  input  [1:0]  _EVAL_101,
  input         _EVAL_102,
  output [2:0]  _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  input  [3:0]  _EVAL_106,
  input         _EVAL_107,
  input         _EVAL_108
);
  wire [3:0] RationalCrossingSource__EVAL;
  wire [1:0] RationalCrossingSource__EVAL_0;
  wire  RationalCrossingSource__EVAL_1;
  wire [7:0] RationalCrossingSource__EVAL_2;
  wire [3:0] RationalCrossingSource__EVAL_3;
  wire [3:0] RationalCrossingSource__EVAL_4;
  wire [2:0] RationalCrossingSource__EVAL_5;
  wire [63:0] RationalCrossingSource__EVAL_6;
  wire [3:0] RationalCrossingSource__EVAL_7;
  wire [7:0] RationalCrossingSource__EVAL_8;
  wire  RationalCrossingSource__EVAL_9;
  wire [2:0] RationalCrossingSource__EVAL_10;
  wire [2:0] RationalCrossingSource__EVAL_11;
  wire  RationalCrossingSource__EVAL_12;
  wire [31:0] RationalCrossingSource__EVAL_13;
  wire [31:0] RationalCrossingSource__EVAL_14;
  wire  RationalCrossingSource__EVAL_15;
  wire [63:0] RationalCrossingSource__EVAL_16;
  wire  RationalCrossingSource__EVAL_17;
  wire [2:0] RationalCrossingSource__EVAL_18;
  wire  RationalCrossingSource__EVAL_19;
  wire  RationalCrossingSource__EVAL_20;
  wire [2:0] RationalCrossingSource__EVAL_21;
  wire  RationalCrossingSource__EVAL_22;
  wire [63:0] RationalCrossingSource__EVAL_23;
  wire [2:0] RationalCrossingSource__EVAL_24;
  wire  RationalCrossingSource__EVAL_25;
  wire [31:0] RationalCrossingSource__EVAL_26;
  wire [3:0] RationalCrossingSource__EVAL_27;
  wire [7:0] RationalCrossingSource__EVAL_28;
  wire [1:0] RationalCrossingSource__EVAL_29;
  wire [3:0] RationalCrossingSource__EVAL_30;
  wire  RationalCrossingSink_1__EVAL;
  wire [1:0] RationalCrossingSink_1__EVAL_0;
  wire  RationalCrossingSink_1__EVAL_1;
  wire [1:0] RationalCrossingSink_1__EVAL_2;
  wire [1:0] RationalCrossingSink_1__EVAL_3;
  wire  RationalCrossingSink_1__EVAL_4;
  wire [1:0] RationalCrossingSink_1__EVAL_5;
  wire [1:0] RationalCrossingSink_1__EVAL_6;
  wire  RationalCrossingSink_1__EVAL_7;
  wire [31:0] RationalCrossingSink_1__EVAL_8;
  wire [31:0] RationalCrossingSink_1__EVAL_9;
  wire [31:0] RationalCrossingSink_1__EVAL_10;
  wire  RationalCrossingSink_1__EVAL_11;
  wire  RationalCrossingSink_1__EVAL_12;
  wire [3:0] RationalCrossingSource_1__EVAL;
  wire [31:0] RationalCrossingSource_1__EVAL_0;
  wire  RationalCrossingSource_1__EVAL_1;
  wire [2:0] RationalCrossingSource_1__EVAL_2;
  wire [63:0] RationalCrossingSource_1__EVAL_3;
  wire [3:0] RationalCrossingSource_1__EVAL_4;
  wire [2:0] RationalCrossingSource_1__EVAL_5;
  wire  RationalCrossingSource_1__EVAL_6;
  wire  RationalCrossingSource_1__EVAL_7;
  wire [31:0] RationalCrossingSource_1__EVAL_8;
  wire  RationalCrossingSource_1__EVAL_9;
  wire [31:0] RationalCrossingSource_1__EVAL_10;
  wire [3:0] RationalCrossingSource_1__EVAL_11;
  wire  RationalCrossingSource_1__EVAL_12;
  wire [3:0] RationalCrossingSource_1__EVAL_13;
  wire [2:0] RationalCrossingSource_1__EVAL_14;
  wire  RationalCrossingSource_1__EVAL_15;
  wire [2:0] RationalCrossingSource_1__EVAL_16;
  wire [3:0] RationalCrossingSource_1__EVAL_17;
  wire  RationalCrossingSource_1__EVAL_18;
  wire [2:0] RationalCrossingSource_1__EVAL_19;
  wire [1:0] RationalCrossingSource_1__EVAL_20;
  wire [3:0] RationalCrossingSource_1__EVAL_21;
  wire  RationalCrossingSource_1__EVAL_22;
  wire [63:0] RationalCrossingSource_1__EVAL_23;
  wire [63:0] RationalCrossingSource_1__EVAL_24;
  wire  RationalCrossingSource_1__EVAL_25;
  wire [1:0] RationalCrossingSource_1__EVAL_26;
  wire [2:0] RationalCrossingSource_1__EVAL_27;
  wire  RationalCrossingSink__EVAL;
  wire [3:0] RationalCrossingSink__EVAL_0;
  wire [1:0] RationalCrossingSink__EVAL_1;
  wire [63:0] RationalCrossingSink__EVAL_2;
  wire  RationalCrossingSink__EVAL_3;
  wire  RationalCrossingSink__EVAL_4;
  wire  RationalCrossingSink__EVAL_5;
  wire  RationalCrossingSink__EVAL_6;
  wire [63:0] RationalCrossingSink__EVAL_7;
  wire [2:0] RationalCrossingSink__EVAL_8;
  wire  RationalCrossingSink__EVAL_9;
  wire  RationalCrossingSink__EVAL_10;
  wire [63:0] RationalCrossingSink__EVAL_11;
  wire [2:0] RationalCrossingSink__EVAL_12;
  wire  RationalCrossingSink__EVAL_13;
  wire [1:0] RationalCrossingSink__EVAL_14;
  wire  RationalCrossingSink__EVAL_15;
  wire [1:0] RationalCrossingSink__EVAL_16;
  wire [3:0] RationalCrossingSink__EVAL_17;
  wire  RationalCrossingSink__EVAL_18;
  wire  RationalCrossingSink__EVAL_19;
  wire  RationalCrossingSink__EVAL_20;
  wire [1:0] RationalCrossingSink__EVAL_21;
  wire [3:0] RationalCrossingSink__EVAL_22;
  wire  RationalCrossingSink__EVAL_23;
  wire [3:0] RationalCrossingSink__EVAL_24;
  wire [2:0] RationalCrossingSink__EVAL_25;
  wire [1:0] RationalCrossingSink__EVAL_26;
  wire [3:0] RationalCrossingSink__EVAL_27;
  wire  RationalCrossingSink__EVAL_28;
  wire  RationalCrossingSink__EVAL_29;
  wire [3:0] RationalCrossingSink__EVAL_30;
  wire  RationalCrossingSource_2__EVAL;
  wire  RationalCrossingSource_2__EVAL_0;
  wire  RationalCrossingSource_2__EVAL_1;
  wire  RationalCrossingSource_2__EVAL_2;
  wire  RationalCrossingSource_2__EVAL_3;
  wire  RationalCrossingSource_2__EVAL_4;
  wire  RationalCrossingSource_2__EVAL_5;
  wire  RationalCrossingSource_2__EVAL_6;
  wire [1:0] RationalCrossingSource_2__EVAL_7;
  wire  RationalCrossingSource_2__EVAL_8;
  wire [1:0] RationalCrossingSource_2__EVAL_9;
  SiFive__EVAL_268 RationalCrossingSource (
    ._EVAL(RationalCrossingSource__EVAL),
    ._EVAL_0(RationalCrossingSource__EVAL_0),
    ._EVAL_1(RationalCrossingSource__EVAL_1),
    ._EVAL_2(RationalCrossingSource__EVAL_2),
    ._EVAL_3(RationalCrossingSource__EVAL_3),
    ._EVAL_4(RationalCrossingSource__EVAL_4),
    ._EVAL_5(RationalCrossingSource__EVAL_5),
    ._EVAL_6(RationalCrossingSource__EVAL_6),
    ._EVAL_7(RationalCrossingSource__EVAL_7),
    ._EVAL_8(RationalCrossingSource__EVAL_8),
    ._EVAL_9(RationalCrossingSource__EVAL_9),
    ._EVAL_10(RationalCrossingSource__EVAL_10),
    ._EVAL_11(RationalCrossingSource__EVAL_11),
    ._EVAL_12(RationalCrossingSource__EVAL_12),
    ._EVAL_13(RationalCrossingSource__EVAL_13),
    ._EVAL_14(RationalCrossingSource__EVAL_14),
    ._EVAL_15(RationalCrossingSource__EVAL_15),
    ._EVAL_16(RationalCrossingSource__EVAL_16),
    ._EVAL_17(RationalCrossingSource__EVAL_17),
    ._EVAL_18(RationalCrossingSource__EVAL_18),
    ._EVAL_19(RationalCrossingSource__EVAL_19),
    ._EVAL_20(RationalCrossingSource__EVAL_20),
    ._EVAL_21(RationalCrossingSource__EVAL_21),
    ._EVAL_22(RationalCrossingSource__EVAL_22),
    ._EVAL_23(RationalCrossingSource__EVAL_23),
    ._EVAL_24(RationalCrossingSource__EVAL_24),
    ._EVAL_25(RationalCrossingSource__EVAL_25),
    ._EVAL_26(RationalCrossingSource__EVAL_26),
    ._EVAL_27(RationalCrossingSource__EVAL_27),
    ._EVAL_28(RationalCrossingSource__EVAL_28),
    ._EVAL_29(RationalCrossingSource__EVAL_29),
    ._EVAL_30(RationalCrossingSource__EVAL_30)
  );
  SiFive__EVAL_270 RationalCrossingSink_1 (
    ._EVAL(RationalCrossingSink_1__EVAL),
    ._EVAL_0(RationalCrossingSink_1__EVAL_0),
    ._EVAL_1(RationalCrossingSink_1__EVAL_1),
    ._EVAL_2(RationalCrossingSink_1__EVAL_2),
    ._EVAL_3(RationalCrossingSink_1__EVAL_3),
    ._EVAL_4(RationalCrossingSink_1__EVAL_4),
    ._EVAL_5(RationalCrossingSink_1__EVAL_5),
    ._EVAL_6(RationalCrossingSink_1__EVAL_6),
    ._EVAL_7(RationalCrossingSink_1__EVAL_7),
    ._EVAL_8(RationalCrossingSink_1__EVAL_8),
    ._EVAL_9(RationalCrossingSink_1__EVAL_9),
    ._EVAL_10(RationalCrossingSink_1__EVAL_10),
    ._EVAL_11(RationalCrossingSink_1__EVAL_11),
    ._EVAL_12(RationalCrossingSink_1__EVAL_12)
  );
  SiFive__EVAL_271 RationalCrossingSource_1 (
    ._EVAL(RationalCrossingSource_1__EVAL),
    ._EVAL_0(RationalCrossingSource_1__EVAL_0),
    ._EVAL_1(RationalCrossingSource_1__EVAL_1),
    ._EVAL_2(RationalCrossingSource_1__EVAL_2),
    ._EVAL_3(RationalCrossingSource_1__EVAL_3),
    ._EVAL_4(RationalCrossingSource_1__EVAL_4),
    ._EVAL_5(RationalCrossingSource_1__EVAL_5),
    ._EVAL_6(RationalCrossingSource_1__EVAL_6),
    ._EVAL_7(RationalCrossingSource_1__EVAL_7),
    ._EVAL_8(RationalCrossingSource_1__EVAL_8),
    ._EVAL_9(RationalCrossingSource_1__EVAL_9),
    ._EVAL_10(RationalCrossingSource_1__EVAL_10),
    ._EVAL_11(RationalCrossingSource_1__EVAL_11),
    ._EVAL_12(RationalCrossingSource_1__EVAL_12),
    ._EVAL_13(RationalCrossingSource_1__EVAL_13),
    ._EVAL_14(RationalCrossingSource_1__EVAL_14),
    ._EVAL_15(RationalCrossingSource_1__EVAL_15),
    ._EVAL_16(RationalCrossingSource_1__EVAL_16),
    ._EVAL_17(RationalCrossingSource_1__EVAL_17),
    ._EVAL_18(RationalCrossingSource_1__EVAL_18),
    ._EVAL_19(RationalCrossingSource_1__EVAL_19),
    ._EVAL_20(RationalCrossingSource_1__EVAL_20),
    ._EVAL_21(RationalCrossingSource_1__EVAL_21),
    ._EVAL_22(RationalCrossingSource_1__EVAL_22),
    ._EVAL_23(RationalCrossingSource_1__EVAL_23),
    ._EVAL_24(RationalCrossingSource_1__EVAL_24),
    ._EVAL_25(RationalCrossingSource_1__EVAL_25),
    ._EVAL_26(RationalCrossingSource_1__EVAL_26),
    ._EVAL_27(RationalCrossingSource_1__EVAL_27)
  );
  SiFive__EVAL_269 RationalCrossingSink (
    ._EVAL(RationalCrossingSink__EVAL),
    ._EVAL_0(RationalCrossingSink__EVAL_0),
    ._EVAL_1(RationalCrossingSink__EVAL_1),
    ._EVAL_2(RationalCrossingSink__EVAL_2),
    ._EVAL_3(RationalCrossingSink__EVAL_3),
    ._EVAL_4(RationalCrossingSink__EVAL_4),
    ._EVAL_5(RationalCrossingSink__EVAL_5),
    ._EVAL_6(RationalCrossingSink__EVAL_6),
    ._EVAL_7(RationalCrossingSink__EVAL_7),
    ._EVAL_8(RationalCrossingSink__EVAL_8),
    ._EVAL_9(RationalCrossingSink__EVAL_9),
    ._EVAL_10(RationalCrossingSink__EVAL_10),
    ._EVAL_11(RationalCrossingSink__EVAL_11),
    ._EVAL_12(RationalCrossingSink__EVAL_12),
    ._EVAL_13(RationalCrossingSink__EVAL_13),
    ._EVAL_14(RationalCrossingSink__EVAL_14),
    ._EVAL_15(RationalCrossingSink__EVAL_15),
    ._EVAL_16(RationalCrossingSink__EVAL_16),
    ._EVAL_17(RationalCrossingSink__EVAL_17),
    ._EVAL_18(RationalCrossingSink__EVAL_18),
    ._EVAL_19(RationalCrossingSink__EVAL_19),
    ._EVAL_20(RationalCrossingSink__EVAL_20),
    ._EVAL_21(RationalCrossingSink__EVAL_21),
    ._EVAL_22(RationalCrossingSink__EVAL_22),
    ._EVAL_23(RationalCrossingSink__EVAL_23),
    ._EVAL_24(RationalCrossingSink__EVAL_24),
    ._EVAL_25(RationalCrossingSink__EVAL_25),
    ._EVAL_26(RationalCrossingSink__EVAL_26),
    ._EVAL_27(RationalCrossingSink__EVAL_27),
    ._EVAL_28(RationalCrossingSink__EVAL_28),
    ._EVAL_29(RationalCrossingSink__EVAL_29),
    ._EVAL_30(RationalCrossingSink__EVAL_30)
  );
  SiFive__EVAL_272 RationalCrossingSource_2 (
    ._EVAL(RationalCrossingSource_2__EVAL),
    ._EVAL_0(RationalCrossingSource_2__EVAL_0),
    ._EVAL_1(RationalCrossingSource_2__EVAL_1),
    ._EVAL_2(RationalCrossingSource_2__EVAL_2),
    ._EVAL_3(RationalCrossingSource_2__EVAL_3),
    ._EVAL_4(RationalCrossingSource_2__EVAL_4),
    ._EVAL_5(RationalCrossingSource_2__EVAL_5),
    ._EVAL_6(RationalCrossingSource_2__EVAL_6),
    ._EVAL_7(RationalCrossingSource_2__EVAL_7),
    ._EVAL_8(RationalCrossingSource_2__EVAL_8),
    ._EVAL_9(RationalCrossingSource_2__EVAL_9)
  );
  assign RationalCrossingSink__EVAL_2 = _EVAL_15;
  assign _EVAL_80 = RationalCrossingSource__EVAL_15;
  assign RationalCrossingSink__EVAL_24 = _EVAL_11;
  assign _EVAL_6 = RationalCrossingSource_1__EVAL_3;
  assign _EVAL_57 = RationalCrossingSource_2__EVAL_9;
  assign RationalCrossingSource_2__EVAL_7 = _EVAL_93;
  assign RationalCrossingSink__EVAL_5 = _EVAL_75;
  assign RationalCrossingSource_2__EVAL_1 = _EVAL_44;
  assign _EVAL_45 = RationalCrossingSink__EVAL_21;
  assign _EVAL_36 = RationalCrossingSource_1__EVAL_14;
  assign _EVAL_46 = RationalCrossingSource__EVAL_11;
  assign _EVAL_63 = RationalCrossingSource_1__EVAL_21;
  assign RationalCrossingSink_1__EVAL_8 = _EVAL_33;
  assign _EVAL_90 = RationalCrossingSink__EVAL_27;
  assign _EVAL_40 = RationalCrossingSource__EVAL_28;
  assign _EVAL_1 = RationalCrossingSource_1__EVAL_9;
  assign _EVAL_18 = RationalCrossingSink_1__EVAL_2;
  assign RationalCrossingSink_1__EVAL_11 = _EVAL_42;
  assign _EVAL_73 = RationalCrossingSink__EVAL_20;
  assign _EVAL_0 = RationalCrossingSource__EVAL_13;
  assign _EVAL_38 = RationalCrossingSink_1__EVAL_4;
  assign RationalCrossingSink__EVAL_13 = _EVAL_105;
  assign _EVAL_59 = RationalCrossingSource_2__EVAL_4;
  assign RationalCrossingSource__EVAL_24 = _EVAL_69;
  assign _EVAL_97 = RationalCrossingSource_1__EVAL_27;
  assign RationalCrossingSink__EVAL_4 = _EVAL_7;
  assign _EVAL_16 = RationalCrossingSource_2__EVAL;
  assign RationalCrossingSource__EVAL_14 = _EVAL_71;
  assign RationalCrossingSink_1__EVAL_7 = _EVAL_13;
  assign _EVAL_98 = RationalCrossingSource__EVAL_10;
  assign _EVAL_91 = RationalCrossingSink__EVAL_8;
  assign RationalCrossingSource_1__EVAL_20 = _EVAL_50;
  assign RationalCrossingSink__EVAL_15 = _EVAL_77;
  assign _EVAL_2 = RationalCrossingSource_1__EVAL_19;
  assign RationalCrossingSource__EVAL_27 = _EVAL_106;
  assign RationalCrossingSink__EVAL_11 = _EVAL_35;
  assign RationalCrossingSource__EVAL_2 = _EVAL_100;
  assign RationalCrossingSource_1__EVAL_22 = _EVAL_42;
  assign RationalCrossingSink__EVAL_30 = _EVAL_21;
  assign _EVAL_39 = RationalCrossingSource__EVAL_22;
  assign _EVAL_51 = RationalCrossingSource_1__EVAL_26;
  assign _EVAL_94 = RationalCrossingSource_1__EVAL_1;
  assign _EVAL_87 = RationalCrossingSink__EVAL_9;
  assign _EVAL_28 = RationalCrossingSource_1__EVAL_18;
  assign RationalCrossingSink__EVAL_0 = _EVAL_34;
  assign RationalCrossingSink_1__EVAL_12 = _EVAL_7;
  assign RationalCrossingSource__EVAL_0 = _EVAL_41;
  assign _EVAL_47 = RationalCrossingSource__EVAL_9;
  assign RationalCrossingSink__EVAL_25 = _EVAL_54;
  assign _EVAL_76 = RationalCrossingSink__EVAL_7;
  assign RationalCrossingSource_1__EVAL_11 = _EVAL_22;
  assign RationalCrossingSource_2__EVAL_6 = _EVAL_7;
  assign RationalCrossingSource_1__EVAL_24 = _EVAL_89;
  assign _EVAL_32 = RationalCrossingSource__EVAL_12;
  assign _EVAL_83 = RationalCrossingSink_1__EVAL_1;
  assign _EVAL_64 = RationalCrossingSource_1__EVAL;
  assign RationalCrossingSource_2__EVAL_2 = _EVAL_4;
  assign _EVAL_8 = RationalCrossingSource__EVAL_7;
  assign RationalCrossingSource__EVAL_17 = _EVAL_42;
  assign _EVAL_5 = RationalCrossingSource__EVAL_30;
  assign RationalCrossingSource_1__EVAL_4 = _EVAL_26;
  assign _EVAL = RationalCrossingSource_1__EVAL_23;
  assign _EVAL_53 = RationalCrossingSink__EVAL_3;
  assign RationalCrossingSource_1__EVAL_15 = _EVAL_7;
  assign _EVAL_72 = RationalCrossingSink__EVAL_19;
  assign RationalCrossingSink__EVAL_1 = _EVAL_66;
  assign RationalCrossingSink__EVAL_14 = _EVAL_101;
  assign RationalCrossingSink_1__EVAL_3 = _EVAL_24;
  assign _EVAL_37 = RationalCrossingSource__EVAL_18;
  assign RationalCrossingSource__EVAL_20 = _EVAL_78;
  assign _EVAL_95 = RationalCrossingSource_1__EVAL_0;
  assign RationalCrossingSource_1__EVAL_16 = _EVAL_82;
  assign RationalCrossingSource_1__EVAL_5 = _EVAL_56;
  assign _EVAL_25 = RationalCrossingSink__EVAL_17;
  assign _EVAL_99 = RationalCrossingSource__EVAL_29;
  assign _EVAL_43 = RationalCrossingSource_2__EVAL_5;
  assign RationalCrossingSource__EVAL_25 = _EVAL_29;
  assign _EVAL_85 = RationalCrossingSource__EVAL_3;
  assign _EVAL_31 = RationalCrossingSource__EVAL_8;
  assign RationalCrossingSink_1__EVAL = _EVAL_96;
  assign RationalCrossingSink__EVAL_10 = _EVAL_108;
  assign RationalCrossingSource_1__EVAL_8 = _EVAL_62;
  assign RationalCrossingSink__EVAL_16 = _EVAL_70;
  assign _EVAL_65 = RationalCrossingSink__EVAL_26;
  assign RationalCrossingSource_2__EVAL_8 = _EVAL_42;
  assign _EVAL_48 = RationalCrossingSource__EVAL;
  assign RationalCrossingSink__EVAL_22 = _EVAL_88;
  assign RationalCrossingSource__EVAL_16 = _EVAL_60;
  assign _EVAL_49 = RationalCrossingSink_1__EVAL_9;
  assign RationalCrossingSink_1__EVAL_10 = _EVAL_68;
  assign RationalCrossingSource_2__EVAL_0 = _EVAL_67;
  assign RationalCrossingSource_1__EVAL_7 = _EVAL_27;
  assign RationalCrossingSink__EVAL_6 = _EVAL_61;
  assign _EVAL_10 = RationalCrossingSink__EVAL_28;
  assign RationalCrossingSource__EVAL_4 = _EVAL_12;
  assign _EVAL_103 = RationalCrossingSource_1__EVAL_2;
  assign _EVAL_19 = RationalCrossingSource_1__EVAL_10;
  assign _EVAL_55 = RationalCrossingSource_2__EVAL_3;
  assign RationalCrossingSink__EVAL = _EVAL_107;
  assign RationalCrossingSource_1__EVAL_12 = _EVAL_104;
  assign _EVAL_58 = RationalCrossingSource_1__EVAL_25;
  assign _EVAL_20 = RationalCrossingSource_1__EVAL_13;
  assign _EVAL_9 = RationalCrossingSink_1__EVAL_0;
  assign RationalCrossingSink__EVAL_29 = _EVAL_3;
  assign RationalCrossingSink_1__EVAL_6 = _EVAL_52;
  assign RationalCrossingSource__EVAL_19 = _EVAL_23;
  assign RationalCrossingSink__EVAL_23 = _EVAL_102;
  assign RationalCrossingSink__EVAL_18 = _EVAL_42;
  assign _EVAL_30 = RationalCrossingSource__EVAL_6;
  assign RationalCrossingSource__EVAL_1 = _EVAL_7;
  assign _EVAL_92 = RationalCrossingSource_1__EVAL_17;
  assign RationalCrossingSink_1__EVAL_5 = _EVAL_86;
  assign RationalCrossingSource_1__EVAL_6 = _EVAL_17;
  assign _EVAL_79 = RationalCrossingSource__EVAL_26;
  assign RationalCrossingSink__EVAL_12 = _EVAL_84;
  assign _EVAL_14 = RationalCrossingSource__EVAL_23;
  assign _EVAL_81 = RationalCrossingSource__EVAL_5;
  assign RationalCrossingSource__EVAL_21 = _EVAL_74;
endmodule
