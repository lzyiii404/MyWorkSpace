//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_55_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_26;
  reg [31:0] _RAND_0;
  reg [1:0] _EVAL_47;
  reg [31:0] _RAND_1;
  reg  _EVAL_80;
  reg [31:0] _RAND_2;
  reg  _EVAL_90;
  reg [31:0] _RAND_3;
  reg  _EVAL_106;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_112;
  reg [31:0] _RAND_5;
  reg [3:0] _EVAL_133;
  reg [31:0] _RAND_6;
  reg [5:0] _EVAL_142;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_151;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_184;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_205;
  reg [31:0] _RAND_10;
  reg [5:0] _EVAL_274;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_276;
  reg [31:0] _RAND_12;
  reg [3:0] _EVAL_283;
  reg [31:0] _RAND_13;
  wire  _EVAL_265;
  wire [31:0] _EVAL_40;
  wire [32:0] _EVAL_194;
  wire  _EVAL_297;
  wire [31:0] _EVAL_71;
  wire [32:0] _EVAL_37;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_207;
  wire  _EVAL_141;
  wire  _EVAL_247;
  wire  _EVAL_239;
  wire  _EVAL_206;
  wire  _EVAL_291;
  wire  _EVAL_255;
  wire  _EVAL_219;
  wire [31:0] _EVAL_246;
  wire [32:0] _EVAL_270;
  wire [31:0] _EVAL_234;
  wire [32:0] _EVAL_91;
  wire [32:0] _EVAL_69;
  wire [32:0] _EVAL_52;
  wire  _EVAL_114;
  wire  _EVAL_64;
  wire  _EVAL_231;
  wire  _EVAL_168;
  wire  _EVAL_147;
  wire  _EVAL_182;
  wire  _EVAL_271;
  wire [31:0] _EVAL_235;
  wire [32:0] _EVAL_216;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_82;
  wire  _EVAL_214;
  wire [32:0] _EVAL_36;
  wire [32:0] _EVAL_158;
  wire  _EVAL_43;
  wire  _EVAL_242;
  wire  _EVAL_169;
  wire [32:0] _EVAL_289;
  wire [32:0] _EVAL_107;
  wire [32:0] _EVAL_27;
  wire  _EVAL_99;
  wire  _EVAL_252;
  wire [32:0] _EVAL_157;
  wire [32:0] _EVAL_46;
  wire  _EVAL_61;
  wire  _EVAL_58;
  wire [31:0] _EVAL_129;
  wire [32:0] _EVAL_211;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_108;
  wire  _EVAL_163;
  wire  _EVAL_17;
  wire [31:0] _EVAL_199;
  wire [32:0] _EVAL_266;
  wire [32:0] _EVAL_28;
  wire [32:0] _EVAL_115;
  wire  _EVAL_109;
  wire  _EVAL_128;
  wire  _EVAL_229;
  wire  _EVAL_227;
  wire  _EVAL_156;
  wire  _EVAL_19;
  wire  _EVAL_93;
  wire  _EVAL_179;
  wire  _EVAL_44;
  wire  _EVAL_264;
  wire  _EVAL_189;
  wire  _EVAL_237;
  wire  _EVAL_135;
  wire  _EVAL_224;
  wire  _EVAL_86;
  wire [1:0] _EVAL_200;
  wire [1:0] _EVAL_225;
  wire  _EVAL_118;
  wire  _EVAL_127;
  wire  _EVAL_191;
  wire  _EVAL_290;
  wire  _EVAL_20;
  wire  _EVAL_164;
  wire  _EVAL_134;
  wire  _EVAL_113;
  wire [22:0] _EVAL_195;
  wire [7:0] _EVAL_49;
  wire [7:0] _EVAL_212;
  wire [31:0] _EVAL_145;
  wire [31:0] _EVAL_153;
  wire  _EVAL_119;
  wire  _EVAL_137;
  wire  _EVAL_175;
  wire [31:0] _EVAL_176;
  wire [32:0] _EVAL_57;
  wire [32:0] _EVAL_97;
  wire [32:0] _EVAL_161;
  wire  _EVAL_240;
  wire  _EVAL_67;
  wire  _EVAL_60;
  wire  _EVAL_32;
  wire  _EVAL_16;
  wire  _EVAL_38;
  wire  _EVAL_122;
  wire  _EVAL_24;
  wire  _EVAL_102;
  wire  _EVAL_186;
  wire  _EVAL_250;
  wire  _EVAL_256;
  wire  _EVAL_117;
  wire  _EVAL_279;
  wire  _EVAL_209;
  wire  _EVAL_293;
  wire  _EVAL_166;
  wire  _EVAL_197;
  wire  _EVAL_146;
  wire  _EVAL_196;
  wire  _EVAL_73;
  wire  _EVAL_173;
  wire  _EVAL_59;
  wire  _EVAL_183;
  wire  _EVAL_50;
  wire  _EVAL_272;
  wire  _EVAL_103;
  wire  _EVAL_261;
  wire  _EVAL_138;
  wire  _EVAL_45;
  wire  _EVAL_143;
  wire [3:0] _EVAL_192;
  wire [3:0] _EVAL_81;
  wire [3:0] _EVAL_178;
  wire  _EVAL_204;
  wire  _EVAL_53;
  wire  _EVAL_213;
  wire  _EVAL_177;
  wire  _EVAL_268;
  wire [1:0] _EVAL_188;
  wire  _EVAL_66;
  wire  _EVAL_154;
  wire  _EVAL_125;
  wire  _EVAL_78;
  wire [1:0] _EVAL_273;
  wire  _EVAL_42;
  wire  _EVAL_22;
  wire  _EVAL_139;
  wire  _EVAL_35;
  wire  _EVAL_172;
  wire  _EVAL_136;
  wire  _EVAL_94;
  wire [22:0] _EVAL_126;
  wire [7:0] _EVAL_217;
  wire [7:0] _EVAL_121;
  wire [5:0] _EVAL_55;
  wire  _EVAL_187;
  wire  _EVAL_221;
  wire [5:0] _EVAL_244;
  wire  _EVAL_30;
  wire  _EVAL_111;
  wire  _EVAL_23;
  wire  _EVAL_248;
  wire  _EVAL_241;
  wire  _EVAL_124;
  wire  _EVAL_31;
  wire  _EVAL_34;
  wire  _EVAL_98;
  wire  _EVAL_101;
  wire  _EVAL_29;
  wire  _EVAL_243;
  wire  _EVAL_190;
  wire  _EVAL_77;
  wire  _EVAL_167;
  wire  _EVAL_292;
  wire  _EVAL_159;
  wire  _EVAL_170;
  wire  _EVAL_269;
  wire  _EVAL_155;
  wire  _EVAL_54;
  wire  _EVAL_132;
  wire [31:0] _EVAL_180;
  wire  _EVAL_120;
  wire  _EVAL_181;
  wire [5:0] _EVAL_25;
  wire  _EVAL_284;
  wire  _EVAL_294;
  wire  _EVAL_56;
  wire  _EVAL_33;
  wire  _EVAL_280;
  wire  _EVAL_236;
  wire  _EVAL_198;
  wire  _EVAL_65;
  wire  _EVAL_72;
  wire [5:0] _EVAL_249;
  wire [5:0] _EVAL_228;
  wire  _EVAL_257;
  wire  _EVAL_41;
  wire  _EVAL_149;
  wire  _EVAL_70;
  wire  _EVAL_286;
  wire  _EVAL_89;
  wire  _EVAL_203;
  wire  _EVAL_278;
  wire  _EVAL_185;
  wire  _EVAL_105;
  wire  _EVAL_87;
  wire  _EVAL_51;
  wire  _EVAL_275;
  wire  _EVAL_100;
  wire  _EVAL_123;
  wire  _EVAL_152;
  wire  _EVAL_74;
  wire  _EVAL_220;
  wire  _EVAL_63;
  wire  _EVAL_296;
  wire  _EVAL_232;
  wire  _EVAL_131;
  wire [5:0] _EVAL_18;
  wire  _EVAL_287;
  wire  _EVAL_174;
  wire  _EVAL_21;
  wire [3:0] _EVAL_208;
  wire  _EVAL_68;
  wire  _EVAL_193;
  wire  _EVAL_295;
  wire  _EVAL_165;
  wire  _EVAL_76;
  wire  _EVAL_222;
  wire  _EVAL_39;
  wire  _EVAL_263;
  wire  _EVAL_202;
  wire  _EVAL_233;
  wire  _EVAL_201;
  wire  _EVAL_226;
  wire  _EVAL_259;
  wire  _EVAL_288;
  wire  _EVAL_160;
  wire  _EVAL_85;
  wire  _EVAL_95;
  wire  _EVAL_223;
  wire  _EVAL_277;
  wire  _EVAL_62;
  wire  _EVAL_254;
  wire  _EVAL_260;
  wire  _EVAL_140;
  wire  _EVAL_116;
  wire  _EVAL_253;
  wire  _EVAL_251;
  wire  _EVAL_258;
  wire  _EVAL_92;
  wire  _EVAL_84;
  wire  _EVAL_110;
  wire  _EVAL_79;
  wire  _EVAL_245;
  wire  _EVAL_285;
  wire  _EVAL_48;
  wire  _EVAL_218;
  wire  _EVAL_215;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_265 = _EVAL_14 == _EVAL_276;
  assign _EVAL_40 = _EVAL_14 ^ 32'h1800000;
  assign _EVAL_194 = {1'b0,$signed(_EVAL_40)};
  assign _EVAL_297 = _EVAL_10 <= 4'h6;
  assign _EVAL_71 = _EVAL_14 ^ 32'h80000000;
  assign _EVAL_37 = {1'b0,$signed(_EVAL_71)};
  assign _EVAL_130 = $signed(_EVAL_37) & $signed(-33'sh20000);
  assign _EVAL_207 = $signed(_EVAL_130);
  assign _EVAL_141 = $signed(_EVAL_207) == $signed(33'sh0);
  assign _EVAL_247 = _EVAL_297 & _EVAL_141;
  assign _EVAL_239 = _EVAL_247 | _EVAL_6;
  assign _EVAL_206 = _EVAL_239 == 1'h0;
  assign _EVAL_291 = _EVAL_0 == _EVAL_90;
  assign _EVAL_255 = _EVAL_291 | _EVAL_6;
  assign _EVAL_219 = _EVAL_255 == 1'h0;
  assign _EVAL_246 = _EVAL_14 ^ 32'hc000000;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_246)};
  assign _EVAL_234 = _EVAL_14 ^ 32'h2000000;
  assign _EVAL_91 = {1'b0,$signed(_EVAL_234)};
  assign _EVAL_69 = $signed(_EVAL_91) & $signed(-33'sh10000);
  assign _EVAL_52 = $signed(_EVAL_69);
  assign _EVAL_114 = $signed(_EVAL_52) == $signed(33'sh0);
  assign _EVAL_64 = _EVAL_106 == 1'h0;
  assign _EVAL_231 = _EVAL_64 | _EVAL_6;
  assign _EVAL_168 = _EVAL_11 & _EVAL_9;
  assign _EVAL_147 = _EVAL_205 == 6'h0;
  assign _EVAL_182 = _EVAL_168 & _EVAL_147;
  assign _EVAL_271 = _EVAL_10 <= 4'h2;
  assign _EVAL_235 = _EVAL_14 ^ 32'h3000;
  assign _EVAL_216 = {1'b0,$signed(_EVAL_235)};
  assign _EVAL_150 = $signed(_EVAL_216) & $signed(-33'sh1000);
  assign _EVAL_82 = $signed(_EVAL_150);
  assign _EVAL_214 = $signed(_EVAL_82) == $signed(33'sh0);
  assign _EVAL_36 = $signed(_EVAL_270) & $signed(-33'sh4000000);
  assign _EVAL_158 = $signed(_EVAL_36);
  assign _EVAL_43 = $signed(_EVAL_158) == $signed(33'sh0);
  assign _EVAL_242 = _EVAL_214 | _EVAL_43;
  assign _EVAL_169 = _EVAL_242 | _EVAL_114;
  assign _EVAL_289 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_107 = $signed(_EVAL_289) & $signed(-33'sh5000);
  assign _EVAL_27 = $signed(_EVAL_107);
  assign _EVAL_99 = $signed(_EVAL_27) == $signed(33'sh0);
  assign _EVAL_252 = _EVAL_169 | _EVAL_99;
  assign _EVAL_157 = $signed(_EVAL_194) & $signed(-33'sh8000);
  assign _EVAL_46 = $signed(_EVAL_157);
  assign _EVAL_61 = $signed(_EVAL_46) == $signed(33'sh0);
  assign _EVAL_58 = _EVAL_252 | _EVAL_61;
  assign _EVAL_129 = _EVAL_14 ^ 32'h1900000;
  assign _EVAL_211 = {1'b0,$signed(_EVAL_129)};
  assign _EVAL_104 = $signed(_EVAL_211) & $signed(-33'sh2000);
  assign _EVAL_108 = $signed(_EVAL_104);
  assign _EVAL_163 = $signed(_EVAL_108) == $signed(33'sh0);
  assign _EVAL_17 = _EVAL_58 | _EVAL_163;
  assign _EVAL_199 = _EVAL_14 ^ 32'h20000000;
  assign _EVAL_266 = {1'b0,$signed(_EVAL_199)};
  assign _EVAL_28 = $signed(_EVAL_266) & $signed(-33'sh2000);
  assign _EVAL_115 = $signed(_EVAL_28);
  assign _EVAL_109 = $signed(_EVAL_115) == $signed(33'sh0);
  assign _EVAL_128 = _EVAL_17 | _EVAL_109;
  assign _EVAL_229 = _EVAL_271 & _EVAL_128;
  assign _EVAL_227 = _EVAL_229 | _EVAL_6;
  assign _EVAL_156 = _EVAL_227 == 1'h0;
  assign _EVAL_19 = _EVAL_274 == 6'h0;
  assign _EVAL_93 = _EVAL_14[1];
  assign _EVAL_179 = _EVAL_93 == 1'h0;
  assign _EVAL_44 = _EVAL_3 == 3'h6;
  assign _EVAL_264 = _EVAL_7 & _EVAL_44;
  assign _EVAL_189 = _EVAL_142 == 6'h0;
  assign _EVAL_237 = _EVAL_10 <= 4'h8;
  assign _EVAL_135 = _EVAL_237 & _EVAL_214;
  assign _EVAL_224 = _EVAL_10 >= 4'h2;
  assign _EVAL_86 = _EVAL_10[0];
  assign _EVAL_200 = 2'h1 << _EVAL_86;
  assign _EVAL_225 = _EVAL_200 | 2'h1;
  assign _EVAL_118 = _EVAL_225[1];
  assign _EVAL_127 = _EVAL_118 & _EVAL_93;
  assign _EVAL_191 = _EVAL_224 | _EVAL_127;
  assign _EVAL_290 = _EVAL_225[0];
  assign _EVAL_20 = _EVAL_14[0];
  assign _EVAL_164 = _EVAL_93 & _EVAL_20;
  assign _EVAL_134 = _EVAL_290 & _EVAL_164;
  assign _EVAL_113 = _EVAL_191 | _EVAL_134;
  assign _EVAL_195 = 23'hff << _EVAL_10;
  assign _EVAL_49 = _EVAL_195[7:0];
  assign _EVAL_212 = ~ _EVAL_49;
  assign _EVAL_145 = {{24'd0}, _EVAL_212};
  assign _EVAL_153 = _EVAL_14 & _EVAL_145;
  assign _EVAL_119 = _EVAL_153 == 32'h0;
  assign _EVAL_137 = _EVAL_119 | _EVAL_6;
  assign _EVAL_175 = _EVAL_137 == 1'h0;
  assign _EVAL_176 = _EVAL_14 ^ 32'h40000000;
  assign _EVAL_57 = {1'b0,$signed(_EVAL_176)};
  assign _EVAL_97 = $signed(_EVAL_57) & $signed(-33'sh2000);
  assign _EVAL_161 = $signed(_EVAL_97);
  assign _EVAL_240 = $signed(_EVAL_161) == $signed(33'sh0);
  assign _EVAL_67 = _EVAL_240 | _EVAL_141;
  assign _EVAL_60 = _EVAL_67 | _EVAL_43;
  assign _EVAL_32 = _EVAL_60 | _EVAL_114;
  assign _EVAL_16 = _EVAL_32 | _EVAL_99;
  assign _EVAL_38 = _EVAL_16 | _EVAL_61;
  assign _EVAL_122 = _EVAL_38 | _EVAL_163;
  assign _EVAL_24 = _EVAL_122 | _EVAL_109;
  assign _EVAL_102 = _EVAL_297 & _EVAL_24;
  assign _EVAL_186 = _EVAL_102 | _EVAL_135;
  assign _EVAL_250 = _EVAL_186 | _EVAL_6;
  assign _EVAL_256 = plusarg_reader_out == 32'h0;
  assign _EVAL_117 = _EVAL_64 | _EVAL_256;
  assign _EVAL_279 = _EVAL_26 < plusarg_reader_out;
  assign _EVAL_209 = _EVAL_117 | _EVAL_279;
  assign _EVAL_293 = _EVAL_209 | _EVAL_6;
  assign _EVAL_166 = _EVAL_293 == 1'h0;
  assign _EVAL_197 = _EVAL_0 == 1'h0;
  assign _EVAL_146 = _EVAL_197 | _EVAL_13;
  assign _EVAL_196 = _EVAL_20 == 1'h0;
  assign _EVAL_73 = _EVAL_93 & _EVAL_196;
  assign _EVAL_173 = _EVAL_290 & _EVAL_73;
  assign _EVAL_59 = _EVAL_191 | _EVAL_173;
  assign _EVAL_183 = _EVAL_118 & _EVAL_179;
  assign _EVAL_50 = _EVAL_224 | _EVAL_183;
  assign _EVAL_272 = _EVAL_179 & _EVAL_20;
  assign _EVAL_103 = _EVAL_290 & _EVAL_272;
  assign _EVAL_261 = _EVAL_50 | _EVAL_103;
  assign _EVAL_138 = _EVAL_179 & _EVAL_196;
  assign _EVAL_45 = _EVAL_290 & _EVAL_138;
  assign _EVAL_143 = _EVAL_50 | _EVAL_45;
  assign _EVAL_192 = {_EVAL_113,_EVAL_59,_EVAL_261,_EVAL_143};
  assign _EVAL_81 = ~ _EVAL_192;
  assign _EVAL_178 = _EVAL_12 & _EVAL_81;
  assign _EVAL_204 = _EVAL_10 == _EVAL_283;
  assign _EVAL_53 = _EVAL_204 | _EVAL_6;
  assign _EVAL_213 = _EVAL_8 & _EVAL_7;
  assign _EVAL_177 = _EVAL_184 == 6'h0;
  assign _EVAL_268 = _EVAL_213 & _EVAL_177;
  assign _EVAL_188 = _EVAL_268 ? 2'h1 : 2'h0;
  assign _EVAL_66 = _EVAL_188[0];
  assign _EVAL_154 = _EVAL_1 == 3'h6;
  assign _EVAL_125 = _EVAL_154 == 1'h0;
  assign _EVAL_78 = _EVAL_182 & _EVAL_125;
  assign _EVAL_273 = _EVAL_78 ? 2'h1 : 2'h0;
  assign _EVAL_42 = _EVAL_273[0];
  assign _EVAL_22 = _EVAL_66 != _EVAL_42;
  assign _EVAL_139 = _EVAL_66 == 1'h0;
  assign _EVAL_35 = _EVAL_22 | _EVAL_139;
  assign _EVAL_172 = _EVAL_35 | _EVAL_6;
  assign _EVAL_136 = _EVAL_172 == 1'h0;
  assign _EVAL_94 = _EVAL_1[0];
  assign _EVAL_126 = 23'hff << _EVAL_4;
  assign _EVAL_217 = _EVAL_126[7:0];
  assign _EVAL_121 = ~ _EVAL_217;
  assign _EVAL_55 = _EVAL_121[7:2];
  assign _EVAL_187 = _EVAL_1 == 3'h4;
  assign _EVAL_221 = _EVAL_9 & _EVAL_187;
  assign _EVAL_244 = _EVAL_205 - 6'h1;
  assign _EVAL_30 = _EVAL_9 & _EVAL_154;
  assign _EVAL_111 = _EVAL_2 != 2'h2;
  assign _EVAL_23 = _EVAL_111 | _EVAL_6;
  assign _EVAL_248 = _EVAL_23 == 1'h0;
  assign _EVAL_241 = _EVAL_3 == 3'h5;
  assign _EVAL_124 = _EVAL_4 == _EVAL_133;
  assign _EVAL_31 = _EVAL_124 | _EVAL_6;
  assign _EVAL_34 = _EVAL_31 == 1'h0;
  assign _EVAL_98 = _EVAL_3 == _EVAL_151;
  assign _EVAL_101 = _EVAL_98 | _EVAL_6;
  assign _EVAL_29 = _EVAL_101 == 1'h0;
  assign _EVAL_243 = _EVAL_3 == 3'h1;
  assign _EVAL_190 = _EVAL_7 & _EVAL_243;
  assign _EVAL_77 = _EVAL_1 == _EVAL_112;
  assign _EVAL_167 = _EVAL_77 | _EVAL_6;
  assign _EVAL_292 = _EVAL_3 == 3'h0;
  assign _EVAL_159 = _EVAL_7 & _EVAL_292;
  assign _EVAL_170 = _EVAL_4 >= 4'h2;
  assign _EVAL_269 = _EVAL_178 == 4'h0;
  assign _EVAL_155 = _EVAL_269 | _EVAL_6;
  assign _EVAL_54 = _EVAL_2 <= 2'h2;
  assign _EVAL_132 = _EVAL_54 | _EVAL_6;
  assign _EVAL_180 = _EVAL_26 + 32'h1;
  assign _EVAL_120 = _EVAL_265 | _EVAL_6;
  assign _EVAL_181 = _EVAL_120 == 1'h0;
  assign _EVAL_25 = _EVAL_184 - 6'h1;
  assign _EVAL_284 = _EVAL_106 | _EVAL_66;
  assign _EVAL_294 = ~ _EVAL_42;
  assign _EVAL_56 = _EVAL_284 & _EVAL_294;
  assign _EVAL_33 = _EVAL_19 == 1'h0;
  assign _EVAL_280 = _EVAL_9 & _EVAL_33;
  assign _EVAL_236 = _EVAL_3 == 3'h3;
  assign _EVAL_198 = _EVAL_7 & _EVAL_236;
  assign _EVAL_65 = _EVAL_3[2];
  assign _EVAL_72 = _EVAL_65 == 1'h0;
  assign _EVAL_249 = _EVAL_212[7:2];
  assign _EVAL_228 = _EVAL_142 - 6'h1;
  assign _EVAL_257 = _EVAL_146 | _EVAL_6;
  assign _EVAL_41 = _EVAL_3 == 3'h7;
  assign _EVAL_149 = _EVAL_7 & _EVAL_41;
  assign _EVAL_70 = _EVAL_170 | _EVAL_6;
  assign _EVAL_286 = _EVAL_70 == 1'h0;
  assign _EVAL_89 = _EVAL_7 & _EVAL_241;
  assign _EVAL_203 = _EVAL_168 & _EVAL_19;
  assign _EVAL_278 = _EVAL_155 == 1'h0;
  assign _EVAL_185 = _EVAL_1 == 3'h1;
  assign _EVAL_105 = _EVAL_9 & _EVAL_185;
  assign _EVAL_87 = _EVAL_6 == 1'h0;
  assign _EVAL_51 = _EVAL_2 == _EVAL_47;
  assign _EVAL_275 = _EVAL_51 | _EVAL_6;
  assign _EVAL_100 = _EVAL_275 == 1'h0;
  assign _EVAL_123 = _EVAL_167 == 1'h0;
  assign _EVAL_152 = _EVAL_213 & _EVAL_189;
  assign _EVAL_74 = _EVAL_1 <= 3'h6;
  assign _EVAL_220 = _EVAL_12 == _EVAL_192;
  assign _EVAL_63 = _EVAL_220 | _EVAL_6;
  assign _EVAL_296 = _EVAL_63 == 1'h0;
  assign _EVAL_232 = _EVAL_1 == 3'h5;
  assign _EVAL_131 = _EVAL_9 & _EVAL_232;
  assign _EVAL_18 = _EVAL_274 - 6'h1;
  assign _EVAL_287 = _EVAL_13 == 1'h0;
  assign _EVAL_174 = _EVAL_287 | _EVAL_6;
  assign _EVAL_21 = _EVAL_174 == 1'h0;
  assign _EVAL_208 = ~ _EVAL_12;
  assign _EVAL_68 = _EVAL_208 == 4'h0;
  assign _EVAL_193 = _EVAL_250 == 1'h0;
  assign _EVAL_295 = _EVAL_1 == 3'h0;
  assign _EVAL_165 = _EVAL_9 & _EVAL_295;
  assign _EVAL_76 = _EVAL_224 | _EVAL_6;
  assign _EVAL_222 = _EVAL_76 == 1'h0;
  assign _EVAL_39 = _EVAL_53 == 1'h0;
  assign _EVAL_263 = _EVAL_1 == 3'h2;
  assign _EVAL_202 = _EVAL_9 & _EVAL_263;
  assign _EVAL_233 = _EVAL_66 | _EVAL_106;
  assign _EVAL_201 = _EVAL_233 | _EVAL_6;
  assign _EVAL_226 = _EVAL_201 == 1'h0;
  assign _EVAL_259 = _EVAL_257 == 1'h0;
  assign _EVAL_288 = _EVAL_3 == 3'h4;
  assign _EVAL_160 = _EVAL_7 & _EVAL_288;
  assign _EVAL_85 = _EVAL_197 | _EVAL_6;
  assign _EVAL_95 = _EVAL_85 == 1'h0;
  assign _EVAL_223 = _EVAL_231 == 1'h0;
  assign _EVAL_277 = _EVAL_5 == _EVAL_80;
  assign _EVAL_62 = _EVAL_277 | _EVAL_6;
  assign _EVAL_254 = _EVAL_3 == 3'h2;
  assign _EVAL_260 = _EVAL_213 | _EVAL_168;
  assign _EVAL_140 = _EVAL_2 == 2'h0;
  assign _EVAL_116 = _EVAL_68 | _EVAL_6;
  assign _EVAL_253 = _EVAL_189 == 1'h0;
  assign _EVAL_251 = _EVAL_7 & _EVAL_253;
  assign _EVAL_258 = _EVAL_132 == 1'h0;
  assign _EVAL_92 = _EVAL_116 == 1'h0;
  assign _EVAL_84 = _EVAL_62 == 1'h0;
  assign _EVAL_110 = _EVAL_135 | _EVAL_6;
  assign _EVAL_79 = _EVAL_7 & _EVAL_254;
  assign _EVAL_245 = _EVAL_74 | _EVAL_6;
  assign _EVAL_285 = _EVAL_140 | _EVAL_6;
  assign _EVAL_48 = _EVAL_285 == 1'h0;
  assign _EVAL_218 = _EVAL_245 == 1'h0;
  assign _EVAL_215 = _EVAL_110 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_47 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_80 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_90 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_106 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_112 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_133 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_142 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_151 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_184 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_205 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_274 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_276 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_283 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_6) begin
      _EVAL_26 <= 32'h0;
    end else begin
      if (_EVAL_260) begin
        _EVAL_26 <= 32'h0;
      end else begin
        _EVAL_26 <= _EVAL_180;
      end
    end
    if (_EVAL_203) begin
      _EVAL_47 <= _EVAL_2;
    end
    if (_EVAL_203) begin
      _EVAL_80 <= _EVAL_5;
    end
    if (_EVAL_203) begin
      _EVAL_90 <= _EVAL_0;
    end
    if (_EVAL_6) begin
      _EVAL_106 <= 1'h0;
    end else begin
      _EVAL_106 <= _EVAL_56;
    end
    if (_EVAL_203) begin
      _EVAL_112 <= _EVAL_1;
    end
    if (_EVAL_203) begin
      _EVAL_133 <= _EVAL_4;
    end
    if (_EVAL_6) begin
      _EVAL_142 <= 6'h0;
    end else begin
      if (_EVAL_213) begin
        if (_EVAL_189) begin
          if (_EVAL_72) begin
            _EVAL_142 <= _EVAL_249;
          end else begin
            _EVAL_142 <= 6'h0;
          end
        end else begin
          _EVAL_142 <= _EVAL_228;
        end
      end
    end
    if (_EVAL_152) begin
      _EVAL_151 <= _EVAL_3;
    end
    if (_EVAL_6) begin
      _EVAL_184 <= 6'h0;
    end else begin
      if (_EVAL_213) begin
        if (_EVAL_177) begin
          if (_EVAL_72) begin
            _EVAL_184 <= _EVAL_249;
          end else begin
            _EVAL_184 <= 6'h0;
          end
        end else begin
          _EVAL_184 <= _EVAL_25;
        end
      end
    end
    if (_EVAL_6) begin
      _EVAL_205 <= 6'h0;
    end else begin
      if (_EVAL_168) begin
        if (_EVAL_147) begin
          if (_EVAL_94) begin
            _EVAL_205 <= _EVAL_55;
          end else begin
            _EVAL_205 <= 6'h0;
          end
        end else begin
          _EVAL_205 <= _EVAL_244;
        end
      end
    end
    if (_EVAL_6) begin
      _EVAL_274 <= 6'h0;
    end else begin
      if (_EVAL_168) begin
        if (_EVAL_19) begin
          if (_EVAL_94) begin
            _EVAL_274 <= _EVAL_55;
          end else begin
            _EVAL_274 <= 6'h0;
          end
        end else begin
          _EVAL_274 <= _EVAL_18;
        end
      end
    end
    if (_EVAL_152) begin
      _EVAL_276 <= _EVAL_14;
    end
    if (_EVAL_152) begin
      _EVAL_283 <= _EVAL_10;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95e9d07f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de5fb75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24b6391b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a52e9692)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff2f4e8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(914904b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a18274)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af9e2719)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ae13398)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fd58b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4908a73e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5653cfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(722ff522)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55b4a6be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eeeaea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a088dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfe0d95c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbf976fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc062825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93b2ddc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1a88ea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14046c46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(940d985)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23623c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11a4969f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aef5224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f090a66c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b8ec764)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57deab67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53e48445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3846b53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1a881fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b965e8f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e75eaf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de71977a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8454b83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2888a2d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e73eba88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb2ddbfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae93c6e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ce61f95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a7cdb85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9dce93c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(930bfb2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e85d929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3543dbb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a68f62de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95854ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c405d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a10a365d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfff346b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dc0031e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(654bea29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e33293f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7fb7cf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79d02293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8f4e96b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65bb7172)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcf67d29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fb2649)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
