//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_148_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [24:0] _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [6:0]  _EVAL_17,
  input  [6:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_58;
  reg [31:0] _RAND_0;
  reg [72:0] _EVAL_87;
  reg [95:0] _RAND_1;
  reg [24:0] _EVAL_94;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_97;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_98;
  reg [31:0] _RAND_4;
  reg [6:0] _EVAL_110;
  reg [31:0] _RAND_5;
  reg  _EVAL_164;
  reg [31:0] _RAND_6;
  reg [1:0] _EVAL_175;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_187;
  reg [31:0] _RAND_8;
  reg [6:0] _EVAL_196;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_199;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_212;
  reg [31:0] _RAND_11;
  reg [3:0] _EVAL_219;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_230;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_247;
  reg [31:0] _RAND_14;
  reg  _EVAL_271;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_272;
  reg [31:0] _RAND_16;
  wire [2:0] _EVAL_233;
  wire  _EVAL_99;
  wire  _EVAL_210;
  wire  _EVAL_317;
  wire [3:0] _EVAL_266;
  wire  _EVAL_72;
  wire  _EVAL_120;
  wire  _EVAL_45;
  wire  _EVAL_31;
  wire  _EVAL_328;
  wire [12:0] _EVAL_332;
  wire [3:0] _EVAL_284;
  wire  _EVAL_217;
  wire  _EVAL_198;
  wire  _EVAL_306;
  wire  _EVAL_270;
  wire  _EVAL_37;
  wire  _EVAL_65;
  wire  _EVAL_23;
  wire  _EVAL_150;
  wire  _EVAL_197;
  wire  _EVAL_229;
  wire  _EVAL_127;
  wire  _EVAL_308;
  wire  _EVAL_131;
  wire  _EVAL_203;
  wire  _EVAL_40;
  wire [127:0] _EVAL_243;
  wire [127:0] _EVAL_228;
  wire [72:0] _EVAL_81;
  wire [72:0] _EVAL_154;
  wire [72:0] _EVAL_141;
  wire  _EVAL_77;
  wire  _EVAL_255;
  wire  _EVAL_331;
  wire [1:0] _EVAL_290;
  wire [1:0] _EVAL_119;
  wire  _EVAL_237;
  wire [72:0] _EVAL_252;
  wire  _EVAL_100;
  wire [5:0] _EVAL_167;
  wire [5:0] _EVAL_78;
  wire  _EVAL_181;
  wire  _EVAL_310;
  wire  _EVAL_265;
  wire  _EVAL_121;
  wire  _EVAL_329;
  wire  _EVAL_33;
  wire  _EVAL_301;
  wire  _EVAL_137;
  wire  _EVAL_295;
  wire  _EVAL_244;
  wire  _EVAL_202;
  wire  _EVAL_263;
  wire  _EVAL_171;
  wire  _EVAL_83;
  wire [3:0] _EVAL_223;
  wire [3:0] _EVAL_103;
  wire  _EVAL_142;
  wire  _EVAL_236;
  wire  _EVAL_186;
  wire  _EVAL_231;
  wire  _EVAL_159;
  wire  _EVAL_279;
  wire  _EVAL_213;
  wire  _EVAL_89;
  wire  _EVAL_157;
  wire [3:0] _EVAL_122;
  wire  _EVAL_240;
  wire  _EVAL_124;
  wire [3:0] _EVAL_225;
  wire  _EVAL_273;
  wire  _EVAL_62;
  wire  _EVAL_205;
  wire  _EVAL_267;
  wire  _EVAL_262;
  wire  _EVAL_117;
  wire  _EVAL_126;
  wire [24:0] _EVAL_291;
  wire [25:0] _EVAL_115;
  wire [25:0] _EVAL_118;
  wire [25:0] _EVAL_74;
  wire  _EVAL_50;
  wire  _EVAL_38;
  wire  _EVAL_112;
  wire  _EVAL_315;
  wire  _EVAL_44;
  wire  _EVAL_52;
  wire  _EVAL_177;
  wire  _EVAL_153;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_285;
  wire [127:0] _EVAL_298;
  wire [127:0] _EVAL_313;
  wire [72:0] _EVAL_151;
  wire  _EVAL_275;
  wire  _EVAL_192;
  wire  _EVAL_302;
  wire  _EVAL_325;
  wire  _EVAL_46;
  wire [24:0] _EVAL_254;
  wire [25:0] _EVAL_54;
  wire [25:0] _EVAL_235;
  wire [25:0] _EVAL_80;
  wire  _EVAL_145;
  wire  _EVAL_114;
  wire  _EVAL_304;
  wire  _EVAL_85;
  wire  _EVAL_162;
  wire  _EVAL_91;
  wire  _EVAL_30;
  wire  _EVAL_278;
  wire  _EVAL_195;
  wire  _EVAL_220;
  wire  _EVAL_260;
  wire  _EVAL_297;
  wire  _EVAL_204;
  wire  _EVAL_253;
  wire  _EVAL_49;
  wire  _EVAL_241;
  wire  _EVAL_32;
  wire  _EVAL_289;
  wire  _EVAL_128;
  wire  _EVAL_173;
  wire  _EVAL_283;
  wire  _EVAL_19;
  wire  _EVAL_138;
  wire  _EVAL_152;
  wire [2:0] _EVAL_56;
  wire  _EVAL_327;
  wire  _EVAL_143;
  wire  _EVAL_206;
  wire  _EVAL_277;
  wire  _EVAL_51;
  wire  _EVAL_324;
  wire  _EVAL_43;
  wire  _EVAL_169;
  wire  _EVAL_84;
  wire  _EVAL_256;
  wire  _EVAL_268;
  wire  _EVAL_221;
  wire  _EVAL_147;
  wire  _EVAL_200;
  wire  _EVAL_39;
  wire  _EVAL_155;
  wire  _EVAL_48;
  wire  _EVAL_227;
  wire  _EVAL_184;
  wire  _EVAL_209;
  wire  _EVAL_264;
  wire [3:0] _EVAL_75;
  wire  _EVAL_148;
  wire  _EVAL_201;
  wire  _EVAL_276;
  wire  _EVAL_70;
  wire  _EVAL_165;
  wire  _EVAL_180;
  wire  _EVAL_320;
  wire  _EVAL_79;
  wire  _EVAL_73;
  wire  _EVAL_189;
  wire  _EVAL_34;
  wire  _EVAL_326;
  wire  _EVAL_149;
  wire  _EVAL_163;
  wire  _EVAL_96;
  wire  _EVAL_68;
  wire  _EVAL_288;
  wire  _EVAL_242;
  wire  _EVAL_67;
  wire  _EVAL_20;
  wire  _EVAL_222;
  wire  _EVAL_111;
  wire  _EVAL_211;
  wire  _EVAL_125;
  wire  _EVAL_214;
  wire  _EVAL_25;
  wire  _EVAL_269;
  wire [12:0] _EVAL_323;
  wire [5:0] _EVAL_322;
  wire [5:0] _EVAL_238;
  wire [3:0] _EVAL_274;
  wire  _EVAL_57;
  wire  _EVAL_286;
  wire  _EVAL_135;
  wire [24:0] _EVAL_105;
  wire [24:0] _EVAL_109;
  wire  _EVAL_41;
  wire  _EVAL_193;
  wire [3:0] _EVAL_282;
  wire  _EVAL_64;
  wire  _EVAL_224;
  wire  _EVAL_232;
  wire  _EVAL_249;
  wire  _EVAL_166;
  wire  _EVAL_71;
  wire  _EVAL_42;
  wire  _EVAL_129;
  wire  _EVAL_82;
  wire  _EVAL_136;
  wire  _EVAL_293;
  wire  _EVAL_296;
  wire [3:0] _EVAL_107;
  wire [3:0] _EVAL_226;
  wire [3:0] _EVAL_208;
  wire  _EVAL_146;
  wire  _EVAL_134;
  wire  _EVAL_95;
  wire  _EVAL_251;
  wire  _EVAL_101;
  wire  _EVAL_190;
  wire  _EVAL_144;
  wire  _EVAL_133;
  wire  _EVAL_104;
  wire  _EVAL_132;
  wire  _EVAL_287;
  wire  _EVAL_215;
  wire  _EVAL_330;
  wire  _EVAL_88;
  wire  _EVAL_170;
  wire  _EVAL_130;
  wire  _EVAL_218;
  wire  _EVAL_292;
  wire  _EVAL_257;
  wire  _EVAL_113;
  wire [72:0] _EVAL_280;
  wire  _EVAL_185;
  wire  _EVAL_311;
  wire  _EVAL_76;
  wire  _EVAL_108;
  wire  _EVAL_305;
  wire  _EVAL_36;
  wire [31:0] _EVAL_47;
  wire  _EVAL_281;
  wire  _EVAL_24;
  wire  _EVAL_248;
  wire  _EVAL_172;
  wire  _EVAL_60;
  wire  _EVAL_294;
  wire  _EVAL_21;
  wire  _EVAL_161;
  wire  _EVAL_250;
  wire  _EVAL_27;
  wire  _EVAL_299;
  wire  _EVAL_55;
  wire  _EVAL_312;
  wire  _EVAL_307;
  wire  _EVAL_174;
  wire  _EVAL_59;
  wire  _EVAL_92;
  wire  _EVAL_318;
  wire  _EVAL_194;
  wire  _EVAL_182;
  wire  _EVAL_160;
  wire  _EVAL_183;
  wire  _EVAL_28;
  wire  _EVAL_188;
  wire  _EVAL_245;
  wire  _EVAL_156;
  wire  _EVAL_63;
  wire  _EVAL_246;
  wire  _EVAL_178;
  wire  _EVAL_207;
  wire  _EVAL_66;
  wire  _EVAL_26;
  wire  _EVAL_303;
  wire  _EVAL_261;
  wire [72:0] _EVAL_300;
  wire  _EVAL_319;
  wire  _EVAL_158;
  wire  _EVAL_90;
  wire  _EVAL_258;
  wire  _EVAL_234;
  wire  _EVAL_86;
  wire  _EVAL_93;
  wire  _EVAL_22;
  wire [72:0] _EVAL_314;
  wire  _EVAL_123;
  wire  _EVAL_168;
  wire  _EVAL_116;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_233 = _EVAL_18[2:0];
  assign _EVAL_99 = _EVAL_219 == 4'h0;
  assign _EVAL_210 = _EVAL_99 == 1'h0;
  assign _EVAL_317 = _EVAL_9 & _EVAL_210;
  assign _EVAL_266 = _EVAL_17[6:3];
  assign _EVAL_72 = _EVAL_266 == 4'h0;
  assign _EVAL_120 = _EVAL_266 == 4'h3;
  assign _EVAL_45 = _EVAL_7[0];
  assign _EVAL_31 = _EVAL_45 == 1'h0;
  assign _EVAL_328 = _EVAL_10 == 3'h4;
  assign _EVAL_332 = 13'h3f << _EVAL_2;
  assign _EVAL_284 = ~ _EVAL_12;
  assign _EVAL_217 = _EVAL_284 == 4'h0;
  assign _EVAL_198 = _EVAL_15 == 1'h0;
  assign _EVAL_306 = _EVAL_198 | _EVAL_6;
  assign _EVAL_270 = _EVAL_306 == 1'h0;
  assign _EVAL_37 = _EVAL_5 == 3'h6;
  assign _EVAL_65 = _EVAL & _EVAL_37;
  assign _EVAL_23 = _EVAL_2 >= 3'h2;
  assign _EVAL_150 = _EVAL_23 | _EVAL_6;
  assign _EVAL_197 = _EVAL_14 <= 3'h2;
  assign _EVAL_229 = _EVAL_197 | _EVAL_6;
  assign _EVAL_127 = _EVAL_229 == 1'h0;
  assign _EVAL_308 = _EVAL_17 == 7'h48;
  assign _EVAL_131 = _EVAL_0 & _EVAL;
  assign _EVAL_203 = _EVAL_272 == 4'h0;
  assign _EVAL_40 = _EVAL_131 & _EVAL_203;
  assign _EVAL_243 = 128'h1 << _EVAL_18;
  assign _EVAL_228 = _EVAL_40 ? _EVAL_243 : 128'h0;
  assign _EVAL_81 = _EVAL_228[72:0];
  assign _EVAL_154 = _EVAL_81 | _EVAL_87;
  assign _EVAL_141 = _EVAL_154 >> _EVAL_17;
  assign _EVAL_77 = _EVAL_141[0];
  assign _EVAL_255 = _EVAL_77 | _EVAL_6;
  assign _EVAL_331 = _EVAL_13[0];
  assign _EVAL_290 = 2'h1 << _EVAL_331;
  assign _EVAL_119 = _EVAL_290 | 2'h1;
  assign _EVAL_237 = _EVAL_119[1];
  assign _EVAL_252 = _EVAL_87 >> _EVAL_18;
  assign _EVAL_100 = 3'h1 <= _EVAL_233;
  assign _EVAL_167 = _EVAL_332[5:0];
  assign _EVAL_78 = ~ _EVAL_167;
  assign _EVAL_181 = _EVAL_16 == _EVAL_164;
  assign _EVAL_310 = _EVAL_181 | _EVAL_6;
  assign _EVAL_265 = _EVAL_252[0];
  assign _EVAL_121 = _EVAL_265 == 1'h0;
  assign _EVAL_329 = _EVAL_121 | _EVAL_6;
  assign _EVAL_33 = _EVAL_329 == 1'h0;
  assign _EVAL_301 = _EVAL_4 == 1'h0;
  assign _EVAL_137 = _EVAL_301 | _EVAL_6;
  assign _EVAL_295 = _EVAL_137 == 1'h0;
  assign _EVAL_244 = _EVAL_98 == 4'h0;
  assign _EVAL_202 = _EVAL_1 & _EVAL_9;
  assign _EVAL_263 = _EVAL_187 == 4'h0;
  assign _EVAL_171 = _EVAL_202 & _EVAL_263;
  assign _EVAL_83 = _EVAL_10[0];
  assign _EVAL_223 = _EVAL_78[5:2];
  assign _EVAL_103 = _EVAL_187 - 4'h1;
  assign _EVAL_142 = _EVAL_18 == 7'h40;
  assign _EVAL_236 = 3'h6 == _EVAL_13;
  assign _EVAL_186 = _EVAL_142 ? _EVAL_236 : 1'h0;
  assign _EVAL_231 = _EVAL_186 | _EVAL_6;
  assign _EVAL_159 = _EVAL_119[0];
  assign _EVAL_279 = _EVAL_7[1];
  assign _EVAL_213 = _EVAL_279 == 1'h0;
  assign _EVAL_89 = _EVAL_213 & _EVAL_31;
  assign _EVAL_157 = _EVAL_159 & _EVAL_89;
  assign _EVAL_122 = _EVAL_219 - 4'h1;
  assign _EVAL_240 = _EVAL_10 == 3'h6;
  assign _EVAL_124 = _EVAL_9 & _EVAL_240;
  assign _EVAL_225 = _EVAL_18[6:3];
  assign _EVAL_273 = _EVAL_4 == _EVAL_271;
  assign _EVAL_62 = _EVAL_7 == _EVAL_94;
  assign _EVAL_205 = _EVAL_213 & _EVAL_45;
  assign _EVAL_267 = _EVAL_237 & _EVAL_213;
  assign _EVAL_262 = _EVAL_14 == _EVAL_247;
  assign _EVAL_117 = _EVAL_262 | _EVAL_6;
  assign _EVAL_126 = _EVAL_117 == 1'h0;
  assign _EVAL_291 = _EVAL_7 ^ 25'h1900000;
  assign _EVAL_115 = {1'b0,$signed(_EVAL_291)};
  assign _EVAL_118 = $signed(_EVAL_115) & $signed(-26'sh2000);
  assign _EVAL_74 = $signed(_EVAL_118);
  assign _EVAL_50 = $signed(_EVAL_74) == $signed(26'sh0);
  assign _EVAL_38 = _EVAL_5 == 3'h4;
  assign _EVAL_112 = _EVAL & _EVAL_38;
  assign _EVAL_315 = _EVAL_2 == _EVAL_97;
  assign _EVAL_44 = _EVAL_315 | _EVAL_6;
  assign _EVAL_52 = _EVAL_44 == 1'h0;
  assign _EVAL_177 = _EVAL_14 == 3'h0;
  assign _EVAL_153 = _EVAL_177 | _EVAL_6;
  assign _EVAL_139 = _EVAL_5 == 3'h1;
  assign _EVAL_140 = _EVAL_240 == 1'h0;
  assign _EVAL_285 = _EVAL_171 & _EVAL_140;
  assign _EVAL_298 = 128'h1 << _EVAL_17;
  assign _EVAL_313 = _EVAL_285 ? _EVAL_298 : 128'h0;
  assign _EVAL_151 = _EVAL_313[72:0];
  assign _EVAL_275 = _EVAL_13 >= 3'h2;
  assign _EVAL_192 = _EVAL_237 & _EVAL_279;
  assign _EVAL_302 = _EVAL_275 | _EVAL_192;
  assign _EVAL_325 = _EVAL_225 == 4'h1;
  assign _EVAL_46 = _EVAL_18 == 7'h48;
  assign _EVAL_254 = _EVAL_7 ^ 25'h1800000;
  assign _EVAL_54 = {1'b0,$signed(_EVAL_254)};
  assign _EVAL_235 = $signed(_EVAL_54) & $signed(-26'sh8000);
  assign _EVAL_80 = $signed(_EVAL_235);
  assign _EVAL_145 = $signed(_EVAL_80) == $signed(26'sh0);
  assign _EVAL_114 = _EVAL_46 | _EVAL_142;
  assign _EVAL_304 = _EVAL_225 == 4'h8;
  assign _EVAL_85 = _EVAL_304 & _EVAL_100;
  assign _EVAL_162 = _EVAL_114 | _EVAL_85;
  assign _EVAL_91 = _EVAL_18 == 7'h20;
  assign _EVAL_30 = _EVAL_162 | _EVAL_91;
  assign _EVAL_278 = _EVAL_225 == 4'h0;
  assign _EVAL_195 = _EVAL_30 | _EVAL_278;
  assign _EVAL_220 = _EVAL_195 | _EVAL_325;
  assign _EVAL_260 = _EVAL_5 == 3'h2;
  assign _EVAL_297 = _EVAL_10 == 3'h1;
  assign _EVAL_204 = _EVAL_8 == _EVAL_175;
  assign _EVAL_253 = _EVAL_204 | _EVAL_6;
  assign _EVAL_49 = _EVAL_253 == 1'h0;
  assign _EVAL_241 = _EVAL_301 | _EVAL_3;
  assign _EVAL_32 = _EVAL_241 | _EVAL_6;
  assign _EVAL_289 = _EVAL_32 == 1'h0;
  assign _EVAL_128 = _EVAL_14 != 3'h0;
  assign _EVAL_173 = _EVAL_10 == _EVAL_199;
  assign _EVAL_283 = _EVAL_173 | _EVAL_6;
  assign _EVAL_19 = _EVAL_17 == 7'h40;
  assign _EVAL_138 = _EVAL_308 | _EVAL_19;
  assign _EVAL_152 = _EVAL_266 == 4'h8;
  assign _EVAL_56 = _EVAL_17[2:0];
  assign _EVAL_327 = 3'h1 <= _EVAL_56;
  assign _EVAL_143 = _EVAL_152 & _EVAL_327;
  assign _EVAL_206 = _EVAL_138 | _EVAL_143;
  assign _EVAL_277 = _EVAL_17 == 7'h20;
  assign _EVAL_51 = _EVAL_206 | _EVAL_277;
  assign _EVAL_324 = _EVAL_275 | _EVAL_267;
  assign _EVAL_43 = _EVAL_283 == 1'h0;
  assign _EVAL_169 = _EVAL_51 | _EVAL_72;
  assign _EVAL_84 = _EVAL_266 == 4'h1;
  assign _EVAL_256 = _EVAL_169 | _EVAL_84;
  assign _EVAL_268 = _EVAL_266 == 4'h2;
  assign _EVAL_221 = _EVAL_256 | _EVAL_268;
  assign _EVAL_147 = _EVAL_279 & _EVAL_45;
  assign _EVAL_200 = _EVAL_159 & _EVAL_147;
  assign _EVAL_39 = _EVAL_302 | _EVAL_200;
  assign _EVAL_155 = _EVAL_279 & _EVAL_31;
  assign _EVAL_48 = _EVAL_159 & _EVAL_155;
  assign _EVAL_227 = _EVAL_302 | _EVAL_48;
  assign _EVAL_184 = _EVAL_159 & _EVAL_205;
  assign _EVAL_209 = _EVAL_324 | _EVAL_184;
  assign _EVAL_264 = _EVAL_324 | _EVAL_157;
  assign _EVAL_75 = {_EVAL_39,_EVAL_227,_EVAL_209,_EVAL_264};
  assign _EVAL_148 = _EVAL_12 == _EVAL_75;
  assign _EVAL_201 = _EVAL_148 | _EVAL_6;
  assign _EVAL_276 = _EVAL_201 == 1'h0;
  assign _EVAL_70 = _EVAL_18 == _EVAL_110;
  assign _EVAL_165 = _EVAL_70 | _EVAL_6;
  assign _EVAL_180 = _EVAL_165 == 1'h0;
  assign _EVAL_320 = _EVAL_13 == _EVAL_212;
  assign _EVAL_79 = _EVAL_320 | _EVAL_6;
  assign _EVAL_73 = _EVAL_231 == 1'h0;
  assign _EVAL_189 = _EVAL_10 == 3'h5;
  assign _EVAL_34 = _EVAL_9 & _EVAL_189;
  assign _EVAL_326 = _EVAL_5 == 3'h7;
  assign _EVAL_149 = _EVAL_10 == 3'h0;
  assign _EVAL_163 = _EVAL_9 & _EVAL_149;
  assign _EVAL_96 = _EVAL_145 | _EVAL_50;
  assign _EVAL_68 = _EVAL_225 == 4'h3;
  assign _EVAL_288 = _EVAL_153 == 1'h0;
  assign _EVAL_242 = _EVAL_5 == _EVAL_230;
  assign _EVAL_67 = _EVAL_242 | _EVAL_6;
  assign _EVAL_20 = _EVAL_13 <= 3'h6;
  assign _EVAL_222 = _EVAL_20 & _EVAL_96;
  assign _EVAL_111 = _EVAL_222 | _EVAL_6;
  assign _EVAL_211 = _EVAL_202 & _EVAL_99;
  assign _EVAL_125 = _EVAL_10 == 3'h2;
  assign _EVAL_214 = _EVAL_8 == 2'h0;
  assign _EVAL_25 = _EVAL_214 | _EVAL_6;
  assign _EVAL_269 = _EVAL_25 == 1'h0;
  assign _EVAL_323 = 13'h3f << _EVAL_13;
  assign _EVAL_322 = _EVAL_323[5:0];
  assign _EVAL_238 = ~ _EVAL_322;
  assign _EVAL_274 = _EVAL_238[5:2];
  assign _EVAL_57 = _EVAL_9 & _EVAL_328;
  assign _EVAL_286 = _EVAL_275 | _EVAL_6;
  assign _EVAL_135 = _EVAL & _EVAL_260;
  assign _EVAL_105 = {{19'd0}, _EVAL_238};
  assign _EVAL_109 = _EVAL_7 & _EVAL_105;
  assign _EVAL_41 = _EVAL_109 == 25'h0;
  assign _EVAL_193 = _EVAL_41 | _EVAL_6;
  assign _EVAL_282 = _EVAL_272 - 4'h1;
  assign _EVAL_64 = _EVAL_3 == 1'h0;
  assign _EVAL_224 = _EVAL_64 | _EVAL_6;
  assign _EVAL_232 = _EVAL_224 == 1'h0;
  assign _EVAL_249 = _EVAL_221 | _EVAL_120;
  assign _EVAL_166 = _EVAL_249 | _EVAL_6;
  assign _EVAL_71 = _EVAL_8 <= 2'h2;
  assign _EVAL_42 = _EVAL_71 | _EVAL_6;
  assign _EVAL_129 = _EVAL_42 == 1'h0;
  assign _EVAL_82 = _EVAL_5[2];
  assign _EVAL_136 = _EVAL_82 == 1'h0;
  assign _EVAL_293 = _EVAL_10 <= 3'h6;
  assign _EVAL_296 = _EVAL_293 | _EVAL_6;
  assign _EVAL_107 = _EVAL_98 - 4'h1;
  assign _EVAL_226 = ~ _EVAL_75;
  assign _EVAL_208 = _EVAL_12 & _EVAL_226;
  assign _EVAL_146 = _EVAL_208 == 4'h0;
  assign _EVAL_134 = _EVAL_81 != 73'h0;
  assign _EVAL_95 = _EVAL & _EVAL_139;
  assign _EVAL_251 = _EVAL_8 != 2'h2;
  assign _EVAL_101 = _EVAL_251 | _EVAL_6;
  assign _EVAL_190 = _EVAL_14 <= 3'h3;
  assign _EVAL_144 = _EVAL_190 | _EVAL_6;
  assign _EVAL_133 = _EVAL_58 < plusarg_reader_out;
  assign _EVAL_104 = _EVAL_5 == 3'h3;
  assign _EVAL_132 = _EVAL & _EVAL_104;
  assign _EVAL_287 = _EVAL_87 != 73'h0;
  assign _EVAL_215 = _EVAL_287 == 1'h0;
  assign _EVAL_330 = plusarg_reader_out == 32'h0;
  assign _EVAL_88 = _EVAL_215 | _EVAL_330;
  assign _EVAL_170 = _EVAL_88 | _EVAL_133;
  assign _EVAL_130 = _EVAL_170 | _EVAL_6;
  assign _EVAL_218 = _EVAL_17 == _EVAL_196;
  assign _EVAL_292 = _EVAL_218 | _EVAL_6;
  assign _EVAL_257 = _EVAL_292 == 1'h0;
  assign _EVAL_113 = _EVAL_5 == 3'h0;
  assign _EVAL_280 = _EVAL_87 | _EVAL_81;
  assign _EVAL_185 = _EVAL_146 | _EVAL_6;
  assign _EVAL_311 = _EVAL_185 == 1'h0;
  assign _EVAL_76 = _EVAL_286 == 1'h0;
  assign _EVAL_108 = _EVAL_128 | _EVAL_6;
  assign _EVAL_305 = _EVAL_108 == 1'h0;
  assign _EVAL_36 = _EVAL_131 & _EVAL_244;
  assign _EVAL_47 = _EVAL_58 + 32'h1;
  assign _EVAL_281 = _EVAL_244 == 1'h0;
  assign _EVAL_24 = _EVAL & _EVAL_281;
  assign _EVAL_248 = _EVAL_111 == 1'h0;
  assign _EVAL_172 = _EVAL_296 == 1'h0;
  assign _EVAL_60 = _EVAL_225 == 4'h2;
  assign _EVAL_294 = _EVAL_220 | _EVAL_60;
  assign _EVAL_21 = _EVAL_5 == 3'h5;
  assign _EVAL_161 = _EVAL_131 | _EVAL_202;
  assign _EVAL_250 = _EVAL_81 != _EVAL_151;
  assign _EVAL_27 = _EVAL_144 == 1'h0;
  assign _EVAL_299 = _EVAL_217 | _EVAL_6;
  assign _EVAL_55 = _EVAL_299 == 1'h0;
  assign _EVAL_312 = _EVAL_294 | _EVAL_68;
  assign _EVAL_307 = _EVAL_310 == 1'h0;
  assign _EVAL_174 = _EVAL_14 <= 3'h4;
  assign _EVAL_59 = _EVAL_174 | _EVAL_6;
  assign _EVAL_92 = _EVAL_101 == 1'h0;
  assign _EVAL_318 = _EVAL_134 == 1'h0;
  assign _EVAL_194 = _EVAL_250 | _EVAL_318;
  assign _EVAL_182 = _EVAL_194 | _EVAL_6;
  assign _EVAL_160 = _EVAL_182 == 1'h0;
  assign _EVAL_183 = _EVAL_59 == 1'h0;
  assign _EVAL_28 = _EVAL_166 == 1'h0;
  assign _EVAL_188 = _EVAL_79 == 1'h0;
  assign _EVAL_245 = _EVAL & _EVAL_326;
  assign _EVAL_156 = _EVAL & _EVAL_113;
  assign _EVAL_63 = _EVAL_312 | _EVAL_6;
  assign _EVAL_246 = _EVAL_62 | _EVAL_6;
  assign _EVAL_178 = _EVAL_246 == 1'h0;
  assign _EVAL_207 = _EVAL_193 == 1'h0;
  assign _EVAL_66 = _EVAL_255 == 1'h0;
  assign _EVAL_26 = _EVAL_63 == 1'h0;
  assign _EVAL_303 = _EVAL_150 == 1'h0;
  assign _EVAL_261 = _EVAL_9 & _EVAL_125;
  assign _EVAL_300 = ~ _EVAL_151;
  assign _EVAL_319 = _EVAL & _EVAL_21;
  assign _EVAL_158 = _EVAL_13 <= 3'h2;
  assign _EVAL_90 = _EVAL_158 & _EVAL_50;
  assign _EVAL_258 = _EVAL_90 | _EVAL_6;
  assign _EVAL_234 = _EVAL_6 == 1'h0;
  assign _EVAL_86 = _EVAL_273 | _EVAL_6;
  assign _EVAL_93 = _EVAL_67 == 1'h0;
  assign _EVAL_22 = _EVAL_86 == 1'h0;
  assign _EVAL_314 = _EVAL_280 & _EVAL_300;
  assign _EVAL_123 = _EVAL_9 & _EVAL_297;
  assign _EVAL_168 = _EVAL_258 == 1'h0;
  assign _EVAL_116 = _EVAL_130 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_58 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _EVAL_87 = _RAND_1[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_94 = _RAND_2[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_97 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_98 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_110 = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_164 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_175 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_187 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_196 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_199 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_212 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_219 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_230 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_247 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_271 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_272 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_11) begin
    if (_EVAL_6) begin
      _EVAL_58 <= 32'h0;
    end else begin
      if (_EVAL_161) begin
        _EVAL_58 <= 32'h0;
      end else begin
        _EVAL_58 <= _EVAL_47;
      end
    end
    if (_EVAL_6) begin
      _EVAL_87 <= 73'h0;
    end else begin
      _EVAL_87 <= _EVAL_314;
    end
    if (_EVAL_36) begin
      _EVAL_94 <= _EVAL_7;
    end
    if (_EVAL_211) begin
      _EVAL_97 <= _EVAL_2;
    end
    if (_EVAL_6) begin
      _EVAL_98 <= 4'h0;
    end else begin
      if (_EVAL_131) begin
        if (_EVAL_244) begin
          if (_EVAL_136) begin
            _EVAL_98 <= _EVAL_274;
          end else begin
            _EVAL_98 <= 4'h0;
          end
        end else begin
          _EVAL_98 <= _EVAL_107;
        end
      end
    end
    if (_EVAL_36) begin
      _EVAL_110 <= _EVAL_18;
    end
    if (_EVAL_211) begin
      _EVAL_164 <= _EVAL_16;
    end
    if (_EVAL_211) begin
      _EVAL_175 <= _EVAL_8;
    end
    if (_EVAL_6) begin
      _EVAL_187 <= 4'h0;
    end else begin
      if (_EVAL_202) begin
        if (_EVAL_263) begin
          if (_EVAL_83) begin
            _EVAL_187 <= _EVAL_223;
          end else begin
            _EVAL_187 <= 4'h0;
          end
        end else begin
          _EVAL_187 <= _EVAL_103;
        end
      end
    end
    if (_EVAL_211) begin
      _EVAL_196 <= _EVAL_17;
    end
    if (_EVAL_211) begin
      _EVAL_199 <= _EVAL_10;
    end
    if (_EVAL_36) begin
      _EVAL_212 <= _EVAL_13;
    end
    if (_EVAL_6) begin
      _EVAL_219 <= 4'h0;
    end else begin
      if (_EVAL_202) begin
        if (_EVAL_99) begin
          if (_EVAL_83) begin
            _EVAL_219 <= _EVAL_223;
          end else begin
            _EVAL_219 <= 4'h0;
          end
        end else begin
          _EVAL_219 <= _EVAL_122;
        end
      end
    end
    if (_EVAL_36) begin
      _EVAL_230 <= _EVAL_5;
    end
    if (_EVAL_36) begin
      _EVAL_247 <= _EVAL_14;
    end
    if (_EVAL_211) begin
      _EVAL_271 <= _EVAL_4;
    end
    if (_EVAL_6) begin
      _EVAL_272 <= 4'h0;
    end else begin
      if (_EVAL_131) begin
        if (_EVAL_203) begin
          if (_EVAL_136) begin
            _EVAL_272 <= _EVAL_274;
          end else begin
            _EVAL_272 <= 4'h0;
          end
        end else begin
          _EVAL_272 <= _EVAL_282;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(900d8f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78e4708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb58796b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f08e778)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7a0e97b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e26c1521)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62fa97ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37a930b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5fb7687)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93b44785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42775c86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40172fba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5098de0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b893664)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4d18eeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f7d0ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ea80fb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60a3085e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc50c033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd8327df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9da6f7f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd36a0ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9488be2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4564e862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97376226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1095087b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb9c92c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28a6271d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8250cfad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78f3c8ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d04a1682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ec6c09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f594552)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(731c267d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13bb53b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c84e5e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a71d8963)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6607e5bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae04f495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b161441a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57715daf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67e45a31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5104d01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9346153a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d72030)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c93aa4b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(535879f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea2e5f5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(491243ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d61ebd59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bca0c8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(677c8bc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f214e06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d531d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f140984)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(119e7d7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(447052b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(964debb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64b8b9df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57f529fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(797331cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dae68f70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(550997c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ea2f406)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c905613e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3442cf59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a14748d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b47cd8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(815b2e65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41978167)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9869586d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d775b7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61081fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7da68dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7567ddc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e510f11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db63fb20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fb7a9c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5fe6894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a49409a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea848012)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2448be5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2378f270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f48d6cf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(682a0470)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7baaeaf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df195cc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66d531c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86eea0df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff60c09c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(395adcb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87dd01ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(442f234b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53e91ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d05ae034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
