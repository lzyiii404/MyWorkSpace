//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_196_assert(
  input        _EVAL,
  input        _EVAL_0,
  input  [1:0] _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input        _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8,
  input  [3:0] _EVAL_9,
  input  [2:0] _EVAL_10,
  input  [8:0] _EVAL_11,
  input  [2:0] _EVAL_12,
  input        _EVAL_13,
  input  [1:0] _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_22;
  reg [31:0] _RAND_0;
  reg  _EVAL_26;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_27;
  reg [31:0] _RAND_2;
  reg  _EVAL_47;
  reg [31:0] _RAND_3;
  reg [8:0] _EVAL_59;
  reg [31:0] _RAND_4;
  reg  _EVAL_96;
  reg [31:0] _RAND_5;
  reg [1:0] _EVAL_100;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_128;
  reg [31:0] _RAND_7;
  reg  _EVAL_137;
  reg [31:0] _RAND_8;
  reg  _EVAL_138;
  reg [31:0] _RAND_9;
  reg  _EVAL_154;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_166;
  reg [31:0] _RAND_11;
  reg  _EVAL_198;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_210;
  reg [31:0] _RAND_13;
  wire  _EVAL_169;
  wire  _EVAL_109;
  wire  _EVAL_126;
  wire  _EVAL_200;
  wire [8:0] _EVAL_66;
  wire [9:0] _EVAL_212;
  wire [9:0] _EVAL_55;
  wire [9:0] _EVAL_120;
  wire [8:0] _EVAL_181;
  wire [9:0] _EVAL_153;
  wire  _EVAL_53;
  wire  _EVAL_165;
  wire  _EVAL_60;
  wire [8:0] _EVAL_88;
  wire [9:0] _EVAL_167;
  wire  _EVAL_83;
  wire [8:0] _EVAL_106;
  wire [9:0] _EVAL_49;
  wire [9:0] _EVAL_84;
  wire [9:0] _EVAL_168;
  wire  _EVAL_51;
  wire  _EVAL_97;
  wire  _EVAL_73;
  wire  _EVAL_40;
  wire  _EVAL_18;
  wire  _EVAL_107;
  wire  _EVAL_91;
  wire  _EVAL_104;
  wire [1:0] _EVAL_194;
  wire  _EVAL_216;
  wire  _EVAL_180;
  wire [9:0] _EVAL_102;
  wire [9:0] _EVAL_130;
  wire  _EVAL_95;
  wire  _EVAL_150;
  wire [3:0] _EVAL_58;
  wire  _EVAL_25;
  wire  _EVAL_121;
  wire  _EVAL_193;
  wire  _EVAL_75;
  wire  _EVAL_131;
  wire  _EVAL_206;
  wire  _EVAL_72;
  wire  _EVAL_70;
  wire  _EVAL_151;
  wire  _EVAL_119;
  wire  _EVAL_20;
  wire  _EVAL_108;
  wire  _EVAL_33;
  wire  _EVAL_175;
  wire  _EVAL_207;
  wire  _EVAL_144;
  wire  _EVAL_172;
  wire  _EVAL_162;
  wire  _EVAL_99;
  wire  _EVAL_39;
  wire  _EVAL_15;
  wire  _EVAL_57;
  wire  _EVAL_134;
  wire  _EVAL_182;
  wire [1:0] _EVAL_203;
  wire [9:0] _EVAL_63;
  wire [9:0] _EVAL_202;
  wire  _EVAL_184;
  wire  _EVAL_110;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_48;
  wire  _EVAL_118;
  wire  _EVAL_146;
  wire [1:0] _EVAL_103;
  wire  _EVAL_142;
  wire  _EVAL_129;
  wire  _EVAL_204;
  wire  _EVAL_38;
  wire  _EVAL_78;
  wire [8:0] _EVAL_67;
  wire [9:0] _EVAL_141;
  wire [9:0] _EVAL_89;
  wire [31:0] _EVAL_29;
  wire [9:0] _EVAL_179;
  wire [9:0] _EVAL_116;
  wire  _EVAL_201;
  wire  _EVAL_173;
  wire  _EVAL_136;
  wire  _EVAL_90;
  wire  _EVAL_35;
  wire  _EVAL_214;
  wire  _EVAL_105;
  wire  _EVAL_30;
  wire  _EVAL_186;
  wire  _EVAL_195;
  wire  _EVAL_24;
  wire [9:0] _EVAL_133;
  wire  _EVAL_43;
  wire  _EVAL_147;
  wire  _EVAL_76;
  wire  _EVAL_113;
  wire  _EVAL_125;
  wire [8:0] _EVAL_170;
  wire  _EVAL_46;
  wire  _EVAL_19;
  wire  _EVAL_161;
  wire  _EVAL_117;
  wire  _EVAL_44;
  wire  _EVAL_187;
  wire  _EVAL_163;
  wire  _EVAL_211;
  wire  _EVAL_171;
  wire  _EVAL_188;
  wire  _EVAL_196;
  wire  _EVAL_189;
  wire  _EVAL_215;
  wire  _EVAL_16;
  wire  _EVAL_139;
  wire  _EVAL_82;
  wire  _EVAL_37;
  wire  _EVAL_71;
  wire  _EVAL_23;
  wire  _EVAL_80;
  wire  _EVAL_77;
  wire  _EVAL_32;
  wire  _EVAL_122;
  wire  _EVAL_56;
  wire  _EVAL_152;
  wire  _EVAL_101;
  wire  _EVAL_68;
  wire  _EVAL_65;
  wire  _EVAL_94;
  wire  _EVAL_155;
  wire  _EVAL_50;
  wire [9:0] _EVAL_114;
  wire  _EVAL_124;
  wire  _EVAL_17;
  wire  _EVAL_36;
  wire  _EVAL_69;
  wire  _EVAL_111;
  wire  _EVAL_190;
  wire  _EVAL_205;
  wire  _EVAL_176;
  wire  _EVAL_199;
  wire  _EVAL_164;
  wire  _EVAL_178;
  wire  _EVAL_143;
  wire  _EVAL_34;
  wire  _EVAL_174;
  wire  _EVAL_115;
  wire  _EVAL_209;
  wire  _EVAL_45;
  wire  _EVAL_92;
  wire  _EVAL_213;
  wire  _EVAL_28;
  wire  _EVAL_93;
  wire  _EVAL_149;
  wire  _EVAL_160;
  wire  _EVAL_123;
  wire  _EVAL_52;
  wire  _EVAL_62;
  wire  _EVAL_31;
  wire  _EVAL_135;
  wire  _EVAL_157;
  wire  _EVAL_145;
  wire  _EVAL_192;
  wire  _EVAL_148;
  wire  _EVAL_183;
  wire  _EVAL_112;
  wire  _EVAL_217;
  wire  _EVAL_21;
  wire  _EVAL_191;
  wire  _EVAL_54;
  wire  _EVAL_64;
  wire  _EVAL_79;
  wire  _EVAL_140;
  wire  _EVAL_156;
  wire  _EVAL_74;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_169 = _EVAL_26 == 1'h0;
  assign _EVAL_109 = _EVAL_169 == 1'h0;
  assign _EVAL_126 = _EVAL_12 == 3'h0;
  assign _EVAL_200 = _EVAL_5 & _EVAL_126;
  assign _EVAL_66 = _EVAL_11 ^ 9'h44;
  assign _EVAL_212 = {1'b0,$signed(_EVAL_66)};
  assign _EVAL_55 = $signed(_EVAL_212) & $signed(-10'sh4);
  assign _EVAL_120 = $signed(_EVAL_55);
  assign _EVAL_181 = _EVAL_11 ^ 9'h60;
  assign _EVAL_153 = {1'b0,$signed(_EVAL_181)};
  assign _EVAL_53 = _EVAL_6 & _EVAL_2;
  assign _EVAL_165 = _EVAL_137 == 1'h0;
  assign _EVAL_60 = _EVAL_137 - 1'h1;
  assign _EVAL_88 = _EVAL_11 ^ 9'h48;
  assign _EVAL_167 = {1'b0,$signed(_EVAL_88)};
  assign _EVAL_83 = _EVAL_12 == _EVAL_27;
  assign _EVAL_106 = _EVAL_11 ^ 9'h100;
  assign _EVAL_49 = {1'b0,$signed(_EVAL_106)};
  assign _EVAL_84 = $signed(_EVAL_49) & $signed(-10'sh100);
  assign _EVAL_168 = $signed(_EVAL_84);
  assign _EVAL_51 = _EVAL_1 == _EVAL_100;
  assign _EVAL_97 = _EVAL_51 | _EVAL_8;
  assign _EVAL_73 = _EVAL_97 == 1'h0;
  assign _EVAL_40 = _EVAL_12 == 3'h7;
  assign _EVAL_18 = _EVAL_5 & _EVAL_40;
  assign _EVAL_107 = _EVAL_4 & _EVAL_5;
  assign _EVAL_91 = _EVAL_138 == 1'h0;
  assign _EVAL_104 = _EVAL_107 & _EVAL_91;
  assign _EVAL_194 = _EVAL_104 ? 2'h1 : 2'h0;
  assign _EVAL_216 = _EVAL_0 == _EVAL_47;
  assign _EVAL_180 = _EVAL_216 | _EVAL_8;
  assign _EVAL_102 = {1'b0,$signed(_EVAL_11)};
  assign _EVAL_130 = $signed(_EVAL_102) & $signed(-10'sh40);
  assign _EVAL_95 = _EVAL_53 & _EVAL_165;
  assign _EVAL_150 = plusarg_reader_out == 32'h0;
  assign _EVAL_58 = ~ _EVAL_9;
  assign _EVAL_25 = _EVAL_58 == 4'h0;
  assign _EVAL_121 = _EVAL_25 | _EVAL_8;
  assign _EVAL_193 = _EVAL == _EVAL_198;
  assign _EVAL_75 = _EVAL_26 - 1'h1;
  assign _EVAL_131 = _EVAL_12 == 3'h6;
  assign _EVAL_206 = _EVAL_138 - 1'h1;
  assign _EVAL_72 = _EVAL_12 == 3'h5;
  assign _EVAL_70 = _EVAL_14 <= 2'h2;
  assign _EVAL_151 = _EVAL_70 | _EVAL_8;
  assign _EVAL_119 = _EVAL_7 == 1'h0;
  assign _EVAL_20 = _EVAL_119 | _EVAL_8;
  assign _EVAL_108 = _EVAL_0 == 1'h0;
  assign _EVAL_33 = _EVAL_108 | _EVAL_13;
  assign _EVAL_175 = _EVAL_33 | _EVAL_8;
  assign _EVAL_207 = _EVAL_12 == 3'h3;
  assign _EVAL_144 = _EVAL_9 == 4'hf;
  assign _EVAL_172 = _EVAL_144 | _EVAL_8;
  assign _EVAL_162 = _EVAL_172 == 1'h0;
  assign _EVAL_99 = $signed(_EVAL_168) == $signed(10'sh0);
  assign _EVAL_39 = _EVAL_107 | _EVAL_53;
  assign _EVAL_15 = _EVAL_194[0];
  assign _EVAL_57 = _EVAL_22 | _EVAL_15;
  assign _EVAL_134 = _EVAL_20 == 1'h0;
  assign _EVAL_182 = _EVAL_1 >= 2'h2;
  assign _EVAL_203 = 2'h1 << _EVAL_7;
  assign _EVAL_63 = $signed(_EVAL_153) & $signed(-10'sh20);
  assign _EVAL_202 = $signed(_EVAL_63);
  assign _EVAL_184 = $signed(_EVAL_202) == $signed(10'sh0);
  assign _EVAL_110 = _EVAL_12 == 3'h4;
  assign _EVAL_86 = _EVAL_10 == 3'h0;
  assign _EVAL_87 = _EVAL_182 | _EVAL_8;
  assign _EVAL_48 = _EVAL_10 == 3'h6;
  assign _EVAL_118 = _EVAL_48 == 1'h0;
  assign _EVAL_146 = _EVAL_95 & _EVAL_118;
  assign _EVAL_103 = _EVAL_146 ? _EVAL_203 : 2'h0;
  assign _EVAL_142 = _EVAL_103[0];
  assign _EVAL_129 = _EVAL_15 != _EVAL_142;
  assign _EVAL_204 = _EVAL_15 == 1'h0;
  assign _EVAL_38 = _EVAL_129 | _EVAL_204;
  assign _EVAL_78 = _EVAL_38 | _EVAL_8;
  assign _EVAL_67 = _EVAL_11 ^ 9'h80;
  assign _EVAL_141 = {1'b0,$signed(_EVAL_67)};
  assign _EVAL_89 = $signed(_EVAL_141) & $signed(-10'sh80);
  assign _EVAL_29 = _EVAL_166 + 32'h1;
  assign _EVAL_179 = $signed(_EVAL_167) & $signed(-10'sh18);
  assign _EVAL_116 = $signed(_EVAL_179);
  assign _EVAL_201 = $signed(_EVAL_116) == $signed(10'sh0);
  assign _EVAL_173 = _EVAL_13 == 1'h0;
  assign _EVAL_136 = _EVAL_173 | _EVAL_8;
  assign _EVAL_90 = _EVAL_193 | _EVAL_8;
  assign _EVAL_35 = _EVAL_175 == 1'h0;
  assign _EVAL_214 = _EVAL_154 == 1'h0;
  assign _EVAL_105 = _EVAL_214 == 1'h0;
  assign _EVAL_30 = _EVAL_2 & _EVAL_105;
  assign _EVAL_186 = _EVAL_14 == 2'h0;
  assign _EVAL_195 = _EVAL_154 - 1'h1;
  assign _EVAL_24 = _EVAL_22 == 1'h0;
  assign _EVAL_133 = $signed(_EVAL_130);
  assign _EVAL_43 = $signed(_EVAL_133) == $signed(10'sh0);
  assign _EVAL_147 = $signed(_EVAL_120) == $signed(10'sh0);
  assign _EVAL_76 = _EVAL_43 | _EVAL_147;
  assign _EVAL_113 = _EVAL_10 <= 3'h6;
  assign _EVAL_125 = _EVAL_113 | _EVAL_8;
  assign _EVAL_170 = _EVAL_11 & 9'h3;
  assign _EVAL_46 = _EVAL_90 == 1'h0;
  assign _EVAL_19 = _EVAL_83 | _EVAL_8;
  assign _EVAL_161 = _EVAL_78 == 1'h0;
  assign _EVAL_117 = _EVAL_10 == 3'h1;
  assign _EVAL_44 = _EVAL_136 == 1'h0;
  assign _EVAL_187 = _EVAL_7 == _EVAL_96;
  assign _EVAL_163 = _EVAL_187 | _EVAL_8;
  assign _EVAL_211 = _EVAL_163 == 1'h0;
  assign _EVAL_171 = _EVAL_10 == _EVAL_128;
  assign _EVAL_188 = _EVAL_5 & _EVAL_207;
  assign _EVAL_196 = _EVAL_151 == 1'h0;
  assign _EVAL_189 = _EVAL_10 == 3'h5;
  assign _EVAL_215 = _EVAL_2 & _EVAL_189;
  assign _EVAL_16 = _EVAL_24 | _EVAL_150;
  assign _EVAL_139 = _EVAL_166 < plusarg_reader_out;
  assign _EVAL_82 = _EVAL_16 | _EVAL_139;
  assign _EVAL_37 = _EVAL_82 | _EVAL_8;
  assign _EVAL_71 = _EVAL_37 == 1'h0;
  assign _EVAL_23 = _EVAL_53 & _EVAL_214;
  assign _EVAL_80 = _EVAL_186 | _EVAL_8;
  assign _EVAL_77 = _EVAL_80 == 1'h0;
  assign _EVAL_32 = _EVAL_87 == 1'h0;
  assign _EVAL_122 = _EVAL_170 == 9'h0;
  assign _EVAL_56 = _EVAL_122 | _EVAL_8;
  assign _EVAL_152 = _EVAL_12 == 3'h1;
  assign _EVAL_101 = _EVAL_5 & _EVAL_109;
  assign _EVAL_68 = ~ _EVAL_142;
  assign _EVAL_65 = _EVAL_57 & _EVAL_68;
  assign _EVAL_94 = _EVAL_14 == _EVAL_210;
  assign _EVAL_155 = _EVAL_76 | _EVAL_201;
  assign _EVAL_50 = _EVAL_155 | _EVAL_184;
  assign _EVAL_114 = $signed(_EVAL_89);
  assign _EVAL_124 = $signed(_EVAL_114) == $signed(10'sh0);
  assign _EVAL_17 = _EVAL_50 | _EVAL_124;
  assign _EVAL_36 = _EVAL_17 | _EVAL_99;
  assign _EVAL_69 = _EVAL_36 | _EVAL_8;
  assign _EVAL_111 = _EVAL_24 | _EVAL_8;
  assign _EVAL_190 = _EVAL_111 == 1'h0;
  assign _EVAL_205 = _EVAL_8 == 1'h0;
  assign _EVAL_176 = _EVAL_10 == 3'h2;
  assign _EVAL_199 = _EVAL_180 == 1'h0;
  assign _EVAL_164 = _EVAL_14 != 2'h2;
  assign _EVAL_178 = _EVAL_164 | _EVAL_8;
  assign _EVAL_143 = _EVAL_178 == 1'h0;
  assign _EVAL_34 = _EVAL_5 & _EVAL_72;
  assign _EVAL_174 = _EVAL_15 | _EVAL_22;
  assign _EVAL_115 = _EVAL_174 >> _EVAL_7;
  assign _EVAL_209 = _EVAL_115 | _EVAL_8;
  assign _EVAL_45 = _EVAL_2 & _EVAL_48;
  assign _EVAL_92 = _EVAL_108 | _EVAL_8;
  assign _EVAL_213 = _EVAL_125 == 1'h0;
  assign _EVAL_28 = _EVAL_56 == 1'h0;
  assign _EVAL_93 = _EVAL_94 | _EVAL_8;
  assign _EVAL_149 = _EVAL_93 == 1'h0;
  assign _EVAL_160 = _EVAL_2 & _EVAL_117;
  assign _EVAL_123 = _EVAL_11 == _EVAL_59;
  assign _EVAL_52 = _EVAL_10 == 3'h4;
  assign _EVAL_62 = _EVAL_2 & _EVAL_52;
  assign _EVAL_31 = _EVAL_209 == 1'h0;
  assign _EVAL_135 = _EVAL_69 == 1'h0;
  assign _EVAL_157 = _EVAL_12 == 3'h2;
  assign _EVAL_145 = _EVAL_107 & _EVAL_169;
  assign _EVAL_192 = _EVAL_92 == 1'h0;
  assign _EVAL_148 = _EVAL_5 & _EVAL_152;
  assign _EVAL_183 = _EVAL_2 & _EVAL_176;
  assign _EVAL_112 = _EVAL_123 | _EVAL_8;
  assign _EVAL_217 = _EVAL_112 == 1'h0;
  assign _EVAL_21 = _EVAL_171 | _EVAL_8;
  assign _EVAL_191 = _EVAL_21 == 1'h0;
  assign _EVAL_54 = _EVAL_5 & _EVAL_131;
  assign _EVAL_64 = _EVAL_121 == 1'h0;
  assign _EVAL_79 = _EVAL_2 & _EVAL_86;
  assign _EVAL_140 = _EVAL_5 & _EVAL_110;
  assign _EVAL_156 = _EVAL_5 & _EVAL_157;
  assign _EVAL_74 = _EVAL_19 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_26 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_27 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_47 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_59 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_96 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_100 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_128 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_137 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_138 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_154 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_166 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_198 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_210 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_8) begin
      _EVAL_22 <= 1'h0;
    end else begin
      _EVAL_22 <= _EVAL_65;
    end
    if (_EVAL_8) begin
      _EVAL_26 <= 1'h0;
    end else begin
      if (_EVAL_107) begin
        if (_EVAL_169) begin
          _EVAL_26 <= 1'h0;
        end else begin
          _EVAL_26 <= _EVAL_75;
        end
      end
    end
    if (_EVAL_145) begin
      _EVAL_27 <= _EVAL_12;
    end
    if (_EVAL_23) begin
      _EVAL_47 <= _EVAL_0;
    end
    if (_EVAL_145) begin
      _EVAL_59 <= _EVAL_11;
    end
    if (_EVAL_23) begin
      _EVAL_96 <= _EVAL_7;
    end
    if (_EVAL_23) begin
      _EVAL_100 <= _EVAL_1;
    end
    if (_EVAL_23) begin
      _EVAL_128 <= _EVAL_10;
    end
    if (_EVAL_8) begin
      _EVAL_137 <= 1'h0;
    end else begin
      if (_EVAL_53) begin
        if (_EVAL_165) begin
          _EVAL_137 <= 1'h0;
        end else begin
          _EVAL_137 <= _EVAL_60;
        end
      end
    end
    if (_EVAL_8) begin
      _EVAL_138 <= 1'h0;
    end else begin
      if (_EVAL_107) begin
        if (_EVAL_91) begin
          _EVAL_138 <= 1'h0;
        end else begin
          _EVAL_138 <= _EVAL_206;
        end
      end
    end
    if (_EVAL_8) begin
      _EVAL_154 <= 1'h0;
    end else begin
      if (_EVAL_53) begin
        if (_EVAL_214) begin
          _EVAL_154 <= 1'h0;
        end else begin
          _EVAL_154 <= _EVAL_195;
        end
      end
    end
    if (_EVAL_8) begin
      _EVAL_166 <= 32'h0;
    end else begin
      if (_EVAL_39) begin
        _EVAL_166 <= 32'h0;
      end else begin
        _EVAL_166 <= _EVAL_29;
      end
    end
    if (_EVAL_23) begin
      _EVAL_198 <= _EVAL;
    end
    if (_EVAL_23) begin
      _EVAL_210 <= _EVAL_14;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5136ab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d65add17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(665a6d76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7245680c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17ec1de3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(371eba89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a85a0f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65ef3e71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(434a4a9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4dd1f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73c0d2fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e84b852)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1151c93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e8ff417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f51c64d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c145ee8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a748a3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d39705ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918329e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3be82c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed9588df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d336bb23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(128376a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d604558a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6bffdb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30613e4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc8633e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41a6e8fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f2c64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcbdbba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69caab5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47be705d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d2b57cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e4efdf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47e86156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e27472b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25d9265c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e038368e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb30eae3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c61b00c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b829e3a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(973f8bca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e73c99a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d231a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(164798cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(168274a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21708521)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85ecb399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b206431d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a712dab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35292fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(817516cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0fa85b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5853330)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830257b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df424449)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f66de93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7c265e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(566e7c2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8d2f142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95508e80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb0e06db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d8388c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e64f7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe56442)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ffa2d3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dae2ef7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3aa61cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1936c7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b19cf6d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
