//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_129(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  output [31:0] _EVAL_1,
  input  [13:0] _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input  [3:0]  _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  output        _EVAL_12,
  input  [2:0]  _EVAL_13,
  output [6:0]  _EVAL_14,
  output [3:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  output [1:0]  _EVAL_18,
  input  [6:0]  _EVAL_19
);
  wire [6:0] buffer__EVAL;
  wire [13:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire [3:0] buffer__EVAL_2;
  wire [2:0] buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [2:0] buffer__EVAL_6;
  wire [3:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [2:0] buffer__EVAL_10;
  wire [2:0] buffer__EVAL_11;
  wire [31:0] buffer__EVAL_12;
  wire [2:0] buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire [1:0] buffer__EVAL_16;
  wire [3:0] buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire [3:0] buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire [6:0] buffer__EVAL_21;
  wire [2:0] buffer__EVAL_22;
  wire [6:0] buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire [6:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire [3:0] buffer__EVAL_29;
  wire [3:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [13:0] buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire  error__EVAL;
  wire [6:0] error__EVAL_0;
  wire  error__EVAL_1;
  wire [2:0] error__EVAL_2;
  wire  error__EVAL_3;
  wire [3:0] error__EVAL_4;
  wire [6:0] error__EVAL_5;
  wire [2:0] error__EVAL_6;
  wire  error__EVAL_7;
  wire  error__EVAL_8;
  wire  error__EVAL_9;
  wire [3:0] error__EVAL_10;
  wire [13:0] error__EVAL_11;
  wire [3:0] error__EVAL_12;
  wire  error__EVAL_13;
  wire [2:0] error__EVAL_14;
  wire  error__EVAL_15;
  SiFive__EVAL_128 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34)
  );
  SiFive__EVAL_125 error (
    ._EVAL(error__EVAL),
    ._EVAL_0(error__EVAL_0),
    ._EVAL_1(error__EVAL_1),
    ._EVAL_2(error__EVAL_2),
    ._EVAL_3(error__EVAL_3),
    ._EVAL_4(error__EVAL_4),
    ._EVAL_5(error__EVAL_5),
    ._EVAL_6(error__EVAL_6),
    ._EVAL_7(error__EVAL_7),
    ._EVAL_8(error__EVAL_8),
    ._EVAL_9(error__EVAL_9),
    ._EVAL_10(error__EVAL_10),
    ._EVAL_11(error__EVAL_11),
    ._EVAL_12(error__EVAL_12),
    ._EVAL_13(error__EVAL_13),
    ._EVAL_14(error__EVAL_14),
    ._EVAL_15(error__EVAL_15)
  );
  assign _EVAL_7 = buffer__EVAL_14;
  assign error__EVAL_2 = buffer__EVAL_11;
  assign _EVAL_1 = buffer__EVAL_12;
  assign error__EVAL = buffer__EVAL_1;
  assign buffer__EVAL_5 = _EVAL_0;
  assign buffer__EVAL_22 = _EVAL_11;
  assign buffer__EVAL_10 = _EVAL_13;
  assign buffer__EVAL_0 = _EVAL_2;
  assign buffer__EVAL_4 = _EVAL_3;
  assign _EVAL_8 = buffer__EVAL_34;
  assign buffer__EVAL_20 = _EVAL_9;
  assign error__EVAL_11 = buffer__EVAL_33;
  assign _EVAL = buffer__EVAL_13;
  assign buffer__EVAL_19 = error__EVAL_12;
  assign _EVAL_4 = buffer__EVAL_28;
  assign error__EVAL_4 = buffer__EVAL_17;
  assign buffer__EVAL_9 = _EVAL_10;
  assign buffer__EVAL_3 = error__EVAL_14;
  assign buffer__EVAL_24 = _EVAL_17;
  assign error__EVAL_7 = buffer__EVAL_32;
  assign error__EVAL_0 = buffer__EVAL_23;
  assign _EVAL_18 = buffer__EVAL_16;
  assign buffer__EVAL_21 = error__EVAL_5;
  assign _EVAL_15 = buffer__EVAL_29;
  assign buffer__EVAL_27 = _EVAL_19;
  assign _EVAL_6 = buffer__EVAL_25;
  assign error__EVAL_10 = buffer__EVAL_7;
  assign buffer__EVAL_15 = error__EVAL_13;
  assign error__EVAL_6 = buffer__EVAL_6;
  assign error__EVAL_15 = _EVAL_17;
  assign error__EVAL_3 = buffer__EVAL_31;
  assign buffer__EVAL_8 = error__EVAL_9;
  assign error__EVAL_8 = _EVAL_10;
  assign buffer__EVAL_30 = _EVAL_16;
  assign buffer__EVAL_2 = _EVAL_5;
  assign buffer__EVAL_26 = error__EVAL_1;
  assign _EVAL_14 = buffer__EVAL;
  assign _EVAL_12 = buffer__EVAL_18;
endmodule
