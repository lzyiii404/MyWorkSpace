//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_192(
  input         _EVAL,
  input  [31:0] _EVAL_0,
  output [31:0] _EVAL_1,
  input         _EVAL_2
);
  wire  reg_30_d;
  wire  reg_30_q;
  wire  reg_30_en;
  wire  reg_30_clk;
  wire  reg_30_rst;
  wire  reg_20_d;
  wire  reg_20_q;
  wire  reg_20_en;
  wire  reg_20_clk;
  wire  reg_20_rst;
  wire  reg_2_d;
  wire  reg_2_q;
  wire  reg_2_en;
  wire  reg_2_clk;
  wire  reg_2_rst;
  wire  reg_28_d;
  wire  reg_28_q;
  wire  reg_28_en;
  wire  reg_28_clk;
  wire  reg_28_rst;
  wire  reg_23_d;
  wire  reg_23_q;
  wire  reg_23_en;
  wire  reg_23_clk;
  wire  reg_23_rst;
  wire  reg_12_d;
  wire  reg_12_q;
  wire  reg_12_en;
  wire  reg_12_clk;
  wire  reg_12_rst;
  wire  reg_9_d;
  wire  reg_9_q;
  wire  reg_9_en;
  wire  reg_9_clk;
  wire  reg_9_rst;
  wire  reg_31_d;
  wire  reg_31_q;
  wire  reg_31_en;
  wire  reg_31_clk;
  wire  reg_31_rst;
  wire  reg_18_d;
  wire  reg_18_q;
  wire  reg_18_en;
  wire  reg_18_clk;
  wire  reg_18_rst;
  wire  reg_27_d;
  wire  reg_27_q;
  wire  reg_27_en;
  wire  reg_27_clk;
  wire  reg_27_rst;
  wire  reg_24_d;
  wire  reg_24_q;
  wire  reg_24_en;
  wire  reg_24_clk;
  wire  reg_24_rst;
  wire  reg_8_d;
  wire  reg_8_q;
  wire  reg_8_en;
  wire  reg_8_clk;
  wire  reg_8_rst;
  wire  reg_4_d;
  wire  reg_4_q;
  wire  reg_4_en;
  wire  reg_4_clk;
  wire  reg_4_rst;
  wire  reg_0_d;
  wire  reg_0_q;
  wire  reg_0_en;
  wire  reg_0_clk;
  wire  reg_0_rst;
  wire  reg_7_d;
  wire  reg_7_q;
  wire  reg_7_en;
  wire  reg_7_clk;
  wire  reg_7_rst;
  wire  reg_25_d;
  wire  reg_25_q;
  wire  reg_25_en;
  wire  reg_25_clk;
  wire  reg_25_rst;
  wire  reg_1_d;
  wire  reg_1_q;
  wire  reg_1_en;
  wire  reg_1_clk;
  wire  reg_1_rst;
  wire  reg_5_d;
  wire  reg_5_q;
  wire  reg_5_en;
  wire  reg_5_clk;
  wire  reg_5_rst;
  wire  reg_16_d;
  wire  reg_16_q;
  wire  reg_16_en;
  wire  reg_16_clk;
  wire  reg_16_rst;
  wire  reg_21_d;
  wire  reg_21_q;
  wire  reg_21_en;
  wire  reg_21_clk;
  wire  reg_21_rst;
  wire  reg_29_d;
  wire  reg_29_q;
  wire  reg_29_en;
  wire  reg_29_clk;
  wire  reg_29_rst;
  wire  reg_19_d;
  wire  reg_19_q;
  wire  reg_19_en;
  wire  reg_19_clk;
  wire  reg_19_rst;
  wire  reg_15_d;
  wire  reg_15_q;
  wire  reg_15_en;
  wire  reg_15_clk;
  wire  reg_15_rst;
  wire  reg_6_d;
  wire  reg_6_q;
  wire  reg_6_en;
  wire  reg_6_clk;
  wire  reg_6_rst;
  wire  reg_13_d;
  wire  reg_13_q;
  wire  reg_13_en;
  wire  reg_13_clk;
  wire  reg_13_rst;
  wire  reg_14_d;
  wire  reg_14_q;
  wire  reg_14_en;
  wire  reg_14_clk;
  wire  reg_14_rst;
  wire  reg_3_d;
  wire  reg_3_q;
  wire  reg_3_en;
  wire  reg_3_clk;
  wire  reg_3_rst;
  wire  reg_10_d;
  wire  reg_10_q;
  wire  reg_10_en;
  wire  reg_10_clk;
  wire  reg_10_rst;
  wire  reg_22_d;
  wire  reg_22_q;
  wire  reg_22_en;
  wire  reg_22_clk;
  wire  reg_22_rst;
  wire  reg_11_d;
  wire  reg_11_q;
  wire  reg_11_en;
  wire  reg_11_clk;
  wire  reg_11_rst;
  wire  reg_17_d;
  wire  reg_17_q;
  wire  reg_17_en;
  wire  reg_17_clk;
  wire  reg_17_rst;
  wire  reg_26_d;
  wire  reg_26_q;
  wire  reg_26_en;
  wire  reg_26_clk;
  wire  reg_26_rst;
  wire [7:0] _EVAL_3;
  wire [7:0] _EVAL_6;
  wire [15:0] _EVAL_5;
  wire [15:0] _EVAL_4;
  AsyncResetReg #(.RESET_VALUE(0)) reg_30 (
    .d(reg_30_d),
    .q(reg_30_q),
    .en(reg_30_en),
    .clk(reg_30_clk),
    .rst(reg_30_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_20 (
    .d(reg_20_d),
    .q(reg_20_q),
    .en(reg_20_en),
    .clk(reg_20_clk),
    .rst(reg_20_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_2 (
    .d(reg_2_d),
    .q(reg_2_q),
    .en(reg_2_en),
    .clk(reg_2_clk),
    .rst(reg_2_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_28 (
    .d(reg_28_d),
    .q(reg_28_q),
    .en(reg_28_en),
    .clk(reg_28_clk),
    .rst(reg_28_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_23 (
    .d(reg_23_d),
    .q(reg_23_q),
    .en(reg_23_en),
    .clk(reg_23_clk),
    .rst(reg_23_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_12 (
    .d(reg_12_d),
    .q(reg_12_q),
    .en(reg_12_en),
    .clk(reg_12_clk),
    .rst(reg_12_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_9 (
    .d(reg_9_d),
    .q(reg_9_q),
    .en(reg_9_en),
    .clk(reg_9_clk),
    .rst(reg_9_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_31 (
    .d(reg_31_d),
    .q(reg_31_q),
    .en(reg_31_en),
    .clk(reg_31_clk),
    .rst(reg_31_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_18 (
    .d(reg_18_d),
    .q(reg_18_q),
    .en(reg_18_en),
    .clk(reg_18_clk),
    .rst(reg_18_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_27 (
    .d(reg_27_d),
    .q(reg_27_q),
    .en(reg_27_en),
    .clk(reg_27_clk),
    .rst(reg_27_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_24 (
    .d(reg_24_d),
    .q(reg_24_q),
    .en(reg_24_en),
    .clk(reg_24_clk),
    .rst(reg_24_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_8 (
    .d(reg_8_d),
    .q(reg_8_q),
    .en(reg_8_en),
    .clk(reg_8_clk),
    .rst(reg_8_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_4 (
    .d(reg_4_d),
    .q(reg_4_q),
    .en(reg_4_en),
    .clk(reg_4_clk),
    .rst(reg_4_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_0 (
    .d(reg_0_d),
    .q(reg_0_q),
    .en(reg_0_en),
    .clk(reg_0_clk),
    .rst(reg_0_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_7 (
    .d(reg_7_d),
    .q(reg_7_q),
    .en(reg_7_en),
    .clk(reg_7_clk),
    .rst(reg_7_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_25 (
    .d(reg_25_d),
    .q(reg_25_q),
    .en(reg_25_en),
    .clk(reg_25_clk),
    .rst(reg_25_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_1 (
    .d(reg_1_d),
    .q(reg_1_q),
    .en(reg_1_en),
    .clk(reg_1_clk),
    .rst(reg_1_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_5 (
    .d(reg_5_d),
    .q(reg_5_q),
    .en(reg_5_en),
    .clk(reg_5_clk),
    .rst(reg_5_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_16 (
    .d(reg_16_d),
    .q(reg_16_q),
    .en(reg_16_en),
    .clk(reg_16_clk),
    .rst(reg_16_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_21 (
    .d(reg_21_d),
    .q(reg_21_q),
    .en(reg_21_en),
    .clk(reg_21_clk),
    .rst(reg_21_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_29 (
    .d(reg_29_d),
    .q(reg_29_q),
    .en(reg_29_en),
    .clk(reg_29_clk),
    .rst(reg_29_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_19 (
    .d(reg_19_d),
    .q(reg_19_q),
    .en(reg_19_en),
    .clk(reg_19_clk),
    .rst(reg_19_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_15 (
    .d(reg_15_d),
    .q(reg_15_q),
    .en(reg_15_en),
    .clk(reg_15_clk),
    .rst(reg_15_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_6 (
    .d(reg_6_d),
    .q(reg_6_q),
    .en(reg_6_en),
    .clk(reg_6_clk),
    .rst(reg_6_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_13 (
    .d(reg_13_d),
    .q(reg_13_q),
    .en(reg_13_en),
    .clk(reg_13_clk),
    .rst(reg_13_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_14 (
    .d(reg_14_d),
    .q(reg_14_q),
    .en(reg_14_en),
    .clk(reg_14_clk),
    .rst(reg_14_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_3 (
    .d(reg_3_d),
    .q(reg_3_q),
    .en(reg_3_en),
    .clk(reg_3_clk),
    .rst(reg_3_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_10 (
    .d(reg_10_d),
    .q(reg_10_q),
    .en(reg_10_en),
    .clk(reg_10_clk),
    .rst(reg_10_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_22 (
    .d(reg_22_d),
    .q(reg_22_q),
    .en(reg_22_en),
    .clk(reg_22_clk),
    .rst(reg_22_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_11 (
    .d(reg_11_d),
    .q(reg_11_q),
    .en(reg_11_en),
    .clk(reg_11_clk),
    .rst(reg_11_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_17 (
    .d(reg_17_d),
    .q(reg_17_q),
    .en(reg_17_en),
    .clk(reg_17_clk),
    .rst(reg_17_rst)
  );
  AsyncResetReg #(.RESET_VALUE(0)) reg_26 (
    .d(reg_26_d),
    .q(reg_26_q),
    .en(reg_26_en),
    .clk(reg_26_clk),
    .rst(reg_26_rst)
  );
  assign _EVAL_3 = {reg_7_q,reg_6_q,reg_5_q,reg_4_q,reg_3_q,reg_2_q,reg_1_q,reg_0_q};
  assign _EVAL_6 = {reg_23_q,reg_22_q,reg_21_q,reg_20_q,reg_19_q,reg_18_q,reg_17_q,reg_16_q};
  assign _EVAL_5 = {reg_15_q,reg_14_q,reg_13_q,reg_12_q,reg_11_q,reg_10_q,reg_9_q,reg_8_q,_EVAL_3};
  assign _EVAL_4 = {reg_31_q,reg_30_q,reg_29_q,reg_28_q,reg_27_q,reg_26_q,reg_25_q,reg_24_q,_EVAL_6};
  assign reg_31_d = _EVAL_0[31];
  assign reg_6_rst = _EVAL_2;
  assign reg_14_en = 1'h1;
  assign reg_9_rst = _EVAL_2;
  assign reg_28_en = 1'h1;
  assign reg_12_en = 1'h1;
  assign reg_11_en = 1'h1;
  assign reg_13_d = _EVAL_0[13];
  assign reg_25_d = _EVAL_0[25];
  assign reg_18_clk = _EVAL;
  assign reg_5_clk = _EVAL;
  assign reg_21_en = 1'h1;
  assign reg_1_clk = _EVAL;
  assign reg_25_rst = _EVAL_2;
  assign reg_10_rst = _EVAL_2;
  assign reg_1_en = 1'h1;
  assign reg_0_rst = _EVAL_2;
  assign reg_1_rst = _EVAL_2;
  assign reg_16_clk = _EVAL;
  assign reg_6_en = 1'h1;
  assign reg_4_clk = _EVAL;
  assign reg_27_clk = _EVAL;
  assign reg_17_d = _EVAL_0[17];
  assign reg_16_rst = _EVAL_2;
  assign reg_21_rst = _EVAL_2;
  assign reg_17_en = 1'h1;
  assign reg_10_clk = _EVAL;
  assign reg_13_clk = _EVAL;
  assign reg_17_clk = _EVAL;
  assign reg_4_en = 1'h1;
  assign reg_25_en = 1'h1;
  assign reg_28_d = _EVAL_0[28];
  assign reg_20_d = _EVAL_0[20];
  assign reg_1_d = _EVAL_0[1];
  assign reg_24_clk = _EVAL;
  assign reg_11_clk = _EVAL;
  assign reg_5_rst = _EVAL_2;
  assign reg_26_clk = _EVAL;
  assign reg_6_d = _EVAL_0[6];
  assign reg_20_en = 1'h1;
  assign reg_30_d = _EVAL_0[30];
  assign reg_23_clk = _EVAL;
  assign reg_26_d = _EVAL_0[26];
  assign reg_2_rst = _EVAL_2;
  assign reg_4_rst = _EVAL_2;
  assign reg_31_rst = _EVAL_2;
  assign reg_28_clk = _EVAL;
  assign reg_7_en = 1'h1;
  assign reg_21_clk = _EVAL;
  assign reg_3_en = 1'h1;
  assign reg_30_en = 1'h1;
  assign reg_15_rst = _EVAL_2;
  assign reg_7_d = _EVAL_0[7];
  assign reg_29_en = 1'h1;
  assign reg_20_rst = _EVAL_2;
  assign reg_0_clk = _EVAL;
  assign reg_13_en = 1'h1;
  assign reg_0_d = _EVAL_0[0];
  assign reg_16_en = 1'h1;
  assign reg_28_rst = _EVAL_2;
  assign reg_2_clk = _EVAL;
  assign reg_4_d = _EVAL_0[4];
  assign reg_0_en = 1'h1;
  assign reg_10_d = _EVAL_0[10];
  assign reg_21_d = _EVAL_0[21];
  assign reg_12_d = _EVAL_0[12];
  assign reg_6_clk = _EVAL;
  assign reg_15_en = 1'h1;
  assign reg_12_clk = _EVAL;
  assign reg_27_d = _EVAL_0[27];
  assign reg_26_en = 1'h1;
  assign reg_23_d = _EVAL_0[23];
  assign reg_30_rst = _EVAL_2;
  assign reg_9_clk = _EVAL;
  assign reg_18_en = 1'h1;
  assign reg_8_clk = _EVAL;
  assign reg_27_en = 1'h1;
  assign reg_7_clk = _EVAL;
  assign reg_29_clk = _EVAL;
  assign reg_22_clk = _EVAL;
  assign reg_10_en = 1'h1;
  assign reg_17_rst = _EVAL_2;
  assign reg_3_rst = _EVAL_2;
  assign reg_24_en = 1'h1;
  assign reg_16_d = _EVAL_0[16];
  assign reg_24_rst = _EVAL_2;
  assign reg_3_clk = _EVAL;
  assign reg_5_d = _EVAL_0[5];
  assign reg_29_d = _EVAL_0[29];
  assign reg_8_rst = _EVAL_2;
  assign reg_31_en = 1'h1;
  assign reg_14_clk = _EVAL;
  assign reg_9_d = _EVAL_0[9];
  assign reg_23_en = 1'h1;
  assign reg_18_rst = _EVAL_2;
  assign reg_11_d = _EVAL_0[11];
  assign reg_8_d = _EVAL_0[8];
  assign reg_13_rst = _EVAL_2;
  assign reg_18_d = _EVAL_0[18];
  assign reg_24_d = _EVAL_0[24];
  assign reg_14_rst = _EVAL_2;
  assign reg_22_d = _EVAL_0[22];
  assign reg_19_rst = _EVAL_2;
  assign reg_23_rst = _EVAL_2;
  assign _EVAL_1 = {_EVAL_4,_EVAL_5};
  assign reg_30_clk = _EVAL;
  assign reg_11_rst = _EVAL_2;
  assign reg_29_rst = _EVAL_2;
  assign reg_27_rst = _EVAL_2;
  assign reg_19_d = _EVAL_0[19];
  assign reg_3_d = _EVAL_0[3];
  assign reg_5_en = 1'h1;
  assign reg_19_clk = _EVAL;
  assign reg_12_rst = _EVAL_2;
  assign reg_15_d = _EVAL_0[15];
  assign reg_26_rst = _EVAL_2;
  assign reg_19_en = 1'h1;
  assign reg_25_clk = _EVAL;
  assign reg_15_clk = _EVAL;
  assign reg_8_en = 1'h1;
  assign reg_2_d = _EVAL_0[2];
  assign reg_2_en = 1'h1;
  assign reg_22_rst = _EVAL_2;
  assign reg_20_clk = _EVAL;
  assign reg_22_en = 1'h1;
  assign reg_14_d = _EVAL_0[14];
  assign reg_9_en = 1'h1;
  assign reg_7_rst = _EVAL_2;
  assign reg_31_clk = _EVAL;
endmodule
