//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_256(
  input         _EVAL,
  input  [31:0] _EVAL_0,
  input  [29:0] _EVAL_1,
  input         _EVAL_2,
  input  [31:0] _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [1:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [29:0] _EVAL_13,
  input         _EVAL_14,
  input  [31:0] _EVAL_15,
  input  [31:0] _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input  [31:0] _EVAL_19,
  input  [29:0] _EVAL_20,
  input  [1:0]  _EVAL_21,
  input  [29:0] _EVAL_22,
  input         _EVAL_23,
  input  [1:0]  _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input  [29:0] _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input  [1:0]  _EVAL_33,
  input  [1:0]  _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input  [31:0] _EVAL_37,
  input         _EVAL_38,
  input  [1:0]  _EVAL_39,
  input         _EVAL_40,
  input  [1:0]  _EVAL_41,
  output        _EVAL_42,
  input  [29:0] _EVAL_43,
  input  [1:0]  _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input  [29:0] _EVAL_48,
  input  [31:0] _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input  [1:0]  _EVAL_54,
  input         _EVAL_55,
  input  [31:0] _EVAL_56,
  input  [29:0] _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60
);
  wire  _EVAL_229;
  wire [31:0] _EVAL_261;
  wire [31:0] _EVAL_62;
  wire [31:0] _EVAL_130;
  wire [31:0] _EVAL_297;
  wire  _EVAL_88;
  wire  _EVAL_225;
  wire [31:0] _EVAL_116;
  wire [31:0] _EVAL_162;
  wire [31:0] _EVAL_154;
  wire [31:0] _EVAL_276;
  wire  _EVAL_263;
  wire  _EVAL_124;
  wire  _EVAL_384;
  wire [31:0] _EVAL_210;
  wire [31:0] _EVAL_298;
  wire [31:0] _EVAL_142;
  wire [31:0] _EVAL_191;
  wire [31:0] _EVAL_273;
  wire [31:0] _EVAL_82;
  wire [31:0] _EVAL_156;
  wire [31:0] _EVAL_107;
  wire  _EVAL_205;
  wire  _EVAL_143;
  wire  _EVAL_146;
  wire [31:0] _EVAL_284;
  wire [31:0] _EVAL_63;
  wire [31:0] _EVAL_105;
  wire [31:0] _EVAL_207;
  wire  _EVAL_360;
  wire  _EVAL_258;
  wire [31:0] _EVAL_322;
  wire [31:0] _EVAL_372;
  wire [31:0] _EVAL_94;
  wire [31:0] _EVAL_131;
  wire  _EVAL_69;
  wire  _EVAL_362;
  wire  _EVAL_219;
  wire [31:0] _EVAL_113;
  wire [31:0] _EVAL_109;
  wire [31:0] _EVAL_202;
  wire  _EVAL_153;
  wire [31:0] _EVAL_280;
  wire [31:0] _EVAL_274;
  wire [31:0] _EVAL_317;
  wire [31:0] _EVAL_86;
  wire [31:0] _EVAL_260;
  wire [31:0] _EVAL_245;
  wire [31:0] _EVAL_222;
  wire  _EVAL_287;
  wire  _EVAL_91;
  wire  _EVAL_349;
  wire  _EVAL_85;
  wire  _EVAL_294;
  wire [31:0] _EVAL_252;
  wire [31:0] _EVAL_377;
  wire [31:0] _EVAL_122;
  wire  _EVAL_251;
  wire  _EVAL_366;
  wire  _EVAL_140;
  wire  _EVAL_329;
  wire  _EVAL_333;
  wire  _EVAL_343;
  wire  _EVAL_358;
  wire  _EVAL_254;
  wire [31:0] _EVAL_72;
  wire [31:0] _EVAL_83;
  wire [31:0] _EVAL_311;
  wire [31:0] _EVAL_168;
  wire [31:0] _EVAL_70;
  wire [31:0] _EVAL_316;
  wire [31:0] _EVAL_357;
  wire  _EVAL_272;
  wire  _EVAL_78;
  wire [31:0] _EVAL_215;
  wire [31:0] _EVAL_315;
  wire  _EVAL_64;
  wire  _EVAL_250;
  wire  _EVAL_267;
  wire  _EVAL_230;
  wire  _EVAL_313;
  wire  _EVAL_312;
  wire  _EVAL_266;
  wire  _EVAL_233;
  wire  _EVAL_161;
  wire  _EVAL_314;
  wire  _EVAL_217;
  wire [31:0] _EVAL_73;
  wire [31:0] _EVAL_378;
  wire [31:0] _EVAL_231;
  wire  _EVAL_151;
  wire  _EVAL_283;
  wire  _EVAL_242;
  wire  _EVAL_376;
  wire  _EVAL_108;
  wire  _EVAL_76;
  wire [31:0] _EVAL_354;
  wire [31:0] _EVAL_320;
  wire  _EVAL_98;
  wire  _EVAL_193;
  wire  _EVAL_211;
  wire  _EVAL_334;
  wire  _EVAL_212;
  wire  _EVAL_160;
  wire  _EVAL_184;
  wire  _EVAL_293;
  wire  _EVAL_353;
  wire  _EVAL_323;
  wire  _EVAL_253;
  wire  _EVAL_326;
  wire  _EVAL_183;
  wire [31:0] _EVAL_179;
  wire [31:0] _EVAL_148;
  wire  _EVAL_145;
  wire  _EVAL_147;
  wire  _EVAL_227;
  wire  _EVAL_114;
  wire  _EVAL_125;
  wire  _EVAL_80;
  wire  _EVAL_203;
  wire  _EVAL_190;
  wire  _EVAL_303;
  wire  _EVAL_68;
  wire  _EVAL_321;
  wire  _EVAL_213;
  wire  _EVAL_99;
  wire  _EVAL_339;
  wire  _EVAL_369;
  wire  _EVAL_169;
  wire  _EVAL_310;
  wire  _EVAL_218;
  wire  _EVAL_338;
  wire  _EVAL_368;
  wire  _EVAL_359;
  wire [31:0] _EVAL_155;
  wire [31:0] _EVAL_241;
  wire [31:0] _EVAL_188;
  wire  _EVAL_336;
  wire  _EVAL_352;
  wire  _EVAL_170;
  wire  _EVAL_281;
  wire  _EVAL_111;
  wire  _EVAL_356;
  wire  _EVAL_302;
  wire  _EVAL_237;
  wire  _EVAL_270;
  wire  _EVAL_185;
  wire  _EVAL_363;
  wire  _EVAL_223;
  wire  _EVAL_126;
  wire  _EVAL_285;
  wire  _EVAL_244;
  wire  _EVAL_118;
  wire  _EVAL_269;
  wire  _EVAL_84;
  wire  _EVAL_259;
  wire  _EVAL_71;
  wire  _EVAL_288;
  wire  _EVAL_381;
  wire  _EVAL_163;
  wire  _EVAL_374;
  wire  _EVAL_286;
  wire  _EVAL_290;
  wire  _EVAL_97;
  wire  _EVAL_373;
  assign _EVAL_229 = _EVAL_9[0];
  assign _EVAL_261 = {_EVAL_48, 2'h0};
  assign _EVAL_62 = ~ _EVAL_261;
  assign _EVAL_130 = _EVAL_62 | 32'h3f;
  assign _EVAL_297 = ~ _EVAL_130;
  assign _EVAL_88 = _EVAL_56 < _EVAL_297;
  assign _EVAL_225 = _EVAL_88 == 1'h0;
  assign _EVAL_116 = {_EVAL_22, 2'h0};
  assign _EVAL_162 = ~ _EVAL_116;
  assign _EVAL_154 = _EVAL_162 | 32'h3f;
  assign _EVAL_276 = ~ _EVAL_154;
  assign _EVAL_263 = _EVAL_56 < _EVAL_276;
  assign _EVAL_124 = _EVAL_225 & _EVAL_263;
  assign _EVAL_384 = _EVAL_229 & _EVAL_124;
  assign _EVAL_210 = {_EVAL_1, 2'h0};
  assign _EVAL_298 = ~ _EVAL_210;
  assign _EVAL_142 = _EVAL_298 | 32'h3f;
  assign _EVAL_191 = ~ _EVAL_142;
  assign _EVAL_273 = {_EVAL_13, 2'h0};
  assign _EVAL_82 = ~ _EVAL_273;
  assign _EVAL_156 = _EVAL_82 | 32'h3f;
  assign _EVAL_107 = ~ _EVAL_156;
  assign _EVAL_205 = _EVAL_56 < _EVAL_107;
  assign _EVAL_143 = _EVAL_205 == 1'h0;
  assign _EVAL_146 = _EVAL_24[0];
  assign _EVAL_284 = {_EVAL_43, 2'h0};
  assign _EVAL_63 = ~ _EVAL_284;
  assign _EVAL_105 = _EVAL_63 | 32'h3f;
  assign _EVAL_207 = ~ _EVAL_105;
  assign _EVAL_360 = _EVAL_56 < _EVAL_207;
  assign _EVAL_258 = _EVAL_360 == 1'h0;
  assign _EVAL_322 = {_EVAL_27, 2'h0};
  assign _EVAL_372 = ~ _EVAL_322;
  assign _EVAL_94 = _EVAL_372 | 32'h3f;
  assign _EVAL_131 = ~ _EVAL_94;
  assign _EVAL_69 = _EVAL_56 < _EVAL_131;
  assign _EVAL_362 = _EVAL_258 & _EVAL_69;
  assign _EVAL_219 = _EVAL_146 & _EVAL_362;
  assign _EVAL_113 = _EVAL_56 ^ _EVAL_297;
  assign _EVAL_109 = ~ _EVAL_19;
  assign _EVAL_202 = _EVAL_113 & _EVAL_109;
  assign _EVAL_153 = _EVAL_34[1];
  assign _EVAL_280 = _EVAL_56 ^ _EVAL_207;
  assign _EVAL_274 = _EVAL_56 ^ _EVAL_191;
  assign _EVAL_317 = ~ _EVAL_0;
  assign _EVAL_86 = {_EVAL_20, 2'h0};
  assign _EVAL_260 = ~ _EVAL_86;
  assign _EVAL_245 = _EVAL_260 | 32'h3f;
  assign _EVAL_222 = ~ _EVAL_245;
  assign _EVAL_287 = _EVAL_56 < _EVAL_222;
  assign _EVAL_91 = _EVAL_33 > 2'h1;
  assign _EVAL_349 = _EVAL_36 == 1'h0;
  assign _EVAL_85 = _EVAL_91 & _EVAL_349;
  assign _EVAL_294 = _EVAL_10 | _EVAL_85;
  assign _EVAL_252 = _EVAL_56 ^ _EVAL_222;
  assign _EVAL_377 = ~ _EVAL_49;
  assign _EVAL_122 = _EVAL_252 & _EVAL_377;
  assign _EVAL_251 = _EVAL_122 == 32'h0;
  assign _EVAL_366 = _EVAL_34[0];
  assign _EVAL_140 = _EVAL_143 & _EVAL_287;
  assign _EVAL_329 = _EVAL_366 & _EVAL_140;
  assign _EVAL_333 = _EVAL_153 ? _EVAL_251 : _EVAL_329;
  assign _EVAL_343 = _EVAL_45 == 1'h0;
  assign _EVAL_358 = _EVAL_91 & _EVAL_343;
  assign _EVAL_254 = _EVAL | _EVAL_358;
  assign _EVAL_72 = {_EVAL_57, 2'h0};
  assign _EVAL_83 = ~ _EVAL_72;
  assign _EVAL_311 = _EVAL_83 | 32'h3f;
  assign _EVAL_168 = ~ _EVAL_311;
  assign _EVAL_70 = _EVAL_56 ^ _EVAL_168;
  assign _EVAL_316 = ~ _EVAL_37;
  assign _EVAL_357 = _EVAL_70 & _EVAL_316;
  assign _EVAL_272 = _EVAL_357 == 32'h0;
  assign _EVAL_78 = _EVAL_44[1];
  assign _EVAL_215 = ~ _EVAL_12;
  assign _EVAL_315 = _EVAL_280 & _EVAL_215;
  assign _EVAL_64 = _EVAL_315 == 32'h0;
  assign _EVAL_250 = _EVAL_44[0];
  assign _EVAL_267 = _EVAL_56 < _EVAL_168;
  assign _EVAL_230 = _EVAL_267 == 1'h0;
  assign _EVAL_313 = _EVAL_230 & _EVAL_360;
  assign _EVAL_312 = _EVAL_250 & _EVAL_313;
  assign _EVAL_266 = _EVAL_78 ? _EVAL_64 : _EVAL_312;
  assign _EVAL_233 = _EVAL_4 == 1'h0;
  assign _EVAL_161 = _EVAL_91 & _EVAL_233;
  assign _EVAL_314 = _EVAL_50 | _EVAL_161;
  assign _EVAL_217 = _EVAL_24[1];
  assign _EVAL_73 = _EVAL_56 ^ _EVAL_131;
  assign _EVAL_378 = ~ _EVAL_3;
  assign _EVAL_231 = _EVAL_73 & _EVAL_378;
  assign _EVAL_151 = _EVAL_231 == 32'h0;
  assign _EVAL_283 = _EVAL_217 ? _EVAL_151 : _EVAL_219;
  assign _EVAL_242 = _EVAL_59 == 1'h0;
  assign _EVAL_376 = _EVAL_91 & _EVAL_242;
  assign _EVAL_108 = _EVAL_40 | _EVAL_376;
  assign _EVAL_76 = _EVAL_39[1];
  assign _EVAL_354 = _EVAL_56 ^ _EVAL_107;
  assign _EVAL_320 = _EVAL_354 & _EVAL_317;
  assign _EVAL_98 = _EVAL_320 == 32'h0;
  assign _EVAL_193 = _EVAL_39[0];
  assign _EVAL_211 = _EVAL_69 == 1'h0;
  assign _EVAL_334 = _EVAL_211 & _EVAL_205;
  assign _EVAL_212 = _EVAL_193 & _EVAL_334;
  assign _EVAL_160 = _EVAL_76 ? _EVAL_98 : _EVAL_212;
  assign _EVAL_184 = _EVAL_55 == 1'h0;
  assign _EVAL_293 = _EVAL_91 & _EVAL_184;
  assign _EVAL_353 = _EVAL_46 | _EVAL_293;
  assign _EVAL_323 = _EVAL_60 == 1'h0;
  assign _EVAL_253 = _EVAL_91 & _EVAL_323;
  assign _EVAL_326 = _EVAL_52 | _EVAL_253;
  assign _EVAL_183 = _EVAL_41[1];
  assign _EVAL_179 = ~ _EVAL_16;
  assign _EVAL_148 = _EVAL_274 & _EVAL_179;
  assign _EVAL_145 = _EVAL_148 == 32'h0;
  assign _EVAL_147 = _EVAL_41[0];
  assign _EVAL_227 = _EVAL_287 == 1'h0;
  assign _EVAL_114 = _EVAL_56 < _EVAL_191;
  assign _EVAL_125 = _EVAL_227 & _EVAL_114;
  assign _EVAL_80 = _EVAL_147 & _EVAL_125;
  assign _EVAL_203 = _EVAL_183 ? _EVAL_145 : _EVAL_80;
  assign _EVAL_190 = _EVAL_53 == 1'h0;
  assign _EVAL_303 = _EVAL_91 & _EVAL_190;
  assign _EVAL_68 = _EVAL_47 | _EVAL_303;
  assign _EVAL_321 = _EVAL_21[1];
  assign _EVAL_213 = _EVAL_202 == 32'h0;
  assign _EVAL_99 = _EVAL_21[0];
  assign _EVAL_339 = _EVAL_114 == 1'h0;
  assign _EVAL_369 = _EVAL_339 & _EVAL_88;
  assign _EVAL_169 = _EVAL_99 & _EVAL_369;
  assign _EVAL_310 = _EVAL_321 ? _EVAL_213 : _EVAL_169;
  assign _EVAL_218 = _EVAL_35 == 1'h0;
  assign _EVAL_338 = _EVAL_91 & _EVAL_218;
  assign _EVAL_368 = _EVAL_58 | _EVAL_338;
  assign _EVAL_359 = _EVAL_9[1];
  assign _EVAL_155 = _EVAL_56 ^ _EVAL_276;
  assign _EVAL_241 = ~ _EVAL_15;
  assign _EVAL_188 = _EVAL_155 & _EVAL_241;
  assign _EVAL_336 = _EVAL_188 == 32'h0;
  assign _EVAL_352 = _EVAL_359 ? _EVAL_336 : _EVAL_384;
  assign _EVAL_170 = _EVAL_23 | _EVAL_358;
  assign _EVAL_281 = _EVAL_352 ? _EVAL_170 : _EVAL_91;
  assign _EVAL_111 = _EVAL_310 ? _EVAL_368 : _EVAL_281;
  assign _EVAL_356 = _EVAL_203 ? _EVAL_68 : _EVAL_111;
  assign _EVAL_302 = _EVAL_333 ? _EVAL_326 : _EVAL_356;
  assign _EVAL_237 = _EVAL_160 ? _EVAL_353 : _EVAL_302;
  assign _EVAL_270 = _EVAL_283 ? _EVAL_108 : _EVAL_237;
  assign _EVAL_185 = _EVAL_266 ? _EVAL_314 : _EVAL_270;
  assign _EVAL_363 = _EVAL_54[1];
  assign _EVAL_223 = _EVAL_54[0];
  assign _EVAL_126 = _EVAL_223 & _EVAL_267;
  assign _EVAL_285 = _EVAL_363 ? _EVAL_272 : _EVAL_126;
  assign _EVAL_244 = _EVAL_14 | _EVAL_85;
  assign _EVAL_118 = _EVAL_30 | _EVAL_253;
  assign _EVAL_269 = _EVAL_51 | _EVAL_338;
  assign _EVAL_84 = _EVAL_5 | _EVAL_161;
  assign _EVAL_259 = _EVAL_8 | _EVAL_376;
  assign _EVAL_71 = _EVAL_26 | _EVAL_293;
  assign _EVAL_288 = _EVAL_25 | _EVAL_303;
  assign _EVAL_381 = _EVAL_352 ? _EVAL_254 : _EVAL_91;
  assign _EVAL_163 = _EVAL_310 ? _EVAL_269 : _EVAL_381;
  assign _EVAL_374 = _EVAL_203 ? _EVAL_288 : _EVAL_163;
  assign _EVAL_286 = _EVAL_333 ? _EVAL_118 : _EVAL_374;
  assign _EVAL_290 = _EVAL_160 ? _EVAL_71 : _EVAL_286;
  assign _EVAL_97 = _EVAL_283 ? _EVAL_259 : _EVAL_290;
  assign _EVAL_373 = _EVAL_266 ? _EVAL_84 : _EVAL_97;
  assign _EVAL_6 = _EVAL_285 ? _EVAL_244 : _EVAL_373;
  assign _EVAL_42 = _EVAL_285 ? _EVAL_294 : _EVAL_185;
endmodule
