//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_186_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [11:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [11:0] _EVAL_8,
  input         _EVAL_9,
  input  [25:0] _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_36;
  reg [31:0] _RAND_0;
  reg [1:0] _EVAL_39;
  reg [31:0] _RAND_1;
  reg  _EVAL_49;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_95;
  reg [31:0] _RAND_3;
  reg [2335:0] _EVAL_118;
  reg [2335:0] _RAND_4;
  reg [11:0] _EVAL_119;
  reg [31:0] _RAND_5;
  reg [1:0] _EVAL_131;
  reg [31:0] _RAND_6;
  reg  _EVAL_132;
  reg [31:0] _RAND_7;
  reg  _EVAL_133;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_146;
  reg [31:0] _RAND_9;
  reg [25:0] _EVAL_154;
  reg [31:0] _RAND_10;
  reg [11:0] _EVAL_179;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_195;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_226;
  reg [31:0] _RAND_13;
  wire  _EVAL_83;
  wire  _EVAL_174;
  wire  _EVAL_161;
  wire  _EVAL_211;
  wire [31:0] _EVAL_199;
  wire  _EVAL_59;
  wire  _EVAL_123;
  wire  _EVAL_99;
  wire  _EVAL_70;
  wire  _EVAL_109;
  wire  _EVAL_157;
  wire  _EVAL_160;
  wire [4095:0] _EVAL_152;
  wire [4095:0] _EVAL_94;
  wire [2335:0] _EVAL_34;
  wire [2335:0] _EVAL_97;
  wire  _EVAL_126;
  wire  _EVAL_37;
  wire  _EVAL_80;
  wire  _EVAL_200;
  wire  _EVAL_44;
  wire [4095:0] _EVAL_127;
  wire [4095:0] _EVAL_167;
  wire [2335:0] _EVAL_55;
  wire [2335:0] _EVAL_107;
  wire [2335:0] _EVAL_155;
  wire  _EVAL_184;
  wire  _EVAL_181;
  wire  _EVAL_104;
  wire  _EVAL_50;
  wire  _EVAL_166;
  wire  _EVAL_61;
  wire  _EVAL_110;
  wire  _EVAL_210;
  wire  _EVAL_203;
  wire [2335:0] _EVAL_29;
  wire [2335:0] _EVAL_105;
  wire  _EVAL_222;
  wire  _EVAL_74;
  wire  _EVAL_89;
  wire  _EVAL_145;
  wire  _EVAL_51;
  wire  _EVAL_28;
  wire  _EVAL_27;
  wire  _EVAL_21;
  wire  _EVAL_180;
  wire  _EVAL_147;
  wire  _EVAL_122;
  wire  _EVAL_142;
  wire  _EVAL_90;
  wire  _EVAL_116;
  wire [1:0] _EVAL_73;
  wire [1:0] _EVAL_188;
  wire  _EVAL_86;
  wire  _EVAL_189;
  wire  _EVAL_112;
  wire  _EVAL_40;
  wire  _EVAL_35;
  wire  _EVAL_148;
  wire  _EVAL_204;
  wire  _EVAL_197;
  wire  _EVAL_92;
  wire  _EVAL_164;
  wire  _EVAL_196;
  wire  _EVAL_212;
  wire  _EVAL_88;
  wire  _EVAL_129;
  wire  _EVAL_182;
  wire  _EVAL_232;
  wire  _EVAL_162;
  wire  _EVAL_111;
  wire  _EVAL_98;
  wire  _EVAL_24;
  wire  _EVAL_87;
  wire  _EVAL_228;
  wire [3:0] _EVAL_143;
  wire  _EVAL_18;
  wire  _EVAL_135;
  wire  _EVAL_52;
  wire  _EVAL_32;
  wire  _EVAL_170;
  wire  _EVAL_202;
  wire  _EVAL_163;
  wire [25:0] _EVAL_186;
  wire [26:0] _EVAL_65;
  wire  _EVAL_91;
  wire  _EVAL_45;
  wire  _EVAL_227;
  wire  _EVAL_121;
  wire  _EVAL_38;
  wire [3:0] _EVAL_23;
  wire [3:0] _EVAL_125;
  wire  _EVAL_77;
  wire  _EVAL_140;
  wire  _EVAL_151;
  wire  _EVAL_84;
  wire  _EVAL_224;
  wire  _EVAL_43;
  wire [4:0] _EVAL_205;
  wire [1:0] _EVAL_207;
  wire [1:0] _EVAL_169;
  wire  _EVAL_221;
  wire  _EVAL_48;
  wire [3:0] _EVAL_120;
  wire  _EVAL_63;
  wire  _EVAL_150;
  wire  _EVAL_225;
  wire  _EVAL_183;
  wire  _EVAL_191;
  wire  _EVAL_100;
  wire [25:0] _EVAL_115;
  wire [25:0] _EVAL_153;
  wire  _EVAL_79;
  wire  _EVAL_114;
  wire  _EVAL_198;
  wire  _EVAL_54;
  wire  _EVAL_217;
  wire  _EVAL_141;
  wire  _EVAL_193;
  wire  _EVAL_57;
  wire  _EVAL_214;
  wire  _EVAL_22;
  wire  _EVAL_144;
  wire  _EVAL_185;
  wire  _EVAL_78;
  wire  _EVAL_139;
  wire  _EVAL_201;
  wire  _EVAL_159;
  wire  _EVAL_75;
  wire [26:0] _EVAL_58;
  wire [26:0] _EVAL_76;
  wire  _EVAL_209;
  wire  _EVAL_15;
  wire  _EVAL_82;
  wire  _EVAL_103;
  wire  _EVAL_229;
  wire  _EVAL_171;
  wire  _EVAL_71;
  wire  _EVAL_194;
  wire  _EVAL_108;
  wire  _EVAL_128;
  wire  _EVAL_165;
  wire  _EVAL_85;
  wire  _EVAL_20;
  wire [2335:0] _EVAL_230;
  wire  _EVAL_208;
  wire  _EVAL_66;
  wire  _EVAL_60;
  wire  _EVAL_219;
  wire  _EVAL_113;
  wire  _EVAL_30;
  wire  _EVAL_173;
  wire  _EVAL_47;
  wire  _EVAL_190;
  wire  _EVAL_138;
  wire  _EVAL_223;
  wire  _EVAL_192;
  wire  _EVAL_72;
  wire  _EVAL_187;
  wire  _EVAL_25;
  wire  _EVAL_68;
  wire  _EVAL_137;
  wire  _EVAL_149;
  wire  _EVAL_33;
  wire  _EVAL_64;
  wire  _EVAL_158;
  wire  _EVAL_117;
  wire  _EVAL_130;
  wire  _EVAL_218;
  wire  _EVAL_134;
  wire  _EVAL_101;
  wire  _EVAL_124;
  wire  _EVAL_176;
  wire  _EVAL_213;
  wire  _EVAL_19;
  wire  _EVAL_220;
  wire  _EVAL_26;
  wire  _EVAL_17;
  wire  _EVAL_31;
  wire  _EVAL_168;
  wire  _EVAL_53;
  wire  _EVAL_106;
  wire  _EVAL_16;
  wire  _EVAL_156;
  wire  _EVAL_206;
  wire  _EVAL_81;
  wire  _EVAL_172;
  wire  _EVAL_136;
  wire  _EVAL_177;
  wire  _EVAL_46;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_83 = _EVAL_13 & _EVAL_14;
  assign _EVAL_174 = _EVAL_7 & _EVAL;
  assign _EVAL_161 = _EVAL_83 | _EVAL_174;
  assign _EVAL_211 = _EVAL_226 < plusarg_reader_out;
  assign _EVAL_199 = _EVAL_226 + 32'h1;
  assign _EVAL_59 = _EVAL_11 == _EVAL_195;
  assign _EVAL_123 = _EVAL_59 | _EVAL_5;
  assign _EVAL_99 = _EVAL_3 <= 3'h2;
  assign _EVAL_70 = _EVAL_99 | _EVAL_5;
  assign _EVAL_109 = _EVAL_70 == 1'h0;
  assign _EVAL_157 = _EVAL_133 == 1'h0;
  assign _EVAL_160 = _EVAL_83 & _EVAL_157;
  assign _EVAL_152 = 4096'h1 << _EVAL_8;
  assign _EVAL_94 = _EVAL_160 ? _EVAL_152 : 4096'h0;
  assign _EVAL_34 = _EVAL_94[2335:0];
  assign _EVAL_97 = _EVAL_118 | _EVAL_34;
  assign _EVAL_126 = _EVAL_49 == 1'h0;
  assign _EVAL_37 = _EVAL_174 & _EVAL_126;
  assign _EVAL_80 = _EVAL_2 == 3'h6;
  assign _EVAL_200 = _EVAL_80 == 1'h0;
  assign _EVAL_44 = _EVAL_37 & _EVAL_200;
  assign _EVAL_127 = 4096'h1 << _EVAL_4;
  assign _EVAL_167 = _EVAL_44 ? _EVAL_127 : 4096'h0;
  assign _EVAL_55 = _EVAL_167[2335:0];
  assign _EVAL_107 = ~ _EVAL_55;
  assign _EVAL_155 = _EVAL_97 & _EVAL_107;
  assign _EVAL_184 = _EVAL_11 == 3'h3;
  assign _EVAL_181 = _EVAL_0 == _EVAL_39;
  assign _EVAL_104 = _EVAL_181 | _EVAL_5;
  assign _EVAL_50 = _EVAL_104 == 1'h0;
  assign _EVAL_166 = _EVAL_0[0];
  assign _EVAL_61 = _EVAL_11 == 3'h2;
  assign _EVAL_110 = _EVAL_14 & _EVAL_61;
  assign _EVAL_210 = _EVAL_36 == 1'h0;
  assign _EVAL_203 = _EVAL_36 - 1'h1;
  assign _EVAL_29 = _EVAL_34 | _EVAL_118;
  assign _EVAL_105 = _EVAL_29 >> _EVAL_4;
  assign _EVAL_222 = _EVAL_105[0];
  assign _EVAL_74 = _EVAL_222 | _EVAL_5;
  assign _EVAL_89 = _EVAL_74 == 1'h0;
  assign _EVAL_145 = _EVAL_4 <= 12'h91f;
  assign _EVAL_51 = _EVAL_145 | _EVAL_5;
  assign _EVAL_28 = _EVAL_51 == 1'h0;
  assign _EVAL_27 = _EVAL_3 <= 3'h3;
  assign _EVAL_21 = _EVAL_3 != 3'h0;
  assign _EVAL_180 = _EVAL_21 | _EVAL_5;
  assign _EVAL_147 = _EVAL_180 == 1'h0;
  assign _EVAL_122 = _EVAL_2 == _EVAL_95;
  assign _EVAL_142 = _EVAL_11 == 3'h1;
  assign _EVAL_90 = _EVAL_14 & _EVAL_142;
  assign _EVAL_116 = _EVAL_0 >= 2'h2;
  assign _EVAL_73 = 2'h1 << _EVAL_166;
  assign _EVAL_188 = _EVAL_73 | 2'h1;
  assign _EVAL_86 = _EVAL_188[1];
  assign _EVAL_189 = _EVAL_10[1];
  assign _EVAL_112 = _EVAL_86 & _EVAL_189;
  assign _EVAL_40 = _EVAL_116 | _EVAL_112;
  assign _EVAL_35 = _EVAL_188[0];
  assign _EVAL_148 = _EVAL_10[0];
  assign _EVAL_204 = _EVAL_189 & _EVAL_148;
  assign _EVAL_197 = _EVAL_35 & _EVAL_204;
  assign _EVAL_92 = _EVAL_40 | _EVAL_197;
  assign _EVAL_164 = _EVAL_148 == 1'h0;
  assign _EVAL_196 = _EVAL_189 & _EVAL_164;
  assign _EVAL_212 = _EVAL_35 & _EVAL_196;
  assign _EVAL_88 = _EVAL_40 | _EVAL_212;
  assign _EVAL_129 = _EVAL_189 == 1'h0;
  assign _EVAL_182 = _EVAL_86 & _EVAL_129;
  assign _EVAL_232 = _EVAL_116 | _EVAL_182;
  assign _EVAL_162 = _EVAL_129 & _EVAL_148;
  assign _EVAL_111 = _EVAL_35 & _EVAL_162;
  assign _EVAL_98 = _EVAL_232 | _EVAL_111;
  assign _EVAL_24 = _EVAL_129 & _EVAL_164;
  assign _EVAL_87 = _EVAL_35 & _EVAL_24;
  assign _EVAL_228 = _EVAL_232 | _EVAL_87;
  assign _EVAL_143 = {_EVAL_92,_EVAL_88,_EVAL_98,_EVAL_228};
  assign _EVAL_18 = _EVAL_1 == _EVAL_143;
  assign _EVAL_135 = _EVAL_9 == 1'h0;
  assign _EVAL_52 = _EVAL_135 | _EVAL_5;
  assign _EVAL_32 = _EVAL_0 <= 2'h2;
  assign _EVAL_170 = _EVAL_3 == 3'h0;
  assign _EVAL_202 = _EVAL_170 | _EVAL_5;
  assign _EVAL_163 = _EVAL_202 == 1'h0;
  assign _EVAL_186 = _EVAL_10 ^ 26'h2000000;
  assign _EVAL_65 = {1'b0,$signed(_EVAL_186)};
  assign _EVAL_91 = _EVAL_8 <= 12'h91f;
  assign _EVAL_45 = _EVAL_91 | _EVAL_5;
  assign _EVAL_227 = _EVAL_45 == 1'h0;
  assign _EVAL_121 = _EVAL_11 == 3'h7;
  assign _EVAL_38 = _EVAL_14 & _EVAL_121;
  assign _EVAL_23 = ~ _EVAL_143;
  assign _EVAL_125 = _EVAL_1 & _EVAL_23;
  assign _EVAL_77 = _EVAL_2 == 3'h5;
  assign _EVAL_140 = _EVAL & _EVAL_77;
  assign _EVAL_151 = _EVAL_3 == _EVAL_146;
  assign _EVAL_84 = _EVAL_12 >= 2'h2;
  assign _EVAL_224 = _EVAL_84 | _EVAL_5;
  assign _EVAL_43 = _EVAL_224 == 1'h0;
  assign _EVAL_205 = 5'h3 << _EVAL_0;
  assign _EVAL_207 = _EVAL_205[1:0];
  assign _EVAL_169 = ~ _EVAL_207;
  assign _EVAL_221 = _EVAL_132 == 1'h0;
  assign _EVAL_48 = _EVAL_174 & _EVAL_221;
  assign _EVAL_120 = ~ _EVAL_1;
  assign _EVAL_63 = _EVAL_120 == 4'h0;
  assign _EVAL_150 = _EVAL_63 | _EVAL_5;
  assign _EVAL_225 = _EVAL_150 == 1'h0;
  assign _EVAL_183 = _EVAL_2 == 3'h1;
  assign _EVAL_191 = _EVAL_3 <= 3'h4;
  assign _EVAL_100 = _EVAL_11 == 3'h5;
  assign _EVAL_115 = {{24'd0}, _EVAL_169};
  assign _EVAL_153 = _EVAL_10 & _EVAL_115;
  assign _EVAL_79 = _EVAL_8 == _EVAL_179;
  assign _EVAL_114 = _EVAL_79 | _EVAL_5;
  assign _EVAL_198 = _EVAL_114 == 1'h0;
  assign _EVAL_54 = _EVAL_2 == 3'h0;
  assign _EVAL_217 = _EVAL & _EVAL_54;
  assign _EVAL_141 = _EVAL & _EVAL_80;
  assign _EVAL_193 = _EVAL_132 - 1'h1;
  assign _EVAL_57 = _EVAL_191 | _EVAL_5;
  assign _EVAL_214 = _EVAL_125 == 4'h0;
  assign _EVAL_22 = _EVAL_214 | _EVAL_5;
  assign _EVAL_144 = _EVAL_22 == 1'h0;
  assign _EVAL_185 = _EVAL_133 - 1'h1;
  assign _EVAL_78 = _EVAL_210 == 1'h0;
  assign _EVAL_139 = _EVAL_27 | _EVAL_5;
  assign _EVAL_201 = _EVAL_12 == _EVAL_131;
  assign _EVAL_159 = _EVAL_201 | _EVAL_5;
  assign _EVAL_75 = _EVAL_159 == 1'h0;
  assign _EVAL_58 = $signed(_EVAL_65) & $signed(-27'sh10000);
  assign _EVAL_76 = $signed(_EVAL_58);
  assign _EVAL_209 = $signed(_EVAL_76) == $signed(27'sh0);
  assign _EVAL_15 = _EVAL_32 & _EVAL_209;
  assign _EVAL_82 = _EVAL_15 | _EVAL_5;
  assign _EVAL_103 = _EVAL_82 == 1'h0;
  assign _EVAL_229 = _EVAL_10 == _EVAL_154;
  assign _EVAL_171 = _EVAL_229 | _EVAL_5;
  assign _EVAL_71 = _EVAL_171 == 1'h0;
  assign _EVAL_194 = _EVAL_2 == 3'h2;
  assign _EVAL_108 = _EVAL & _EVAL_194;
  assign _EVAL_128 = _EVAL_2 <= 3'h6;
  assign _EVAL_165 = _EVAL_128 | _EVAL_5;
  assign _EVAL_85 = _EVAL_165 == 1'h0;
  assign _EVAL_20 = _EVAL_2 == 3'h4;
  assign _EVAL_230 = _EVAL_118 >> _EVAL_8;
  assign _EVAL_208 = _EVAL_230[0];
  assign _EVAL_66 = _EVAL_118 != 2336'h0;
  assign _EVAL_60 = _EVAL_66 == 1'h0;
  assign _EVAL_219 = _EVAL_221 == 1'h0;
  assign _EVAL_113 = _EVAL_208 == 1'h0;
  assign _EVAL_30 = _EVAL_11 == 3'h4;
  assign _EVAL_173 = _EVAL_14 & _EVAL_30;
  assign _EVAL_47 = _EVAL_153 == 26'h0;
  assign _EVAL_190 = plusarg_reader_out == 32'h0;
  assign _EVAL_138 = _EVAL_60 | _EVAL_190;
  assign _EVAL_223 = _EVAL_11 == 3'h0;
  assign _EVAL_192 = _EVAL_14 & _EVAL_223;
  assign _EVAL_72 = _EVAL_49 - 1'h1;
  assign _EVAL_187 = _EVAL_123 == 1'h0;
  assign _EVAL_25 = _EVAL_122 | _EVAL_5;
  assign _EVAL_68 = _EVAL_25 == 1'h0;
  assign _EVAL_137 = _EVAL_4 == _EVAL_119;
  assign _EVAL_149 = _EVAL_14 & _EVAL_78;
  assign _EVAL_33 = _EVAL_18 | _EVAL_5;
  assign _EVAL_64 = _EVAL_33 == 1'h0;
  assign _EVAL_158 = _EVAL_11 == 3'h6;
  assign _EVAL_117 = _EVAL_137 | _EVAL_5;
  assign _EVAL_130 = _EVAL_117 == 1'h0;
  assign _EVAL_218 = _EVAL_57 == 1'h0;
  assign _EVAL_134 = _EVAL_138 | _EVAL_211;
  assign _EVAL_101 = _EVAL_134 | _EVAL_5;
  assign _EVAL_124 = _EVAL & _EVAL_183;
  assign _EVAL_176 = _EVAL_113 | _EVAL_5;
  assign _EVAL_213 = _EVAL_176 == 1'h0;
  assign _EVAL_19 = _EVAL_14 & _EVAL_158;
  assign _EVAL_220 = _EVAL_5 == 1'h0;
  assign _EVAL_26 = _EVAL_139 == 1'h0;
  assign _EVAL_17 = _EVAL & _EVAL_20;
  assign _EVAL_31 = _EVAL & _EVAL_219;
  assign _EVAL_168 = _EVAL_116 | _EVAL_5;
  assign _EVAL_53 = _EVAL_168 == 1'h0;
  assign _EVAL_106 = _EVAL_47 | _EVAL_5;
  assign _EVAL_16 = _EVAL_106 == 1'h0;
  assign _EVAL_156 = _EVAL_14 & _EVAL_100;
  assign _EVAL_206 = _EVAL_52 == 1'h0;
  assign _EVAL_81 = _EVAL_14 & _EVAL_184;
  assign _EVAL_172 = _EVAL_151 | _EVAL_5;
  assign _EVAL_136 = _EVAL_101 == 1'h0;
  assign _EVAL_177 = _EVAL_172 == 1'h0;
  assign _EVAL_46 = _EVAL_83 & _EVAL_210;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_36 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_39 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_49 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_95 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {73{`RANDOM}};
  _EVAL_118 = _RAND_4[2335:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_119 = _RAND_5[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_131 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_132 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_133 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_146 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_154 = _RAND_10[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_179 = _RAND_11[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_195 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_226 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_6) begin
    if (_EVAL_5) begin
      _EVAL_36 <= 1'h0;
    end else begin
      if (_EVAL_83) begin
        if (_EVAL_210) begin
          _EVAL_36 <= 1'h0;
        end else begin
          _EVAL_36 <= _EVAL_203;
        end
      end
    end
    if (_EVAL_46) begin
      _EVAL_39 <= _EVAL_0;
    end
    if (_EVAL_5) begin
      _EVAL_49 <= 1'h0;
    end else begin
      if (_EVAL_174) begin
        if (_EVAL_126) begin
          _EVAL_49 <= 1'h0;
        end else begin
          _EVAL_49 <= _EVAL_72;
        end
      end
    end
    if (_EVAL_48) begin
      _EVAL_95 <= _EVAL_2;
    end
    if (_EVAL_5) begin
      _EVAL_118 <= 2336'h0;
    end else begin
      _EVAL_118 <= _EVAL_155;
    end
    if (_EVAL_48) begin
      _EVAL_119 <= _EVAL_4;
    end
    if (_EVAL_48) begin
      _EVAL_131 <= _EVAL_12;
    end
    if (_EVAL_5) begin
      _EVAL_132 <= 1'h0;
    end else begin
      if (_EVAL_174) begin
        if (_EVAL_221) begin
          _EVAL_132 <= 1'h0;
        end else begin
          _EVAL_132 <= _EVAL_193;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_133 <= 1'h0;
    end else begin
      if (_EVAL_83) begin
        if (_EVAL_157) begin
          _EVAL_133 <= 1'h0;
        end else begin
          _EVAL_133 <= _EVAL_185;
        end
      end
    end
    if (_EVAL_46) begin
      _EVAL_146 <= _EVAL_3;
    end
    if (_EVAL_46) begin
      _EVAL_154 <= _EVAL_10;
    end
    if (_EVAL_46) begin
      _EVAL_179 <= _EVAL_8;
    end
    if (_EVAL_46) begin
      _EVAL_195 <= _EVAL_11;
    end
    if (_EVAL_5) begin
      _EVAL_226 <= 32'h0;
    end else begin
      if (_EVAL_161) begin
        _EVAL_226 <= 32'h0;
      end else begin
        _EVAL_226 <= _EVAL_199;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c449091)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4efed878)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60fd7c25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69d41dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14e2f350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37730a8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96274fa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5185208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e013b5e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb2bd77a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a661060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baa0350f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de9d6f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a4268c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d01bea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db43c511)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab395ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6402889b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfb81090)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7e21bcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f40ec1a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac154cdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee00e844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c27938d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b217e8ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93e31beb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fa87ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7388bf00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc7233e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f9622ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88094bbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1334fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5639dc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3eea9ee1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f54c4c73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(879452a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8577f3c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9803939a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2c57440)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c2e8448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c3e1934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1f916d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90396575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(201fb6f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(985a103d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e7fda5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7dc8374)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d050aaa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(649534d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f05cec9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9016)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb9c9161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c623b40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(371f8fa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31e4f3b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7751c23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e14713c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62fffe28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16b9b574)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c213697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc780a12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21fd42f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34393ad9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d8e5a88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a3c9b66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6676c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ced76a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27c0c9e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16558a59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923bae2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2289885)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
