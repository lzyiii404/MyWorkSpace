//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_238(
  output [2:0]  _EVAL,
  output [63:0] _EVAL_0,
  input         _EVAL_1,
  output [2:0]  _EVAL_2,
  input  [6:0]  _EVAL_3,
  input  [24:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  output [7:0]  _EVAL_6,
  output [2:0]  _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  output [24:0] _EVAL_14,
  output [6:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [3:0]  _EVAL_17,
  output [6:0]  _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input  [6:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  input  [63:0] _EVAL_23,
  input  [31:0] _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  output        _EVAL_27,
  output [31:0] _EVAL_28
);
  wire  Repeater__EVAL;
  wire [2:0] Repeater__EVAL_0;
  wire [2:0] Repeater__EVAL_1;
  wire  Repeater__EVAL_2;
  wire [63:0] Repeater__EVAL_3;
  wire [6:0] Repeater__EVAL_4;
  wire [2:0] Repeater__EVAL_5;
  wire [63:0] Repeater__EVAL_6;
  wire  Repeater__EVAL_7;
  wire [2:0] Repeater__EVAL_8;
  wire  Repeater__EVAL_9;
  wire  Repeater__EVAL_10;
  wire  Repeater__EVAL_11;
  wire [6:0] Repeater__EVAL_12;
  wire  Repeater__EVAL_13;
  reg  _EVAL_44;
  reg [31:0] _RAND_0;
  reg  _EVAL_49;
  reg [31:0] _RAND_1;
  reg  _EVAL_51;
  reg [31:0] _RAND_2;
  reg  _EVAL_52;
  reg [31:0] _RAND_3;
  reg  _EVAL_53;
  reg [31:0] _RAND_4;
  reg  _EVAL_54;
  reg [31:0] _RAND_5;
  reg  _EVAL_69;
  reg [31:0] _RAND_6;
  reg  _EVAL_76;
  reg [31:0] _RAND_7;
  reg  _EVAL_78;
  reg [31:0] _RAND_8;
  reg  _EVAL_80;
  reg [31:0] _RAND_9;
  reg  _EVAL_87;
  reg [31:0] _RAND_10;
  reg  _EVAL_90;
  reg [31:0] _RAND_11;
  reg  _EVAL_91;
  reg [31:0] _RAND_12;
  reg  _EVAL_98;
  reg [31:0] _RAND_13;
  reg  _EVAL_103;
  reg [31:0] _RAND_14;
  reg  _EVAL_104;
  reg [31:0] _RAND_15;
  reg [31:0] _EVAL_114;
  reg [31:0] _RAND_16;
  reg  _EVAL_115;
  reg [31:0] _RAND_17;
  reg [3:0] _EVAL_116;
  reg [31:0] _RAND_18;
  reg  _EVAL_118;
  reg [31:0] _RAND_19;
  reg  _EVAL_127;
  reg [31:0] _RAND_20;
  reg  _EVAL_142;
  reg [31:0] _RAND_21;
  reg  _EVAL_147;
  reg [31:0] _RAND_22;
  reg  _EVAL_153;
  reg [31:0] _RAND_23;
  reg  _EVAL_154;
  reg [31:0] _RAND_24;
  reg  _EVAL_155;
  reg [31:0] _RAND_25;
  reg  _EVAL_165;
  reg [31:0] _RAND_26;
  reg  _EVAL_182;
  reg [31:0] _RAND_27;
  reg  _EVAL_194;
  reg [31:0] _RAND_28;
  reg  _EVAL_198;
  reg [31:0] _RAND_29;
  reg  _EVAL_203;
  reg [31:0] _RAND_30;
  reg  _EVAL_204;
  reg [31:0] _RAND_31;
  reg  _EVAL_211;
  reg [31:0] _RAND_32;
  reg  _EVAL_214;
  reg [31:0] _RAND_33;
  reg  _EVAL_227;
  reg [31:0] _RAND_34;
  reg  _EVAL_243;
  reg [31:0] _RAND_35;
  reg  _EVAL_244;
  reg [31:0] _RAND_36;
  reg  _EVAL_253;
  reg [31:0] _RAND_37;
  reg  _EVAL_255;
  reg [31:0] _RAND_38;
  reg  _EVAL_258;
  reg [31:0] _RAND_39;
  reg  _EVAL_274;
  reg [31:0] _RAND_40;
  reg  _EVAL_280;
  reg [31:0] _RAND_41;
  reg  _EVAL_281;
  reg [31:0] _RAND_42;
  reg  _EVAL_287;
  reg [31:0] _RAND_43;
  reg  _EVAL_291;
  reg [31:0] _RAND_44;
  reg  _EVAL_292;
  reg [31:0] _RAND_45;
  reg  _EVAL_294;
  reg [31:0] _RAND_46;
  wire  _EVAL_117;
  wire  _EVAL_235;
  wire  _EVAL_66;
  wire  _EVAL_30;
  wire  _EVAL_137;
  wire  _EVAL_285;
  wire  _EVAL_202;
  wire  _EVAL_133;
  wire [9:0] _EVAL_93;
  wire [2:0] _EVAL_172;
  wire [2:0] _EVAL_171;
  wire  _EVAL_184;
  wire  _EVAL_231;
  wire  _EVAL_180;
  wire  _EVAL_224;
  wire  _EVAL_175;
  wire  _EVAL_106;
  wire [6:0] _EVAL_36;
  wire  _EVAL_208;
  wire  _EVAL_277;
  wire  _EVAL_110;
  wire  _EVAL_77;
  wire  _EVAL_257;
  wire  _EVAL_239;
  wire  _EVAL_60;
  wire  _EVAL_176;
  wire  _EVAL_72;
  wire  _EVAL_65;
  wire  _EVAL_206;
  wire  _EVAL_57;
  wire  _EVAL_275;
  wire  _EVAL_31;
  wire  _EVAL_75;
  wire  _EVAL_29;
  wire  _EVAL_141;
  wire  _EVAL_125;
  wire  _EVAL_158;
  wire  _EVAL_283;
  wire  _EVAL_174;
  wire  _EVAL_156;
  wire  _EVAL_201;
  wire  _EVAL_225;
  wire  _EVAL_48;
  wire  _EVAL_178;
  wire  _EVAL_113;
  wire  _EVAL_242;
  wire  _EVAL_237;
  wire  _EVAL_268;
  wire  _EVAL_261;
  wire  _EVAL_265;
  wire  _EVAL_102;
  wire  _EVAL_168;
  wire  _EVAL_228;
  wire  _EVAL_139;
  wire  _EVAL_162;
  wire  _EVAL_215;
  wire  _EVAL_73;
  wire  _EVAL_121;
  wire  _EVAL_124;
  wire  _EVAL_33;
  wire [1:0] _EVAL_240;
  wire [3:0] _EVAL_190;
  wire [2:0] _EVAL_39;
  wire [2:0] _EVAL_68;
  wire  _EVAL_143;
  wire  _EVAL_160;
  wire  _EVAL_167;
  wire  _EVAL_286;
  wire  _EVAL_67;
  wire  _EVAL_83;
  wire  _EVAL_256;
  wire  _EVAL_212;
  wire  _EVAL_181;
  wire  _EVAL_59;
  wire  _EVAL_238;
  wire  _EVAL_157;
  wire  _EVAL_97;
  wire  _EVAL_135;
  wire  _EVAL_186;
  wire  _EVAL_272;
  wire  _EVAL_84;
  wire  _EVAL_267;
  wire  _EVAL_74;
  wire  _EVAL_159;
  wire  _EVAL_79;
  wire  _EVAL_63;
  wire  _EVAL_112;
  wire  _EVAL_144;
  wire  _EVAL_131;
  wire  _EVAL_119;
  wire  _EVAL_134;
  wire  _EVAL_138;
  wire  _EVAL_164;
  wire  _EVAL_282;
  wire  _EVAL_289;
  wire  _EVAL_226;
  wire  _EVAL_32;
  wire  _EVAL_136;
  wire  _EVAL_290;
  wire  _EVAL_185;
  wire  _EVAL_266;
  wire  _EVAL_34;
  wire  _EVAL_50;
  wire  _EVAL_229;
  wire [31:0] _EVAL_234;
  wire [31:0] _EVAL_187;
  wire [63:0] _EVAL_88;
  wire [31:0] _EVAL_233;
  wire  _EVAL_205;
  wire  _EVAL_220;
  wire [3:0] _EVAL_99;
  wire  _EVAL_279;
  wire  _EVAL_61;
  wire  _EVAL_195;
  wire [2:0] _EVAL_92;
  wire [9:0] _EVAL_236;
  wire [2:0] _EVAL_62;
  wire [2:0] _EVAL_183;
  wire  _EVAL_192;
  wire  _EVAL_170;
  wire [2:0] _EVAL_241;
  wire  _EVAL_58;
  wire  _EVAL_123;
  wire  _EVAL_161;
  wire  _EVAL_56;
  wire  _EVAL_188;
  wire  _EVAL_64;
  wire  _EVAL_140;
  wire  _EVAL_70;
  wire  _EVAL_149;
  wire  _EVAL_284;
  wire  _EVAL_271;
  wire  _EVAL_100;
  wire  _EVAL_199;
  wire  _EVAL_55;
  wire  _EVAL_38;
  wire  _EVAL_96;
  wire  _EVAL_105;
  wire  _EVAL_130;
  wire  _EVAL_166;
  wire  _EVAL_108;
  wire  _EVAL_259;
  wire  _EVAL_107;
  wire  _EVAL_218;
  wire  _EVAL_230;
  wire  _EVAL_94;
  wire  _EVAL_210;
  wire  _EVAL_42;
  wire  _EVAL_260;
  wire  _EVAL_196;
  wire  _EVAL_81;
  wire  _EVAL_132;
  wire  _EVAL_95;
  wire  _EVAL_221;
  wire  _EVAL_145;
  wire  _EVAL_173;
  wire  _EVAL_47;
  wire  _EVAL_247;
  wire  _EVAL_246;
  wire  _EVAL_191;
  wire  _EVAL_263;
  wire [7:0] _EVAL_209;
  wire  _EVAL_71;
  wire [31:0] _EVAL_273;
  wire [7:0] _EVAL_177;
  wire [7:0] _EVAL_86;
  wire  _EVAL_248;
  wire  _EVAL_43;
  wire  _EVAL_41;
  wire [31:0] _EVAL_293;
  wire  _EVAL_252;
  SiFive__EVAL_237 Repeater (
    ._EVAL(Repeater__EVAL),
    ._EVAL_0(Repeater__EVAL_0),
    ._EVAL_1(Repeater__EVAL_1),
    ._EVAL_2(Repeater__EVAL_2),
    ._EVAL_3(Repeater__EVAL_3),
    ._EVAL_4(Repeater__EVAL_4),
    ._EVAL_5(Repeater__EVAL_5),
    ._EVAL_6(Repeater__EVAL_6),
    ._EVAL_7(Repeater__EVAL_7),
    ._EVAL_8(Repeater__EVAL_8),
    ._EVAL_9(Repeater__EVAL_9),
    ._EVAL_10(Repeater__EVAL_10),
    ._EVAL_11(Repeater__EVAL_11),
    ._EVAL_12(Repeater__EVAL_12),
    ._EVAL_13(Repeater__EVAL_13)
  );
  assign _EVAL_117 = _EVAL_4[2];
  assign _EVAL_235 = _EVAL_4[1];
  assign _EVAL_66 = _EVAL_117 & _EVAL_235;
  assign _EVAL_30 = _EVAL_4[0];
  assign _EVAL_137 = _EVAL_30 == 1'h0;
  assign _EVAL_285 = _EVAL_66 & _EVAL_137;
  assign _EVAL_202 = _EVAL_5[2];
  assign _EVAL_133 = _EVAL_202 == 1'h0;
  assign _EVAL_93 = 10'h7 << _EVAL_16;
  assign _EVAL_172 = _EVAL_93[2:0];
  assign _EVAL_171 = ~ _EVAL_172;
  assign _EVAL_184 = _EVAL_171[2:2];
  assign _EVAL_231 = _EVAL_227 == _EVAL_184;
  assign _EVAL_180 = _EVAL_133 == 1'h0;
  assign _EVAL_224 = _EVAL_231 | _EVAL_180;
  assign _EVAL_175 = _EVAL_224 == 1'h0;
  assign _EVAL_106 = _EVAL_26 | _EVAL_175;
  assign _EVAL_36 = Repeater__EVAL_4;
  assign _EVAL_208 = 7'h1 == _EVAL_36 ? _EVAL_90 : _EVAL_153;
  assign _EVAL_277 = 7'h2 == _EVAL_36 ? _EVAL_78 : _EVAL_208;
  assign _EVAL_110 = 7'h3 == _EVAL_36 ? _EVAL_76 : _EVAL_277;
  assign _EVAL_77 = 7'h4 == _EVAL_36 ? _EVAL_54 : _EVAL_110;
  assign _EVAL_257 = 7'h5 == _EVAL_36 ? _EVAL_182 : _EVAL_77;
  assign _EVAL_239 = 7'h6 == _EVAL_36 ? _EVAL_294 : _EVAL_257;
  assign _EVAL_60 = 7'h7 == _EVAL_36 ? _EVAL_253 : _EVAL_239;
  assign _EVAL_176 = 7'h8 == _EVAL_36 ? _EVAL_154 : _EVAL_60;
  assign _EVAL_72 = 7'h9 == _EVAL_36 ? _EVAL_214 : _EVAL_176;
  assign _EVAL_65 = 7'ha == _EVAL_36 ? _EVAL_44 : _EVAL_72;
  assign _EVAL_206 = 7'hb == _EVAL_36 ? _EVAL_103 : _EVAL_65;
  assign _EVAL_57 = 7'hc == _EVAL_36 ? _EVAL_142 : _EVAL_206;
  assign _EVAL_275 = 7'hd == _EVAL_36 ? _EVAL_280 : _EVAL_57;
  assign _EVAL_31 = 7'he == _EVAL_36 ? _EVAL_91 : _EVAL_275;
  assign _EVAL_75 = 7'hf == _EVAL_36 ? _EVAL_127 : _EVAL_31;
  assign _EVAL_29 = 7'h10 == _EVAL_36 ? _EVAL_287 : _EVAL_75;
  assign _EVAL_141 = 7'h11 == _EVAL_36 ? _EVAL_255 : _EVAL_29;
  assign _EVAL_125 = 7'h12 == _EVAL_36 ? _EVAL_258 : _EVAL_141;
  assign _EVAL_158 = 7'h13 == _EVAL_36 ? _EVAL_281 : _EVAL_125;
  assign _EVAL_283 = 7'h14 == _EVAL_36 ? _EVAL_115 : _EVAL_158;
  assign _EVAL_174 = 7'h15 == _EVAL_36 ? _EVAL_98 : _EVAL_283;
  assign _EVAL_156 = 7'h16 == _EVAL_36 ? _EVAL_244 : _EVAL_174;
  assign _EVAL_201 = 7'h17 == _EVAL_36 ? _EVAL_165 : _EVAL_156;
  assign _EVAL_225 = 7'h18 == _EVAL_36 ? _EVAL_155 : _EVAL_201;
  assign _EVAL_48 = 7'h19 == _EVAL_36 ? _EVAL_292 : _EVAL_225;
  assign _EVAL_178 = 7'h1a == _EVAL_36 ? _EVAL_147 : _EVAL_48;
  assign _EVAL_113 = 7'h1b == _EVAL_36 ? _EVAL_211 : _EVAL_178;
  assign _EVAL_242 = 7'h1c == _EVAL_36 ? _EVAL_69 : _EVAL_113;
  assign _EVAL_237 = 7'h1d == _EVAL_36 ? _EVAL_194 : _EVAL_242;
  assign _EVAL_268 = 7'h1e == _EVAL_36 ? _EVAL_118 : _EVAL_237;
  assign _EVAL_261 = 7'h1f == _EVAL_36 ? _EVAL_87 : _EVAL_268;
  assign _EVAL_265 = 7'h20 == _EVAL_36 ? _EVAL_49 : _EVAL_261;
  assign _EVAL_102 = 7'h21 == _EVAL_36 ? 1'h0 : _EVAL_265;
  assign _EVAL_168 = 7'h22 == _EVAL_36 ? 1'h0 : _EVAL_102;
  assign _EVAL_228 = 7'h23 == _EVAL_36 ? 1'h0 : _EVAL_168;
  assign _EVAL_139 = 7'h24 == _EVAL_36 ? 1'h0 : _EVAL_228;
  assign _EVAL_162 = 7'h25 == _EVAL_36 ? 1'h0 : _EVAL_139;
  assign _EVAL_215 = 7'h26 == _EVAL_36 ? 1'h0 : _EVAL_162;
  assign _EVAL_73 = 7'h27 == _EVAL_36 ? 1'h0 : _EVAL_215;
  assign _EVAL_121 = 7'h28 == _EVAL_36 ? 1'h0 : _EVAL_73;
  assign _EVAL_124 = 7'h29 == _EVAL_36 ? 1'h0 : _EVAL_121;
  assign _EVAL_33 = 7'h2a == _EVAL_36 ? 1'h0 : _EVAL_124;
  assign _EVAL_240 = _EVAL_16[1:0];
  assign _EVAL_190 = 4'h1 << _EVAL_240;
  assign _EVAL_39 = _EVAL_190[2:0];
  assign _EVAL_68 = _EVAL_39 | 3'h1;
  assign _EVAL_143 = _EVAL_68[2];
  assign _EVAL_160 = _EVAL_16 >= 3'h3;
  assign _EVAL_167 = _EVAL_143 & _EVAL_117;
  assign _EVAL_286 = _EVAL_160 | _EVAL_167;
  assign _EVAL_67 = _EVAL_51 + 1'h1;
  assign _EVAL_83 = 7'h2b == _EVAL_36 ? 1'h0 : _EVAL_33;
  assign _EVAL_256 = 7'h2c == _EVAL_36 ? 1'h0 : _EVAL_83;
  assign _EVAL_212 = 7'h2d == _EVAL_36 ? 1'h0 : _EVAL_256;
  assign _EVAL_181 = 7'h2e == _EVAL_36 ? 1'h0 : _EVAL_212;
  assign _EVAL_59 = 7'h2f == _EVAL_36 ? 1'h0 : _EVAL_181;
  assign _EVAL_238 = 7'h30 == _EVAL_36 ? 1'h0 : _EVAL_59;
  assign _EVAL_157 = 7'h31 == _EVAL_36 ? 1'h0 : _EVAL_238;
  assign _EVAL_97 = 7'h32 == _EVAL_36 ? 1'h0 : _EVAL_157;
  assign _EVAL_135 = 7'h33 == _EVAL_36 ? 1'h0 : _EVAL_97;
  assign _EVAL_186 = 7'h34 == _EVAL_36 ? 1'h0 : _EVAL_135;
  assign _EVAL_272 = 7'h35 == _EVAL_36 ? 1'h0 : _EVAL_186;
  assign _EVAL_84 = 7'h36 == _EVAL_36 ? 1'h0 : _EVAL_272;
  assign _EVAL_267 = 7'h37 == _EVAL_36 ? 1'h0 : _EVAL_84;
  assign _EVAL_74 = 7'h38 == _EVAL_36 ? 1'h0 : _EVAL_267;
  assign _EVAL_159 = 7'h39 == _EVAL_36 ? 1'h0 : _EVAL_74;
  assign _EVAL_79 = 7'h3a == _EVAL_36 ? 1'h0 : _EVAL_159;
  assign _EVAL_63 = 7'h3b == _EVAL_36 ? 1'h0 : _EVAL_79;
  assign _EVAL_112 = 7'h3c == _EVAL_36 ? 1'h0 : _EVAL_63;
  assign _EVAL_144 = 7'h3d == _EVAL_36 ? 1'h0 : _EVAL_112;
  assign _EVAL_131 = 7'h3e == _EVAL_36 ? 1'h0 : _EVAL_144;
  assign _EVAL_119 = 7'h3f == _EVAL_36 ? 1'h0 : _EVAL_131;
  assign _EVAL_134 = 7'h40 == _EVAL_36 ? _EVAL_198 : _EVAL_119;
  assign _EVAL_138 = 7'h41 == _EVAL_36 ? _EVAL_52 : _EVAL_134;
  assign _EVAL_164 = 7'h42 == _EVAL_36 ? _EVAL_203 : _EVAL_138;
  assign _EVAL_282 = 7'h43 == _EVAL_36 ? _EVAL_243 : _EVAL_164;
  assign _EVAL_289 = 7'h44 == _EVAL_36 ? _EVAL_104 : _EVAL_282;
  assign _EVAL_226 = Repeater__EVAL_7;
  assign _EVAL_32 = _EVAL_117 == 1'h0;
  assign _EVAL_136 = _EVAL_143 & _EVAL_32;
  assign _EVAL_290 = _EVAL_68[1];
  assign _EVAL_185 = _EVAL_235 == 1'h0;
  assign _EVAL_266 = _EVAL_32 & _EVAL_185;
  assign _EVAL_34 = _EVAL_290 & _EVAL_266;
  assign _EVAL_50 = _EVAL_106 & _EVAL_11;
  assign _EVAL_229 = _EVAL_227 + 1'h1;
  assign _EVAL_234 = Repeater__EVAL_3[63:32];
  assign _EVAL_187 = _EVAL_23[31:0];
  assign _EVAL_88 = {_EVAL_234,_EVAL_187};
  assign _EVAL_233 = _EVAL_88[63:32];
  assign _EVAL_205 = _EVAL_227 & _EVAL_184;
  assign _EVAL_220 = _EVAL_205 == 1'h0;
  assign _EVAL_99 = _EVAL_220 ? _EVAL_17 : _EVAL_116;
  assign _EVAL_279 = _EVAL_117 & _EVAL_185;
  assign _EVAL_61 = _EVAL_290 & _EVAL_279;
  assign _EVAL_195 = _EVAL_286 | _EVAL_61;
  assign _EVAL_92 = Repeater__EVAL_5;
  assign _EVAL_236 = 10'h7 << _EVAL_92;
  assign _EVAL_62 = _EVAL_236[2:0];
  assign _EVAL_183 = ~ _EVAL_62;
  assign _EVAL_192 = _EVAL_183[2:2];
  assign _EVAL_170 = _EVAL_51 == _EVAL_192;
  assign _EVAL_241 = Repeater__EVAL_1;
  assign _EVAL_58 = _EVAL_241[0];
  assign _EVAL_123 = _EVAL_58 == 1'h0;
  assign _EVAL_161 = _EVAL_170 | _EVAL_123;
  assign _EVAL_56 = _EVAL_32 & _EVAL_235;
  assign _EVAL_188 = _EVAL_56 & _EVAL_30;
  assign _EVAL_64 = _EVAL_68[0];
  assign _EVAL_140 = _EVAL_290 & _EVAL_56;
  assign _EVAL_70 = _EVAL_66 & _EVAL_30;
  assign _EVAL_149 = _EVAL_51 == 1'h0;
  assign _EVAL_284 = 7'h45 == _EVAL_36 ? _EVAL_53 : _EVAL_289;
  assign _EVAL_271 = 7'h46 == _EVAL_36 ? _EVAL_80 : _EVAL_284;
  assign _EVAL_100 = 7'h47 == _EVAL_36 ? _EVAL_204 : _EVAL_271;
  assign _EVAL_199 = 7'h48 == _EVAL_36 ? _EVAL_291 : _EVAL_100;
  assign _EVAL_55 = _EVAL_149 ? _EVAL_199 : _EVAL_274;
  assign _EVAL_38 = _EVAL_290 & _EVAL_66;
  assign _EVAL_96 = _EVAL_286 | _EVAL_38;
  assign _EVAL_105 = _EVAL_64 & _EVAL_285;
  assign _EVAL_130 = _EVAL_96 | _EVAL_105;
  assign _EVAL_166 = _EVAL_266 & _EVAL_137;
  assign _EVAL_108 = _EVAL_64 & _EVAL_166;
  assign _EVAL_259 = _EVAL_279 & _EVAL_137;
  assign _EVAL_107 = _EVAL_160 | _EVAL_136;
  assign _EVAL_218 = _EVAL_107 | _EVAL_140;
  assign _EVAL_230 = _EVAL_107 | _EVAL_34;
  assign _EVAL_94 = _EVAL_230 | _EVAL_108;
  assign _EVAL_210 = _EVAL_64 & _EVAL_188;
  assign _EVAL_42 = _EVAL_64 & _EVAL_70;
  assign _EVAL_260 = _EVAL_96 | _EVAL_42;
  assign _EVAL_196 = _EVAL_279 & _EVAL_30;
  assign _EVAL_81 = _EVAL_64 & _EVAL_196;
  assign _EVAL_132 = _EVAL_195 | _EVAL_81;
  assign _EVAL_95 = _EVAL_64 & _EVAL_259;
  assign _EVAL_221 = _EVAL_195 | _EVAL_95;
  assign _EVAL_145 = _EVAL_218 | _EVAL_210;
  assign _EVAL_173 = _EVAL_56 & _EVAL_137;
  assign _EVAL_47 = _EVAL_64 & _EVAL_173;
  assign _EVAL_247 = _EVAL_218 | _EVAL_47;
  assign _EVAL_246 = _EVAL_266 & _EVAL_30;
  assign _EVAL_191 = _EVAL_64 & _EVAL_246;
  assign _EVAL_263 = _EVAL_230 | _EVAL_191;
  assign _EVAL_209 = {_EVAL_260,_EVAL_130,_EVAL_132,_EVAL_221,_EVAL_145,_EVAL_247,_EVAL_263,_EVAL_94};
  assign _EVAL_71 = _EVAL_20 & _EVAL_226;
  assign _EVAL_273 = _EVAL_88[31:0];
  assign _EVAL_177 = {_EVAL_17,_EVAL_99};
  assign _EVAL_86 = _EVAL_133 ? _EVAL_177 : 8'hff;
  assign _EVAL_248 = ~ _EVAL_192;
  assign _EVAL_43 = _EVAL_55 & _EVAL_248;
  assign _EVAL_41 = _EVAL_43 | _EVAL_51;
  assign _EVAL_293 = _EVAL_220 ? _EVAL_24 : _EVAL_114;
  assign _EVAL_252 = _EVAL_50 & _EVAL_175;
  assign _EVAL_27 = Repeater__EVAL_11;
  assign _EVAL_10 = Repeater__EVAL_7;
  assign Repeater__EVAL_2 = _EVAL_20;
  assign _EVAL_8 = _EVAL_26 | _EVAL_175;
  assign _EVAL_6 = _EVAL_209 & _EVAL_86;
  assign Repeater__EVAL_6 = _EVAL_23;
  assign _EVAL_15 = _EVAL_21;
  assign _EVAL_0 = {_EVAL_24,_EVAL_293};
  assign _EVAL = Repeater__EVAL_1;
  assign _EVAL_18 = Repeater__EVAL_4;
  assign Repeater__EVAL_12 = _EVAL_3;
  assign Repeater__EVAL_8 = _EVAL_25;
  assign Repeater__EVAL_0 = _EVAL_13;
  assign _EVAL_22 = Repeater__EVAL_5;
  assign _EVAL_28 = _EVAL_41 ? _EVAL_233 : _EVAL_273;
  assign Repeater__EVAL_13 = _EVAL_161 == 1'h0;
  assign Repeater__EVAL_10 = _EVAL_12;
  assign _EVAL_2 = _EVAL_16;
  assign _EVAL_14 = _EVAL_4;
  assign Repeater__EVAL_9 = _EVAL_1;
  assign _EVAL_7 = _EVAL_5;
  assign _EVAL_19 = _EVAL_11 & _EVAL_224;
  assign Repeater__EVAL = _EVAL_9;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_44 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_49 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_51 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_52 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_53 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_54 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_69 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_76 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_78 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_80 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_87 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_90 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_91 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_98 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_103 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_104 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_114 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_115 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_116 = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_118 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_127 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_142 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_147 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_153 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_154 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_155 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_165 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_182 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_194 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_198 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_203 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_204 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_211 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_214 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_227 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_243 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_244 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_253 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_255 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_258 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_274 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_280 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_281 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_287 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_291 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_292 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_294 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_9) begin
    if (_EVAL_50) begin
      if (7'ha == _EVAL_21) begin
        _EVAL_44 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h20 == _EVAL_21) begin
        _EVAL_49 <= _EVAL_117;
      end
    end
    if (_EVAL_12) begin
      _EVAL_51 <= 1'h0;
    end else begin
      if (_EVAL_71) begin
        if (_EVAL_161) begin
          _EVAL_51 <= 1'h0;
        end else begin
          _EVAL_51 <= _EVAL_67;
        end
      end
    end
    if (_EVAL_50) begin
      if (7'h41 == _EVAL_21) begin
        _EVAL_52 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h45 == _EVAL_21) begin
        _EVAL_53 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h4 == _EVAL_21) begin
        _EVAL_54 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h1c == _EVAL_21) begin
        _EVAL_69 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h3 == _EVAL_21) begin
        _EVAL_76 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h2 == _EVAL_21) begin
        _EVAL_78 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h46 == _EVAL_21) begin
        _EVAL_80 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h1f == _EVAL_21) begin
        _EVAL_87 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h1 == _EVAL_21) begin
        _EVAL_90 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'he == _EVAL_21) begin
        _EVAL_91 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h15 == _EVAL_21) begin
        _EVAL_98 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'hb == _EVAL_21) begin
        _EVAL_103 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h44 == _EVAL_21) begin
        _EVAL_104 <= _EVAL_117;
      end
    end
    if (_EVAL_252) begin
      if (_EVAL_220) begin
        _EVAL_114 <= _EVAL_24;
      end
    end
    if (_EVAL_50) begin
      if (7'h14 == _EVAL_21) begin
        _EVAL_115 <= _EVAL_117;
      end
    end
    if (_EVAL_252) begin
      if (_EVAL_220) begin
        _EVAL_116 <= _EVAL_17;
      end
    end
    if (_EVAL_50) begin
      if (7'h1e == _EVAL_21) begin
        _EVAL_118 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'hf == _EVAL_21) begin
        _EVAL_127 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'hc == _EVAL_21) begin
        _EVAL_142 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h1a == _EVAL_21) begin
        _EVAL_147 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h0 == _EVAL_21) begin
        _EVAL_153 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h8 == _EVAL_21) begin
        _EVAL_154 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h18 == _EVAL_21) begin
        _EVAL_155 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h17 == _EVAL_21) begin
        _EVAL_165 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h5 == _EVAL_21) begin
        _EVAL_182 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h1d == _EVAL_21) begin
        _EVAL_194 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h40 == _EVAL_21) begin
        _EVAL_198 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h42 == _EVAL_21) begin
        _EVAL_203 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h47 == _EVAL_21) begin
        _EVAL_204 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h1b == _EVAL_21) begin
        _EVAL_211 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h9 == _EVAL_21) begin
        _EVAL_214 <= _EVAL_117;
      end
    end
    if (_EVAL_12) begin
      _EVAL_227 <= 1'h0;
    end else begin
      if (_EVAL_50) begin
        if (_EVAL_224) begin
          _EVAL_227 <= 1'h0;
        end else begin
          _EVAL_227 <= _EVAL_229;
        end
      end
    end
    if (_EVAL_50) begin
      if (7'h43 == _EVAL_21) begin
        _EVAL_243 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h16 == _EVAL_21) begin
        _EVAL_244 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h7 == _EVAL_21) begin
        _EVAL_253 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h11 == _EVAL_21) begin
        _EVAL_255 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h12 == _EVAL_21) begin
        _EVAL_258 <= _EVAL_117;
      end
    end
    if (_EVAL_149) begin
      if (7'h48 == _EVAL_36) begin
        _EVAL_274 <= _EVAL_291;
      end else begin
        if (7'h47 == _EVAL_36) begin
          _EVAL_274 <= _EVAL_204;
        end else begin
          if (7'h46 == _EVAL_36) begin
            _EVAL_274 <= _EVAL_80;
          end else begin
            if (7'h45 == _EVAL_36) begin
              _EVAL_274 <= _EVAL_53;
            end else begin
              if (7'h44 == _EVAL_36) begin
                _EVAL_274 <= _EVAL_104;
              end else begin
                if (7'h43 == _EVAL_36) begin
                  _EVAL_274 <= _EVAL_243;
                end else begin
                  if (7'h42 == _EVAL_36) begin
                    _EVAL_274 <= _EVAL_203;
                  end else begin
                    if (7'h41 == _EVAL_36) begin
                      _EVAL_274 <= _EVAL_52;
                    end else begin
                      if (7'h40 == _EVAL_36) begin
                        _EVAL_274 <= _EVAL_198;
                      end else begin
                        if (7'h3f == _EVAL_36) begin
                          _EVAL_274 <= 1'h0;
                        end else begin
                          if (7'h3e == _EVAL_36) begin
                            _EVAL_274 <= 1'h0;
                          end else begin
                            if (7'h3d == _EVAL_36) begin
                              _EVAL_274 <= 1'h0;
                            end else begin
                              if (7'h3c == _EVAL_36) begin
                                _EVAL_274 <= 1'h0;
                              end else begin
                                if (7'h3b == _EVAL_36) begin
                                  _EVAL_274 <= 1'h0;
                                end else begin
                                  if (7'h3a == _EVAL_36) begin
                                    _EVAL_274 <= 1'h0;
                                  end else begin
                                    if (7'h39 == _EVAL_36) begin
                                      _EVAL_274 <= 1'h0;
                                    end else begin
                                      if (7'h38 == _EVAL_36) begin
                                        _EVAL_274 <= 1'h0;
                                      end else begin
                                        if (7'h37 == _EVAL_36) begin
                                          _EVAL_274 <= 1'h0;
                                        end else begin
                                          if (7'h36 == _EVAL_36) begin
                                            _EVAL_274 <= 1'h0;
                                          end else begin
                                            if (7'h35 == _EVAL_36) begin
                                              _EVAL_274 <= 1'h0;
                                            end else begin
                                              if (7'h34 == _EVAL_36) begin
                                                _EVAL_274 <= 1'h0;
                                              end else begin
                                                if (7'h33 == _EVAL_36) begin
                                                  _EVAL_274 <= 1'h0;
                                                end else begin
                                                  if (7'h32 == _EVAL_36) begin
                                                    _EVAL_274 <= 1'h0;
                                                  end else begin
                                                    if (7'h31 == _EVAL_36) begin
                                                      _EVAL_274 <= 1'h0;
                                                    end else begin
                                                      if (7'h30 == _EVAL_36) begin
                                                        _EVAL_274 <= 1'h0;
                                                      end else begin
                                                        if (7'h2f == _EVAL_36) begin
                                                          _EVAL_274 <= 1'h0;
                                                        end else begin
                                                          if (7'h2e == _EVAL_36) begin
                                                            _EVAL_274 <= 1'h0;
                                                          end else begin
                                                            if (7'h2d == _EVAL_36) begin
                                                              _EVAL_274 <= 1'h0;
                                                            end else begin
                                                              if (7'h2c == _EVAL_36) begin
                                                                _EVAL_274 <= 1'h0;
                                                              end else begin
                                                                if (7'h2b == _EVAL_36) begin
                                                                  _EVAL_274 <= 1'h0;
                                                                end else begin
                                                                  if (7'h2a == _EVAL_36) begin
                                                                    _EVAL_274 <= 1'h0;
                                                                  end else begin
                                                                    if (7'h29 == _EVAL_36) begin
                                                                      _EVAL_274 <= 1'h0;
                                                                    end else begin
                                                                      if (7'h28 == _EVAL_36) begin
                                                                        _EVAL_274 <= 1'h0;
                                                                      end else begin
                                                                        if (7'h27 == _EVAL_36) begin
                                                                          _EVAL_274 <= 1'h0;
                                                                        end else begin
                                                                          if (7'h26 == _EVAL_36) begin
                                                                            _EVAL_274 <= 1'h0;
                                                                          end else begin
                                                                            if (7'h25 == _EVAL_36) begin
                                                                              _EVAL_274 <= 1'h0;
                                                                            end else begin
                                                                              if (7'h24 == _EVAL_36) begin
                                                                                _EVAL_274 <= 1'h0;
                                                                              end else begin
                                                                                if (7'h23 == _EVAL_36) begin
                                                                                  _EVAL_274 <= 1'h0;
                                                                                end else begin
                                                                                  if (7'h22 == _EVAL_36) begin
                                                                                    _EVAL_274 <= 1'h0;
                                                                                  end else begin
                                                                                    if (7'h21 == _EVAL_36) begin
                                                                                      _EVAL_274 <= 1'h0;
                                                                                    end else begin
                                                                                      if (7'h20 == _EVAL_36) begin
                                                                                        _EVAL_274 <= _EVAL_49;
                                                                                      end else begin
                                                                                        if (7'h1f == _EVAL_36) begin
                                                                                          _EVAL_274 <= _EVAL_87;
                                                                                        end else begin
                                                                                          if (7'h1e == _EVAL_36) begin
                                                                                            _EVAL_274 <= _EVAL_118;
                                                                                          end else begin
                                                                                            if (7'h1d == _EVAL_36) begin
                                                                                              _EVAL_274 <= _EVAL_194;
                                                                                            end else begin
                                                                                              if (7'h1c == _EVAL_36) begin
                                                                                                _EVAL_274 <= _EVAL_69;
                                                                                              end else begin
                                                                                                if (7'h1b == _EVAL_36) begin
                                                                                                  _EVAL_274 <= _EVAL_211;
                                                                                                end else begin
                                                                                                  if (7'h1a == _EVAL_36) begin
                                                                                                    _EVAL_274 <= _EVAL_147;
                                                                                                  end else begin
                                                                                                    if (7'h19 == _EVAL_36) begin
                                                                                                      _EVAL_274 <= _EVAL_292;
                                                                                                    end else begin
                                                                                                      if (7'h18 == _EVAL_36) begin
                                                                                                        _EVAL_274 <= _EVAL_155;
                                                                                                      end else begin
                                                                                                        if (7'h17 == _EVAL_36) begin
                                                                                                          _EVAL_274 <= _EVAL_165;
                                                                                                        end else begin
                                                                                                          if (7'h16 == _EVAL_36) begin
                                                                                                            _EVAL_274 <= _EVAL_244;
                                                                                                          end else begin
                                                                                                            if (7'h15 == _EVAL_36) begin
                                                                                                              _EVAL_274 <= _EVAL_98;
                                                                                                            end else begin
                                                                                                              if (7'h14 == _EVAL_36) begin
                                                                                                                _EVAL_274 <= _EVAL_115;
                                                                                                              end else begin
                                                                                                                if (7'h13 == _EVAL_36) begin
                                                                                                                  _EVAL_274 <= _EVAL_281;
                                                                                                                end else begin
                                                                                                                  if (7'h12 == _EVAL_36) begin
                                                                                                                    _EVAL_274 <= _EVAL_258;
                                                                                                                  end else begin
                                                                                                                    if (7'h11 == _EVAL_36) begin
                                                                                                                      _EVAL_274 <= _EVAL_255;
                                                                                                                    end else begin
                                                                                                                      if (7'h10 == _EVAL_36) begin
                                                                                                                        _EVAL_274 <= _EVAL_287;
                                                                                                                      end else begin
                                                                                                                        if (7'hf == _EVAL_36) begin
                                                                                                                          _EVAL_274 <= _EVAL_127;
                                                                                                                        end else begin
                                                                                                                          if (7'he == _EVAL_36) begin
                                                                                                                            _EVAL_274 <= _EVAL_91;
                                                                                                                          end else begin
                                                                                                                            if (7'hd == _EVAL_36) begin
                                                                                                                              _EVAL_274 <= _EVAL_280;
                                                                                                                            end else begin
                                                                                                                              if (7'hc == _EVAL_36) begin
                                                                                                                                _EVAL_274 <= _EVAL_142;
                                                                                                                              end else begin
                                                                                                                                if (7'hb == _EVAL_36) begin
                                                                                                                                  _EVAL_274 <= _EVAL_103;
                                                                                                                                end else begin
                                                                                                                                  if (7'ha == _EVAL_36) begin
                                                                                                                                    _EVAL_274 <= _EVAL_44;
                                                                                                                                  end else begin
                                                                                                                                    if (7'h9 == _EVAL_36) begin
                                                                                                                                      _EVAL_274 <= _EVAL_214;
                                                                                                                                    end else begin
                                                                                                                                      if (7'h8 == _EVAL_36) begin
                                                                                                                                        _EVAL_274 <= _EVAL_154;
                                                                                                                                      end else begin
                                                                                                                                        if (7'h7 == _EVAL_36) begin
                                                                                                                                          _EVAL_274 <= _EVAL_253;
                                                                                                                                        end else begin
                                                                                                                                          if (7'h6 == _EVAL_36) begin
                                                                                                                                            _EVAL_274 <= _EVAL_294;
                                                                                                                                          end else begin
                                                                                                                                            if (7'h5 == _EVAL_36) begin
                                                                                                                                              _EVAL_274 <= _EVAL_182;
                                                                                                                                            end else begin
                                                                                                                                              if (7'h4 == _EVAL_36) begin
                                                                                                                                                _EVAL_274 <= _EVAL_54;
                                                                                                                                              end else begin
                                                                                                                                                if (7'h3 == _EVAL_36) begin
                                                                                                                                                  _EVAL_274 <= _EVAL_76;
                                                                                                                                                end else begin
                                                                                                                                                  if (7'h2 == _EVAL_36) begin
                                                                                                                                                    _EVAL_274 <= _EVAL_78;
                                                                                                                                                  end else begin
                                                                                                                                                    if (7'h1 == _EVAL_36) begin
                                                                                                                                                      _EVAL_274 <= _EVAL_90;
                                                                                                                                                    end else begin
                                                                                                                                                      _EVAL_274 <= _EVAL_153;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_50) begin
      if (7'hd == _EVAL_21) begin
        _EVAL_280 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h13 == _EVAL_21) begin
        _EVAL_281 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h10 == _EVAL_21) begin
        _EVAL_287 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h48 == _EVAL_21) begin
        _EVAL_291 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h19 == _EVAL_21) begin
        _EVAL_292 <= _EVAL_117;
      end
    end
    if (_EVAL_50) begin
      if (7'h6 == _EVAL_21) begin
        _EVAL_294 <= _EVAL_117;
      end
    end
  end
endmodule
