//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_130_assert(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [27:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [6:0]  _EVAL_8,
  input  [6:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [72:0] _EVAL_38;
  reg [95:0] _RAND_0;
  reg [27:0] _EVAL_44;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_117;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_124;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_133;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_144;
  reg [31:0] _RAND_5;
  reg [6:0] _EVAL_198;
  reg [31:0] _RAND_6;
  reg [6:0] _EVAL_204;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_209;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_228;
  reg [31:0] _RAND_9;
  reg [31:0] _EVAL_235;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_254;
  reg [31:0] _RAND_11;
  reg [3:0] _EVAL_286;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_287;
  reg [31:0] _RAND_13;
  wire  _EVAL_188;
  wire  _EVAL_282;
  wire  _EVAL_266;
  wire [12:0] _EVAL_248;
  wire [5:0] _EVAL_269;
  wire [5:0] _EVAL_241;
  wire [3:0] _EVAL_160;
  wire  _EVAL_103;
  wire  _EVAL_113;
  wire  _EVAL_118;
  wire  _EVAL_141;
  wire  _EVAL_120;
  wire  _EVAL_201;
  wire  _EVAL_104;
  wire  _EVAL_108;
  wire  _EVAL_157;
  wire  _EVAL_86;
  wire  _EVAL_191;
  wire  _EVAL_202;
  wire [31:0] _EVAL_55;
  wire  _EVAL_142;
  wire  _EVAL_46;
  wire  _EVAL_162;
  wire  _EVAL_255;
  wire  _EVAL_181;
  wire [3:0] _EVAL_213;
  wire  _EVAL_262;
  wire [2:0] _EVAL_26;
  wire  _EVAL_130;
  wire  _EVAL_21;
  wire  _EVAL_159;
  wire  _EVAL_154;
  wire  _EVAL_219;
  wire  _EVAL_132;
  wire  _EVAL_170;
  wire  _EVAL_183;
  wire  _EVAL_275;
  wire  _EVAL_40;
  wire  _EVAL_166;
  wire  _EVAL_33;
  wire  _EVAL_182;
  wire  _EVAL_83;
  wire  _EVAL_123;
  wire  _EVAL_62;
  wire  _EVAL_152;
  wire  _EVAL_242;
  wire  _EVAL_131;
  wire [27:0] _EVAL_177;
  wire [27:0] _EVAL_91;
  wire  _EVAL_85;
  wire [3:0] _EVAL_51;
  wire  _EVAL_127;
  wire  _EVAL_121;
  wire [1:0] _EVAL_52;
  wire [1:0] _EVAL_64;
  wire  _EVAL_110;
  wire  _EVAL_47;
  wire  _EVAL_99;
  wire  _EVAL_218;
  wire  _EVAL_258;
  wire  _EVAL_185;
  wire  _EVAL_259;
  wire  _EVAL_116;
  wire [3:0] _EVAL_70;
  wire  _EVAL_176;
  wire  _EVAL_109;
  wire  _EVAL_216;
  wire  _EVAL_54;
  wire  _EVAL_264;
  wire  _EVAL_25;
  wire  _EVAL_252;
  wire  _EVAL_97;
  wire  _EVAL_236;
  wire  _EVAL_39;
  wire  _EVAL_73;
  wire  _EVAL_164;
  wire  _EVAL_207;
  wire  _EVAL_283;
  wire  _EVAL_178;
  wire  _EVAL_126;
  wire  _EVAL_245;
  wire  _EVAL_59;
  wire  _EVAL_221;
  wire  _EVAL_153;
  wire  _EVAL_187;
  wire  _EVAL_172;
  wire  _EVAL_143;
  wire  _EVAL_71;
  wire  _EVAL_76;
  wire [3:0] _EVAL_88;
  wire [3:0] _EVAL_173;
  wire [3:0] _EVAL_224;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_261;
  wire  _EVAL_56;
  wire  _EVAL_156;
  wire  _EVAL_145;
  wire  _EVAL_30;
  wire  _EVAL_23;
  wire [2:0] _EVAL_107;
  wire  _EVAL_273;
  wire  _EVAL_253;
  wire  _EVAL_122;
  wire  _EVAL_281;
  wire  _EVAL_89;
  wire  _EVAL_134;
  wire  _EVAL_36;
  wire  _EVAL_227;
  wire  _EVAL_214;
  wire  _EVAL_135;
  wire  _EVAL_238;
  wire  _EVAL_230;
  wire  _EVAL_151;
  wire  _EVAL_257;
  wire  _EVAL_244;
  wire  _EVAL_226;
  wire [12:0] _EVAL_93;
  wire [5:0] _EVAL_284;
  wire [5:0] _EVAL_63;
  wire [3:0] _EVAL_174;
  wire [3:0] _EVAL_24;
  wire  _EVAL_17;
  wire  _EVAL_140;
  wire  _EVAL_60;
  wire  _EVAL_288;
  wire  _EVAL_280;
  wire  _EVAL_50;
  wire  _EVAL_77;
  wire  _EVAL_267;
  wire  _EVAL_58;
  wire  _EVAL_20;
  wire [127:0] _EVAL_171;
  wire [127:0] _EVAL_210;
  wire [72:0] _EVAL_66;
  wire [72:0] _EVAL_84;
  wire [72:0] _EVAL_277;
  wire  _EVAL_37;
  wire  _EVAL_94;
  wire [127:0] _EVAL_41;
  wire [127:0] _EVAL_270;
  wire [72:0] _EVAL_112;
  wire  _EVAL_92;
  wire  _EVAL_212;
  wire  _EVAL_203;
  wire  _EVAL_278;
  wire  _EVAL_69;
  wire  _EVAL_175;
  wire  _EVAL_81;
  wire  _EVAL_197;
  wire [27:0] _EVAL_48;
  wire [72:0] _EVAL_279;
  wire  _EVAL_82;
  wire  _EVAL_150;
  wire  _EVAL_193;
  wire  _EVAL_95;
  wire [28:0] _EVAL_87;
  wire [28:0] _EVAL_106;
  wire [28:0] _EVAL_146;
  wire  _EVAL_67;
  wire  _EVAL_158;
  wire  _EVAL_222;
  wire  _EVAL_234;
  wire  _EVAL_272;
  wire  _EVAL_240;
  wire  _EVAL_32;
  wire  _EVAL_239;
  wire  _EVAL_163;
  wire  _EVAL_29;
  wire  _EVAL_229;
  wire  _EVAL_196;
  wire [72:0] _EVAL_225;
  wire [72:0] _EVAL_43;
  wire [72:0] _EVAL_190;
  wire  _EVAL_79;
  wire  _EVAL_90;
  wire  _EVAL_249;
  wire  _EVAL_167;
  wire  _EVAL_31;
  wire  _EVAL_208;
  wire  _EVAL_80;
  wire  _EVAL_215;
  wire  _EVAL_199;
  wire  _EVAL_165;
  wire  _EVAL_194;
  wire [3:0] _EVAL_195;
  wire [3:0] _EVAL_206;
  wire  _EVAL_28;
  wire  _EVAL_78;
  wire  _EVAL_205;
  wire  _EVAL_128;
  wire  _EVAL_276;
  wire  _EVAL_75;
  wire  _EVAL_200;
  wire  _EVAL_22;
  wire  _EVAL_136;
  wire  _EVAL_102;
  wire  _EVAL_100;
  wire  _EVAL_139;
  wire  _EVAL_45;
  wire  _EVAL_98;
  wire  _EVAL_161;
  wire  _EVAL_256;
  wire  _EVAL_250;
  wire  _EVAL_148;
  wire  _EVAL_211;
  wire  _EVAL_155;
  wire  _EVAL_168;
  wire  _EVAL_179;
  wire  _EVAL_19;
  wire  _EVAL_263;
  wire  _EVAL_260;
  wire  _EVAL_251;
  wire  _EVAL_180;
  wire  _EVAL_217;
  wire  _EVAL_265;
  wire  _EVAL_111;
  wire  _EVAL_114;
  wire  _EVAL_247;
  wire  _EVAL_105;
  wire  _EVAL_57;
  wire  _EVAL_101;
  wire  _EVAL_268;
  wire  _EVAL_68;
  wire  _EVAL_237;
  wire  _EVAL_189;
  wire  _EVAL_65;
  wire  _EVAL_149;
  wire  _EVAL_147;
  wire  _EVAL_137;
  wire  _EVAL_186;
  wire [3:0] _EVAL_274;
  wire  _EVAL_115;
  wire  _EVAL_192;
  wire  _EVAL_285;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_184;
  wire  _EVAL_138;
  wire  _EVAL_233;
  wire  _EVAL_42;
  wire  _EVAL_271;
  wire  _EVAL_53;
  wire  _EVAL_49;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_188 = _EVAL_0 == 3'h1;
  assign _EVAL_282 = _EVAL_0[2];
  assign _EVAL_266 = _EVAL_282 == 1'h0;
  assign _EVAL_248 = 13'h3f << _EVAL_1;
  assign _EVAL_269 = _EVAL_248[5:0];
  assign _EVAL_241 = ~ _EVAL_269;
  assign _EVAL_160 = _EVAL_241[5:2];
  assign _EVAL_103 = _EVAL_14 == 3'h4;
  assign _EVAL_113 = _EVAL_6 & _EVAL_103;
  assign _EVAL_118 = _EVAL_0 == 3'h5;
  assign _EVAL_141 = _EVAL_12 <= 3'h3;
  assign _EVAL_120 = _EVAL_38 != 73'h0;
  assign _EVAL_201 = _EVAL_120 == 1'h0;
  assign _EVAL_104 = _EVAL_12 == 3'h0;
  assign _EVAL_108 = _EVAL_104 | _EVAL_7;
  assign _EVAL_157 = _EVAL_108 == 1'h0;
  assign _EVAL_86 = _EVAL_3 & _EVAL_13;
  assign _EVAL_191 = _EVAL_5 & _EVAL_6;
  assign _EVAL_202 = _EVAL_86 | _EVAL_191;
  assign _EVAL_55 = _EVAL_235 + 32'h1;
  assign _EVAL_142 = _EVAL_0 == 3'h0;
  assign _EVAL_46 = _EVAL_13 & _EVAL_142;
  assign _EVAL_162 = _EVAL_9 == 7'h48;
  assign _EVAL_255 = _EVAL_9 == 7'h40;
  assign _EVAL_181 = _EVAL_162 | _EVAL_255;
  assign _EVAL_213 = _EVAL_9[6:3];
  assign _EVAL_262 = _EVAL_213 == 4'h8;
  assign _EVAL_26 = _EVAL_9[2:0];
  assign _EVAL_130 = 3'h1 <= _EVAL_26;
  assign _EVAL_21 = _EVAL_262 & _EVAL_130;
  assign _EVAL_159 = _EVAL_181 | _EVAL_21;
  assign _EVAL_154 = _EVAL_9 == 7'h20;
  assign _EVAL_219 = _EVAL_159 | _EVAL_154;
  assign _EVAL_132 = _EVAL_213 == 4'h0;
  assign _EVAL_170 = _EVAL_219 | _EVAL_132;
  assign _EVAL_183 = _EVAL_213 == 4'h1;
  assign _EVAL_275 = _EVAL_170 | _EVAL_183;
  assign _EVAL_40 = _EVAL_213 == 4'h2;
  assign _EVAL_166 = _EVAL_275 | _EVAL_40;
  assign _EVAL_33 = _EVAL_213 == 4'h3;
  assign _EVAL_182 = _EVAL_166 | _EVAL_33;
  assign _EVAL_83 = _EVAL_182 | _EVAL_7;
  assign _EVAL_123 = _EVAL_209 == 4'h0;
  assign _EVAL_62 = _EVAL_191 & _EVAL_123;
  assign _EVAL_152 = _EVAL_14 == 3'h6;
  assign _EVAL_242 = _EVAL_152 == 1'h0;
  assign _EVAL_131 = _EVAL_62 & _EVAL_242;
  assign _EVAL_177 = {{22'd0}, _EVAL_241};
  assign _EVAL_91 = _EVAL_2 & _EVAL_177;
  assign _EVAL_85 = _EVAL_91 == 28'h0;
  assign _EVAL_51 = _EVAL_209 - 4'h1;
  assign _EVAL_127 = _EVAL_12 != 3'h0;
  assign _EVAL_121 = _EVAL_1[0];
  assign _EVAL_52 = 2'h1 << _EVAL_121;
  assign _EVAL_64 = _EVAL_52 | 2'h1;
  assign _EVAL_110 = _EVAL_64[0];
  assign _EVAL_47 = _EVAL_2[1];
  assign _EVAL_99 = _EVAL_47 == 1'h0;
  assign _EVAL_218 = _EVAL_2[0];
  assign _EVAL_258 = _EVAL_99 & _EVAL_218;
  assign _EVAL_185 = _EVAL_110 & _EVAL_258;
  assign _EVAL_259 = _EVAL_47 & _EVAL_218;
  assign _EVAL_116 = _EVAL_110 & _EVAL_259;
  assign _EVAL_70 = _EVAL_8[6:3];
  assign _EVAL_176 = _EVAL_70 == 4'h3;
  assign _EVAL_109 = _EVAL_70 == 4'h2;
  assign _EVAL_216 = _EVAL_286 == 4'h0;
  assign _EVAL_54 = _EVAL_216 == 1'h0;
  assign _EVAL_264 = _EVAL_0 == 3'h6;
  assign _EVAL_25 = _EVAL_13 & _EVAL_264;
  assign _EVAL_252 = _EVAL_9 == _EVAL_204;
  assign _EVAL_97 = _EVAL_252 | _EVAL_7;
  assign _EVAL_236 = _EVAL_97 == 1'h0;
  assign _EVAL_39 = _EVAL_70 == 4'h0;
  assign _EVAL_73 = _EVAL_1 >= 3'h2;
  assign _EVAL_164 = _EVAL_64[1];
  assign _EVAL_207 = _EVAL_164 & _EVAL_47;
  assign _EVAL_283 = _EVAL_73 | _EVAL_207;
  assign _EVAL_178 = _EVAL_283 | _EVAL_116;
  assign _EVAL_126 = _EVAL_218 == 1'h0;
  assign _EVAL_245 = _EVAL_47 & _EVAL_126;
  assign _EVAL_59 = _EVAL_110 & _EVAL_245;
  assign _EVAL_221 = _EVAL_283 | _EVAL_59;
  assign _EVAL_153 = _EVAL_164 & _EVAL_99;
  assign _EVAL_187 = _EVAL_73 | _EVAL_153;
  assign _EVAL_172 = _EVAL_187 | _EVAL_185;
  assign _EVAL_143 = _EVAL_99 & _EVAL_126;
  assign _EVAL_71 = _EVAL_110 & _EVAL_143;
  assign _EVAL_76 = _EVAL_187 | _EVAL_71;
  assign _EVAL_88 = {_EVAL_178,_EVAL_221,_EVAL_172,_EVAL_76};
  assign _EVAL_173 = ~ _EVAL_88;
  assign _EVAL_224 = _EVAL_10 & _EVAL_173;
  assign _EVAL_34 = _EVAL_10 == _EVAL_88;
  assign _EVAL_35 = _EVAL_34 | _EVAL_7;
  assign _EVAL_261 = _EVAL_14 == 3'h2;
  assign _EVAL_56 = _EVAL_14 <= 3'h6;
  assign _EVAL_156 = _EVAL_8 == 7'h48;
  assign _EVAL_145 = _EVAL_8 == 7'h40;
  assign _EVAL_30 = _EVAL_156 | _EVAL_145;
  assign _EVAL_23 = _EVAL_70 == 4'h8;
  assign _EVAL_107 = _EVAL_8[2:0];
  assign _EVAL_273 = 3'h1 <= _EVAL_107;
  assign _EVAL_253 = _EVAL_23 & _EVAL_273;
  assign _EVAL_122 = _EVAL_30 | _EVAL_253;
  assign _EVAL_281 = _EVAL_8 == 7'h20;
  assign _EVAL_89 = _EVAL_122 | _EVAL_281;
  assign _EVAL_134 = _EVAL_89 | _EVAL_39;
  assign _EVAL_36 = _EVAL_70 == 4'h1;
  assign _EVAL_227 = _EVAL_134 | _EVAL_36;
  assign _EVAL_214 = _EVAL_227 | _EVAL_109;
  assign _EVAL_135 = _EVAL_214 | _EVAL_176;
  assign _EVAL_238 = _EVAL_141 | _EVAL_7;
  assign _EVAL_230 = _EVAL_12 == _EVAL_254;
  assign _EVAL_151 = _EVAL_230 | _EVAL_7;
  assign _EVAL_257 = _EVAL_14 == 3'h5;
  assign _EVAL_244 = _EVAL_6 & _EVAL_257;
  assign _EVAL_226 = _EVAL_14[0];
  assign _EVAL_93 = 13'h3f << _EVAL;
  assign _EVAL_284 = _EVAL_93[5:0];
  assign _EVAL_63 = ~ _EVAL_284;
  assign _EVAL_174 = _EVAL_63[5:2];
  assign _EVAL_24 = _EVAL_286 - 4'h1;
  assign _EVAL_17 = _EVAL_1 <= 3'h6;
  assign _EVAL_140 = 3'h6 == _EVAL_1;
  assign _EVAL_60 = _EVAL_145 ? _EVAL_140 : 1'h0;
  assign _EVAL_288 = plusarg_reader_out == 32'h0;
  assign _EVAL_280 = _EVAL_201 | _EVAL_288;
  assign _EVAL_50 = _EVAL_235 < plusarg_reader_out;
  assign _EVAL_77 = _EVAL_280 | _EVAL_50;
  assign _EVAL_267 = _EVAL_77 | _EVAL_7;
  assign _EVAL_58 = _EVAL_144 == 4'h0;
  assign _EVAL_20 = _EVAL_86 & _EVAL_58;
  assign _EVAL_171 = 128'h1 << _EVAL_8;
  assign _EVAL_210 = _EVAL_20 ? _EVAL_171 : 128'h0;
  assign _EVAL_66 = _EVAL_210[72:0];
  assign _EVAL_84 = _EVAL_66 | _EVAL_38;
  assign _EVAL_277 = _EVAL_84 >> _EVAL_9;
  assign _EVAL_37 = _EVAL_277[0];
  assign _EVAL_94 = _EVAL_37 | _EVAL_7;
  assign _EVAL_41 = 128'h1 << _EVAL_9;
  assign _EVAL_270 = _EVAL_131 ? _EVAL_41 : 128'h0;
  assign _EVAL_112 = _EVAL_270[72:0];
  assign _EVAL_92 = _EVAL_66 != _EVAL_112;
  assign _EVAL_212 = _EVAL_66 != 73'h0;
  assign _EVAL_203 = _EVAL_212 == 1'h0;
  assign _EVAL_278 = _EVAL_92 | _EVAL_203;
  assign _EVAL_69 = _EVAL_278 | _EVAL_7;
  assign _EVAL_175 = _EVAL_69 == 1'h0;
  assign _EVAL_81 = _EVAL_6 & _EVAL_261;
  assign _EVAL_197 = _EVAL_13 & _EVAL_188;
  assign _EVAL_48 = _EVAL_2 ^ 28'hc000000;
  assign _EVAL_279 = _EVAL_38 >> _EVAL_8;
  assign _EVAL_82 = _EVAL_279[0];
  assign _EVAL_150 = _EVAL_82 == 1'h0;
  assign _EVAL_193 = _EVAL_150 | _EVAL_7;
  assign _EVAL_95 = _EVAL_193 == 1'h0;
  assign _EVAL_87 = {1'b0,$signed(_EVAL_48)};
  assign _EVAL_106 = $signed(_EVAL_87) & $signed(-29'sh4000000);
  assign _EVAL_146 = $signed(_EVAL_106);
  assign _EVAL_67 = $signed(_EVAL_146) == $signed(29'sh0);
  assign _EVAL_158 = _EVAL_0 == 3'h2;
  assign _EVAL_222 = _EVAL_11 == 1'h0;
  assign _EVAL_234 = _EVAL_73 | _EVAL_7;
  assign _EVAL_272 = _EVAL_234 == 1'h0;
  assign _EVAL_240 = _EVAL_135 | _EVAL_7;
  assign _EVAL_32 = _EVAL_240 == 1'h0;
  assign _EVAL_239 = _EVAL_12 <= 3'h4;
  assign _EVAL_163 = _EVAL_239 | _EVAL_7;
  assign _EVAL_29 = _EVAL_56 | _EVAL_7;
  assign _EVAL_229 = _EVAL_29 == 1'h0;
  assign _EVAL_196 = _EVAL_0 == 3'h3;
  assign _EVAL_225 = _EVAL_38 | _EVAL_66;
  assign _EVAL_43 = ~ _EVAL_112;
  assign _EVAL_190 = _EVAL_225 & _EVAL_43;
  assign _EVAL_79 = _EVAL_14 == 3'h0;
  assign _EVAL_90 = _EVAL_6 & _EVAL_79;
  assign _EVAL_249 = _EVAL_12 <= 3'h2;
  assign _EVAL_167 = _EVAL_249 | _EVAL_7;
  assign _EVAL_31 = _EVAL_60 | _EVAL_7;
  assign _EVAL_208 = _EVAL_17 & _EVAL_67;
  assign _EVAL_80 = _EVAL_208 | _EVAL_7;
  assign _EVAL_215 = _EVAL_2 == _EVAL_44;
  assign _EVAL_199 = _EVAL_267 == 1'h0;
  assign _EVAL_165 = _EVAL_222 | _EVAL_7;
  assign _EVAL_194 = _EVAL >= 3'h2;
  assign _EVAL_195 = _EVAL_144 - 4'h1;
  assign _EVAL_206 = ~ _EVAL_10;
  assign _EVAL_28 = _EVAL_206 == 4'h0;
  assign _EVAL_78 = _EVAL_191 & _EVAL_216;
  assign _EVAL_205 = _EVAL_31 == 1'h0;
  assign _EVAL_128 = _EVAL_124 == 4'h0;
  assign _EVAL_276 = _EVAL_128 == 1'h0;
  assign _EVAL_75 = _EVAL_85 | _EVAL_7;
  assign _EVAL_200 = _EVAL_215 | _EVAL_7;
  assign _EVAL_22 = _EVAL_200 == 1'h0;
  assign _EVAL_136 = _EVAL_224 == 4'h0;
  assign _EVAL_102 = _EVAL_136 | _EVAL_7;
  assign _EVAL_100 = _EVAL_165 == 1'h0;
  assign _EVAL_139 = _EVAL_14 == 3'h1;
  assign _EVAL_45 = _EVAL_6 & _EVAL_152;
  assign _EVAL_98 = _EVAL_75 == 1'h0;
  assign _EVAL_161 = _EVAL_8 == _EVAL_198;
  assign _EVAL_256 = _EVAL_161 | _EVAL_7;
  assign _EVAL_250 = _EVAL == _EVAL_133;
  assign _EVAL_148 = _EVAL_0 == 3'h4;
  assign _EVAL_211 = _EVAL_0 == 3'h7;
  assign _EVAL_155 = _EVAL_0 == _EVAL_287;
  assign _EVAL_168 = _EVAL_155 | _EVAL_7;
  assign _EVAL_179 = _EVAL_13 & _EVAL_148;
  assign _EVAL_19 = _EVAL_80 == 1'h0;
  assign _EVAL_263 = _EVAL_250 | _EVAL_7;
  assign _EVAL_260 = _EVAL_263 == 1'h0;
  assign _EVAL_251 = _EVAL_1 == _EVAL_228;
  assign _EVAL_180 = _EVAL_251 | _EVAL_7;
  assign _EVAL_217 = _EVAL_168 == 1'h0;
  assign _EVAL_265 = _EVAL_151 == 1'h0;
  assign _EVAL_111 = _EVAL_28 | _EVAL_7;
  assign _EVAL_114 = _EVAL_13 & _EVAL_118;
  assign _EVAL_247 = _EVAL_167 == 1'h0;
  assign _EVAL_105 = _EVAL_6 & _EVAL_54;
  assign _EVAL_57 = _EVAL_7 == 1'h0;
  assign _EVAL_101 = _EVAL_13 & _EVAL_276;
  assign _EVAL_268 = _EVAL_13 & _EVAL_196;
  assign _EVAL_68 = _EVAL_180 == 1'h0;
  assign _EVAL_237 = _EVAL_238 == 1'h0;
  assign _EVAL_189 = _EVAL_35 == 1'h0;
  assign _EVAL_65 = _EVAL_127 | _EVAL_7;
  assign _EVAL_149 = _EVAL_65 == 1'h0;
  assign _EVAL_147 = _EVAL_194 | _EVAL_7;
  assign _EVAL_137 = _EVAL_147 == 1'h0;
  assign _EVAL_186 = _EVAL_83 == 1'h0;
  assign _EVAL_274 = _EVAL_124 - 4'h1;
  assign _EVAL_115 = _EVAL_14 == _EVAL_117;
  assign _EVAL_192 = _EVAL_86 & _EVAL_128;
  assign _EVAL_285 = _EVAL_94 == 1'h0;
  assign _EVAL_72 = _EVAL_115 | _EVAL_7;
  assign _EVAL_74 = _EVAL_102 == 1'h0;
  assign _EVAL_184 = _EVAL_13 & _EVAL_211;
  assign _EVAL_138 = _EVAL_13 & _EVAL_158;
  assign _EVAL_233 = _EVAL_163 == 1'h0;
  assign _EVAL_42 = _EVAL_6 & _EVAL_139;
  assign _EVAL_271 = _EVAL_111 == 1'h0;
  assign _EVAL_53 = _EVAL_72 == 1'h0;
  assign _EVAL_49 = _EVAL_256 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  _EVAL_38 = _RAND_0[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_44 = _RAND_1[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_117 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_124 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_133 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_144 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_198 = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_204 = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_209 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_228 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_235 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_254 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_286 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_287 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_7) begin
      _EVAL_38 <= 73'h0;
    end else begin
      _EVAL_38 <= _EVAL_190;
    end
    if (_EVAL_192) begin
      _EVAL_44 <= _EVAL_2;
    end
    if (_EVAL_78) begin
      _EVAL_117 <= _EVAL_14;
    end
    if (_EVAL_7) begin
      _EVAL_124 <= 4'h0;
    end else begin
      if (_EVAL_86) begin
        if (_EVAL_128) begin
          if (_EVAL_266) begin
            _EVAL_124 <= _EVAL_160;
          end else begin
            _EVAL_124 <= 4'h0;
          end
        end else begin
          _EVAL_124 <= _EVAL_274;
        end
      end
    end
    if (_EVAL_78) begin
      _EVAL_133 <= _EVAL;
    end
    if (_EVAL_7) begin
      _EVAL_144 <= 4'h0;
    end else begin
      if (_EVAL_86) begin
        if (_EVAL_58) begin
          if (_EVAL_266) begin
            _EVAL_144 <= _EVAL_160;
          end else begin
            _EVAL_144 <= 4'h0;
          end
        end else begin
          _EVAL_144 <= _EVAL_195;
        end
      end
    end
    if (_EVAL_192) begin
      _EVAL_198 <= _EVAL_8;
    end
    if (_EVAL_78) begin
      _EVAL_204 <= _EVAL_9;
    end
    if (_EVAL_7) begin
      _EVAL_209 <= 4'h0;
    end else begin
      if (_EVAL_191) begin
        if (_EVAL_123) begin
          if (_EVAL_226) begin
            _EVAL_209 <= _EVAL_174;
          end else begin
            _EVAL_209 <= 4'h0;
          end
        end else begin
          _EVAL_209 <= _EVAL_51;
        end
      end
    end
    if (_EVAL_192) begin
      _EVAL_228 <= _EVAL_1;
    end
    if (_EVAL_7) begin
      _EVAL_235 <= 32'h0;
    end else begin
      if (_EVAL_202) begin
        _EVAL_235 <= 32'h0;
      end else begin
        _EVAL_235 <= _EVAL_55;
      end
    end
    if (_EVAL_192) begin
      _EVAL_254 <= _EVAL_12;
    end
    if (_EVAL_7) begin
      _EVAL_286 <= 4'h0;
    end else begin
      if (_EVAL_191) begin
        if (_EVAL_216) begin
          if (_EVAL_226) begin
            _EVAL_286 <= _EVAL_174;
          end else begin
            _EVAL_286 <= 4'h0;
          end
        end else begin
          _EVAL_286 <= _EVAL_24;
        end
      end
    end
    if (_EVAL_192) begin
      _EVAL_287 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e37f725)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9044f576)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81a5269f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c844bcdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b2e7e28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d05d8812)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf2fbf05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80ae187e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11ef4d21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53cb8465)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1eb8d67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a74bb991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b92cc26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19cf74e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1da22fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84a81312)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9aab613)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a36adb5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3615785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(532cdd7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd2f0060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfdbd1b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d02a754e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6224381)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d557f10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5164bd99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dc86dbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2725ecc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54146dc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e7b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d17d59f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bda73412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f7a9669)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bb5e64d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e8927dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(850d3984)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e92a7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0576dd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33b0eb13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c108b7e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fedd04ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(388ada6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3faedc1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c460fcb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83279c8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a49e6fd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9db6495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(439d4e91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dbc2447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a79f75a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0d32d33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98cce06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d31027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df6c0ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19cad84b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1777fc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf92a907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(746cb02d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cfaffff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7dbf7f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ea2bb7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23099bc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2532c1fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678c13da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1788a378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceb0c77b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4793818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dcca396)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c10a690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b42af990)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1a31e0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79c52aa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
