//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_92(
  output        _EVAL,
  input         _EVAL_0,
  output [3:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  output [3:0]  _EVAL_4,
  output        _EVAL_5,
  output [3:0]  _EVAL_6,
  output [63:0] _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  output [3:0]  _EVAL_12,
  output [31:0] _EVAL_13,
  input         _EVAL_14,
  output [2:0]  _EVAL_15,
  output [7:0]  _EVAL_16,
  input         _EVAL_17,
  output [4:0]  _EVAL_18,
  input         _EVAL_19,
  output [3:0]  _EVAL_20,
  output        _EVAL_21,
  input  [3:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  input  [1:0]  _EVAL_24,
  input  [3:0]  _EVAL_25,
  output        _EVAL_26,
  input  [3:0]  _EVAL_27,
  output [31:0] _EVAL_28,
  output        _EVAL_29,
  input  [63:0] _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input  [2:0]  _EVAL_33,
  input  [1:0]  _EVAL_34,
  output [2:0]  _EVAL_35,
  input  [7:0]  _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  input  [1:0]  _EVAL_39,
  output        _EVAL_40,
  output        _EVAL_41,
  output [3:0]  _EVAL_42,
  output [1:0]  _EVAL_43,
  input         _EVAL_44,
  output        _EVAL_45,
  input  [3:0]  _EVAL_46,
  input         _EVAL_47,
  output [7:0]  _EVAL_48,
  input         _EVAL_49,
  input  [31:0] _EVAL_50,
  output [1:0]  _EVAL_51,
  input  [7:0]  _EVAL_52,
  input  [3:0]  _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input  [63:0] _EVAL_56,
  output [2:0]  _EVAL_57,
  input  [3:0]  _EVAL_58,
  output [1:0]  _EVAL_59,
  output        _EVAL_60,
  input  [7:0]  _EVAL_61,
  output        _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  output [4:0]  _EVAL_65,
  output        _EVAL_66,
  output [3:0]  _EVAL_67,
  output [2:0]  _EVAL_68,
  output [63:0] _EVAL_69,
  input  [4:0]  _EVAL_70,
  input  [2:0]  _EVAL_71,
  output        _EVAL_72,
  input  [2:0]  _EVAL_73,
  input  [4:0]  _EVAL_74,
  output [1:0]  _EVAL_75,
  output [3:0]  _EVAL_76,
  input  [3:0]  _EVAL_77,
  input  [31:0] _EVAL_78,
  input         _EVAL_79,
  output [7:0]  _EVAL_80
);
  wire [4:0] Queue_2__EVAL;
  wire  Queue_2__EVAL_0;
  wire  Queue_2__EVAL_1;
  wire  Queue_2__EVAL_2;
  wire  Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire  Queue_2__EVAL_5;
  wire [4:0] Queue_2__EVAL_6;
  wire [4:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire [4:0] Queue_1__EVAL_6;
  wire [4:0] Queue_3__EVAL;
  wire  Queue_3__EVAL_0;
  wire  Queue_3__EVAL_1;
  wire  Queue_3__EVAL_2;
  wire  Queue_3__EVAL_3;
  wire  Queue_3__EVAL_4;
  wire  Queue_3__EVAL_5;
  wire [4:0] Queue_3__EVAL_6;
  wire [4:0] Queue__EVAL;
  wire  Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire [4:0] Queue__EVAL_6;
  wire  _EVAL_159;
  wire [15:0] _EVAL_185;
  wire  _EVAL_200;
  wire [4:0] _EVAL_195;
  wire [4:0] _EVAL_89;
  wire [4:0] _EVAL_106;
  wire [4:0] _EVAL_191;
  wire [4:0] _EVAL_151;
  wire [4:0] _EVAL_85;
  wire [4:0] _EVAL_103;
  wire [4:0] _EVAL_186;
  wire [4:0] _EVAL_161;
  wire [4:0] _EVAL_118;
  wire [4:0] _EVAL_91;
  wire [15:0] _EVAL_92;
  wire  _EVAL_127;
  wire  _EVAL_177;
  wire  _EVAL_187;
  wire  _EVAL_121;
  wire  _EVAL_140;
  wire  _EVAL_108;
  wire  _EVAL_107;
  wire  _EVAL_173;
  wire  _EVAL_171;
  wire  _EVAL_148;
  wire  _EVAL_88;
  wire [4:0] _EVAL_167;
  wire [4:0] _EVAL_204;
  wire [4:0] _EVAL_137;
  wire [4:0] _EVAL_158;
  wire [4:0] _EVAL_194;
  wire [4:0] _EVAL_144;
  wire [4:0] _EVAL_122;
  wire [4:0] _EVAL_124;
  wire [4:0] _EVAL_112;
  wire [4:0] _EVAL_199;
  wire [4:0] _EVAL_170;
  wire [4:0] _EVAL_160;
  wire [4:0] _EVAL_206;
  wire [4:0] _EVAL_193;
  wire [4:0] _EVAL_97;
  wire  _EVAL_132;
  wire  _EVAL_142;
  wire  _EVAL_138;
  wire  _EVAL_94;
  wire  _EVAL_135;
  wire  _EVAL_147;
  wire  _EVAL_156;
  wire  _EVAL_174;
  wire  _EVAL_169;
  wire  _EVAL_166;
  wire [4:0] _EVAL_152;
  wire  _EVAL_192;
  wire  _EVAL_115;
  wire  _EVAL_202;
  wire  _EVAL_81;
  wire  _EVAL_84;
  wire  _EVAL_164;
  wire [15:0] _EVAL_150;
  wire  _EVAL_126;
  wire  _EVAL_180;
  wire  _EVAL_198;
  wire  _EVAL_183;
  wire  _EVAL_130;
  wire [15:0] _EVAL_176;
  wire  _EVAL_120;
  wire  _EVAL_172;
  wire  _EVAL_146;
  wire  _EVAL_197;
  wire  _EVAL_104;
  wire  _EVAL_203;
  wire  _EVAL_157;
  wire  _EVAL_111;
  wire  _EVAL_128;
  wire  _EVAL_143;
  wire  _EVAL_101;
  wire  _EVAL_82;
  wire [4:0] _EVAL_196;
  wire [4:0] _EVAL_181;
  wire [4:0] _EVAL_99;
  wire [4:0] _EVAL_113;
  wire [4:0] _EVAL_123;
  wire  _EVAL_155;
  wire  _EVAL_139;
  SiFive__EVAL_91 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6)
  );
  SiFive__EVAL_91 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6)
  );
  SiFive__EVAL_91 Queue_3 (
    ._EVAL(Queue_3__EVAL),
    ._EVAL_0(Queue_3__EVAL_0),
    ._EVAL_1(Queue_3__EVAL_1),
    ._EVAL_2(Queue_3__EVAL_2),
    ._EVAL_3(Queue_3__EVAL_3),
    ._EVAL_4(Queue_3__EVAL_4),
    ._EVAL_5(Queue_3__EVAL_5),
    ._EVAL_6(Queue_3__EVAL_6)
  );
  SiFive__EVAL_91 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6)
  );
  assign _EVAL_159 = _EVAL_44 & _EVAL_19;
  assign _EVAL_185 = 16'h1 << _EVAL_53;
  assign _EVAL_200 = _EVAL_185[1];
  assign _EVAL_195 = Queue_3__EVAL;
  assign _EVAL_89 = Queue_2__EVAL;
  assign _EVAL_106 = 4'h1 == _EVAL_25 ? _EVAL_195 : _EVAL_89;
  assign _EVAL_191 = 4'h2 == _EVAL_25 ? 5'h0 : _EVAL_106;
  assign _EVAL_151 = 4'h3 == _EVAL_25 ? 5'h0 : _EVAL_191;
  assign _EVAL_85 = 4'h4 == _EVAL_25 ? 5'h0 : _EVAL_151;
  assign _EVAL_103 = 4'h5 == _EVAL_25 ? 5'h0 : _EVAL_85;
  assign _EVAL_186 = 4'h6 == _EVAL_25 ? 5'h0 : _EVAL_103;
  assign _EVAL_161 = 4'h7 == _EVAL_25 ? 5'h0 : _EVAL_186;
  assign _EVAL_118 = 4'h8 == _EVAL_25 ? 5'h0 : _EVAL_161;
  assign _EVAL_91 = 4'h9 == _EVAL_25 ? 5'h0 : _EVAL_118;
  assign _EVAL_92 = 16'h1 << _EVAL_25;
  assign _EVAL_127 = _EVAL_92[1];
  assign _EVAL_177 = Queue_3__EVAL_2;
  assign _EVAL_187 = Queue_2__EVAL_2;
  assign _EVAL_121 = 4'h1 == _EVAL_77 ? _EVAL_177 : _EVAL_187;
  assign _EVAL_140 = 4'h2 == _EVAL_77 ? 1'h0 : _EVAL_121;
  assign _EVAL_108 = 4'h3 == _EVAL_77 ? 1'h0 : _EVAL_140;
  assign _EVAL_107 = 4'h4 == _EVAL_77 ? 1'h0 : _EVAL_108;
  assign _EVAL_173 = 4'h5 == _EVAL_77 ? 1'h0 : _EVAL_107;
  assign _EVAL_171 = 4'h6 == _EVAL_77 ? 1'h0 : _EVAL_173;
  assign _EVAL_148 = 4'h7 == _EVAL_77 ? 1'h0 : _EVAL_171;
  assign _EVAL_88 = 4'h8 == _EVAL_77 ? 1'h0 : _EVAL_148;
  assign _EVAL_167 = Queue_1__EVAL;
  assign _EVAL_204 = Queue__EVAL;
  assign _EVAL_137 = 4'h1 == _EVAL_53 ? _EVAL_167 : _EVAL_204;
  assign _EVAL_158 = 4'h2 == _EVAL_53 ? 5'h0 : _EVAL_137;
  assign _EVAL_194 = 4'h3 == _EVAL_53 ? 5'h0 : _EVAL_158;
  assign _EVAL_144 = 4'h4 == _EVAL_53 ? 5'h0 : _EVAL_194;
  assign _EVAL_122 = 4'h5 == _EVAL_53 ? 5'h0 : _EVAL_144;
  assign _EVAL_124 = 4'h6 == _EVAL_53 ? 5'h0 : _EVAL_122;
  assign _EVAL_112 = 4'h7 == _EVAL_53 ? 5'h0 : _EVAL_124;
  assign _EVAL_199 = 4'h8 == _EVAL_53 ? 5'h0 : _EVAL_112;
  assign _EVAL_170 = 4'h9 == _EVAL_53 ? 5'h0 : _EVAL_199;
  assign _EVAL_160 = 4'ha == _EVAL_53 ? 5'h0 : _EVAL_170;
  assign _EVAL_206 = 4'hb == _EVAL_53 ? 5'h0 : _EVAL_160;
  assign _EVAL_193 = 4'hc == _EVAL_53 ? 5'h0 : _EVAL_206;
  assign _EVAL_97 = 4'hd == _EVAL_53 ? 5'h0 : _EVAL_193;
  assign _EVAL_132 = Queue_1__EVAL_2;
  assign _EVAL_142 = Queue__EVAL_2;
  assign _EVAL_138 = 4'h1 == _EVAL_58 ? _EVAL_132 : _EVAL_142;
  assign _EVAL_94 = 4'h2 == _EVAL_58 ? 1'h0 : _EVAL_138;
  assign _EVAL_135 = 4'h3 == _EVAL_58 ? 1'h0 : _EVAL_94;
  assign _EVAL_147 = 4'h4 == _EVAL_58 ? 1'h0 : _EVAL_135;
  assign _EVAL_156 = 4'h5 == _EVAL_58 ? 1'h0 : _EVAL_147;
  assign _EVAL_174 = 4'h6 == _EVAL_58 ? 1'h0 : _EVAL_156;
  assign _EVAL_169 = 4'h7 == _EVAL_58 ? 1'h0 : _EVAL_174;
  assign _EVAL_166 = 4'h8 == _EVAL_58 ? 1'h0 : _EVAL_169;
  assign _EVAL_152 = 4'he == _EVAL_53 ? 5'h0 : _EVAL_97;
  assign _EVAL_192 = _EVAL_32 & _EVAL_17;
  assign _EVAL_115 = _EVAL_185[0];
  assign _EVAL_202 = _EVAL_192 & _EVAL_115;
  assign _EVAL_81 = 4'h9 == _EVAL_58 ? 1'h0 : _EVAL_166;
  assign _EVAL_84 = 4'ha == _EVAL_58 ? 1'h0 : _EVAL_81;
  assign _EVAL_164 = 4'hb == _EVAL_58 ? 1'h0 : _EVAL_84;
  assign _EVAL_150 = 16'h1 << _EVAL_77;
  assign _EVAL_126 = _EVAL_150[1];
  assign _EVAL_180 = 4'hc == _EVAL_58 ? 1'h0 : _EVAL_164;
  assign _EVAL_198 = 4'hd == _EVAL_58 ? 1'h0 : _EVAL_180;
  assign _EVAL_183 = 4'he == _EVAL_58 ? 1'h0 : _EVAL_198;
  assign _EVAL_130 = 4'hf == _EVAL_58 ? 1'h0 : _EVAL_183;
  assign _EVAL_176 = 16'h1 << _EVAL_58;
  assign _EVAL_120 = _EVAL_176[1];
  assign _EVAL_172 = 4'h9 == _EVAL_77 ? 1'h0 : _EVAL_88;
  assign _EVAL_146 = 4'ha == _EVAL_77 ? 1'h0 : _EVAL_172;
  assign _EVAL_197 = _EVAL_8 & _EVAL_31;
  assign _EVAL_104 = 4'hb == _EVAL_77 ? 1'h0 : _EVAL_146;
  assign _EVAL_203 = 4'hc == _EVAL_77 ? 1'h0 : _EVAL_104;
  assign _EVAL_157 = 4'hd == _EVAL_77 ? 1'h0 : _EVAL_203;
  assign _EVAL_111 = 4'he == _EVAL_77 ? 1'h0 : _EVAL_157;
  assign _EVAL_128 = 4'hf == _EVAL_77 ? 1'h0 : _EVAL_111;
  assign _EVAL_143 = _EVAL_14 & _EVAL_10;
  assign _EVAL_101 = _EVAL_92[0];
  assign _EVAL_82 = _EVAL_176[0];
  assign _EVAL_196 = 4'ha == _EVAL_25 ? 5'h0 : _EVAL_91;
  assign _EVAL_181 = 4'hb == _EVAL_25 ? 5'h0 : _EVAL_196;
  assign _EVAL_99 = 4'hc == _EVAL_25 ? 5'h0 : _EVAL_181;
  assign _EVAL_113 = 4'hd == _EVAL_25 ? 5'h0 : _EVAL_99;
  assign _EVAL_123 = 4'he == _EVAL_25 ? 5'h0 : _EVAL_113;
  assign _EVAL_155 = _EVAL_192 & _EVAL_200;
  assign _EVAL_139 = _EVAL_150[0];
  assign _EVAL_80 = _EVAL_52;
  assign _EVAL_69 = _EVAL_30;
  assign Queue_3__EVAL_6 = _EVAL_74;
  assign _EVAL_43 = _EVAL_39;
  assign _EVAL_48 = _EVAL_36;
  assign _EVAL_67 = _EVAL_27;
  assign Queue__EVAL_5 = _EVAL_202 & _EVAL_64;
  assign _EVAL_20 = _EVAL_58;
  assign _EVAL_60 = _EVAL_47;
  assign Queue_1__EVAL_4 = _EVAL_54;
  assign _EVAL_21 = _EVAL_8 & _EVAL_130;
  assign Queue_1__EVAL_6 = _EVAL_70;
  assign Queue__EVAL_6 = _EVAL_70;
  assign Queue_2__EVAL_1 = _EVAL_159 & _EVAL_139;
  assign Queue_2__EVAL_6 = _EVAL_74;
  assign _EVAL_29 = _EVAL_10;
  assign _EVAL_59 = _EVAL_34;
  assign Queue_2__EVAL_0 = _EVAL_79;
  assign Queue_2__EVAL_5 = _EVAL_143 & _EVAL_101;
  assign _EVAL_1 = _EVAL_77;
  assign _EVAL_9 = _EVAL_14;
  assign _EVAL_72 = _EVAL_17;
  assign _EVAL_66 = _EVAL_55;
  assign Queue_3__EVAL_1 = _EVAL_159 & _EVAL_126;
  assign _EVAL_57 = _EVAL_73;
  assign _EVAL_6 = _EVAL_25;
  assign _EVAL_15 = _EVAL_33;
  assign _EVAL_26 = _EVAL_31 & _EVAL_130;
  assign _EVAL_40 = _EVAL_0;
  assign _EVAL = _EVAL_32;
  assign _EVAL_62 = _EVAL_19 & _EVAL_128;
  assign _EVAL_35 = _EVAL_23;
  assign _EVAL_18 = 4'hf == _EVAL_53 ? 5'h0 : _EVAL_152;
  assign _EVAL_41 = _EVAL_3;
  assign _EVAL_5 = _EVAL_64;
  assign _EVAL_42 = _EVAL_11;
  assign _EVAL_45 = _EVAL_49;
  assign Queue__EVAL_1 = _EVAL_197 & _EVAL_82;
  assign _EVAL_7 = _EVAL_56;
  assign _EVAL_12 = _EVAL_22;
  assign _EVAL_13 = _EVAL_50;
  assign _EVAL_28 = _EVAL_78;
  assign _EVAL_16 = _EVAL_61;
  assign _EVAL_75 = _EVAL_24;
  assign _EVAL_4 = _EVAL_53;
  assign _EVAL_76 = _EVAL_46;
  assign _EVAL_38 = _EVAL_44 & _EVAL_128;
  assign Queue_1__EVAL_1 = _EVAL_197 & _EVAL_120;
  assign Queue_3__EVAL_0 = _EVAL_79;
  assign Queue_2__EVAL_4 = _EVAL_54;
  assign Queue__EVAL_4 = _EVAL_54;
  assign Queue_3__EVAL_4 = _EVAL_54;
  assign _EVAL_68 = _EVAL_71;
  assign Queue__EVAL_0 = _EVAL_79;
  assign _EVAL_65 = 4'hf == _EVAL_25 ? 5'h0 : _EVAL_123;
  assign Queue_1__EVAL_5 = _EVAL_155 & _EVAL_64;
  assign _EVAL_37 = _EVAL_63;
  assign Queue_3__EVAL_5 = _EVAL_143 & _EVAL_127;
  assign _EVAL_51 = _EVAL_2;
  assign Queue_1__EVAL_0 = _EVAL_79;
endmodule
