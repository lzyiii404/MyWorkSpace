//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_103(
  output [7:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  output [31:0] _EVAL_4,
  output [63:0] _EVAL_5,
  output [2:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input  [63:0] _EVAL_10,
  input  [7:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  output        _EVAL_15,
  output [63:0] _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  input  [63:0] _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input  [2:0]  _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  output [2:0]  _EVAL_32,
  input         _EVAL_33,
  output        _EVAL_34,
  output [2:0]  _EVAL_35,
  output        _EVAL_36
);
  assign _EVAL_8 = _EVAL_28;
  assign _EVAL_34 = _EVAL_29;
  assign _EVAL_35 = _EVAL_22;
  assign _EVAL_26 = _EVAL_33;
  assign _EVAL_36 = _EVAL_9;
  assign _EVAL_15 = _EVAL_31;
  assign _EVAL_20 = _EVAL_27;
  assign _EVAL_5 = _EVAL_10;
  assign _EVAL_6 = _EVAL_7;
  assign _EVAL_18 = _EVAL_14;
  assign _EVAL_16 = _EVAL_19;
  assign _EVAL_1 = _EVAL_3;
  assign _EVAL = _EVAL_11;
  assign _EVAL_4 = _EVAL_2;
  assign _EVAL_21 = _EVAL_0;
  assign _EVAL_23 = _EVAL_24;
  assign _EVAL_32 = _EVAL_13;
  assign _EVAL_30 = _EVAL_12;
endmodule
