//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_109(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [63:0] _EVAL_3,
  output [2:0]  _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  output [2:0]  _EVAL_8,
  input         _EVAL_9,
  output [2:0]  _EVAL_10,
  output [63:0] _EVAL_11,
  input  [7:0]  _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  output [7:0]  _EVAL_16,
  output        _EVAL_17,
  input  [63:0] _EVAL_18,
  output [2:0]  _EVAL_19,
  input         _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [63:0] _EVAL_22,
  input  [2:0]  _EVAL_23,
  input  [2:0]  _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [31:0] _EVAL_26,
  input  [2:0]  _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36
);
  wire  binder__EVAL;
  wire [2:0] binder__EVAL_0;
  wire [63:0] binder__EVAL_1;
  wire [2:0] binder__EVAL_2;
  wire  binder__EVAL_3;
  wire  binder__EVAL_4;
  wire  binder__EVAL_5;
  wire [31:0] binder__EVAL_6;
  wire [2:0] binder__EVAL_7;
  wire [31:0] binder__EVAL_8;
  wire  binder__EVAL_9;
  wire [2:0] binder__EVAL_10;
  wire [2:0] binder__EVAL_11;
  wire [2:0] binder__EVAL_12;
  wire  binder__EVAL_13;
  wire  binder__EVAL_14;
  wire  binder__EVAL_15;
  wire [2:0] binder__EVAL_16;
  wire [7:0] binder__EVAL_17;
  wire [63:0] binder__EVAL_18;
  wire [2:0] binder__EVAL_19;
  wire  binder__EVAL_20;
  wire  binder__EVAL_21;
  wire  binder__EVAL_22;
  wire  binder__EVAL_23;
  wire [2:0] binder__EVAL_24;
  wire  binder__EVAL_25;
  wire  binder__EVAL_26;
  wire  binder__EVAL_27;
  wire [2:0] binder__EVAL_28;
  wire  binder__EVAL_29;
  wire [63:0] binder__EVAL_30;
  wire [63:0] binder__EVAL_31;
  wire  binder__EVAL_32;
  wire  binder__EVAL_33;
  wire  binder__EVAL_34;
  wire [7:0] binder__EVAL_35;
  wire  binder__EVAL_36;
  SiFive__EVAL_108 binder (
    ._EVAL(binder__EVAL),
    ._EVAL_0(binder__EVAL_0),
    ._EVAL_1(binder__EVAL_1),
    ._EVAL_2(binder__EVAL_2),
    ._EVAL_3(binder__EVAL_3),
    ._EVAL_4(binder__EVAL_4),
    ._EVAL_5(binder__EVAL_5),
    ._EVAL_6(binder__EVAL_6),
    ._EVAL_7(binder__EVAL_7),
    ._EVAL_8(binder__EVAL_8),
    ._EVAL_9(binder__EVAL_9),
    ._EVAL_10(binder__EVAL_10),
    ._EVAL_11(binder__EVAL_11),
    ._EVAL_12(binder__EVAL_12),
    ._EVAL_13(binder__EVAL_13),
    ._EVAL_14(binder__EVAL_14),
    ._EVAL_15(binder__EVAL_15),
    ._EVAL_16(binder__EVAL_16),
    ._EVAL_17(binder__EVAL_17),
    ._EVAL_18(binder__EVAL_18),
    ._EVAL_19(binder__EVAL_19),
    ._EVAL_20(binder__EVAL_20),
    ._EVAL_21(binder__EVAL_21),
    ._EVAL_22(binder__EVAL_22),
    ._EVAL_23(binder__EVAL_23),
    ._EVAL_24(binder__EVAL_24),
    ._EVAL_25(binder__EVAL_25),
    ._EVAL_26(binder__EVAL_26),
    ._EVAL_27(binder__EVAL_27),
    ._EVAL_28(binder__EVAL_28),
    ._EVAL_29(binder__EVAL_29),
    ._EVAL_30(binder__EVAL_30),
    ._EVAL_31(binder__EVAL_31),
    ._EVAL_32(binder__EVAL_32),
    ._EVAL_33(binder__EVAL_33),
    ._EVAL_34(binder__EVAL_34),
    ._EVAL_35(binder__EVAL_35),
    ._EVAL_36(binder__EVAL_36)
  );
  assign binder__EVAL_13 = _EVAL_20;
  assign _EVAL_26 = binder__EVAL_6;
  assign binder__EVAL_8 = _EVAL_2;
  assign binder__EVAL_31 = _EVAL_3;
  assign binder__EVAL_3 = _EVAL_29;
  assign binder__EVAL_1 = _EVAL_18;
  assign _EVAL_10 = binder__EVAL_19;
  assign binder__EVAL_22 = _EVAL_15;
  assign _EVAL_17 = binder__EVAL_27;
  assign _EVAL_14 = binder__EVAL_15;
  assign _EVAL_22 = binder__EVAL_30;
  assign binder__EVAL_35 = _EVAL_12;
  assign binder__EVAL_36 = _EVAL_5;
  assign _EVAL_8 = binder__EVAL_12;
  assign binder__EVAL_11 = _EVAL_25;
  assign _EVAL_30 = binder__EVAL_5;
  assign _EVAL_31 = binder__EVAL_9;
  assign binder__EVAL_16 = _EVAL_24;
  assign binder__EVAL_21 = _EVAL_28;
  assign binder__EVAL_24 = _EVAL_23;
  assign _EVAL_19 = binder__EVAL_10;
  assign binder__EVAL_20 = _EVAL_9;
  assign _EVAL_4 = binder__EVAL_28;
  assign _EVAL_6 = binder__EVAL_14;
  assign binder__EVAL_4 = _EVAL_35;
  assign binder__EVAL_34 = _EVAL_32;
  assign _EVAL_7 = binder__EVAL_29;
  assign _EVAL_11 = binder__EVAL_18;
  assign binder__EVAL_0 = _EVAL_27;
  assign _EVAL = binder__EVAL_7;
  assign binder__EVAL_2 = _EVAL_21;
  assign _EVAL_33 = binder__EVAL_32;
  assign _EVAL_13 = binder__EVAL_23;
  assign binder__EVAL_25 = _EVAL_0;
  assign binder__EVAL_33 = _EVAL_1;
  assign binder__EVAL = _EVAL_36;
  assign _EVAL_34 = binder__EVAL_26;
  assign _EVAL_16 = binder__EVAL_17;
endmodule
