//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_54(
  input         _EVAL,
  output [1:0]  _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output [31:0] _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  output [31:0] _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [31:0] _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output [3:0]  _EVAL_18,
  output [3:0]  _EVAL_19,
  output [2:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  input  [3:0]  _EVAL_22,
  output [31:0] _EVAL_23,
  output [3:0]  _EVAL_24,
  input         _EVAL_25,
  input  [1:0]  _EVAL_26,
  input         _EVAL_27,
  output [2:0]  _EVAL_28,
  input         _EVAL_29,
  input  [31:0] _EVAL_30,
  input         _EVAL_31,
  output        _EVAL_32
);
  assign _EVAL_23 = _EVAL_30;
  assign _EVAL_3 = _EVAL_10;
  assign _EVAL_18 = _EVAL_22;
  assign _EVAL_12 = _EVAL_27;
  assign _EVAL_32 = _EVAL_1;
  assign _EVAL_19 = _EVAL_7;
  assign _EVAL_28 = _EVAL_21;
  assign _EVAL_17 = _EVAL_4;
  assign _EVAL_11 = _EVAL;
  assign _EVAL_16 = _EVAL_14;
  assign _EVAL_20 = _EVAL_9;
  assign _EVAL_5 = _EVAL_25;
  assign _EVAL_24 = _EVAL_8;
  assign _EVAL_2 = _EVAL_31;
  assign _EVAL_6 = _EVAL_13;
  assign _EVAL_0 = _EVAL_26;
endmodule
