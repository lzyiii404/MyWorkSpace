//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_108(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [63:0] _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  output [31:0] _EVAL_6,
  output [2:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  output        _EVAL_9,
  output [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  input  [2:0]  _EVAL_16,
  output [7:0]  _EVAL_17,
  output [63:0] _EVAL_18,
  output [2:0]  _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [2:0]  _EVAL_24,
  input         _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  output [2:0]  _EVAL_28,
  output        _EVAL_29,
  output [63:0] _EVAL_30,
  input  [63:0] _EVAL_31,
  output        _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input  [7:0]  _EVAL_35,
  input         _EVAL_36
);
  assign _EVAL_9 = _EVAL;
  assign _EVAL_12 = _EVAL_24;
  assign _EVAL_10 = _EVAL_0;
  assign _EVAL_7 = _EVAL_16;
  assign _EVAL_32 = _EVAL_33;
  assign _EVAL_18 = _EVAL_1;
  assign _EVAL_5 = _EVAL_22;
  assign _EVAL_6 = _EVAL_8;
  assign _EVAL_26 = _EVAL_13;
  assign _EVAL_28 = _EVAL_11;
  assign _EVAL_19 = _EVAL_2;
  assign _EVAL_29 = _EVAL_21;
  assign _EVAL_23 = _EVAL_25;
  assign _EVAL_15 = _EVAL_4;
  assign _EVAL_14 = _EVAL_3;
  assign _EVAL_30 = _EVAL_31;
  assign _EVAL_27 = _EVAL_20;
  assign _EVAL_17 = _EVAL_35;
endmodule
