//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_173(
  output [31:0] _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  output [3:0]  _EVAL_2,
  output [29:0] _EVAL_3,
  output        _EVAL_4,
  output [31:0] _EVAL_5,
  output [2:0]  _EVAL_6,
  output        _EVAL_7,
  output [6:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  output [6:0]  _EVAL_17,
  input  [6:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  input  [6:0]  _EVAL_20,
  input  [29:0] _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  output [2:0]  _EVAL_28,
  input  [3:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  output [2:0]  _EVAL_31,
  output        _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input  [2:0]  _EVAL_35,
  input         _EVAL_36
);
  assign _EVAL_5 = _EVAL_0;
  assign _EVAL_12 = _EVAL_1;
  assign _EVAL_26 = _EVAL_9;
  assign _EVAL_6 = _EVAL_10;
  assign _EVAL_15 = _EVAL_13;
  assign _EVAL_23 = _EVAL_11;
  assign _EVAL_32 = _EVAL_14;
  assign _EVAL_28 = _EVAL_25;
  assign _EVAL_2 = _EVAL_29;
  assign _EVAL_30 = _EVAL_19;
  assign _EVAL_22 = _EVAL_36;
  assign _EVAL_4 = _EVAL_33;
  assign _EVAL_3 = _EVAL_21;
  assign _EVAL_7 = _EVAL_34;
  assign _EVAL_31 = _EVAL_35;
  assign _EVAL = _EVAL_27;
  assign _EVAL_17 = _EVAL_20;
  assign _EVAL_8 = _EVAL_18;
endmodule
