//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_104_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [31:0] _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [7:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_20;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_27;
  reg [31:0] _RAND_1;
  reg [31:0] _EVAL_58;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_69;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_78;
  reg [31:0] _RAND_4;
  reg  _EVAL_97;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_102;
  reg [31:0] _RAND_6;
  reg  _EVAL_111;
  reg [31:0] _RAND_7;
  reg  _EVAL_187;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_205;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_206;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_220;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_228;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_265;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_276;
  reg [31:0] _RAND_14;
  wire  _EVAL_277;
  wire  _EVAL_110;
  wire [12:0] _EVAL_267;
  wire [5:0] _EVAL_269;
  wire [5:0] _EVAL_250;
  wire [31:0] _EVAL_81;
  wire [31:0] _EVAL_180;
  wire  _EVAL_50;
  wire  _EVAL_17;
  wire  _EVAL_54;
  wire  _EVAL_151;
  wire  _EVAL_62;
  wire  _EVAL_35;
  wire  _EVAL_30;
  wire  _EVAL_281;
  wire  _EVAL_227;
  wire  _EVAL_189;
  wire  _EVAL_106;
  wire  _EVAL_271;
  wire  _EVAL_28;
  wire  _EVAL_258;
  wire  _EVAL_32;
  wire [1:0] _EVAL_134;
  wire [3:0] _EVAL_18;
  wire [2:0] _EVAL_44;
  wire [2:0] _EVAL_113;
  wire  _EVAL_157;
  wire  _EVAL_268;
  wire  _EVAL_76;
  wire  _EVAL_196;
  wire  _EVAL_248;
  wire  _EVAL_83;
  wire [1:0] _EVAL_177;
  wire  _EVAL_215;
  wire  _EVAL_108;
  wire  _EVAL_262;
  wire  _EVAL_25;
  wire  _EVAL_38;
  wire  _EVAL_148;
  wire  _EVAL_133;
  wire  _EVAL_222;
  wire  _EVAL_200;
  wire  _EVAL_139;
  wire  _EVAL_223;
  wire  _EVAL_183;
  wire  _EVAL_199;
  wire  _EVAL_99;
  wire  _EVAL_253;
  wire  _EVAL_242;
  wire  _EVAL_226;
  wire  _EVAL_64;
  wire  _EVAL_89;
  wire  _EVAL_45;
  wire  _EVAL_260;
  wire  _EVAL_105;
  wire  _EVAL_138;
  wire [1:0] _EVAL_202;
  wire [1:0] _EVAL_79;
  wire [1:0] _EVAL_161;
  wire [1:0] _EVAL_165;
  wire  _EVAL_230;
  wire  _EVAL_147;
  wire  _EVAL_121;
  wire  _EVAL_34;
  wire [2:0] _EVAL_254;
  wire [2:0] _EVAL_184;
  wire  _EVAL_149;
  wire  _EVAL_87;
  wire  _EVAL_143;
  wire  _EVAL_72;
  wire  _EVAL_278;
  wire  _EVAL_53;
  wire  _EVAL_95;
  wire  _EVAL_280;
  wire  _EVAL_19;
  wire  _EVAL_31;
  wire  _EVAL_198;
  wire  _EVAL_116;
  wire  _EVAL_245;
  wire  _EVAL_176;
  wire  _EVAL_178;
  wire  _EVAL_244;
  wire  _EVAL_86;
  wire  _EVAL_137;
  wire  _EVAL_235;
  wire  _EVAL_234;
  wire  _EVAL_114;
  wire  _EVAL_48;
  wire  _EVAL_144;
  wire  _EVAL_197;
  wire  _EVAL_193;
  wire  _EVAL_140;
  wire  _EVAL_167;
  wire  _EVAL_104;
  wire  _EVAL_238;
  wire [7:0] _EVAL_66;
  wire [7:0] _EVAL_154;
  wire [7:0] _EVAL_229;
  wire  _EVAL_77;
  wire  _EVAL_24;
  wire  _EVAL_49;
  wire  _EVAL_141;
  wire [7:0] _EVAL_282;
  wire  _EVAL_52;
  wire  _EVAL_168;
  wire  _EVAL_43;
  wire  _EVAL_60;
  wire  _EVAL_98;
  wire  _EVAL_128;
  wire  _EVAL_170;
  wire  _EVAL_93;
  wire  _EVAL_264;
  wire  _EVAL_158;
  wire  _EVAL_231;
  wire [12:0] _EVAL_283;
  wire [5:0] _EVAL_59;
  wire [5:0] _EVAL_246;
  wire  _EVAL_65;
  wire  _EVAL_272;
  wire  _EVAL_150;
  wire  _EVAL_40;
  wire  _EVAL_124;
  wire  _EVAL_204;
  wire  _EVAL_173;
  wire  _EVAL_263;
  wire  _EVAL_243;
  wire  _EVAL_174;
  wire  _EVAL_29;
  wire  _EVAL_125;
  wire  _EVAL_130;
  wire  _EVAL_224;
  wire  _EVAL_36;
  wire  _EVAL_156;
  wire  _EVAL_192;
  wire [1:0] _EVAL_85;
  wire [1:0] _EVAL_225;
  wire  _EVAL_67;
  wire  _EVAL_46;
  wire  _EVAL_233;
  wire  _EVAL_182;
  wire  _EVAL_70;
  wire  _EVAL_162;
  wire  _EVAL_101;
  wire  _EVAL_214;
  wire  _EVAL_266;
  wire  _EVAL_41;
  wire  _EVAL_96;
  wire  _EVAL_47;
  wire  _EVAL_270;
  wire  _EVAL_88;
  wire  _EVAL_33;
  wire  _EVAL_203;
  wire  _EVAL_237;
  wire  _EVAL_82;
  wire  _EVAL_219;
  wire  _EVAL_142;
  wire  _EVAL_160;
  wire [1:0] _EVAL_186;
  wire [2:0] _EVAL_191;
  wire  _EVAL_118;
  wire  _EVAL_100;
  wire  _EVAL_232;
  wire  _EVAL_208;
  wire [31:0] _EVAL_201;
  wire [32:0] _EVAL_152;
  wire [32:0] _EVAL_22;
  wire [32:0] _EVAL_247;
  wire  _EVAL_236;
  wire [2:0] _EVAL_155;
  wire  _EVAL_123;
  wire  _EVAL_127;
  wire  _EVAL_257;
  wire  _EVAL_195;
  wire  _EVAL_117;
  wire  _EVAL_261;
  wire  _EVAL_119;
  wire  _EVAL_194;
  wire  _EVAL_179;
  wire  _EVAL_255;
  wire  _EVAL_251;
  wire  _EVAL_240;
  wire  _EVAL_56;
  wire  _EVAL_241;
  wire  _EVAL_57;
  wire [2:0] _EVAL_256;
  wire  _EVAL_42;
  wire  _EVAL_213;
  wire  _EVAL_84;
  wire  _EVAL_74;
  wire  _EVAL_91;
  wire  _EVAL_159;
  wire  _EVAL_126;
  wire  _EVAL_92;
  wire [1:0] _EVAL_94;
  wire [1:0] _EVAL_132;
  wire  _EVAL_75;
  wire  _EVAL_274;
  wire  _EVAL_211;
  wire  _EVAL_145;
  wire  _EVAL_61;
  wire  _EVAL_249;
  wire  _EVAL_37;
  wire  _EVAL_207;
  wire  _EVAL_120;
  wire  _EVAL_209;
  wire  _EVAL_175;
  wire  _EVAL_210;
  wire  _EVAL_273;
  wire  _EVAL_63;
  wire  _EVAL_136;
  wire  _EVAL_122;
  wire  _EVAL_171;
  wire  _EVAL_153;
  wire  _EVAL_166;
  wire  _EVAL_90;
  wire  _EVAL_163;
  wire  _EVAL_68;
  wire  _EVAL_80;
  wire  _EVAL_279;
  wire [2:0] _EVAL_275;
  wire  _EVAL_164;
  wire  _EVAL_188;
  wire  _EVAL_216;
  wire [31:0] _EVAL_112;
  wire  _EVAL_39;
  wire  _EVAL_73;
  wire  _EVAL_259;
  wire  _EVAL_218;
  wire  _EVAL_55;
  wire  _EVAL_26;
  wire  _EVAL_221;
  wire  _EVAL_71;
  wire  _EVAL_51;
  wire  _EVAL_107;
  wire  _EVAL_212;
  wire  _EVAL_169;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_277 = _EVAL_12[2];
  assign _EVAL_110 = _EVAL_277 == 1'h0;
  assign _EVAL_267 = 13'h3f << _EVAL_10;
  assign _EVAL_269 = _EVAL_267[5:0];
  assign _EVAL_250 = ~ _EVAL_269;
  assign _EVAL_81 = {{26'd0}, _EVAL_250};
  assign _EVAL_180 = _EVAL_11 & _EVAL_81;
  assign _EVAL_50 = _EVAL_180 == 32'h0;
  assign _EVAL_17 = _EVAL_50 | _EVAL_6;
  assign _EVAL_54 = _EVAL_17 == 1'h0;
  assign _EVAL_151 = _EVAL_12 == 3'h3;
  assign _EVAL_62 = _EVAL_4 & _EVAL_151;
  assign _EVAL_35 = _EVAL_12 == 3'h5;
  assign _EVAL_30 = _EVAL_4 & _EVAL_35;
  assign _EVAL_281 = _EVAL_12 == 3'h2;
  assign _EVAL_227 = _EVAL_5 & _EVAL_15;
  assign _EVAL_189 = _EVAL_228 == 3'h0;
  assign _EVAL_106 = _EVAL_227 & _EVAL_189;
  assign _EVAL_271 = _EVAL_7 == 1'h0;
  assign _EVAL_28 = _EVAL_271 | _EVAL_6;
  assign _EVAL_258 = _EVAL_8 != 3'h0;
  assign _EVAL_32 = _EVAL_258 | _EVAL_6;
  assign _EVAL_134 = _EVAL_10[1:0];
  assign _EVAL_18 = 4'h1 << _EVAL_134;
  assign _EVAL_44 = _EVAL_18[2:0];
  assign _EVAL_113 = _EVAL_44 | 3'h1;
  assign _EVAL_157 = _EVAL_113[1];
  assign _EVAL_268 = _EVAL_11[2];
  assign _EVAL_76 = _EVAL_11[1];
  assign _EVAL_196 = _EVAL_76 == 1'h0;
  assign _EVAL_248 = _EVAL_268 & _EVAL_196;
  assign _EVAL_83 = _EVAL_157 & _EVAL_248;
  assign _EVAL_177 = _EVAL_206 >> _EVAL_16;
  assign _EVAL_215 = _EVAL_113[0];
  assign _EVAL_108 = _EVAL_11[0];
  assign _EVAL_262 = _EVAL_248 & _EVAL_108;
  assign _EVAL_25 = _EVAL_215 & _EVAL_262;
  assign _EVAL_38 = _EVAL_268 & _EVAL_76;
  assign _EVAL_148 = _EVAL_38 & _EVAL_108;
  assign _EVAL_133 = _EVAL_8 == _EVAL_205;
  assign _EVAL_222 = _EVAL_133 | _EVAL_6;
  assign _EVAL_200 = _EVAL_268 == 1'h0;
  assign _EVAL_139 = _EVAL_200 & _EVAL_76;
  assign _EVAL_223 = _EVAL_157 & _EVAL_139;
  assign _EVAL_183 = _EVAL_10 >= 3'h3;
  assign _EVAL_199 = _EVAL_113[2];
  assign _EVAL_99 = _EVAL_199 & _EVAL_200;
  assign _EVAL_253 = _EVAL_183 | _EVAL_99;
  assign _EVAL_242 = _EVAL_253 | _EVAL_223;
  assign _EVAL_226 = _EVAL_108 == 1'h0;
  assign _EVAL_64 = _EVAL_139 & _EVAL_226;
  assign _EVAL_89 = _EVAL_215 & _EVAL_64;
  assign _EVAL_45 = _EVAL_242 | _EVAL_89;
  assign _EVAL_260 = _EVAL_2 & _EVAL_4;
  assign _EVAL_105 = _EVAL_78 == 3'h0;
  assign _EVAL_138 = _EVAL_260 & _EVAL_105;
  assign _EVAL_202 = 2'h1 << _EVAL_16;
  assign _EVAL_79 = _EVAL_138 ? _EVAL_202 : 2'h0;
  assign _EVAL_161 = _EVAL_79 | _EVAL_206;
  assign _EVAL_165 = _EVAL_161 >> _EVAL_3;
  assign _EVAL_230 = _EVAL_165[0];
  assign _EVAL_147 = _EVAL_20 == 3'h0;
  assign _EVAL_121 = _EVAL_147 == 1'h0;
  assign _EVAL_34 = _EVAL_15 & _EVAL_121;
  assign _EVAL_254 = _EVAL_250[5:3];
  assign _EVAL_184 = _EVAL_78 - 3'h1;
  assign _EVAL_149 = _EVAL_9 == 3'h6;
  assign _EVAL_87 = _EVAL_149 == 1'h0;
  assign _EVAL_143 = _EVAL_106 & _EVAL_87;
  assign _EVAL_72 = _EVAL_199 & _EVAL_268;
  assign _EVAL_278 = _EVAL_183 | _EVAL_72;
  assign _EVAL_53 = _EVAL_157 & _EVAL_38;
  assign _EVAL_95 = _EVAL_278 | _EVAL_53;
  assign _EVAL_280 = _EVAL_215 & _EVAL_148;
  assign _EVAL_19 = _EVAL_95 | _EVAL_280;
  assign _EVAL_31 = _EVAL_38 & _EVAL_226;
  assign _EVAL_198 = _EVAL_215 & _EVAL_31;
  assign _EVAL_116 = _EVAL_95 | _EVAL_198;
  assign _EVAL_245 = _EVAL_278 | _EVAL_83;
  assign _EVAL_176 = _EVAL_245 | _EVAL_25;
  assign _EVAL_178 = _EVAL_248 & _EVAL_226;
  assign _EVAL_244 = _EVAL_215 & _EVAL_178;
  assign _EVAL_86 = _EVAL_245 | _EVAL_244;
  assign _EVAL_137 = _EVAL_139 & _EVAL_108;
  assign _EVAL_235 = _EVAL_215 & _EVAL_137;
  assign _EVAL_234 = _EVAL_242 | _EVAL_235;
  assign _EVAL_114 = _EVAL_200 & _EVAL_196;
  assign _EVAL_48 = _EVAL_157 & _EVAL_114;
  assign _EVAL_144 = _EVAL_253 | _EVAL_48;
  assign _EVAL_197 = _EVAL_114 & _EVAL_108;
  assign _EVAL_193 = _EVAL_215 & _EVAL_197;
  assign _EVAL_140 = _EVAL_144 | _EVAL_193;
  assign _EVAL_167 = _EVAL_114 & _EVAL_226;
  assign _EVAL_104 = _EVAL_215 & _EVAL_167;
  assign _EVAL_238 = _EVAL_144 | _EVAL_104;
  assign _EVAL_66 = {_EVAL_19,_EVAL_116,_EVAL_176,_EVAL_86,_EVAL_234,_EVAL_45,_EVAL_140,_EVAL_238};
  assign _EVAL_154 = ~ _EVAL_66;
  assign _EVAL_229 = _EVAL_13 & _EVAL_154;
  assign _EVAL_77 = _EVAL_12 == 3'h4;
  assign _EVAL_24 = _EVAL_229 == 8'h0;
  assign _EVAL_49 = _EVAL == 1'h0;
  assign _EVAL_141 = _EVAL_12 == 3'h7;
  assign _EVAL_282 = ~ _EVAL_13;
  assign _EVAL_52 = _EVAL_282 == 8'h0;
  assign _EVAL_168 = _EVAL_183 | _EVAL_6;
  assign _EVAL_43 = _EVAL_168 == 1'h0;
  assign _EVAL_60 = _EVAL_177[0];
  assign _EVAL_98 = _EVAL_60 == 1'h0;
  assign _EVAL_128 = _EVAL_98 | _EVAL_6;
  assign _EVAL_170 = _EVAL_128 == 1'h0;
  assign _EVAL_93 = _EVAL_9[0];
  assign _EVAL_264 = _EVAL_24 | _EVAL_6;
  assign _EVAL_158 = _EVAL_14 >= 3'h3;
  assign _EVAL_231 = _EVAL_158 | _EVAL_6;
  assign _EVAL_283 = 13'h3f << _EVAL_14;
  assign _EVAL_59 = _EVAL_283[5:0];
  assign _EVAL_246 = ~ _EVAL_59;
  assign _EVAL_65 = _EVAL_6 == 1'h0;
  assign _EVAL_272 = _EVAL_102 == 3'h0;
  assign _EVAL_150 = _EVAL_12 == 3'h1;
  assign _EVAL_40 = _EVAL_4 & _EVAL_150;
  assign _EVAL_124 = _EVAL_10 <= 3'h6;
  assign _EVAL_204 = _EVAL_206 != 2'h0;
  assign _EVAL_173 = _EVAL_204 == 1'h0;
  assign _EVAL_263 = plusarg_reader_out == 32'h0;
  assign _EVAL_243 = _EVAL_173 | _EVAL_263;
  assign _EVAL_174 = _EVAL_27 < plusarg_reader_out;
  assign _EVAL_29 = _EVAL_243 | _EVAL_174;
  assign _EVAL_125 = _EVAL_29 | _EVAL_6;
  assign _EVAL_130 = _EVAL_125 == 1'h0;
  assign _EVAL_224 = _EVAL_13 == _EVAL_66;
  assign _EVAL_36 = _EVAL_9 == 3'h0;
  assign _EVAL_156 = _EVAL_15 & _EVAL_36;
  assign _EVAL_192 = _EVAL_9 == 3'h5;
  assign _EVAL_85 = 2'h1 << _EVAL_3;
  assign _EVAL_225 = _EVAL_143 ? _EVAL_85 : 2'h0;
  assign _EVAL_67 = _EVAL_79 != _EVAL_225;
  assign _EVAL_46 = _EVAL_79 != 2'h0;
  assign _EVAL_233 = _EVAL_46 == 1'h0;
  assign _EVAL_182 = _EVAL_260 | _EVAL_227;
  assign _EVAL_70 = _EVAL_8 <= 3'h4;
  assign _EVAL_162 = _EVAL_70 | _EVAL_6;
  assign _EVAL_101 = _EVAL_162 == 1'h0;
  assign _EVAL_214 = _EVAL_67 | _EVAL_233;
  assign _EVAL_266 = _EVAL_214 | _EVAL_6;
  assign _EVAL_41 = _EVAL_272 == 1'h0;
  assign _EVAL_96 = _EVAL_4 & _EVAL_41;
  assign _EVAL_47 = _EVAL_10 == _EVAL_265;
  assign _EVAL_270 = _EVAL_47 | _EVAL_6;
  assign _EVAL_88 = _EVAL_270 == 1'h0;
  assign _EVAL_33 = _EVAL_9 == 3'h1;
  assign _EVAL_203 = _EVAL_15 & _EVAL_33;
  assign _EVAL_237 = _EVAL_16 == _EVAL_97;
  assign _EVAL_82 = _EVAL_237 | _EVAL_6;
  assign _EVAL_219 = _EVAL_82 == 1'h0;
  assign _EVAL_142 = _EVAL_14 == _EVAL_69;
  assign _EVAL_160 = _EVAL_9 == _EVAL_276;
  assign _EVAL_186 = _EVAL_206 | _EVAL_79;
  assign _EVAL_191 = _EVAL_246[5:3];
  assign _EVAL_118 = _EVAL_4 & _EVAL_141;
  assign _EVAL_100 = _EVAL_8 == 3'h0;
  assign _EVAL_232 = _EVAL_11 == _EVAL_58;
  assign _EVAL_208 = _EVAL_232 | _EVAL_6;
  assign _EVAL_201 = _EVAL_11 ^ 32'h80000000;
  assign _EVAL_152 = {1'b0,$signed(_EVAL_201)};
  assign _EVAL_22 = $signed(_EVAL_152) & $signed(-33'sh20000);
  assign _EVAL_247 = $signed(_EVAL_22);
  assign _EVAL_236 = _EVAL_208 == 1'h0;
  assign _EVAL_155 = _EVAL_228 - 3'h1;
  assign _EVAL_123 = _EVAL_15 & _EVAL_149;
  assign _EVAL_127 = _EVAL_9 == 3'h2;
  assign _EVAL_257 = _EVAL_15 & _EVAL_127;
  assign _EVAL_195 = _EVAL_1 == _EVAL_187;
  assign _EVAL_117 = _EVAL_195 | _EVAL_6;
  assign _EVAL_261 = _EVAL_1 == 1'h0;
  assign _EVAL_119 = _EVAL_261 | _EVAL_7;
  assign _EVAL_194 = _EVAL_3 == _EVAL_111;
  assign _EVAL_179 = _EVAL_194 | _EVAL_6;
  assign _EVAL_255 = _EVAL_179 == 1'h0;
  assign _EVAL_251 = _EVAL_12 == 3'h6;
  assign _EVAL_240 = _EVAL_4 & _EVAL_251;
  assign _EVAL_56 = _EVAL_15 & _EVAL_192;
  assign _EVAL_241 = _EVAL_8 <= 3'h3;
  assign _EVAL_57 = _EVAL_241 | _EVAL_6;
  assign _EVAL_256 = _EVAL_102 - 3'h1;
  assign _EVAL_42 = _EVAL_142 | _EVAL_6;
  assign _EVAL_213 = _EVAL_12 == 3'h0;
  assign _EVAL_84 = _EVAL_261 | _EVAL_6;
  assign _EVAL_74 = _EVAL_84 == 1'h0;
  assign _EVAL_91 = $signed(_EVAL_247) == $signed(33'sh0);
  assign _EVAL_159 = _EVAL_124 & _EVAL_91;
  assign _EVAL_126 = _EVAL_159 | _EVAL_6;
  assign _EVAL_92 = _EVAL_126 == 1'h0;
  assign _EVAL_94 = ~ _EVAL_225;
  assign _EVAL_132 = _EVAL_186 & _EVAL_94;
  assign _EVAL_75 = _EVAL_227 & _EVAL_147;
  assign _EVAL_274 = _EVAL_224 | _EVAL_6;
  assign _EVAL_211 = _EVAL_274 == 1'h0;
  assign _EVAL_145 = _EVAL_9 <= 3'h6;
  assign _EVAL_61 = _EVAL_145 | _EVAL_6;
  assign _EVAL_249 = _EVAL_61 == 1'h0;
  assign _EVAL_37 = _EVAL_119 | _EVAL_6;
  assign _EVAL_207 = _EVAL_12 == _EVAL_220;
  assign _EVAL_120 = _EVAL_260 & _EVAL_272;
  assign _EVAL_209 = _EVAL_222 == 1'h0;
  assign _EVAL_175 = _EVAL_4 & _EVAL_213;
  assign _EVAL_210 = _EVAL_52 | _EVAL_6;
  assign _EVAL_273 = _EVAL_210 == 1'h0;
  assign _EVAL_63 = _EVAL_37 == 1'h0;
  assign _EVAL_136 = _EVAL_9 == 3'h4;
  assign _EVAL_122 = _EVAL_15 & _EVAL_136;
  assign _EVAL_171 = _EVAL_207 | _EVAL_6;
  assign _EVAL_153 = _EVAL_117 == 1'h0;
  assign _EVAL_166 = _EVAL_230 | _EVAL_6;
  assign _EVAL_90 = _EVAL_4 & _EVAL_77;
  assign _EVAL_163 = _EVAL_8 <= 3'h2;
  assign _EVAL_68 = _EVAL_163 | _EVAL_6;
  assign _EVAL_80 = _EVAL_49 | _EVAL_6;
  assign _EVAL_279 = _EVAL_80 == 1'h0;
  assign _EVAL_275 = _EVAL_20 - 3'h1;
  assign _EVAL_164 = _EVAL_160 | _EVAL_6;
  assign _EVAL_188 = _EVAL_57 == 1'h0;
  assign _EVAL_216 = _EVAL_100 | _EVAL_6;
  assign _EVAL_112 = _EVAL_27 + 32'h1;
  assign _EVAL_39 = _EVAL_68 == 1'h0;
  assign _EVAL_73 = _EVAL_166 == 1'h0;
  assign _EVAL_259 = _EVAL_4 & _EVAL_281;
  assign _EVAL_218 = _EVAL_216 == 1'h0;
  assign _EVAL_55 = _EVAL_171 == 1'h0;
  assign _EVAL_26 = _EVAL_231 == 1'h0;
  assign _EVAL_221 = _EVAL_266 == 1'h0;
  assign _EVAL_71 = _EVAL_164 == 1'h0;
  assign _EVAL_51 = _EVAL_32 == 1'h0;
  assign _EVAL_107 = _EVAL_42 == 1'h0;
  assign _EVAL_212 = _EVAL_264 == 1'h0;
  assign _EVAL_169 = _EVAL_28 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_27 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_58 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_69 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_78 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_97 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_102 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_111 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_187 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_205 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_206 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_220 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_228 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_265 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_276 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_6) begin
      _EVAL_20 <= 3'h0;
    end else begin
      if (_EVAL_227) begin
        if (_EVAL_147) begin
          if (_EVAL_93) begin
            _EVAL_20 <= _EVAL_191;
          end else begin
            _EVAL_20 <= 3'h0;
          end
        end else begin
          _EVAL_20 <= _EVAL_275;
        end
      end
    end
    if (_EVAL_6) begin
      _EVAL_27 <= 32'h0;
    end else begin
      if (_EVAL_182) begin
        _EVAL_27 <= 32'h0;
      end else begin
        _EVAL_27 <= _EVAL_112;
      end
    end
    if (_EVAL_120) begin
      _EVAL_58 <= _EVAL_11;
    end
    if (_EVAL_75) begin
      _EVAL_69 <= _EVAL_14;
    end
    if (_EVAL_6) begin
      _EVAL_78 <= 3'h0;
    end else begin
      if (_EVAL_260) begin
        if (_EVAL_105) begin
          if (_EVAL_110) begin
            _EVAL_78 <= _EVAL_254;
          end else begin
            _EVAL_78 <= 3'h0;
          end
        end else begin
          _EVAL_78 <= _EVAL_184;
        end
      end
    end
    if (_EVAL_120) begin
      _EVAL_97 <= _EVAL_16;
    end
    if (_EVAL_6) begin
      _EVAL_102 <= 3'h0;
    end else begin
      if (_EVAL_260) begin
        if (_EVAL_272) begin
          if (_EVAL_110) begin
            _EVAL_102 <= _EVAL_254;
          end else begin
            _EVAL_102 <= 3'h0;
          end
        end else begin
          _EVAL_102 <= _EVAL_256;
        end
      end
    end
    if (_EVAL_75) begin
      _EVAL_111 <= _EVAL_3;
    end
    if (_EVAL_75) begin
      _EVAL_187 <= _EVAL_1;
    end
    if (_EVAL_120) begin
      _EVAL_205 <= _EVAL_8;
    end
    if (_EVAL_6) begin
      _EVAL_206 <= 2'h0;
    end else begin
      _EVAL_206 <= _EVAL_132;
    end
    if (_EVAL_120) begin
      _EVAL_220 <= _EVAL_12;
    end
    if (_EVAL_6) begin
      _EVAL_228 <= 3'h0;
    end else begin
      if (_EVAL_227) begin
        if (_EVAL_189) begin
          if (_EVAL_93) begin
            _EVAL_228 <= _EVAL_191;
          end else begin
            _EVAL_228 <= 3'h0;
          end
        end else begin
          _EVAL_228 <= _EVAL_155;
        end
      end
    end
    if (_EVAL_120) begin
      _EVAL_265 <= _EVAL_10;
    end
    if (_EVAL_75) begin
      _EVAL_276 <= _EVAL_9;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d634fe93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(116da6e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(418b0996)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(231cddd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37e4cdf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31104fd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ab9c392)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(758b9f68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17667086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11203ddc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eb918d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba26f7a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1ed4dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b47d8b16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c518a577)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c06bbaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54242d54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80f56e66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3012273e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85fce7d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48157ae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(934fad6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adc455b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86e2d58d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c5c36d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e44bd62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec88a2f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(552149fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6f69e8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(886973c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a01bd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5bc068b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9854642d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcb92cea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7d34e93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45151c4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c21bc8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e00fe89e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddc25e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8c66200)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c87b737a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9221d02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a73bc4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f100a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b1ed499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91aa36f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a44b1a66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a77ffdc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53ba47d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a919416)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4197c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2464a4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26327e4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c93d73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6493ce7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26efc925)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66f40114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc8f28c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(648002c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b39345cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73f13064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6477b1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2d64e6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd50e2e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(354ef866)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eba505e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
