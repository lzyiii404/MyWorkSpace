//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_303(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  input         _EVAL_1,
  output [32:0] _EVAL_2,
  output [6:0]  _EVAL_3,
  output        _EVAL_4,
  input  [4:0]  _EVAL_5,
  input  [32:0] _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output [31:0] _EVAL_9,
  output [2:0]  _EVAL_10,
  input  [4:0]  _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output [6:0]  _EVAL_17,
  output [4:0]  _EVAL_18,
  input  [32:0] _EVAL_19,
  output        _EVAL_20,
  output [32:0] _EVAL_21,
  output        _EVAL_22,
  output [6:0]  _EVAL_23,
  output        _EVAL_24,
  output [4:0]  _EVAL_25,
  output [4:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [4:0]  _EVAL_28,
  output [4:0]  _EVAL_29,
  output [32:0] _EVAL_30,
  input  [2:0]  _EVAL_31,
  input  [32:0] _EVAL_32,
  input         _EVAL_33,
  output [2:0]  _EVAL_34,
  output [4:0]  _EVAL_35,
  input         _EVAL_36,
  output [4:0]  _EVAL_37,
  input         _EVAL_38,
  output [2:0]  _EVAL_39,
  output        _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  output [4:0]  _EVAL_43,
  output        _EVAL_44,
  output [4:0]  _EVAL_45,
  input         _EVAL_46,
  output [4:0]  _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  input  [6:0]  _EVAL_50,
  output [2:0]  _EVAL_51,
  output        _EVAL_52,
  output        _EVAL_53,
  output [4:0]  _EVAL_54,
  output        _EVAL_55,
  output        _EVAL_56,
  output [4:0]  _EVAL_57,
  input         _EVAL_58,
  output [6:0]  _EVAL_59,
  output [32:0] _EVAL_60
);
  wire  simpleOps__EVAL;
  wire [6:0] simpleOps__EVAL_0;
  wire  simpleOps__EVAL_1;
  wire [31:0] simpleOps__EVAL_2;
  wire [32:0] simpleOps__EVAL_3;
  wire [4:0] simpleOps__EVAL_4;
  wire [31:0] simpleOps__EVAL_5;
  wire  simpleOps__EVAL_6;
  wire [4:0] simpleOps__EVAL_7;
  wire  simpleOps__EVAL_8;
  wire [32:0] simpleOps__EVAL_9;
  wire  simpleOps__EVAL_10;
  wire [32:0] simpleOps__EVAL_11;
  wire [2:0] simpleOps__EVAL_12;
  wire [4:0] divSqrts_0__EVAL;
  wire [2:0] divSqrts_0__EVAL_0;
  wire  divSqrts_0__EVAL_1;
  wire  divSqrts_0__EVAL_2;
  wire  divSqrts_0__EVAL_3;
  wire  divSqrts_0__EVAL_4;
  wire  divSqrts_0__EVAL_5;
  wire  divSqrts_0__EVAL_6;
  wire  divSqrts_0__EVAL_7;
  wire [32:0] divSqrts_0__EVAL_8;
  wire [32:0] divSqrts_0__EVAL_9;
  wire [32:0] divSqrts_0__EVAL_10;
  wire  divSqrts_0__EVAL_11;
  wire [32:0] fmas_0__EVAL;
  wire [4:0] fmas_0__EVAL_0;
  wire [32:0] fmas_0__EVAL_1;
  wire [2:0] fmas_0__EVAL_2;
  wire  fmas_0__EVAL_3;
  wire [32:0] fmas_0__EVAL_4;
  wire  fmas_0__EVAL_5;
  wire  fmas_0__EVAL_6;
  wire  fmas_0__EVAL_7;
  wire [32:0] fmas_0__EVAL_8;
  reg  _EVAL_62;
  reg [31:0] _RAND_0;
  reg  _EVAL_64;
  reg [31:0] _RAND_1;
  reg  _EVAL_67;
  reg [31:0] _RAND_2;
  reg [32:0] _EVAL_75;
  reg [63:0] _RAND_3;
  reg  _EVAL_77;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_80;
  reg [31:0] _RAND_5;
  reg  _EVAL_83;
  reg [31:0] _RAND_6;
  reg [32:0] _EVAL_92;
  reg [63:0] _RAND_7;
  reg [2:0] _EVAL_98;
  reg [31:0] _RAND_8;
  reg [4:0] _EVAL_104;
  reg [31:0] _RAND_9;
  reg [6:0] _EVAL_110;
  reg [31:0] _RAND_10;
  reg  _EVAL_116;
  reg [31:0] _RAND_11;
  reg [6:0] _EVAL_117;
  reg [31:0] _RAND_12;
  reg [32:0] _EVAL_119;
  reg [63:0] _RAND_13;
  reg  _EVAL_125;
  reg [31:0] _RAND_14;
  reg [32:0] _EVAL_127;
  reg [63:0] _RAND_15;
  reg  _EVAL_138;
  reg [31:0] _RAND_16;
  reg  _EVAL_143;
  reg [31:0] _RAND_17;
  reg [32:0] _EVAL_146;
  reg [63:0] _RAND_18;
  reg [4:0] _EVAL_148;
  reg [31:0] _RAND_19;
  reg [4:0] _EVAL_158;
  reg [31:0] _RAND_20;
  reg  _EVAL_160;
  reg [31:0] _RAND_21;
  reg  _EVAL_171;
  reg [31:0] _RAND_22;
  reg [6:0] _EVAL_177;
  reg [31:0] _RAND_23;
  reg  _EVAL_181;
  reg [31:0] _RAND_24;
  reg [6:0] _EVAL_182;
  reg [31:0] _RAND_25;
  reg [4:0] _EVAL_186;
  reg [31:0] _RAND_26;
  reg  _EVAL_188;
  reg [31:0] _RAND_27;
  reg  _EVAL_189;
  reg [31:0] _RAND_28;
  reg  _EVAL_191;
  reg [31:0] _RAND_29;
  reg [32:0] _EVAL_192;
  reg [63:0] _RAND_30;
  reg [4:0] _EVAL_197;
  reg [31:0] _RAND_31;
  reg [4:0] _EVAL_200;
  reg [31:0] _RAND_32;
  reg  _EVAL_216;
  reg [31:0] _RAND_33;
  reg [4:0] _EVAL_219;
  reg [31:0] _RAND_34;
  reg  _EVAL_222;
  reg [31:0] _RAND_35;
  reg  _EVAL_227;
  reg [31:0] _RAND_36;
  reg  _EVAL_232;
  reg [31:0] _RAND_37;
  reg [4:0] _EVAL_233;
  reg [31:0] _RAND_38;
  reg [4:0] _EVAL_234;
  reg [31:0] _RAND_39;
  reg [31:0] _EVAL_246;
  reg [31:0] _RAND_40;
  reg [4:0] _EVAL_249;
  reg [31:0] _RAND_41;
  reg  _EVAL_256;
  reg [31:0] _RAND_42;
  reg  _EVAL_257;
  reg [31:0] _RAND_43;
  reg [4:0] _EVAL_276;
  reg [31:0] _RAND_44;
  wire [4:0] _EVAL_142;
  wire  _EVAL_273;
  wire  _EVAL_243;
  wire  _EVAL_68;
  wire  _EVAL_74;
  wire  _EVAL_145;
  wire  _EVAL_174;
  wire  _EVAL_95;
  wire  _EVAL_82;
  wire  _EVAL_121;
  wire  _EVAL_123;
  wire  _EVAL_91;
  wire  _EVAL_259;
  wire  _EVAL_226;
  wire  _EVAL_268;
  wire  _EVAL_179;
  wire [2:0] _EVAL_248;
  wire  _EVAL_195;
  wire [4:0] _EVAL_81;
  wire  _EVAL_131;
  wire  _EVAL_202;
  wire  _EVAL_220;
  wire  _EVAL_113;
  wire  _EVAL_206;
  wire  _EVAL_203;
  wire  _EVAL_228;
  wire  _EVAL_173;
  wire  _EVAL_212;
  wire  _EVAL_78;
  wire [4:0] _EVAL_163;
  wire [4:0] _EVAL_152;
  wire  _EVAL_198;
  wire  _EVAL_86;
  wire  _EVAL_76;
  wire  _EVAL_251;
  wire  _EVAL_115;
  wire  _EVAL_155;
  wire  _EVAL_275;
  wire [4:0] _EVAL_190;
  wire  _EVAL_109;
  wire  _EVAL_258;
  wire  _EVAL_242;
  wire  _EVAL_204;
  wire  _EVAL_264;
  wire  _EVAL_245;
  wire [4:0] _EVAL_150;
  wire  _EVAL_261;
  wire  _EVAL_221;
  wire  _EVAL_209;
  wire  _EVAL_254;
  wire  _EVAL_112;
  wire [32:0] _EVAL_105;
  wire  _EVAL_154;
  wire  _EVAL_136;
  wire [4:0] _EVAL_96;
  wire  _EVAL_260;
  wire  _EVAL_229;
  wire  _EVAL_201;
  wire  _EVAL_61;
  wire  _EVAL_237;
  wire  _EVAL_99;
  wire  _EVAL_278;
  wire  _EVAL_277;
  wire [4:0] _EVAL_135;
  wire  _EVAL_124;
  wire [4:0] _EVAL_240;
  wire  _EVAL_252;
  wire  _EVAL_175;
  wire  _EVAL_71;
  wire  _EVAL_134;
  wire  _EVAL_137;
  wire  _EVAL_270;
  wire  _EVAL_120;
  wire  _EVAL_97;
  wire  _EVAL_118;
  wire  _EVAL_262;
  wire  _EVAL_250;
  wire  _EVAL_79;
  wire  _EVAL_139;
  wire  _EVAL_132;
  wire [32:0] _EVAL_239;
  wire  _EVAL_73;
  wire  _EVAL_101;
  wire  _EVAL_69;
  wire  _EVAL_238;
  wire  _EVAL_230;
  wire  _EVAL_211;
  wire [32:0] _EVAL_265;
  wire [32:0] _EVAL_207;
  wire  _EVAL_122;
  wire  _EVAL_141;
  wire  _EVAL_111;
  wire [4:0] _EVAL_144;
  wire  _EVAL_130;
  wire  _EVAL_88;
  wire  _EVAL_126;
  wire  _EVAL_225;
  wire  _EVAL_159;
  wire  _EVAL_85;
  wire  _EVAL_102;
  wire  _EVAL_87;
  wire  _EVAL_172;
  wire  _EVAL_185;
  wire  _EVAL_178;
  wire  _EVAL_183;
  wire  _EVAL_210;
  wire  _EVAL_253;
  wire  _EVAL_224;
  wire  _EVAL_149;
  wire  _EVAL_241;
  wire [4:0] _EVAL_165;
  wire  _EVAL_63;
  wire  _EVAL_187;
  wire  _EVAL_176;
  wire  _EVAL_151;
  wire  _EVAL_267;
  wire  _EVAL_90;
  wire  _EVAL_215;
  wire  _EVAL_66;
  wire  _EVAL_269;
  wire  _EVAL_194;
  wire  _EVAL_100;
  wire [2:0] _EVAL_208;
  wire  _EVAL_217;
  wire  _EVAL_271;
  wire  _EVAL_167;
  wire  _EVAL_205;
  wire [1:0] _EVAL_128;
  wire  _EVAL_223;
  wire  _EVAL_114;
  wire  _EVAL_213;
  wire  _EVAL_157;
  wire  _EVAL_214;
  wire [2:0] _EVAL_170;
  wire  _EVAL_193;
  wire  _EVAL_108;
  wire  _EVAL_84;
  wire  _EVAL_164;
  wire  _EVAL_93;
  wire [32:0] _EVAL_236;
  wire [32:0] _EVAL_140;
  wire  _EVAL_162;
  wire  _EVAL_94;
  wire [1:0] _EVAL_279;
  wire  _EVAL_247;
  wire [32:0] _EVAL_70;
  wire  _EVAL_255;
  wire [2:0] _EVAL_156;
  wire  _EVAL_196;
  wire [32:0] _EVAL_106;
  SiFive__EVAL_302 simpleOps (
    ._EVAL(simpleOps__EVAL),
    ._EVAL_0(simpleOps__EVAL_0),
    ._EVAL_1(simpleOps__EVAL_1),
    ._EVAL_2(simpleOps__EVAL_2),
    ._EVAL_3(simpleOps__EVAL_3),
    ._EVAL_4(simpleOps__EVAL_4),
    ._EVAL_5(simpleOps__EVAL_5),
    ._EVAL_6(simpleOps__EVAL_6),
    ._EVAL_7(simpleOps__EVAL_7),
    ._EVAL_8(simpleOps__EVAL_8),
    ._EVAL_9(simpleOps__EVAL_9),
    ._EVAL_10(simpleOps__EVAL_10),
    ._EVAL_11(simpleOps__EVAL_11),
    ._EVAL_12(simpleOps__EVAL_12)
  );
  SiFive__EVAL_296 divSqrts_0 (
    ._EVAL(divSqrts_0__EVAL),
    ._EVAL_0(divSqrts_0__EVAL_0),
    ._EVAL_1(divSqrts_0__EVAL_1),
    ._EVAL_2(divSqrts_0__EVAL_2),
    ._EVAL_3(divSqrts_0__EVAL_3),
    ._EVAL_4(divSqrts_0__EVAL_4),
    ._EVAL_5(divSqrts_0__EVAL_5),
    ._EVAL_6(divSqrts_0__EVAL_6),
    ._EVAL_7(divSqrts_0__EVAL_7),
    ._EVAL_8(divSqrts_0__EVAL_8),
    ._EVAL_9(divSqrts_0__EVAL_9),
    ._EVAL_10(divSqrts_0__EVAL_10),
    ._EVAL_11(divSqrts_0__EVAL_11)
  );
  SiFive__EVAL_293 fmas_0 (
    ._EVAL(fmas_0__EVAL),
    ._EVAL_0(fmas_0__EVAL_0),
    ._EVAL_1(fmas_0__EVAL_1),
    ._EVAL_2(fmas_0__EVAL_2),
    ._EVAL_3(fmas_0__EVAL_3),
    ._EVAL_4(fmas_0__EVAL_4),
    ._EVAL_5(fmas_0__EVAL_5),
    ._EVAL_6(fmas_0__EVAL_6),
    ._EVAL_7(fmas_0__EVAL_7),
    ._EVAL_8(fmas_0__EVAL_8)
  );
  assign _EVAL_142 = _EVAL_59[6:2];
  assign _EVAL_273 = _EVAL_142 == 5'h0;
  assign _EVAL_243 = _EVAL_142 == 5'h1;
  assign _EVAL_68 = _EVAL_273 | _EVAL_243;
  assign _EVAL_74 = _EVAL_44 | _EVAL_68;
  assign _EVAL_145 = _EVAL_142 == 5'h2;
  assign _EVAL_174 = _EVAL_74 | _EVAL_145;
  assign _EVAL_95 = _EVAL_142 == 5'h3;
  assign _EVAL_82 = _EVAL_142 == 5'h7;
  assign _EVAL_121 = _EVAL_95 | _EVAL_82;
  assign _EVAL_123 = _EVAL_142 == 5'hb;
  assign _EVAL_91 = _EVAL_121 | _EVAL_123;
  assign _EVAL_259 = _EVAL_142 == 5'hf;
  assign _EVAL_226 = _EVAL_91 | _EVAL_259;
  assign _EVAL_268 = _EVAL_174 | _EVAL_226;
  assign _EVAL_179 = _EVAL_268 == 1'h0;
  assign _EVAL_248 = {{2'd0}, _EVAL_179};
  assign _EVAL_195 = _EVAL_257 == 1'h0;
  assign _EVAL_81 = _EVAL_110[6:2];
  assign _EVAL_131 = _EVAL_81 == 5'h3;
  assign _EVAL_202 = _EVAL_81 == 5'h7;
  assign _EVAL_220 = _EVAL_131 | _EVAL_202;
  assign _EVAL_113 = _EVAL_81 == 5'hb;
  assign _EVAL_206 = _EVAL_220 | _EVAL_113;
  assign _EVAL_203 = _EVAL_81 == 5'hf;
  assign _EVAL_228 = _EVAL_206 | _EVAL_203;
  assign _EVAL_173 = _EVAL_195 & _EVAL_228;
  assign _EVAL_212 = _EVAL_20 | _EVAL_22;
  assign _EVAL_78 = _EVAL_212 | _EVAL_8;
  assign _EVAL_163 = _EVAL_17[6:2];
  assign _EVAL_152 = _EVAL_117[6:2];
  assign _EVAL_198 = _EVAL_152 == 5'h3;
  assign _EVAL_86 = _EVAL_152 == 5'h7;
  assign _EVAL_76 = _EVAL_198 | _EVAL_86;
  assign _EVAL_251 = _EVAL_152 == 5'hb;
  assign _EVAL_115 = _EVAL_76 | _EVAL_251;
  assign _EVAL_155 = _EVAL_152 == 5'hf;
  assign _EVAL_275 = _EVAL_115 | _EVAL_155;
  assign _EVAL_190 = _EVAL_50[6:2];
  assign _EVAL_109 = _EVAL_190 == 5'h3;
  assign _EVAL_258 = _EVAL_163 == 5'h0;
  assign _EVAL_242 = _EVAL_163 == 5'h1;
  assign _EVAL_204 = _EVAL_258 | _EVAL_242;
  assign _EVAL_264 = _EVAL_7 | _EVAL_204;
  assign _EVAL_245 = _EVAL_13 & _EVAL_4;
  assign _EVAL_150 = _EVAL_3[6:2];
  assign _EVAL_261 = _EVAL_150 == 5'h0;
  assign _EVAL_221 = _EVAL_150 == 5'h1;
  assign _EVAL_209 = _EVAL_261 | _EVAL_221;
  assign _EVAL_254 = _EVAL_14 | _EVAL_209;
  assign _EVAL_112 = _EVAL_104[1];
  assign _EVAL_105 = _EVAL_112 ? 33'h100000000 : 33'h0;
  assign _EVAL_154 = _EVAL_62 == 1'h0;
  assign _EVAL_136 = _EVAL_154 & _EVAL_275;
  assign _EVAL_96 = _EVAL_23[6:2];
  assign _EVAL_260 = _EVAL_96 == 5'h0;
  assign _EVAL_229 = _EVAL_96 == 5'h1;
  assign _EVAL_201 = _EVAL_260 | _EVAL_229;
  assign _EVAL_61 = _EVAL_53 | _EVAL_201;
  assign _EVAL_237 = _EVAL_96 == 5'h2;
  assign _EVAL_99 = _EVAL_61 | _EVAL_237;
  assign _EVAL_278 = _EVAL_189 == 1'h0;
  assign _EVAL_277 = _EVAL_186 != 5'h0;
  assign _EVAL_135 = _EVAL_186 - 5'h1;
  assign _EVAL_124 = _EVAL_64 == 1'h0;
  assign _EVAL_240 = _EVAL_182[6:2];
  assign _EVAL_252 = _EVAL_240 == 5'h3;
  assign _EVAL_175 = _EVAL_240 == 5'h7;
  assign _EVAL_71 = _EVAL_252 | _EVAL_175;
  assign _EVAL_134 = _EVAL_240 == 5'hb;
  assign _EVAL_137 = _EVAL_71 | _EVAL_134;
  assign _EVAL_270 = _EVAL_240 == 5'hf;
  assign _EVAL_120 = _EVAL_137 | _EVAL_270;
  assign _EVAL_97 = _EVAL_124 & _EVAL_120;
  assign _EVAL_118 = _EVAL_227 & _EVAL_97;
  assign _EVAL_262 = _EVAL_118 ? 1'h0 : 1'h1;
  assign _EVAL_250 = divSqrts_0__EVAL_6 & divSqrts_0__EVAL_3;
  assign _EVAL_79 = _EVAL_190 == 5'hb;
  assign _EVAL_139 = _EVAL_58 | _EVAL_38;
  assign _EVAL_132 = _EVAL_190 == 5'h1;
  assign _EVAL_239 = _EVAL_92 ^ _EVAL_192;
  assign _EVAL_73 = _EVAL_190 == 5'h7;
  assign _EVAL_101 = _EVAL_109 | _EVAL_73;
  assign _EVAL_69 = _EVAL_104[0];
  assign _EVAL_238 = _EVAL_240[0];
  assign _EVAL_230 = _EVAL_124 & _EVAL_238;
  assign _EVAL_211 = _EVAL_69 | _EVAL_230;
  assign _EVAL_265 = _EVAL_211 ? 33'h100000000 : 33'h0;
  assign _EVAL_207 = _EVAL_119 ^ _EVAL_265;
  assign _EVAL_122 = _EVAL_190 == 5'h0;
  assign _EVAL_141 = _EVAL_92[23];
  assign _EVAL_111 = _EVAL_256 == 1'h0;
  assign _EVAL_144 = _EVAL_177[6:2];
  assign _EVAL_130 = _EVAL_144 == 5'h3;
  assign _EVAL_88 = _EVAL_144 == 5'h7;
  assign _EVAL_126 = _EVAL_130 | _EVAL_88;
  assign _EVAL_225 = _EVAL_144 == 5'hb;
  assign _EVAL_159 = _EVAL_126 | _EVAL_225;
  assign _EVAL_85 = _EVAL_144 == 5'hf;
  assign _EVAL_102 = _EVAL_159 | _EVAL_85;
  assign _EVAL_87 = _EVAL_111 & _EVAL_102;
  assign _EVAL_172 = _EVAL_77 & _EVAL_87;
  assign _EVAL_185 = _EVAL_160 & _EVAL_173;
  assign _EVAL_178 = _EVAL_185 ? 1'h0 : _EVAL_262;
  assign _EVAL_183 = _EVAL_172 ? 1'h0 : _EVAL_178;
  assign _EVAL_210 = _EVAL_83 == 1'h0;
  assign _EVAL_253 = _EVAL_1 == 1'h0;
  assign _EVAL_224 = _EVAL_160 & _EVAL_253;
  assign _EVAL_149 = _EVAL_116 == 1'h0;
  assign _EVAL_241 = fmas_0__EVAL_5;
  assign _EVAL_165 = _EVAL_241 ? fmas_0__EVAL_0 : _EVAL_197;
  assign _EVAL_63 = _EVAL_122 | _EVAL_132;
  assign _EVAL_187 = _EVAL_58 | _EVAL_63;
  assign _EVAL_176 = _EVAL_190 == 5'h2;
  assign _EVAL_151 = _EVAL_187 | _EVAL_176;
  assign _EVAL_267 = _EVAL_101 | _EVAL_79;
  assign _EVAL_90 = _EVAL_190 == 5'hf;
  assign _EVAL_215 = _EVAL_267 | _EVAL_90;
  assign _EVAL_66 = _EVAL_151 | _EVAL_215;
  assign _EVAL_269 = _EVAL_190[1];
  assign _EVAL_194 = _EVAL_138 == 1'h0;
  assign _EVAL_100 = _EVAL_194 == 1'h0;
  assign _EVAL_208 = _EVAL_174 ? 3'h4 : 3'h0;
  assign _EVAL_217 = _EVAL_58 | _EVAL_269;
  assign _EVAL_271 = _EVAL_151 & _EVAL_217;
  assign _EVAL_167 = _EVAL_150 == 5'h2;
  assign _EVAL_205 = _EVAL_254 | _EVAL_167;
  assign _EVAL_128 = _EVAL_205 ? 2'h3 : 2'h0;
  assign _EVAL_223 = _EVAL_181 & _EVAL_136;
  assign _EVAL_114 = _EVAL_223 ? 1'h0 : _EVAL_183;
  assign _EVAL_213 = _EVAL_41 & _EVAL_49;
  assign _EVAL_157 = _EVAL_213 & _EVAL_4;
  assign _EVAL_214 = divSqrts_0__EVAL_1 & divSqrts_0__EVAL_4;
  assign _EVAL_170 = _EVAL_151 ? 3'h4 : 3'h0;
  assign _EVAL_193 = _EVAL_78 | _EVAL_48;
  assign _EVAL_108 = _EVAL_269 == 1'h0;
  assign _EVAL_84 = _EVAL_58 | _EVAL_108;
  assign _EVAL_164 = _EVAL_151 & _EVAL_84;
  assign _EVAL_93 = _EVAL_163 == 5'h2;
  assign _EVAL_236 = _EVAL_241 ? fmas_0__EVAL_8 : _EVAL_75;
  assign _EVAL_140 = _EVAL_194 ? 33'h0 : _EVAL_239;
  assign _EVAL_162 = _EVAL_58 == 1'h0;
  assign _EVAL_94 = _EVAL_264 | _EVAL_93;
  assign _EVAL_279 = _EVAL_94 ? 2'h2 : 2'h0;
  assign _EVAL_247 = _EVAL_66 == 1'h0;
  assign _EVAL_70 = 33'h100000000 & _EVAL_140;
  assign _EVAL_255 = divSqrts_0__EVAL_4 | _EVAL_13;
  assign _EVAL_156 = {{2'd0}, _EVAL_247};
  assign _EVAL_196 = divSqrts_0__EVAL_6 == 1'h0;
  assign _EVAL_106 = _EVAL_92 ^ _EVAL_105;
  assign _EVAL_16 = _EVAL_125;
  assign _EVAL_44 = _EVAL_64;
  assign _EVAL_25 = _EVAL_276;
  assign _EVAL_26 = _EVAL_234;
  assign _EVAL_40 = _EVAL_255 | _EVAL_193;
  assign _EVAL_8 = _EVAL_77;
  assign divSqrts_0__EVAL_8 = _EVAL_192;
  assign divSqrts_0__EVAL_11 = _EVAL_67 == 1'h0;
  assign _EVAL_0 = _EVAL_156 | _EVAL_170;
  assign _EVAL_60 = simpleOps__EVAL_3;
  assign _EVAL_9 = simpleOps__EVAL_2;
  assign simpleOps__EVAL = _EVAL_67;
  assign _EVAL_47 = _EVAL_171 ? _EVAL_197 : _EVAL_165;
  assign _EVAL_52 = 1'h1;
  assign divSqrts_0__EVAL_1 = _EVAL_181 ? 1'h0 : _EVAL_114;
  assign _EVAL_7 = _EVAL_256;
  assign _EVAL_57 = _EVAL_233;
  assign _EVAL_13 = divSqrts_0__EVAL_3 | _EVAL_196;
  assign simpleOps__EVAL_9 = _EVAL_149 ? 33'he0400000 : _EVAL_92;
  assign _EVAL_20 = _EVAL_227;
  assign _EVAL_56 = _EVAL_232;
  assign _EVAL_51 = {{2'd0}, _EVAL_99};
  assign _EVAL_54 = _EVAL_186;
  assign fmas_0__EVAL_2 = _EVAL_98;
  assign simpleOps__EVAL_1 = _EVAL;
  assign divSqrts_0__EVAL_2 = _EVAL_185 ? _EVAL_1 : 1'h0;
  assign _EVAL_48 = _EVAL_181;
  assign divSqrts_0__EVAL_10 = _EVAL_92;
  assign simpleOps__EVAL_8 = _EVAL_227 & _EVAL_116;
  assign simpleOps__EVAL_4 = _EVAL_148;
  assign _EVAL_2 = _EVAL_127;
  assign _EVAL_4 = _EVAL_162 & _EVAL_215;
  assign _EVAL_43 = _EVAL_219;
  assign fmas_0__EVAL_6 = _EVAL_46;
  assign divSqrts_0__EVAL_7 = _EVAL_46;
  assign _EVAL_42 = _EVAL_222;
  assign fmas_0__EVAL = _EVAL_194 ? 33'h80000000 : _EVAL_106;
  assign _EVAL_34 = {{1'd0}, _EVAL_279};
  assign _EVAL_59 = _EVAL_182;
  assign simpleOps__EVAL_5 = _EVAL_246;
  assign _EVAL_24 = _EVAL_188;
  assign _EVAL_53 = _EVAL_62;
  assign fmas_0__EVAL_3 = _EVAL;
  assign divSqrts_0__EVAL_0 = _EVAL_98;
  assign simpleOps__EVAL_11 = _EVAL_149 ? 33'he0400000 : _EVAL_192;
  assign _EVAL_23 = _EVAL_117;
  assign _EVAL_17 = _EVAL_177;
  assign _EVAL_37 = _EVAL_200;
  assign fmas_0__EVAL_4 = _EVAL_278 ? _EVAL_70 : _EVAL_207;
  assign _EVAL_22 = _EVAL_160;
  assign _EVAL_41 = _EVAL_245 == 1'h0;
  assign fmas_0__EVAL_1 = _EVAL_210 ? 33'h80000000 : _EVAL_192;
  assign _EVAL_35 = _EVAL_249;
  assign simpleOps__EVAL_6 = _EVAL_125;
  assign simpleOps__EVAL_10 = _EVAL_191;
  assign _EVAL_30 = _EVAL_146;
  assign _EVAL_3 = _EVAL_110;
  assign divSqrts_0__EVAL_3 = _EVAL_227 & _EVAL_97;
  assign fmas_0__EVAL_7 = _EVAL_227 & _EVAL_100;
  assign _EVAL_14 = _EVAL_257;
  assign _EVAL_45 = simpleOps__EVAL_7;
  assign _EVAL_29 = _EVAL_158;
  assign simpleOps__EVAL_0 = _EVAL_182;
  assign _EVAL_10 = _EVAL_248 | _EVAL_208;
  assign _EVAL_21 = _EVAL_171 ? _EVAL_75 : _EVAL_236;
  assign _EVAL_12 = _EVAL_143;
  assign _EVAL_55 = _EVAL_216;
  assign simpleOps__EVAL_12 = _EVAL_98;
  assign divSqrts_0__EVAL_5 = _EVAL;
  assign _EVAL_39 = {{1'd0}, _EVAL_128};
  assign _EVAL_18 = _EVAL_80;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_62 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_64 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_67 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  _EVAL_75 = _RAND_3[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_77 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_80 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_83 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _EVAL_92 = _RAND_7[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_98 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_104 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_110 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_116 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_117 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _EVAL_119 = _RAND_13[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_125 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _EVAL_127 = _RAND_15[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_138 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_143 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _EVAL_146 = _RAND_18[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_148 = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_158 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_160 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_171 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_177 = _RAND_23[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_181 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_182 = _RAND_25[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_186 = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_188 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_189 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_191 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _EVAL_192 = _RAND_30[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_197 = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_200 = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_216 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_219 = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_222 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_227 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_232 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_233 = _RAND_38[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_234 = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_246 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_249 = _RAND_41[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_256 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_257 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_276 = _RAND_44[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_77) begin
      _EVAL_62 <= _EVAL_256;
    end
    if (_EVAL_213) begin
      _EVAL_64 <= _EVAL_58;
    end
    if (_EVAL_213) begin
      _EVAL_67 <= _EVAL_38;
    end
    if (_EVAL_214) begin
      _EVAL_75 <= divSqrts_0__EVAL_9;
    end else begin
      if (_EVAL_181) begin
        _EVAL_75 <= _EVAL_2;
      end
    end
    if (_EVAL_46) begin
      _EVAL_77 <= 1'h0;
    end else begin
      _EVAL_77 <= _EVAL_224;
    end
    if (_EVAL_77) begin
      _EVAL_80 <= _EVAL_43;
    end
    if (_EVAL_213) begin
      _EVAL_83 <= _EVAL_271;
    end
    if (_EVAL_213) begin
      if (_EVAL_15) begin
        _EVAL_92 <= _EVAL_6;
      end
    end
    if (_EVAL_213) begin
      _EVAL_98 <= _EVAL_31;
    end
    if (_EVAL_213) begin
      _EVAL_104 <= _EVAL_5;
    end
    if (_EVAL_227) begin
      _EVAL_110 <= _EVAL_182;
    end
    if (_EVAL_213) begin
      _EVAL_116 <= _EVAL_247;
    end
    if (_EVAL_77) begin
      _EVAL_117 <= _EVAL_177;
    end
    if (_EVAL_213) begin
      if (_EVAL_139) begin
        _EVAL_119 <= _EVAL_19;
      end
    end
    if (_EVAL_213) begin
      _EVAL_125 <= _EVAL_36;
    end
    if (_EVAL_77) begin
      _EVAL_127 <= _EVAL_30;
    end
    if (_EVAL_213) begin
      _EVAL_138 <= _EVAL_151;
    end
    if (_EVAL_46) begin
      _EVAL_143 <= 1'h0;
    end else begin
      if (_EVAL_214) begin
        _EVAL_143 <= 1'h1;
      end else begin
        if (_EVAL_181) begin
          if (_EVAL_136) begin
            _EVAL_143 <= 1'h0;
          end else begin
            _EVAL_143 <= _EVAL_181;
          end
        end else begin
          _EVAL_143 <= _EVAL_181;
        end
      end
    end
    if (_EVAL_160) begin
      _EVAL_146 <= _EVAL_60;
    end
    if (_EVAL_213) begin
      _EVAL_148 <= _EVAL_28;
    end
    if (_EVAL_214) begin
      _EVAL_158 <= _EVAL_37;
    end else begin
      if (_EVAL_181) begin
        _EVAL_158 <= _EVAL_276;
      end
    end
    if (_EVAL_46) begin
      _EVAL_160 <= 1'h0;
    end else begin
      _EVAL_160 <= _EVAL_227;
    end
    _EVAL_171 <= divSqrts_0__EVAL_1 & divSqrts_0__EVAL_4;
    if (_EVAL_160) begin
      _EVAL_177 <= _EVAL_110;
    end
    if (_EVAL_46) begin
      _EVAL_181 <= 1'h0;
    end else begin
      _EVAL_181 <= _EVAL_77;
    end
    if (_EVAL_213) begin
      _EVAL_182 <= _EVAL_50;
    end
    if (_EVAL_250) begin
      if (divSqrts_0__EVAL_11) begin
        if (_EVAL_141) begin
          _EVAL_186 <= 5'h18;
        end else begin
          _EVAL_186 <= 5'h19;
        end
      end else begin
        _EVAL_186 <= 5'h1a;
      end
    end else begin
      if (_EVAL_157) begin
        _EVAL_186 <= 5'h1b;
      end else begin
        if (_EVAL_277) begin
          _EVAL_186 <= _EVAL_135;
        end
      end
    end
    if (_EVAL_160) begin
      _EVAL_188 <= _EVAL_232;
    end
    if (_EVAL_213) begin
      _EVAL_189 <= _EVAL_164;
    end
    if (_EVAL_213) begin
      _EVAL_191 <= _EVAL_15;
    end
    if (_EVAL_213) begin
      if (_EVAL_38) begin
        _EVAL_192 <= _EVAL_32;
      end
    end
    if (_EVAL_214) begin
      _EVAL_197 <= divSqrts_0__EVAL;
    end else begin
      if (_EVAL_181) begin
        _EVAL_197 <= _EVAL_18;
      end
    end
    if (_EVAL_157) begin
      _EVAL_200 <= _EVAL_11;
    end
    if (_EVAL_214) begin
      _EVAL_216 <= _EVAL_52;
    end else begin
      if (_EVAL_181) begin
        _EVAL_216 <= _EVAL_222;
      end
    end
    if (_EVAL_160) begin
      _EVAL_219 <= _EVAL_45;
    end
    if (_EVAL_77) begin
      _EVAL_222 <= _EVAL_188;
    end
    _EVAL_227 <= _EVAL_41 & _EVAL_49;
    if (_EVAL_227) begin
      _EVAL_232 <= _EVAL_125;
    end
    if (_EVAL_160) begin
      _EVAL_233 <= _EVAL_234;
    end
    if (_EVAL_227) begin
      _EVAL_234 <= _EVAL_249;
    end
    if (_EVAL_213) begin
      if (_EVAL_33) begin
        _EVAL_246 <= _EVAL_27;
      end
    end
    if (_EVAL_213) begin
      _EVAL_249 <= _EVAL_11;
    end
    if (_EVAL_160) begin
      _EVAL_256 <= _EVAL_257;
    end
    if (_EVAL_227) begin
      _EVAL_257 <= _EVAL_64;
    end
    if (_EVAL_77) begin
      _EVAL_276 <= _EVAL_233;
    end
  end
endmodule
