//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_113_assert(
  input  [2:0]  _EVAL,
  input  [1:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [29:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [6:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [6:0]  _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [6:0] _EVAL_28;
  reg [31:0] _RAND_0;
  reg  _EVAL_31;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_83;
  reg [31:0] _RAND_2;
  reg [29:0] _EVAL_96;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_97;
  reg [31:0] _RAND_4;
  reg [5:0] _EVAL_121;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_166;
  reg [31:0] _RAND_6;
  reg [5:0] _EVAL_212;
  reg [31:0] _RAND_7;
  reg [31:0] _EVAL_214;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_227;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_237;
  reg [31:0] _RAND_10;
  reg [6:0] _EVAL_261;
  reg [31:0] _RAND_11;
  reg [5:0] _EVAL_276;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_324;
  reg [31:0] _RAND_13;
  reg [72:0] _EVAL_350;
  reg [95:0] _RAND_14;
  reg  _EVAL_355;
  reg [31:0] _RAND_15;
  reg [1:0] _EVAL_361;
  reg [31:0] _RAND_16;
  wire  _EVAL_190;
  wire  _EVAL_255;
  wire  _EVAL_133;
  wire [3:0] _EVAL_312;
  wire  _EVAL_198;
  wire [2:0] _EVAL_109;
  wire  _EVAL_29;
  wire  _EVAL_63;
  wire  _EVAL_72;
  wire  _EVAL_36;
  wire  _EVAL_358;
  wire  _EVAL_65;
  wire  _EVAL_293;
  wire  _EVAL_39;
  wire  _EVAL_314;
  wire  _EVAL_100;
  wire  _EVAL_205;
  wire  _EVAL_91;
  wire  _EVAL_254;
  wire [22:0] _EVAL_199;
  wire [7:0] _EVAL_229;
  wire [7:0] _EVAL_107;
  wire [5:0] _EVAL_111;
  wire [5:0] _EVAL_315;
  wire [29:0] _EVAL_154;
  wire [30:0] _EVAL_287;
  wire [30:0] _EVAL_114;
  wire [30:0] _EVAL_363;
  wire  _EVAL_20;
  wire [127:0] _EVAL_175;
  wire [29:0] _EVAL_165;
  wire [30:0] _EVAL_278;
  wire [30:0] _EVAL_23;
  wire [30:0] _EVAL_296;
  wire  _EVAL_171;
  wire [29:0] _EVAL_325;
  wire  _EVAL_176;
  wire  _EVAL_76;
  wire  _EVAL_279;
  wire  _EVAL_351;
  wire  _EVAL_217;
  wire  _EVAL_42;
  wire  _EVAL_232;
  wire  _EVAL_197;
  wire  _EVAL_61;
  wire  _EVAL_290;
  wire [127:0] _EVAL_188;
  wire [72:0] _EVAL_265;
  wire [72:0] _EVAL_334;
  wire [72:0] _EVAL_260;
  wire  _EVAL_174;
  wire  _EVAL_346;
  wire  _EVAL_228;
  wire [22:0] _EVAL_50;
  wire [7:0] _EVAL_366;
  wire [7:0] _EVAL_248;
  wire [5:0] _EVAL_230;
  wire [5:0] _EVAL_353;
  wire  _EVAL_24;
  wire  _EVAL_48;
  wire  _EVAL_289;
  wire [29:0] _EVAL_362;
  wire  _EVAL_368;
  wire [29:0] _EVAL_354;
  wire [30:0] _EVAL_213;
  wire [30:0] _EVAL_84;
  wire [30:0] _EVAL_356;
  wire  _EVAL_85;
  wire  _EVAL_286;
  wire [30:0] _EVAL_115;
  wire [30:0] _EVAL_147;
  wire [30:0] _EVAL_302;
  wire  _EVAL_145;
  wire  _EVAL_123;
  wire [3:0] _EVAL_159;
  wire  _EVAL_195;
  wire [29:0] _EVAL_89;
  wire [30:0] _EVAL_342;
  wire [30:0] _EVAL_273;
  wire [30:0] _EVAL_127;
  wire  _EVAL_196;
  wire  _EVAL_136;
  wire [30:0] _EVAL_86;
  wire [30:0] _EVAL_60;
  wire [30:0] _EVAL_69;
  wire  _EVAL_34;
  wire  _EVAL_371;
  wire [30:0] _EVAL_41;
  wire [30:0] _EVAL_82;
  wire [30:0] _EVAL_93;
  wire  _EVAL_359;
  wire  _EVAL_59;
  wire  _EVAL_87;
  wire  _EVAL_193;
  wire  _EVAL_204;
  wire  _EVAL_219;
  wire  _EVAL_291;
  wire  _EVAL_49;
  wire  _EVAL_277;
  wire  _EVAL_44;
  wire  _EVAL_344;
  wire  _EVAL_95;
  wire  _EVAL_146;
  wire  _EVAL_27;
  wire  _EVAL_235;
  wire  _EVAL_57;
  wire  _EVAL_184;
  wire [72:0] _EVAL_104;
  wire [29:0] _EVAL_112;
  wire [29:0] _EVAL_216;
  wire  _EVAL_304;
  wire  _EVAL_30;
  wire  _EVAL_347;
  wire  _EVAL_222;
  wire  _EVAL_58;
  wire  _EVAL_134;
  wire [127:0] _EVAL_266;
  wire [127:0] _EVAL_340;
  wire [72:0] _EVAL_186;
  wire  _EVAL_337;
  wire  _EVAL_318;
  wire  _EVAL_224;
  wire  _EVAL_321;
  wire  _EVAL_241;
  wire  _EVAL_299;
  wire  _EVAL_38;
  wire  _EVAL_239;
  wire [1:0] _EVAL_345;
  wire [1:0] _EVAL_173;
  wire  _EVAL_256;
  wire  _EVAL_211;
  wire  _EVAL_187;
  wire  _EVAL_294;
  wire  _EVAL_335;
  wire  _EVAL_47;
  wire  _EVAL_52;
  wire  _EVAL_99;
  wire  _EVAL_178;
  wire  _EVAL_162;
  wire  _EVAL_108;
  wire  _EVAL_117;
  wire  _EVAL_66;
  wire  _EVAL_45;
  wire  _EVAL_206;
  wire  _EVAL_240;
  wire  _EVAL_129;
  wire  _EVAL_168;
  wire [3:0] _EVAL_223;
  wire [3:0] _EVAL_333;
  wire [3:0] _EVAL_336;
  wire  _EVAL_179;
  wire  _EVAL_307;
  wire  _EVAL_274;
  wire  _EVAL_236;
  wire  _EVAL_367;
  wire  _EVAL_157;
  wire  _EVAL_226;
  wire  _EVAL_330;
  wire  _EVAL_251;
  wire  _EVAL_282;
  wire [72:0] _EVAL_110;
  wire  _EVAL_267;
  wire  _EVAL_292;
  wire  _EVAL_281;
  wire  _EVAL_221;
  wire  _EVAL_137;
  wire  _EVAL_142;
  wire  _EVAL_308;
  wire  _EVAL_90;
  wire  _EVAL_357;
  wire  _EVAL_349;
  wire  _EVAL_288;
  wire  _EVAL_317;
  wire  _EVAL_189;
  wire  _EVAL_98;
  wire  _EVAL_319;
  wire  _EVAL_126;
  wire  _EVAL_118;
  wire  _EVAL_210;
  wire  _EVAL_155;
  wire  _EVAL_249;
  wire  _EVAL_144;
  wire  _EVAL_306;
  wire  _EVAL_125;
  wire  _EVAL_202;
  wire  _EVAL_139;
  wire  _EVAL_322;
  wire  _EVAL_148;
  wire  _EVAL_339;
  wire  _EVAL_218;
  wire  _EVAL_46;
  wire  _EVAL_243;
  wire  _EVAL_67;
  wire  _EVAL_343;
  wire  _EVAL_183;
  wire  _EVAL_268;
  wire  _EVAL_297;
  wire  _EVAL_113;
  wire  _EVAL_284;
  wire  _EVAL_71;
  wire  _EVAL_338;
  wire  _EVAL_25;
  wire  _EVAL_250;
  wire  _EVAL_94;
  wire  _EVAL_130;
  wire  _EVAL_327;
  wire [72:0] _EVAL_138;
  wire  _EVAL_208;
  wire  _EVAL_56;
  wire  _EVAL_26;
  wire [2:0] _EVAL_140;
  wire [3:0] _EVAL_275;
  wire  _EVAL_231;
  wire  _EVAL_103;
  wire  _EVAL_329;
  wire  _EVAL_215;
  wire  _EVAL_101;
  wire  _EVAL_194;
  wire  _EVAL_102;
  wire  _EVAL_207;
  wire  _EVAL_55;
  wire  _EVAL_180;
  wire  _EVAL_158;
  wire  _EVAL_53;
  wire  _EVAL_19;
  wire  _EVAL_238;
  wire  _EVAL_203;
  wire  _EVAL_106;
  wire  _EVAL_141;
  wire  _EVAL_311;
  wire  _EVAL_264;
  wire  _EVAL_105;
  wire  _EVAL_167;
  wire  _EVAL_182;
  wire  _EVAL_259;
  wire [31:0] _EVAL_160;
  wire  _EVAL_209;
  wire  _EVAL_326;
  wire  _EVAL_242;
  wire  _EVAL_75;
  wire  _EVAL_332;
  wire  _EVAL_119;
  wire  _EVAL_149;
  wire  _EVAL_269;
  wire  _EVAL_246;
  wire  _EVAL_32;
  wire  _EVAL_22;
  wire  _EVAL_170;
  wire [5:0] _EVAL_253;
  wire  _EVAL_247;
  wire  _EVAL_369;
  wire  _EVAL_352;
  wire  _EVAL_77;
  wire  _EVAL_35;
  wire  _EVAL_271;
  wire  _EVAL_177;
  wire  _EVAL_348;
  wire  _EVAL_220;
  wire  _EVAL_128;
  wire  _EVAL_233;
  wire  _EVAL_201;
  wire  _EVAL_152;
  wire  _EVAL_257;
  wire  _EVAL_124;
  wire  _EVAL_305;
  wire  _EVAL_252;
  wire  _EVAL_88;
  wire  _EVAL_64;
  wire  _EVAL_234;
  wire  _EVAL_122;
  wire  _EVAL_51;
  wire  _EVAL_54;
  wire  _EVAL_181;
  wire  _EVAL_331;
  wire  _EVAL_132;
  wire  _EVAL_301;
  wire  _EVAL_298;
  wire  _EVAL_360;
  wire  _EVAL_79;
  wire  _EVAL_68;
  wire  _EVAL_200;
  wire  _EVAL_283;
  wire  _EVAL_40;
  wire  _EVAL_323;
  wire  _EVAL_225;
  wire [5:0] _EVAL_151;
  wire  _EVAL_37;
  wire  _EVAL_78;
  wire  _EVAL_131;
  wire  _EVAL_309;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_43;
  wire  _EVAL_328;
  wire  _EVAL_161;
  wire  _EVAL_262;
  wire  _EVAL_21;
  wire  _EVAL_163;
  wire  _EVAL_74;
  wire  _EVAL_244;
  wire  _EVAL_92;
  wire  _EVAL_185;
  wire  _EVAL_303;
  wire  _EVAL_116;
  wire  _EVAL_143;
  wire  _EVAL_263;
  wire  _EVAL_150;
  wire  _EVAL_270;
  wire  _EVAL_80;
  wire  _EVAL_320;
  wire [72:0] _EVAL_300;
  wire  _EVAL_135;
  wire  _EVAL_70;
  wire  _EVAL_364;
  wire  _EVAL_73;
  wire  _EVAL_153;
  wire  _EVAL_280;
  wire  _EVAL_120;
  wire  _EVAL_164;
  wire  _EVAL_169;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_190 = _EVAL_13 == 7'h48;
  assign _EVAL_255 = _EVAL_13 == 7'h40;
  assign _EVAL_133 = _EVAL_190 | _EVAL_255;
  assign _EVAL_312 = _EVAL_13[6:3];
  assign _EVAL_198 = _EVAL_312 == 4'h8;
  assign _EVAL_109 = _EVAL_13[2:0];
  assign _EVAL_29 = 3'h1 <= _EVAL_109;
  assign _EVAL_63 = _EVAL_198 & _EVAL_29;
  assign _EVAL_72 = _EVAL_133 | _EVAL_63;
  assign _EVAL_36 = _EVAL_13 == 7'h20;
  assign _EVAL_358 = _EVAL_72 | _EVAL_36;
  assign _EVAL_65 = _EVAL_312 == 4'h0;
  assign _EVAL_293 = _EVAL_358 | _EVAL_65;
  assign _EVAL_39 = _EVAL == 3'h0;
  assign _EVAL_314 = _EVAL_1 == 3'h5;
  assign _EVAL_100 = _EVAL_12 & _EVAL_314;
  assign _EVAL_205 = _EVAL_16 == 7'h40;
  assign _EVAL_91 = _EVAL_276 == 6'h0;
  assign _EVAL_254 = _EVAL[0];
  assign _EVAL_199 = 23'hff << _EVAL_7;
  assign _EVAL_229 = _EVAL_199[7:0];
  assign _EVAL_107 = ~ _EVAL_229;
  assign _EVAL_111 = _EVAL_107[7:2];
  assign _EVAL_315 = _EVAL_276 - 6'h1;
  assign _EVAL_154 = _EVAL_2 ^ 30'h3000;
  assign _EVAL_287 = {1'b0,$signed(_EVAL_154)};
  assign _EVAL_114 = $signed(_EVAL_287) & $signed(-31'sh1000);
  assign _EVAL_363 = $signed(_EVAL_114);
  assign _EVAL_20 = $signed(_EVAL_363) == $signed(31'sh0);
  assign _EVAL_175 = 128'h1 << _EVAL_16;
  assign _EVAL_165 = _EVAL_2 ^ 30'hc000000;
  assign _EVAL_278 = {1'b0,$signed(_EVAL_165)};
  assign _EVAL_23 = $signed(_EVAL_278) & $signed(-31'sh4000000);
  assign _EVAL_296 = $signed(_EVAL_23);
  assign _EVAL_171 = $signed(_EVAL_296) == $signed(31'sh0);
  assign _EVAL_325 = _EVAL_2 ^ 30'h20000000;
  assign _EVAL_176 = _EVAL_0 == 2'h0;
  assign _EVAL_76 = _EVAL_176 | _EVAL_4;
  assign _EVAL_279 = _EVAL_76 == 1'h0;
  assign _EVAL_351 = _EVAL_6 <= 4'h8;
  assign _EVAL_217 = _EVAL_10 == _EVAL_324;
  assign _EVAL_42 = _EVAL_217 | _EVAL_4;
  assign _EVAL_232 = _EVAL_42 == 1'h0;
  assign _EVAL_197 = _EVAL_15 & _EVAL_12;
  assign _EVAL_61 = _EVAL_212 == 6'h0;
  assign _EVAL_290 = _EVAL_197 & _EVAL_61;
  assign _EVAL_188 = _EVAL_290 ? _EVAL_175 : 128'h0;
  assign _EVAL_265 = _EVAL_188[72:0];
  assign _EVAL_334 = _EVAL_265 | _EVAL_350;
  assign _EVAL_260 = _EVAL_334 >> _EVAL_13;
  assign _EVAL_174 = _EVAL_260[0];
  assign _EVAL_346 = _EVAL_1[2];
  assign _EVAL_228 = _EVAL_346 == 1'h0;
  assign _EVAL_50 = 23'hff << _EVAL_6;
  assign _EVAL_366 = _EVAL_50[7:0];
  assign _EVAL_248 = ~ _EVAL_366;
  assign _EVAL_230 = _EVAL_248[7:2];
  assign _EVAL_353 = _EVAL_212 - 6'h1;
  assign _EVAL_24 = _EVAL_10 <= 3'h4;
  assign _EVAL_48 = _EVAL_24 | _EVAL_4;
  assign _EVAL_289 = _EVAL_214 < plusarg_reader_out;
  assign _EVAL_362 = _EVAL_2 ^ 30'h1900000;
  assign _EVAL_368 = _EVAL_20 | _EVAL_171;
  assign _EVAL_354 = _EVAL_2 ^ 30'h2000000;
  assign _EVAL_213 = {1'b0,$signed(_EVAL_354)};
  assign _EVAL_84 = $signed(_EVAL_213) & $signed(-31'sh10000);
  assign _EVAL_356 = $signed(_EVAL_84);
  assign _EVAL_85 = $signed(_EVAL_356) == $signed(31'sh0);
  assign _EVAL_286 = _EVAL_368 | _EVAL_85;
  assign _EVAL_115 = {1'b0,$signed(_EVAL_2)};
  assign _EVAL_147 = $signed(_EVAL_115) & $signed(-31'sh5000);
  assign _EVAL_302 = $signed(_EVAL_147);
  assign _EVAL_145 = $signed(_EVAL_302) == $signed(31'sh0);
  assign _EVAL_123 = _EVAL_286 | _EVAL_145;
  assign _EVAL_159 = _EVAL_16[6:3];
  assign _EVAL_195 = _EVAL_159 == 4'h8;
  assign _EVAL_89 = _EVAL_2 ^ 30'h1800000;
  assign _EVAL_342 = {1'b0,$signed(_EVAL_89)};
  assign _EVAL_273 = $signed(_EVAL_342) & $signed(-31'sh8000);
  assign _EVAL_127 = $signed(_EVAL_273);
  assign _EVAL_196 = $signed(_EVAL_127) == $signed(31'sh0);
  assign _EVAL_136 = _EVAL_123 | _EVAL_196;
  assign _EVAL_86 = {1'b0,$signed(_EVAL_362)};
  assign _EVAL_60 = $signed(_EVAL_86) & $signed(-31'sh2000);
  assign _EVAL_69 = $signed(_EVAL_60);
  assign _EVAL_34 = $signed(_EVAL_69) == $signed(31'sh0);
  assign _EVAL_371 = _EVAL_136 | _EVAL_34;
  assign _EVAL_41 = {1'b0,$signed(_EVAL_325)};
  assign _EVAL_82 = $signed(_EVAL_41) & $signed(-31'sh2000);
  assign _EVAL_93 = $signed(_EVAL_82);
  assign _EVAL_359 = $signed(_EVAL_93) == $signed(31'sh0);
  assign _EVAL_59 = _EVAL_371 | _EVAL_359;
  assign _EVAL_87 = _EVAL_2[1];
  assign _EVAL_193 = _EVAL_87 == 1'h0;
  assign _EVAL_204 = _EVAL_2[0];
  assign _EVAL_219 = _EVAL_193 & _EVAL_204;
  assign _EVAL_291 = _EVAL_10 <= 3'h2;
  assign _EVAL_49 = _EVAL_291 | _EVAL_4;
  assign _EVAL_277 = _EVAL_6 <= 4'h2;
  assign _EVAL_44 = _EVAL_277 & _EVAL_59;
  assign _EVAL_344 = _EVAL_44 | _EVAL_4;
  assign _EVAL_95 = _EVAL <= 3'h6;
  assign _EVAL_146 = _EVAL_95 | _EVAL_4;
  assign _EVAL_27 = _EVAL_146 == 1'h0;
  assign _EVAL_235 = _EVAL_1 == 3'h7;
  assign _EVAL_57 = _EVAL_1 == 3'h1;
  assign _EVAL_184 = _EVAL_12 & _EVAL_57;
  assign _EVAL_104 = _EVAL_350 | _EVAL_265;
  assign _EVAL_112 = {{22'd0}, _EVAL_248};
  assign _EVAL_216 = _EVAL_2 & _EVAL_112;
  assign _EVAL_304 = _EVAL_216 == 30'h0;
  assign _EVAL_30 = _EVAL_11 & _EVAL_5;
  assign _EVAL_347 = _EVAL_30 & _EVAL_91;
  assign _EVAL_222 = _EVAL == 3'h6;
  assign _EVAL_58 = _EVAL_222 == 1'h0;
  assign _EVAL_134 = _EVAL_347 & _EVAL_58;
  assign _EVAL_266 = 128'h1 << _EVAL_13;
  assign _EVAL_340 = _EVAL_134 ? _EVAL_266 : 128'h0;
  assign _EVAL_186 = _EVAL_340[72:0];
  assign _EVAL_337 = _EVAL_265 != _EVAL_186;
  assign _EVAL_318 = _EVAL_265 != 73'h0;
  assign _EVAL_224 = _EVAL_318 == 1'h0;
  assign _EVAL_321 = _EVAL_337 | _EVAL_224;
  assign _EVAL_241 = _EVAL_321 | _EVAL_4;
  assign _EVAL_299 = _EVAL_312 == 4'h1;
  assign _EVAL_38 = _EVAL_6 >= 4'h2;
  assign _EVAL_239 = _EVAL_6[0];
  assign _EVAL_345 = 2'h1 << _EVAL_239;
  assign _EVAL_173 = _EVAL_345 | 2'h1;
  assign _EVAL_256 = _EVAL_173[1];
  assign _EVAL_211 = _EVAL_256 & _EVAL_87;
  assign _EVAL_187 = _EVAL_38 | _EVAL_211;
  assign _EVAL_294 = _EVAL_173[0];
  assign _EVAL_335 = _EVAL_87 & _EVAL_204;
  assign _EVAL_47 = _EVAL_294 & _EVAL_335;
  assign _EVAL_52 = _EVAL_187 | _EVAL_47;
  assign _EVAL_99 = _EVAL_204 == 1'h0;
  assign _EVAL_178 = _EVAL_87 & _EVAL_99;
  assign _EVAL_162 = _EVAL_294 & _EVAL_178;
  assign _EVAL_108 = _EVAL_187 | _EVAL_162;
  assign _EVAL_117 = _EVAL_256 & _EVAL_193;
  assign _EVAL_66 = _EVAL_38 | _EVAL_117;
  assign _EVAL_45 = _EVAL_294 & _EVAL_219;
  assign _EVAL_206 = _EVAL_66 | _EVAL_45;
  assign _EVAL_240 = _EVAL_193 & _EVAL_99;
  assign _EVAL_129 = _EVAL_294 & _EVAL_240;
  assign _EVAL_168 = _EVAL_66 | _EVAL_129;
  assign _EVAL_223 = {_EVAL_52,_EVAL_108,_EVAL_206,_EVAL_168};
  assign _EVAL_333 = ~ _EVAL_223;
  assign _EVAL_336 = _EVAL_9 & _EVAL_333;
  assign _EVAL_179 = _EVAL_336 == 4'h0;
  assign _EVAL_307 = _EVAL_350 != 73'h0;
  assign _EVAL_274 = _EVAL_307 == 1'h0;
  assign _EVAL_236 = plusarg_reader_out == 32'h0;
  assign _EVAL_367 = _EVAL_274 | _EVAL_236;
  assign _EVAL_157 = _EVAL_367 | _EVAL_289;
  assign _EVAL_226 = _EVAL_157 | _EVAL_4;
  assign _EVAL_330 = _EVAL_226 == 1'h0;
  assign _EVAL_251 = _EVAL_13 == _EVAL_261;
  assign _EVAL_282 = _EVAL_251 | _EVAL_4;
  assign _EVAL_110 = _EVAL_350 >> _EVAL_16;
  assign _EVAL_267 = _EVAL_110[0];
  assign _EVAL_292 = _EVAL_267 == 1'h0;
  assign _EVAL_281 = _EVAL_292 | _EVAL_4;
  assign _EVAL_221 = _EVAL_281 == 1'h0;
  assign _EVAL_137 = _EVAL_7 >= 4'h2;
  assign _EVAL_142 = _EVAL_137 | _EVAL_4;
  assign _EVAL_308 = _EVAL_142 == 1'h0;
  assign _EVAL_90 = _EVAL_351 & _EVAL_20;
  assign _EVAL_357 = _EVAL_6 <= 4'h6;
  assign _EVAL_349 = _EVAL_171 | _EVAL_85;
  assign _EVAL_288 = _EVAL_349 | _EVAL_145;
  assign _EVAL_317 = _EVAL_288 | _EVAL_196;
  assign _EVAL_189 = _EVAL_317 | _EVAL_34;
  assign _EVAL_98 = _EVAL_189 | _EVAL_359;
  assign _EVAL_319 = _EVAL_357 & _EVAL_98;
  assign _EVAL_126 = _EVAL_90 | _EVAL_319;
  assign _EVAL_118 = _EVAL_126 | _EVAL_4;
  assign _EVAL_210 = _EVAL_118 == 1'h0;
  assign _EVAL_155 = _EVAL_7 == _EVAL_97;
  assign _EVAL_249 = _EVAL_155 | _EVAL_4;
  assign _EVAL_144 = _EVAL_249 == 1'h0;
  assign _EVAL_306 = _EVAL_90 | _EVAL_4;
  assign _EVAL_125 = _EVAL_306 == 1'h0;
  assign _EVAL_202 = 4'h6 == _EVAL_6;
  assign _EVAL_139 = _EVAL_205 ? _EVAL_202 : 1'h0;
  assign _EVAL_322 = _EVAL_9 == _EVAL_223;
  assign _EVAL_148 = _EVAL_322 | _EVAL_4;
  assign _EVAL_339 = _EVAL_5 & _EVAL_39;
  assign _EVAL_218 = _EVAL_83 == 6'h0;
  assign _EVAL_46 = _EVAL_18 == _EVAL_31;
  assign _EVAL_243 = _EVAL_46 | _EVAL_4;
  assign _EVAL_67 = _EVAL_10 <= 3'h3;
  assign _EVAL_343 = _EVAL_67 | _EVAL_4;
  assign _EVAL_183 = _EVAL_343 == 1'h0;
  assign _EVAL_268 = _EVAL_8 == 1'h0;
  assign _EVAL_297 = _EVAL_268 | _EVAL_4;
  assign _EVAL_113 = _EVAL_0 <= 2'h2;
  assign _EVAL_284 = _EVAL_113 | _EVAL_4;
  assign _EVAL_71 = _EVAL_293 | _EVAL_299;
  assign _EVAL_338 = _EVAL_312 == 4'h2;
  assign _EVAL_25 = _EVAL_71 | _EVAL_338;
  assign _EVAL_250 = _EVAL_243 == 1'h0;
  assign _EVAL_94 = _EVAL_14 == _EVAL_355;
  assign _EVAL_130 = _EVAL_94 | _EVAL_4;
  assign _EVAL_327 = _EVAL_130 == 1'h0;
  assign _EVAL_138 = ~ _EVAL_186;
  assign _EVAL_208 = _EVAL_297 == 1'h0;
  assign _EVAL_56 = _EVAL_121 == 6'h0;
  assign _EVAL_26 = _EVAL_56 == 1'h0;
  assign _EVAL_140 = _EVAL_16[2:0];
  assign _EVAL_275 = ~ _EVAL_9;
  assign _EVAL_231 = _EVAL == _EVAL_237;
  assign _EVAL_103 = _EVAL_231 | _EVAL_4;
  assign _EVAL_329 = _EVAL_103 == 1'h0;
  assign _EVAL_215 = _EVAL_0 == _EVAL_361;
  assign _EVAL_101 = _EVAL_215 | _EVAL_4;
  assign _EVAL_194 = _EVAL_101 == 1'h0;
  assign _EVAL_102 = _EVAL_16 == 7'h20;
  assign _EVAL_207 = _EVAL_304 | _EVAL_4;
  assign _EVAL_55 = _EVAL_207 == 1'h0;
  assign _EVAL_180 = _EVAL == 3'h1;
  assign _EVAL_158 = _EVAL_5 & _EVAL_180;
  assign _EVAL_53 = _EVAL_312 == 4'h3;
  assign _EVAL_19 = _EVAL_48 == 1'h0;
  assign _EVAL_238 = 3'h1 <= _EVAL_140;
  assign _EVAL_203 = _EVAL == 3'h5;
  assign _EVAL_106 = _EVAL_16 == 7'h48;
  assign _EVAL_141 = _EVAL_106 | _EVAL_205;
  assign _EVAL_311 = _EVAL_195 & _EVAL_238;
  assign _EVAL_264 = _EVAL_141 | _EVAL_311;
  assign _EVAL_105 = _EVAL_264 | _EVAL_102;
  assign _EVAL_167 = _EVAL_1 == 3'h4;
  assign _EVAL_182 = _EVAL_174 | _EVAL_4;
  assign _EVAL_259 = _EVAL_182 == 1'h0;
  assign _EVAL_160 = _EVAL_214 + 32'h1;
  assign _EVAL_209 = _EVAL_197 | _EVAL_30;
  assign _EVAL_326 = _EVAL_30 & _EVAL_218;
  assign _EVAL_242 = _EVAL_38 | _EVAL_4;
  assign _EVAL_75 = _EVAL_242 == 1'h0;
  assign _EVAL_332 = _EVAL_6 == _EVAL_227;
  assign _EVAL_119 = _EVAL_332 | _EVAL_4;
  assign _EVAL_149 = _EVAL_10 == 3'h0;
  assign _EVAL_269 = _EVAL_149 | _EVAL_4;
  assign _EVAL_246 = _EVAL_16 == _EVAL_28;
  assign _EVAL_32 = _EVAL_246 | _EVAL_4;
  assign _EVAL_22 = _EVAL_2 == _EVAL_96;
  assign _EVAL_170 = _EVAL_22 | _EVAL_4;
  assign _EVAL_253 = _EVAL_121 - 6'h1;
  assign _EVAL_247 = _EVAL_1 == _EVAL_166;
  assign _EVAL_369 = _EVAL_1 == 3'h6;
  assign _EVAL_352 = _EVAL_12 & _EVAL_369;
  assign _EVAL_77 = _EVAL_275 == 4'h0;
  assign _EVAL_35 = _EVAL_77 | _EVAL_4;
  assign _EVAL_271 = _EVAL_35 == 1'h0;
  assign _EVAL_177 = _EVAL_119 == 1'h0;
  assign _EVAL_348 = _EVAL_241 == 1'h0;
  assign _EVAL_220 = _EVAL_170 == 1'h0;
  assign _EVAL_128 = _EVAL_139 | _EVAL_4;
  assign _EVAL_233 = _EVAL_269 == 1'h0;
  assign _EVAL_201 = _EVAL == 3'h4;
  assign _EVAL_152 = _EVAL_12 & _EVAL_26;
  assign _EVAL_257 = _EVAL_14 == 1'h0;
  assign _EVAL_124 = _EVAL_5 & _EVAL_201;
  assign _EVAL_305 = _EVAL_218 == 1'h0;
  assign _EVAL_252 = _EVAL_5 & _EVAL_305;
  assign _EVAL_88 = _EVAL_257 | _EVAL_3;
  assign _EVAL_64 = _EVAL_88 | _EVAL_4;
  assign _EVAL_234 = _EVAL_64 == 1'h0;
  assign _EVAL_122 = _EVAL_344 == 1'h0;
  assign _EVAL_51 = _EVAL_32 == 1'h0;
  assign _EVAL_54 = _EVAL_247 | _EVAL_4;
  assign _EVAL_181 = _EVAL_54 == 1'h0;
  assign _EVAL_331 = _EVAL_5 & _EVAL_222;
  assign _EVAL_132 = _EVAL_284 == 1'h0;
  assign _EVAL_301 = _EVAL_159 == 4'h0;
  assign _EVAL_298 = _EVAL_105 | _EVAL_301;
  assign _EVAL_360 = _EVAL_159 == 4'h1;
  assign _EVAL_79 = _EVAL_1 == 3'h2;
  assign _EVAL_68 = _EVAL_159 == 4'h3;
  assign _EVAL_200 = _EVAL_298 | _EVAL_360;
  assign _EVAL_283 = _EVAL_179 | _EVAL_4;
  assign _EVAL_40 = _EVAL == 3'h2;
  assign _EVAL_323 = _EVAL_5 & _EVAL_40;
  assign _EVAL_225 = _EVAL_25 | _EVAL_53;
  assign _EVAL_151 = _EVAL_83 - 6'h1;
  assign _EVAL_37 = _EVAL_225 | _EVAL_4;
  assign _EVAL_78 = _EVAL_159 == 4'h2;
  assign _EVAL_131 = _EVAL_200 | _EVAL_78;
  assign _EVAL_309 = _EVAL_131 | _EVAL_68;
  assign _EVAL_191 = _EVAL_309 | _EVAL_4;
  assign _EVAL_192 = _EVAL_191 == 1'h0;
  assign _EVAL_43 = _EVAL_49 == 1'h0;
  assign _EVAL_328 = _EVAL_282 == 1'h0;
  assign _EVAL_161 = _EVAL_128 == 1'h0;
  assign _EVAL_262 = _EVAL_3 == 1'h0;
  assign _EVAL_21 = _EVAL_148 == 1'h0;
  assign _EVAL_163 = _EVAL_4 == 1'h0;
  assign _EVAL_74 = _EVAL_262 | _EVAL_4;
  assign _EVAL_244 = _EVAL_10 != 3'h0;
  assign _EVAL_92 = _EVAL_244 | _EVAL_4;
  assign _EVAL_185 = _EVAL_283 == 1'h0;
  assign _EVAL_303 = _EVAL_1 == 3'h3;
  assign _EVAL_116 = _EVAL_12 & _EVAL_235;
  assign _EVAL_143 = _EVAL_0 != 2'h2;
  assign _EVAL_263 = _EVAL_37 == 1'h0;
  assign _EVAL_150 = _EVAL_257 | _EVAL_4;
  assign _EVAL_270 = _EVAL_197 & _EVAL_56;
  assign _EVAL_80 = _EVAL_1 == 3'h0;
  assign _EVAL_320 = _EVAL_12 & _EVAL_80;
  assign _EVAL_300 = _EVAL_104 & _EVAL_138;
  assign _EVAL_135 = _EVAL_150 == 1'h0;
  assign _EVAL_70 = _EVAL_74 == 1'h0;
  assign _EVAL_364 = _EVAL_12 & _EVAL_303;
  assign _EVAL_73 = _EVAL_92 == 1'h0;
  assign _EVAL_153 = _EVAL_12 & _EVAL_79;
  assign _EVAL_280 = _EVAL_143 | _EVAL_4;
  assign _EVAL_120 = _EVAL_280 == 1'h0;
  assign _EVAL_164 = _EVAL_5 & _EVAL_203;
  assign _EVAL_169 = _EVAL_12 & _EVAL_167;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_28 = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_31 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_83 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_96 = _RAND_3[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_97 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_121 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_166 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_212 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_214 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_227 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_237 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_261 = _RAND_11[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_276 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_324 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {3{`RANDOM}};
  _EVAL_350 = _RAND_14[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_355 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_361 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_17) begin
    if (_EVAL_270) begin
      _EVAL_28 <= _EVAL_16;
    end
    if (_EVAL_326) begin
      _EVAL_31 <= _EVAL_18;
    end
    if (_EVAL_4) begin
      _EVAL_83 <= 6'h0;
    end else begin
      if (_EVAL_30) begin
        if (_EVAL_218) begin
          if (_EVAL_254) begin
            _EVAL_83 <= _EVAL_111;
          end else begin
            _EVAL_83 <= 6'h0;
          end
        end else begin
          _EVAL_83 <= _EVAL_151;
        end
      end
    end
    if (_EVAL_270) begin
      _EVAL_96 <= _EVAL_2;
    end
    if (_EVAL_326) begin
      _EVAL_97 <= _EVAL_7;
    end
    if (_EVAL_4) begin
      _EVAL_121 <= 6'h0;
    end else begin
      if (_EVAL_197) begin
        if (_EVAL_56) begin
          if (_EVAL_228) begin
            _EVAL_121 <= _EVAL_230;
          end else begin
            _EVAL_121 <= 6'h0;
          end
        end else begin
          _EVAL_121 <= _EVAL_253;
        end
      end
    end
    if (_EVAL_270) begin
      _EVAL_166 <= _EVAL_1;
    end
    if (_EVAL_4) begin
      _EVAL_212 <= 6'h0;
    end else begin
      if (_EVAL_197) begin
        if (_EVAL_61) begin
          if (_EVAL_228) begin
            _EVAL_212 <= _EVAL_230;
          end else begin
            _EVAL_212 <= 6'h0;
          end
        end else begin
          _EVAL_212 <= _EVAL_353;
        end
      end
    end
    if (_EVAL_4) begin
      _EVAL_214 <= 32'h0;
    end else begin
      if (_EVAL_209) begin
        _EVAL_214 <= 32'h0;
      end else begin
        _EVAL_214 <= _EVAL_160;
      end
    end
    if (_EVAL_270) begin
      _EVAL_227 <= _EVAL_6;
    end
    if (_EVAL_326) begin
      _EVAL_237 <= _EVAL;
    end
    if (_EVAL_326) begin
      _EVAL_261 <= _EVAL_13;
    end
    if (_EVAL_4) begin
      _EVAL_276 <= 6'h0;
    end else begin
      if (_EVAL_30) begin
        if (_EVAL_91) begin
          if (_EVAL_254) begin
            _EVAL_276 <= _EVAL_111;
          end else begin
            _EVAL_276 <= 6'h0;
          end
        end else begin
          _EVAL_276 <= _EVAL_315;
        end
      end
    end
    if (_EVAL_270) begin
      _EVAL_324 <= _EVAL_10;
    end
    if (_EVAL_4) begin
      _EVAL_350 <= 73'h0;
    end else begin
      _EVAL_350 <= _EVAL_300;
    end
    if (_EVAL_326) begin
      _EVAL_355 <= _EVAL_14;
    end
    if (_EVAL_326) begin
      _EVAL_361 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(643d55e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dfa26bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bce2ff8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae54e9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(890de656)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c616e2f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47741d1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07ffc1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7be58c32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e565538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb55d3c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7965fc89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(867c175)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1d8d65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad2c709)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_329) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67aebff8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8cb4ce2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7447ad9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af6f28a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d50cd139)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_329) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da8f7d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3312ddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b22d240)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78d60381)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(927fdd0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e7c430b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4b5b554)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b12738c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(150d7e87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24809aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68b494f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2fb9465)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f85782b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5da0d0bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf32b12b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_328) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e4a2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e795e8e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71456eac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf1807eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(512eb12b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa3ac06a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a61a750)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbbb5865)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7b610fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7645cf76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1febabe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a9d9507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3452e9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fdb4717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c43cbd38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac1ee4e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6958b8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(756ca17b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21b96a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c515b1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10bb6f29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(283a1cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72643eb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65e82d8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8415d2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fd91bbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9826e40b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(183f172a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fc4ce6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecee6dac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33253038)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c715a32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e34e1e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61db8f48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea666531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47ddc33c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ad06dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63d28983)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(763bb36b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee86b6a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d02e2364)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1dce008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed57a4fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c11d162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1b9c822)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51b0c796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bf430c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f373e398)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ba9be45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af5cdabf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_328) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20e7ecf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5d96c8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aef6a83a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db446642)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87d75d49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
