//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_321_assert(
  input         _EVAL,
  input  [8:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [8:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [7:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input  [2:0]  _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_18;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_21;
  reg [31:0] _RAND_1;
  reg [31:0] _EVAL_27;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_36;
  reg [31:0] _RAND_3;
  reg [511:0] _EVAL_41;
  reg [511:0] _RAND_4;
  reg [2:0] _EVAL_77;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_125;
  reg [31:0] _RAND_6;
  reg [8:0] _EVAL_132;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_137;
  reg [31:0] _RAND_8;
  reg [31:0] _EVAL_168;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_181;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_196;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_214;
  reg [31:0] _RAND_12;
  reg  _EVAL_238;
  reg [31:0] _RAND_13;
  reg [8:0] _EVAL_254;
  reg [31:0] _RAND_14;
  wire  _EVAL_147;
  wire  _EVAL_249;
  wire  _EVAL_191;
  wire  _EVAL_102;
  wire  _EVAL_118;
  wire  _EVAL_68;
  wire  _EVAL_282;
  wire  _EVAL_31;
  wire [12:0] _EVAL_101;
  wire [5:0] _EVAL_54;
  wire [5:0] _EVAL_275;
  wire  _EVAL_271;
  wire  _EVAL_247;
  wire  _EVAL_151;
  wire [511:0] _EVAL_35;
  wire [511:0] _EVAL_195;
  wire [511:0] _EVAL_274;
  wire [511:0] _EVAL_146;
  wire  _EVAL_232;
  wire  _EVAL_66;
  wire  _EVAL_246;
  wire [1:0] _EVAL_60;
  wire [3:0] _EVAL_205;
  wire [2:0] _EVAL_261;
  wire [2:0] _EVAL_113;
  wire  _EVAL_23;
  wire  _EVAL_152;
  wire  _EVAL_17;
  wire  _EVAL_33;
  wire  _EVAL_257;
  wire  _EVAL_131;
  wire  _EVAL_30;
  wire  _EVAL_201;
  wire  _EVAL_115;
  wire [2:0] _EVAL_268;
  wire [2:0] _EVAL_142;
  wire  _EVAL_110;
  wire  _EVAL_78;
  wire  _EVAL_166;
  wire  _EVAL_48;
  wire  _EVAL_145;
  wire  _EVAL_126;
  wire  _EVAL_197;
  wire  _EVAL_94;
  wire  _EVAL_230;
  wire  _EVAL_141;
  wire  _EVAL_179;
  wire  _EVAL_186;
  wire  _EVAL_167;
  wire  _EVAL_262;
  wire  _EVAL_207;
  wire  _EVAL_52;
  wire [12:0] _EVAL_194;
  wire [5:0] _EVAL_228;
  wire [5:0] _EVAL_248;
  wire [2:0] _EVAL_114;
  wire [2:0] _EVAL_255;
  wire  _EVAL_171;
  wire  _EVAL_26;
  wire  _EVAL_103;
  wire  _EVAL_22;
  wire  _EVAL_51;
  wire  _EVAL_267;
  wire  _EVAL_128;
  wire  _EVAL_97;
  wire  _EVAL_25;
  wire  _EVAL_225;
  wire  _EVAL_49;
  wire  _EVAL_119;
  wire  _EVAL_34;
  wire  _EVAL_221;
  wire [31:0] _EVAL_74;
  wire [31:0] _EVAL_204;
  wire  _EVAL_192;
  wire  _EVAL_209;
  wire  _EVAL_277;
  wire  _EVAL_50;
  wire  _EVAL_169;
  wire  _EVAL_227;
  wire  _EVAL_283;
  wire  _EVAL_38;
  wire  _EVAL_135;
  wire  _EVAL_158;
  wire  _EVAL_75;
  wire  _EVAL_105;
  wire  _EVAL_29;
  wire  _EVAL_239;
  wire [31:0] _EVAL_272;
  wire [32:0] _EVAL_69;
  wire  _EVAL_140;
  wire  _EVAL_122;
  wire  _EVAL_215;
  wire  _EVAL_59;
  wire  _EVAL_258;
  wire  _EVAL_280;
  wire  _EVAL_63;
  wire [511:0] _EVAL_121;
  wire [511:0] _EVAL_70;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_202;
  wire  _EVAL_86;
  wire  _EVAL_243;
  wire  _EVAL_155;
  wire  _EVAL_20;
  wire  _EVAL_88;
  wire  _EVAL_276;
  wire  _EVAL_153;
  wire [511:0] _EVAL_189;
  wire [2:0] _EVAL_266;
  wire  _EVAL_84;
  wire  _EVAL_174;
  wire  _EVAL_165;
  wire [7:0] _EVAL_172;
  wire  _EVAL_278;
  wire  _EVAL_46;
  wire  _EVAL_129;
  wire  _EVAL_199;
  wire  _EVAL_85;
  wire  _EVAL_245;
  wire  _EVAL_111;
  wire  _EVAL_162;
  wire  _EVAL_244;
  wire  _EVAL_67;
  wire  _EVAL_154;
  wire  _EVAL_62;
  wire  _EVAL_269;
  wire [511:0] _EVAL_53;
  wire  _EVAL_133;
  wire  _EVAL_156;
  wire  _EVAL_109;
  wire  _EVAL_163;
  wire  _EVAL_90;
  wire  _EVAL_24;
  wire  _EVAL_112;
  wire  _EVAL_108;
  wire  _EVAL_58;
  wire  _EVAL_100;
  wire  _EVAL_95;
  wire  _EVAL_270;
  wire  _EVAL_253;
  wire  _EVAL_61;
  wire  _EVAL_149;
  wire  _EVAL_178;
  wire  _EVAL_216;
  wire  _EVAL_99;
  wire  _EVAL_264;
  wire  _EVAL_93;
  wire  _EVAL_182;
  wire  _EVAL_150;
  wire  _EVAL_47;
  wire  _EVAL_226;
  wire  _EVAL_252;
  wire [7:0] _EVAL_183;
  wire [7:0] _EVAL_159;
  wire [7:0] _EVAL_81;
  wire  _EVAL_213;
  wire  _EVAL_265;
  wire  _EVAL_281;
  wire  _EVAL_206;
  wire  _EVAL_208;
  wire  _EVAL_229;
  wire  _EVAL_242;
  wire  _EVAL_79;
  wire  _EVAL_42;
  wire  _EVAL_130;
  wire  _EVAL_104;
  wire  _EVAL_176;
  wire  _EVAL_148;
  wire [2:0] _EVAL_120;
  wire  _EVAL_134;
  wire  _EVAL_138;
  wire  _EVAL_76;
  wire  _EVAL_107;
  wire  _EVAL_175;
  wire  _EVAL_106;
  wire  _EVAL_116;
  wire  _EVAL_211;
  wire  _EVAL_259;
  wire  _EVAL_87;
  wire  _EVAL_44;
  wire  _EVAL_223;
  wire  _EVAL_263;
  wire  _EVAL_37;
  wire  _EVAL_184;
  wire  _EVAL_117;
  wire [32:0] _EVAL_273;
  wire [31:0] _EVAL_73;
  wire  _EVAL_161;
  wire  _EVAL_203;
  wire  _EVAL_32;
  wire [32:0] _EVAL_218;
  wire  _EVAL_256;
  wire  _EVAL_89;
  wire  _EVAL_157;
  wire  _EVAL_40;
  wire  _EVAL_80;
  wire  _EVAL_210;
  wire  _EVAL_173;
  wire  _EVAL_98;
  wire  _EVAL_188;
  wire  _EVAL_164;
  wire  _EVAL_279;
  wire  _EVAL_19;
  wire  _EVAL_224;
  wire [511:0] _EVAL_198;
  wire  _EVAL_143;
  wire  _EVAL_136;
  wire  _EVAL_144;
  wire  _EVAL_233;
  wire  _EVAL_219;
  wire  _EVAL_187;
  wire  _EVAL_92;
  wire  _EVAL_139;
  wire  _EVAL_260;
  wire  _EVAL_193;
  wire  _EVAL_212;
  wire  _EVAL_170;
  wire  _EVAL_45;
  wire  _EVAL_222;
  wire  _EVAL_123;
  wire  _EVAL_217;
  wire  _EVAL_65;
  wire  _EVAL_185;
  wire  _EVAL_231;
  wire  _EVAL_56;
  wire  _EVAL_39;
  wire  _EVAL_43;
  wire  _EVAL_28;
  wire  _EVAL_236;
  wire  _EVAL_64;
  wire  _EVAL_160;
  wire  _EVAL_72;
  wire [511:0] _EVAL_220;
  wire  _EVAL_241;
  wire  _EVAL_91;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_147 = _EVAL_12[2];
  assign _EVAL_249 = _EVAL_12[1];
  assign _EVAL_191 = _EVAL_147 & _EVAL_249;
  assign _EVAL_102 = _EVAL_12[0];
  assign _EVAL_118 = _EVAL_102 == 1'h0;
  assign _EVAL_68 = _EVAL_191 & _EVAL_118;
  assign _EVAL_282 = _EVAL_15 == 1'h0;
  assign _EVAL_31 = _EVAL_12 == _EVAL_27;
  assign _EVAL_101 = 13'h3f << _EVAL_7;
  assign _EVAL_54 = _EVAL_101[5:0];
  assign _EVAL_275 = ~ _EVAL_54;
  assign _EVAL_271 = _EVAL_9 & _EVAL_5;
  assign _EVAL_247 = _EVAL_77 == 3'h0;
  assign _EVAL_151 = _EVAL_271 & _EVAL_247;
  assign _EVAL_35 = 512'h1 << _EVAL_0;
  assign _EVAL_195 = _EVAL_151 ? _EVAL_35 : 512'h0;
  assign _EVAL_274 = _EVAL_195 | _EVAL_41;
  assign _EVAL_146 = _EVAL_274 >> _EVAL_8;
  assign _EVAL_232 = _EVAL_146[0];
  assign _EVAL_66 = _EVAL_232 | _EVAL_15;
  assign _EVAL_246 = _EVAL_66 == 1'h0;
  assign _EVAL_60 = _EVAL_7[1:0];
  assign _EVAL_205 = 4'h1 << _EVAL_60;
  assign _EVAL_261 = _EVAL_205[2:0];
  assign _EVAL_113 = _EVAL_261 | 3'h1;
  assign _EVAL_23 = _EVAL_113[0];
  assign _EVAL_152 = _EVAL_147 == 1'h0;
  assign _EVAL_17 = _EVAL_152 & _EVAL_249;
  assign _EVAL_33 = _EVAL_17 & _EVAL_118;
  assign _EVAL_257 = _EVAL_23 & _EVAL_33;
  assign _EVAL_131 = _EVAL_0 == _EVAL_132;
  assign _EVAL_30 = _EVAL_131 | _EVAL_15;
  assign _EVAL_201 = _EVAL_11[2];
  assign _EVAL_115 = _EVAL_201 == 1'h0;
  assign _EVAL_268 = _EVAL_275[5:3];
  assign _EVAL_142 = _EVAL_196 - 3'h1;
  assign _EVAL_110 = _EVAL_7 <= 3'h6;
  assign _EVAL_78 = _EVAL_7 >= 3'h3;
  assign _EVAL_166 = _EVAL_113[2];
  assign _EVAL_48 = _EVAL_166 & _EVAL_147;
  assign _EVAL_145 = _EVAL_78 | _EVAL_48;
  assign _EVAL_126 = _EVAL_113[1];
  assign _EVAL_197 = _EVAL_249 == 1'h0;
  assign _EVAL_94 = _EVAL_147 & _EVAL_197;
  assign _EVAL_230 = _EVAL_126 & _EVAL_94;
  assign _EVAL_141 = _EVAL_145 | _EVAL_230;
  assign _EVAL_179 = _EVAL_94 & _EVAL_102;
  assign _EVAL_186 = _EVAL_23 & _EVAL_179;
  assign _EVAL_167 = _EVAL_141 | _EVAL_186;
  assign _EVAL_262 = _EVAL_1 & _EVAL_10;
  assign _EVAL_207 = _EVAL_137 == 3'h0;
  assign _EVAL_52 = _EVAL_4[0];
  assign _EVAL_194 = 13'h3f << _EVAL_16;
  assign _EVAL_228 = _EVAL_194[5:0];
  assign _EVAL_248 = ~ _EVAL_228;
  assign _EVAL_114 = _EVAL_248[5:3];
  assign _EVAL_255 = _EVAL_137 - 3'h1;
  assign _EVAL_171 = _EVAL_11 == 3'h7;
  assign _EVAL_26 = _EVAL_5 & _EVAL_171;
  assign _EVAL_103 = _EVAL_16 >= 3'h3;
  assign _EVAL_22 = _EVAL_103 | _EVAL_15;
  assign _EVAL_51 = _EVAL_22 == 1'h0;
  assign _EVAL_267 = _EVAL == 1'h0;
  assign _EVAL_128 = _EVAL_267 | _EVAL_15;
  assign _EVAL_97 = _EVAL_128 == 1'h0;
  assign _EVAL_25 = _EVAL_271 | _EVAL_262;
  assign _EVAL_225 = _EVAL_126 & _EVAL_191;
  assign _EVAL_49 = _EVAL_145 | _EVAL_225;
  assign _EVAL_119 = _EVAL_191 & _EVAL_102;
  assign _EVAL_34 = _EVAL_23 & _EVAL_119;
  assign _EVAL_221 = _EVAL_49 | _EVAL_34;
  assign _EVAL_74 = {{26'd0}, _EVAL_275};
  assign _EVAL_204 = _EVAL_12 & _EVAL_74;
  assign _EVAL_192 = _EVAL_204 == 32'h0;
  assign _EVAL_209 = _EVAL_192 | _EVAL_15;
  assign _EVAL_277 = _EVAL_209 == 1'h0;
  assign _EVAL_50 = _EVAL_8 == _EVAL_254;
  assign _EVAL_169 = _EVAL_50 | _EVAL_15;
  assign _EVAL_227 = _EVAL_14 == 3'h0;
  assign _EVAL_283 = _EVAL_227 | _EVAL_15;
  assign _EVAL_38 = _EVAL_41 != 512'h0;
  assign _EVAL_135 = _EVAL_38 == 1'h0;
  assign _EVAL_158 = plusarg_reader_out == 32'h0;
  assign _EVAL_75 = _EVAL_135 | _EVAL_158;
  assign _EVAL_105 = _EVAL_168 < plusarg_reader_out;
  assign _EVAL_29 = _EVAL_75 | _EVAL_105;
  assign _EVAL_239 = _EVAL_29 | _EVAL_15;
  assign _EVAL_272 = _EVAL_12 ^ 32'h80000000;
  assign _EVAL_69 = {1'b0,$signed(_EVAL_272)};
  assign _EVAL_140 = _EVAL_14 <= 3'h4;
  assign _EVAL_122 = _EVAL_140 | _EVAL_15;
  assign _EVAL_215 = _EVAL_122 == 1'h0;
  assign _EVAL_59 = _EVAL_262 & _EVAL_207;
  assign _EVAL_258 = _EVAL_4 == 3'h6;
  assign _EVAL_280 = _EVAL_258 == 1'h0;
  assign _EVAL_63 = _EVAL_59 & _EVAL_280;
  assign _EVAL_121 = 512'h1 << _EVAL_8;
  assign _EVAL_70 = _EVAL_63 ? _EVAL_121 : 512'h0;
  assign _EVAL_82 = _EVAL_195 != _EVAL_70;
  assign _EVAL_83 = _EVAL_195 != 512'h0;
  assign _EVAL_202 = _EVAL_83 == 1'h0;
  assign _EVAL_86 = _EVAL_82 | _EVAL_202;
  assign _EVAL_243 = _EVAL_86 | _EVAL_15;
  assign _EVAL_155 = _EVAL_243 == 1'h0;
  assign _EVAL_20 = _EVAL_31 | _EVAL_15;
  assign _EVAL_88 = _EVAL_6 == 1'h0;
  assign _EVAL_276 = _EVAL_11 == 3'h1;
  assign _EVAL_153 = _EVAL_5 & _EVAL_276;
  assign _EVAL_189 = ~ _EVAL_70;
  assign _EVAL_266 = _EVAL_77 - 3'h1;
  assign _EVAL_84 = _EVAL_14 != 3'h0;
  assign _EVAL_174 = _EVAL_84 | _EVAL_15;
  assign _EVAL_165 = _EVAL_174 == 1'h0;
  assign _EVAL_172 = ~ _EVAL_13;
  assign _EVAL_278 = _EVAL_16 == _EVAL_181;
  assign _EVAL_46 = _EVAL_278 | _EVAL_15;
  assign _EVAL_129 = _EVAL_11 == _EVAL_21;
  assign _EVAL_199 = _EVAL_129 | _EVAL_15;
  assign _EVAL_85 = _EVAL_199 == 1'h0;
  assign _EVAL_245 = _EVAL_11 == 3'h2;
  assign _EVAL_111 = _EVAL_5 & _EVAL_245;
  assign _EVAL_162 = _EVAL_4 <= 3'h6;
  assign _EVAL_244 = _EVAL_166 & _EVAL_152;
  assign _EVAL_67 = _EVAL_78 | _EVAL_244;
  assign _EVAL_154 = _EVAL_126 & _EVAL_17;
  assign _EVAL_62 = _EVAL_67 | _EVAL_154;
  assign _EVAL_269 = _EVAL_62 | _EVAL_257;
  assign _EVAL_53 = _EVAL_41 >> _EVAL_0;
  assign _EVAL_133 = _EVAL_53[0];
  assign _EVAL_156 = _EVAL_133 == 1'h0;
  assign _EVAL_109 = _EVAL_156 | _EVAL_15;
  assign _EVAL_163 = _EVAL_109 == 1'h0;
  assign _EVAL_90 = _EVAL_17 & _EVAL_102;
  assign _EVAL_24 = _EVAL_14 == _EVAL_214;
  assign _EVAL_112 = _EVAL_24 | _EVAL_15;
  assign _EVAL_108 = _EVAL_7 == _EVAL_125;
  assign _EVAL_58 = _EVAL_162 | _EVAL_15;
  assign _EVAL_100 = _EVAL_23 & _EVAL_68;
  assign _EVAL_95 = _EVAL_49 | _EVAL_100;
  assign _EVAL_270 = _EVAL_94 & _EVAL_118;
  assign _EVAL_253 = _EVAL_23 & _EVAL_270;
  assign _EVAL_61 = _EVAL_141 | _EVAL_253;
  assign _EVAL_149 = _EVAL_23 & _EVAL_90;
  assign _EVAL_178 = _EVAL_62 | _EVAL_149;
  assign _EVAL_216 = _EVAL_152 & _EVAL_197;
  assign _EVAL_99 = _EVAL_126 & _EVAL_216;
  assign _EVAL_264 = _EVAL_67 | _EVAL_99;
  assign _EVAL_93 = _EVAL_216 & _EVAL_102;
  assign _EVAL_182 = _EVAL_23 & _EVAL_93;
  assign _EVAL_150 = _EVAL_264 | _EVAL_182;
  assign _EVAL_47 = _EVAL_216 & _EVAL_118;
  assign _EVAL_226 = _EVAL_23 & _EVAL_47;
  assign _EVAL_252 = _EVAL_264 | _EVAL_226;
  assign _EVAL_183 = {_EVAL_221,_EVAL_95,_EVAL_167,_EVAL_61,_EVAL_178,_EVAL_269,_EVAL_150,_EVAL_252};
  assign _EVAL_159 = ~ _EVAL_183;
  assign _EVAL_81 = _EVAL_13 & _EVAL_159;
  assign _EVAL_213 = _EVAL_11 == 3'h6;
  assign _EVAL_265 = _EVAL_11 == 3'h4;
  assign _EVAL_281 = _EVAL_5 & _EVAL_265;
  assign _EVAL_206 = _EVAL_4 == 3'h2;
  assign _EVAL_208 = _EVAL_10 & _EVAL_206;
  assign _EVAL_229 = _EVAL_4 == 3'h5;
  assign _EVAL_242 = _EVAL_10 & _EVAL_229;
  assign _EVAL_79 = _EVAL_4 == _EVAL_36;
  assign _EVAL_42 = _EVAL_79 | _EVAL_15;
  assign _EVAL_130 = _EVAL_42 == 1'h0;
  assign _EVAL_104 = _EVAL_14 <= 3'h3;
  assign _EVAL_176 = _EVAL_104 | _EVAL_15;
  assign _EVAL_148 = _EVAL_18 == 3'h0;
  assign _EVAL_120 = _EVAL_18 - 3'h1;
  assign _EVAL_134 = _EVAL_148 == 1'h0;
  assign _EVAL_138 = _EVAL_196 == 3'h0;
  assign _EVAL_76 = _EVAL == _EVAL_238;
  assign _EVAL_107 = _EVAL_30 == 1'h0;
  assign _EVAL_175 = _EVAL_11 == 3'h5;
  assign _EVAL_106 = _EVAL_5 & _EVAL_175;
  assign _EVAL_116 = _EVAL_239 == 1'h0;
  assign _EVAL_211 = _EVAL_4 == 3'h4;
  assign _EVAL_259 = _EVAL_10 & _EVAL_211;
  assign _EVAL_87 = _EVAL_88 | _EVAL_15;
  assign _EVAL_44 = _EVAL_87 == 1'h0;
  assign _EVAL_223 = _EVAL_176 == 1'h0;
  assign _EVAL_263 = _EVAL_10 & _EVAL_134;
  assign _EVAL_37 = _EVAL_13 == _EVAL_183;
  assign _EVAL_184 = _EVAL_37 | _EVAL_15;
  assign _EVAL_117 = _EVAL_184 == 1'h0;
  assign _EVAL_273 = $signed(_EVAL_69) & $signed(-33'sh20000);
  assign _EVAL_73 = _EVAL_168 + 32'h1;
  assign _EVAL_161 = _EVAL_4 == 3'h1;
  assign _EVAL_203 = _EVAL_78 | _EVAL_15;
  assign _EVAL_32 = _EVAL_203 == 1'h0;
  assign _EVAL_218 = $signed(_EVAL_273);
  assign _EVAL_256 = _EVAL_11 == 3'h3;
  assign _EVAL_89 = _EVAL_5 & _EVAL_256;
  assign _EVAL_157 = _EVAL_46 == 1'h0;
  assign _EVAL_40 = _EVAL_172 == 8'h0;
  assign _EVAL_80 = _EVAL_40 | _EVAL_15;
  assign _EVAL_210 = _EVAL_112 == 1'h0;
  assign _EVAL_173 = _EVAL_4 == 3'h0;
  assign _EVAL_98 = _EVAL_10 & _EVAL_173;
  assign _EVAL_188 = _EVAL_20 == 1'h0;
  assign _EVAL_164 = $signed(_EVAL_218) == $signed(33'sh0);
  assign _EVAL_279 = _EVAL_138 == 1'h0;
  assign _EVAL_19 = _EVAL_5 & _EVAL_279;
  assign _EVAL_224 = _EVAL_76 | _EVAL_15;
  assign _EVAL_198 = _EVAL_41 | _EVAL_195;
  assign _EVAL_143 = _EVAL_14 <= 3'h2;
  assign _EVAL_136 = _EVAL_143 | _EVAL_15;
  assign _EVAL_144 = _EVAL_108 | _EVAL_15;
  assign _EVAL_233 = _EVAL_144 == 1'h0;
  assign _EVAL_219 = _EVAL_224 == 1'h0;
  assign _EVAL_187 = _EVAL_169 == 1'h0;
  assign _EVAL_92 = _EVAL_10 & _EVAL_258;
  assign _EVAL_139 = _EVAL_10 & _EVAL_161;
  assign _EVAL_260 = _EVAL_110 & _EVAL_164;
  assign _EVAL_193 = _EVAL_260 | _EVAL_15;
  assign _EVAL_212 = _EVAL_193 == 1'h0;
  assign _EVAL_170 = _EVAL_262 & _EVAL_148;
  assign _EVAL_45 = _EVAL_80 == 1'h0;
  assign _EVAL_222 = _EVAL_3 == 1'h0;
  assign _EVAL_123 = _EVAL_222 | _EVAL_15;
  assign _EVAL_217 = _EVAL_11 == 3'h0;
  assign _EVAL_65 = _EVAL_81 == 8'h0;
  assign _EVAL_185 = _EVAL_267 | _EVAL_6;
  assign _EVAL_231 = _EVAL_185 | _EVAL_15;
  assign _EVAL_56 = _EVAL_231 == 1'h0;
  assign _EVAL_39 = _EVAL_65 | _EVAL_15;
  assign _EVAL_43 = _EVAL_271 & _EVAL_138;
  assign _EVAL_28 = _EVAL_283 == 1'h0;
  assign _EVAL_236 = _EVAL_136 == 1'h0;
  assign _EVAL_64 = _EVAL_5 & _EVAL_213;
  assign _EVAL_160 = _EVAL_123 == 1'h0;
  assign _EVAL_72 = _EVAL_58 == 1'h0;
  assign _EVAL_220 = _EVAL_198 & _EVAL_189;
  assign _EVAL_241 = _EVAL_39 == 1'h0;
  assign _EVAL_91 = _EVAL_5 & _EVAL_217;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_18 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_21 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_27 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_36 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {16{`RANDOM}};
  _EVAL_41 = _RAND_4[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_77 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_125 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_132 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_137 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_168 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_181 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_196 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_214 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_238 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_254 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_15) begin
      _EVAL_18 <= 3'h0;
    end else begin
      if (_EVAL_262) begin
        if (_EVAL_148) begin
          if (_EVAL_52) begin
            _EVAL_18 <= _EVAL_114;
          end else begin
            _EVAL_18 <= 3'h0;
          end
        end else begin
          _EVAL_18 <= _EVAL_120;
        end
      end
    end
    if (_EVAL_43) begin
      _EVAL_21 <= _EVAL_11;
    end
    if (_EVAL_43) begin
      _EVAL_27 <= _EVAL_12;
    end
    if (_EVAL_170) begin
      _EVAL_36 <= _EVAL_4;
    end
    if (_EVAL_15) begin
      _EVAL_41 <= 512'h0;
    end else begin
      _EVAL_41 <= _EVAL_220;
    end
    if (_EVAL_15) begin
      _EVAL_77 <= 3'h0;
    end else begin
      if (_EVAL_271) begin
        if (_EVAL_247) begin
          if (_EVAL_115) begin
            _EVAL_77 <= _EVAL_268;
          end else begin
            _EVAL_77 <= 3'h0;
          end
        end else begin
          _EVAL_77 <= _EVAL_266;
        end
      end
    end
    if (_EVAL_43) begin
      _EVAL_125 <= _EVAL_7;
    end
    if (_EVAL_43) begin
      _EVAL_132 <= _EVAL_0;
    end
    if (_EVAL_15) begin
      _EVAL_137 <= 3'h0;
    end else begin
      if (_EVAL_262) begin
        if (_EVAL_207) begin
          if (_EVAL_52) begin
            _EVAL_137 <= _EVAL_114;
          end else begin
            _EVAL_137 <= 3'h0;
          end
        end else begin
          _EVAL_137 <= _EVAL_255;
        end
      end
    end
    if (_EVAL_15) begin
      _EVAL_168 <= 32'h0;
    end else begin
      if (_EVAL_25) begin
        _EVAL_168 <= 32'h0;
      end else begin
        _EVAL_168 <= _EVAL_73;
      end
    end
    if (_EVAL_170) begin
      _EVAL_181 <= _EVAL_16;
    end
    if (_EVAL_15) begin
      _EVAL_196 <= 3'h0;
    end else begin
      if (_EVAL_271) begin
        if (_EVAL_138) begin
          if (_EVAL_115) begin
            _EVAL_196 <= _EVAL_268;
          end else begin
            _EVAL_196 <= 3'h0;
          end
        end else begin
          _EVAL_196 <= _EVAL_142;
        end
      end
    end
    if (_EVAL_43) begin
      _EVAL_214 <= _EVAL_14;
    end
    if (_EVAL_170) begin
      _EVAL_238 <= _EVAL;
    end
    if (_EVAL_170) begin
      _EVAL_254 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f16d540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a96e1d08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90b28326)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64236761)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a132d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87845dc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28b22f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bdf4fab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff30e175)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed1b55cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e4b8b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f81d250f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f559c1b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5132ea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddec9de9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(786fdfdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48bb6716)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c81592c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d4078f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(548ef7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d28e5eaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa3768fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2026dc3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68d97eee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2c0bc61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689a3d34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c866367)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f091508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae376215)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d7666ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71299d9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38f900b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0a08f5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd3ef60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac6784c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aae4385)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aac74ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ac40fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9150265)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf01dc45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d5f8097)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6102b6fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4b85ed6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4807d36d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9803924c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c7d4f03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(144080fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f7d54e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32433cc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d9da04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13e49e14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd69eb2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c5cbb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c164de9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73733854)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(573516fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7865003)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff46aee6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f149e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f546e9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ce0a395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b1356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70df6c84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b98a1f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38d577e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fed13bc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
