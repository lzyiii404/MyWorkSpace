//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_116(
  output [27:0] _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [6:0]  _EVAL_5,
  output [3:0]  _EVAL_6,
  output        _EVAL_7,
  output [2:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [29:0] _EVAL_10,
  input  [2:0]  _EVAL_11,
  output [3:0]  _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input  [6:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  input  [6:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  input  [2:0]  _EVAL_22,
  output [13:0] _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output [6:0]  _EVAL_26,
  input  [2:0]  _EVAL_27,
  output [2:0]  _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  output [2:0]  _EVAL_32,
  input         _EVAL_33,
  output [3:0]  _EVAL_34,
  output [6:0]  _EVAL_35,
  output [6:0]  _EVAL_36,
  output        _EVAL_37,
  output [29:0] _EVAL_38,
  output        _EVAL_39,
  input  [31:0] _EVAL_40,
  output        _EVAL_41,
  output [2:0]  _EVAL_42,
  output [2:0]  _EVAL_43,
  input  [31:0] _EVAL_44,
  input         _EVAL_45,
  input  [6:0]  _EVAL_46,
  output [2:0]  _EVAL_47,
  input  [6:0]  _EVAL_48,
  input         _EVAL_49,
  output [6:0]  _EVAL_50,
  output [2:0]  _EVAL_51,
  input  [31:0] _EVAL_52,
  input  [6:0]  _EVAL_53,
  output [6:0]  _EVAL_54,
  output [14:0] _EVAL_55,
  input  [3:0]  _EVAL_56,
  output        _EVAL_57,
  input  [2:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  output [2:0]  _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  output [31:0] _EVAL_65,
  input         _EVAL_66,
  output        _EVAL_67,
  output [3:0]  _EVAL_68,
  output [3:0]  _EVAL_69,
  input         _EVAL_70,
  output [3:0]  _EVAL_71,
  input         _EVAL_72,
  input         _EVAL_73,
  output [31:0] _EVAL_74,
  input  [6:0]  _EVAL_75,
  input         _EVAL_76,
  input         _EVAL_77,
  output        _EVAL_78,
  output        _EVAL_79,
  output        _EVAL_80,
  input  [31:0] _EVAL_81,
  input         _EVAL_82,
  output [24:0] _EVAL_83,
  input         _EVAL_84,
  output [2:0]  _EVAL_85,
  output [6:0]  _EVAL_86,
  output        _EVAL_87,
  output        _EVAL_88,
  output [1:0]  _EVAL_89,
  output [6:0]  _EVAL_90,
  input  [2:0]  _EVAL_91,
  input         _EVAL_92,
  output [31:0] _EVAL_93,
  output [3:0]  _EVAL_94,
  output [2:0]  _EVAL_95,
  input  [31:0] _EVAL_96,
  output        _EVAL_97,
  output [25:0] _EVAL_98,
  output [3:0]  _EVAL_99,
  output        _EVAL_100,
  input         _EVAL_101,
  input  [2:0]  _EVAL_102,
  output        _EVAL_103,
  output [2:0]  _EVAL_104,
  output [2:0]  _EVAL_105,
  input  [31:0] _EVAL_106,
  input  [2:0]  _EVAL_107,
  input  [6:0]  _EVAL_108,
  output        _EVAL_109,
  output [31:0] _EVAL_110,
  output [2:0]  _EVAL_111,
  output        _EVAL_112,
  input  [3:0]  _EVAL_113,
  output [6:0]  _EVAL_114,
  output [11:0] _EVAL_115,
  input  [2:0]  _EVAL_116,
  output [2:0]  _EVAL_117,
  output        _EVAL_118,
  output [31:0] _EVAL_119,
  output [31:0] _EVAL_120,
  input  [2:0]  _EVAL_121,
  output        _EVAL_122,
  input         _EVAL_123,
  output        _EVAL_124,
  output [2:0]  _EVAL_125,
  output [2:0]  _EVAL_126,
  input  [3:0]  _EVAL_127,
  input         _EVAL_128,
  input         _EVAL_129,
  output        _EVAL_130,
  output        _EVAL_131,
  input  [1:0]  _EVAL_132,
  input  [2:0]  _EVAL_133,
  output        _EVAL_134,
  input  [1:0]  _EVAL_135,
  output [2:0]  _EVAL_136,
  output        _EVAL_137,
  input  [31:0] _EVAL_138,
  input  [2:0]  _EVAL_139,
  output [31:0] _EVAL_140,
  output [2:0]  _EVAL_141
);
  reg  _EVAL_164;
  reg [31:0] _RAND_0;
  reg  _EVAL_206;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_208;
  reg [31:0] _RAND_2;
  reg  _EVAL_212;
  reg [31:0] _RAND_3;
  reg  _EVAL_215;
  reg [31:0] _RAND_4;
  reg  _EVAL_223;
  reg [31:0] _RAND_5;
  reg  _EVAL_255;
  reg [31:0] _RAND_6;
  reg [6:0] _EVAL_393;
  reg [31:0] _RAND_7;
  reg  _EVAL_397;
  reg [31:0] _RAND_8;
  wire [3:0] _EVAL_229;
  wire [20:0] _EVAL_170;
  wire  _EVAL_360;
  wire [22:0] _EVAL_381;
  wire [7:0] _EVAL_155;
  wire [7:0] _EVAL_288;
  wire [5:0] _EVAL_227;
  wire [5:0] _EVAL_260;
  wire  _EVAL_376;
  wire  _EVAL_327;
  wire  _EVAL_326;
  wire [6:0] _EVAL_168;
  wire [6:0] _EVAL_299;
  wire [6:0] _EVAL_400;
  wire [13:0] _EVAL_317;
  wire [12:0] _EVAL_345;
  wire [13:0] _EVAL_281;
  wire [13:0] _EVAL_366;
  wire [11:0] _EVAL_211;
  wire [13:0] _EVAL_198;
  wire [13:0] _EVAL_339;
  wire [9:0] _EVAL_188;
  wire [13:0] _EVAL_395;
  wire [13:0] _EVAL_246;
  wire [12:0] _EVAL_307;
  wire [13:0] _EVAL_262;
  wire [13:0] _EVAL_216;
  wire [13:0] _EVAL_279;
  wire [6:0] _EVAL_259;
  wire [6:0] _EVAL_399;
  wire [6:0] _EVAL_404;
  wire [6:0] _EVAL_294;
  wire  _EVAL_391;
  wire  _EVAL_148;
  wire  _EVAL_387;
  wire [3:0] _EVAL_238;
  wire [20:0] _EVAL_258;
  wire [5:0] _EVAL_414;
  wire [5:0] _EVAL_403;
  wire [3:0] _EVAL_213;
  wire [3:0] _EVAL_250;
  wire [3:0] _EVAL_343;
  wire  _EVAL_225;
  wire [29:0] _EVAL_312;
  wire [30:0] _EVAL_396;
  wire [30:0] _EVAL_243;
  wire [30:0] _EVAL_382;
  wire  _EVAL_301;
  wire  _EVAL_325;
  wire  _EVAL_410;
  wire  _EVAL_207;
  wire  _EVAL_291;
  wire [50:0] _EVAL_192;
  wire [50:0] _EVAL_334;
  wire  _EVAL_329;
  wire  _EVAL_222;
  wire  _EVAL_210;
  wire [3:0] _EVAL_364;
  wire [50:0] _EVAL_303;
  wire [50:0] _EVAL_333;
  wire [50:0] _EVAL_146;
  wire  _EVAL_142;
  wire [50:0] _EVAL_315;
  wire [50:0] _EVAL_306;
  wire [50:0] _EVAL_244;
  wire [6:0] _EVAL_354;
  wire [7:0] _EVAL_236;
  wire [6:0] _EVAL_268;
  wire [6:0] _EVAL_295;
  wire [8:0] _EVAL_256;
  wire [6:0] _EVAL_272;
  wire [6:0] _EVAL_271;
  wire [10:0] _EVAL_214;
  wire [6:0] _EVAL_277;
  wire [6:0] _EVAL_324;
  wire [29:0] _EVAL_199;
  wire [30:0] _EVAL_349;
  wire [30:0] _EVAL_251;
  wire [30:0] _EVAL_356;
  wire  _EVAL_261;
  wire  _EVAL_341;
  wire  _EVAL_323;
  wire [50:0] _EVAL_378;
  wire [50:0] _EVAL_302;
  wire [3:0] _EVAL_369;
  wire [20:0] _EVAL_195;
  wire [5:0] _EVAL_413;
  wire  _EVAL_145;
  wire [20:0] _EVAL_372;
  wire [5:0] _EVAL_411;
  wire [5:0] _EVAL_300;
  wire [3:0] _EVAL_247;
  wire [3:0] _EVAL_157;
  wire [3:0] _EVAL_293;
  wire [5:0] _EVAL_330;
  wire [5:0] _EVAL_384;
  wire [5:0] _EVAL_167;
  wire [5:0] _EVAL_196;
  wire  _EVAL_314;
  wire  _EVAL_270;
  wire  _EVAL_388;
  wire [5:0] _EVAL_368;
  wire [5:0] _EVAL_209;
  wire [3:0] _EVAL_316;
  wire [3:0] _EVAL_370;
  wire [3:0] _EVAL_178;
  wire [5:0] _EVAL_313;
  wire [5:0] _EVAL_161;
  wire  _EVAL_239;
  wire [5:0] _EVAL_180;
  wire [5:0] _EVAL_350;
  wire [3:0] _EVAL_389;
  wire [3:0] _EVAL_169;
  wire [3:0] _EVAL_171;
  wire [5:0] _EVAL_228;
  wire [5:0] _EVAL_187;
  wire  _EVAL_336;
  wire  _EVAL_275;
  wire  _EVAL_357;
  wire [3:0] _EVAL_308;
  wire [20:0] _EVAL_221;
  wire [5:0] _EVAL_398;
  wire [5:0] _EVAL_402;
  wire [3:0] _EVAL_347;
  wire [3:0] _EVAL_184;
  wire [3:0] _EVAL_355;
  wire [5:0] _EVAL_367;
  wire [5:0] _EVAL_264;
  wire  _EVAL_286;
  wire  _EVAL_310;
  wire  _EVAL_280;
  wire [3:0] _EVAL_278;
  wire [20:0] _EVAL_346;
  wire [5:0] _EVAL_219;
  wire [5:0] _EVAL_408;
  wire [3:0] _EVAL_149;
  wire [3:0] _EVAL_379;
  wire [3:0] _EVAL_153;
  wire [5:0] _EVAL_183;
  wire [5:0] _EVAL_189;
  wire [29:0] _EVAL_371;
  wire [30:0] _EVAL_220;
  wire [30:0] _EVAL_224;
  wire [30:0] _EVAL_390;
  wire  _EVAL_337;
  wire  _EVAL_181;
  wire  _EVAL_363;
  wire  _EVAL_186;
  wire  _EVAL_297;
  wire  _EVAL_309;
  wire  _EVAL_358;
  wire  _EVAL_394;
  wire  _EVAL_385;
  wire  _EVAL_159;
  wire [30:0] _EVAL_266;
  wire [30:0] _EVAL_165;
  wire  _EVAL_298;
  wire  _EVAL_267;
  wire  _EVAL_254;
  wire [29:0] _EVAL_252;
  wire [30:0] _EVAL_377;
  wire [30:0] _EVAL_375;
  wire [30:0] _EVAL_241;
  wire [30:0] _EVAL_194;
  wire [30:0] _EVAL_151;
  wire [30:0] _EVAL_190;
  wire  _EVAL_318;
  wire [29:0] _EVAL_147;
  wire  _EVAL_202;
  wire [50:0] _EVAL_292;
  wire [50:0] _EVAL_328;
  wire [50:0] _EVAL_248;
  wire [50:0] _EVAL_175;
  wire  _EVAL_365;
  wire [50:0] _EVAL_380;
  wire [50:0] _EVAL_409;
  wire [50:0] _EVAL_234;
  wire  _EVAL_332;
  wire [50:0] _EVAL_290;
  wire [50:0] _EVAL_179;
  wire [50:0] _EVAL_322;
  wire  _EVAL_320;
  wire [29:0] _EVAL_353;
  wire [30:0] _EVAL_348;
  wire [30:0] _EVAL_163;
  wire [30:0] _EVAL_374;
  wire  _EVAL_158;
  wire  _EVAL_200;
  wire  _EVAL_284;
  wire  _EVAL_257;
  wire  _EVAL_177;
  wire  _EVAL_331;
  wire  _EVAL_182;
  wire  _EVAL_185;
  wire [30:0] _EVAL_150;
  wire [30:0] _EVAL_245;
  wire [30:0] _EVAL_152;
  wire  _EVAL_304;
  wire  _EVAL_237;
  wire  _EVAL_412;
  wire  _EVAL_249;
  wire  _EVAL_173;
  wire  _EVAL_265;
  wire  _EVAL_154;
  wire  _EVAL_406;
  wire  _EVAL_230;
  wire  _EVAL_263;
  wire  _EVAL_218;
  wire  _EVAL_401;
  wire  _EVAL_166;
  wire  _EVAL_340;
  wire  _EVAL_296;
  wire [5:0] _EVAL_335;
  wire [5:0] _EVAL_233;
  wire  _EVAL_285;
  wire  _EVAL_351;
  wire  _EVAL_203;
  wire  _EVAL_226;
  wire  _EVAL_283;
  wire  _EVAL_311;
  wire  _EVAL_217;
  wire  _EVAL_305;
  wire  _EVAL_160;
  assign _EVAL_229 = {{1'd0}, _EVAL_27};
  assign _EVAL_170 = 21'h3f << _EVAL_229;
  assign _EVAL_360 = _EVAL_19[0];
  assign _EVAL_381 = 23'hff << _EVAL_56;
  assign _EVAL_155 = _EVAL_381[7:0];
  assign _EVAL_288 = ~ _EVAL_155;
  assign _EVAL_227 = _EVAL_288[7:2];
  assign _EVAL_260 = _EVAL_360 ? _EVAL_227 : 6'h0;
  assign _EVAL_376 = _EVAL_215 ? _EVAL_128 : 1'h0;
  assign _EVAL_327 = _EVAL_397 ? _EVAL_3 : 1'h0;
  assign _EVAL_326 = _EVAL_376 | _EVAL_327;
  assign _EVAL_168 = {_EVAL_63,_EVAL_70,_EVAL_31,_EVAL_101,_EVAL_17,_EVAL_3,_EVAL_128};
  assign _EVAL_299 = ~ _EVAL_393;
  assign _EVAL_400 = _EVAL_168 & _EVAL_299;
  assign _EVAL_317 = {_EVAL_400,_EVAL_63,_EVAL_70,_EVAL_31,_EVAL_101,_EVAL_17,_EVAL_3,_EVAL_128};
  assign _EVAL_345 = _EVAL_317[13:1];
  assign _EVAL_281 = {{1'd0}, _EVAL_345};
  assign _EVAL_366 = _EVAL_317 | _EVAL_281;
  assign _EVAL_211 = _EVAL_366[13:2];
  assign _EVAL_198 = {{2'd0}, _EVAL_211};
  assign _EVAL_339 = _EVAL_366 | _EVAL_198;
  assign _EVAL_188 = _EVAL_339[13:4];
  assign _EVAL_395 = {{4'd0}, _EVAL_188};
  assign _EVAL_246 = _EVAL_339 | _EVAL_395;
  assign _EVAL_307 = _EVAL_246[13:1];
  assign _EVAL_262 = {{1'd0}, _EVAL_307};
  assign _EVAL_216 = {_EVAL_393, 7'h0};
  assign _EVAL_279 = _EVAL_262 | _EVAL_216;
  assign _EVAL_259 = _EVAL_279[13:7];
  assign _EVAL_399 = _EVAL_279[6:0];
  assign _EVAL_404 = _EVAL_259 & _EVAL_399;
  assign _EVAL_294 = ~ _EVAL_404;
  assign _EVAL_391 = _EVAL_294[2];
  assign _EVAL_148 = _EVAL_391 & _EVAL_17;
  assign _EVAL_387 = _EVAL_2[0];
  assign _EVAL_238 = {{1'd0}, _EVAL_91};
  assign _EVAL_258 = 21'h3f << _EVAL_238;
  assign _EVAL_414 = _EVAL_258[5:0];
  assign _EVAL_403 = ~ _EVAL_414;
  assign _EVAL_213 = _EVAL_403[5:2];
  assign _EVAL_250 = _EVAL_387 ? _EVAL_213 : 4'h0;
  assign _EVAL_343 = _EVAL_148 ? _EVAL_250 : 4'h0;
  assign _EVAL_225 = _EVAL_168 != 7'h0;
  assign _EVAL_312 = _EVAL_10 ^ 30'h1000000;
  assign _EVAL_396 = {1'b0,$signed(_EVAL_312)};
  assign _EVAL_243 = $signed(_EVAL_396) & $signed(31'sh2b004000);
  assign _EVAL_382 = $signed(_EVAL_243);
  assign _EVAL_301 = $signed(_EVAL_382) == $signed(31'sh0);
  assign _EVAL_325 = _EVAL_294[0];
  assign _EVAL_410 = _EVAL_208 == 6'h0;
  assign _EVAL_207 = _EVAL_325 & _EVAL_128;
  assign _EVAL_291 = _EVAL_410 ? _EVAL_207 : _EVAL_215;
  assign _EVAL_192 = {_EVAL_19,_EVAL_135,_EVAL_56,_EVAL_15,_EVAL_60,_EVAL_66,_EVAL_44,_EVAL_84};
  assign _EVAL_334 = _EVAL_291 ? _EVAL_192 : 51'h0;
  assign _EVAL_329 = _EVAL_294[1];
  assign _EVAL_222 = _EVAL_329 & _EVAL_3;
  assign _EVAL_210 = _EVAL_410 ? _EVAL_222 : _EVAL_397;
  assign _EVAL_364 = {{1'd0}, _EVAL_9};
  assign _EVAL_303 = {_EVAL_102,2'h0,_EVAL_364,_EVAL_5,2'h0,_EVAL_81,1'h0};
  assign _EVAL_333 = _EVAL_210 ? _EVAL_303 : 51'h0;
  assign _EVAL_146 = _EVAL_334 | _EVAL_333;
  assign _EVAL_142 = _EVAL_410 ? _EVAL_148 : _EVAL_206;
  assign _EVAL_315 = {_EVAL_2,2'h0,_EVAL_238,_EVAL_48,2'h0,_EVAL_52,1'h0};
  assign _EVAL_306 = _EVAL_142 ? _EVAL_315 : 51'h0;
  assign _EVAL_244 = _EVAL_146 | _EVAL_306;
  assign _EVAL_354 = _EVAL_294 & _EVAL_168;
  assign _EVAL_236 = {_EVAL_354, 1'h0};
  assign _EVAL_268 = _EVAL_236[6:0];
  assign _EVAL_295 = _EVAL_354 | _EVAL_268;
  assign _EVAL_256 = {_EVAL_295, 2'h0};
  assign _EVAL_272 = _EVAL_256[6:0];
  assign _EVAL_271 = _EVAL_295 | _EVAL_272;
  assign _EVAL_214 = {_EVAL_271, 4'h0};
  assign _EVAL_277 = _EVAL_214[6:0];
  assign _EVAL_324 = _EVAL_271 | _EVAL_277;
  assign _EVAL_199 = _EVAL_10 ^ 30'h2000000;
  assign _EVAL_349 = {1'b0,$signed(_EVAL_199)};
  assign _EVAL_251 = $signed(_EVAL_349) & $signed(31'sh2b000000);
  assign _EVAL_356 = $signed(_EVAL_251);
  assign _EVAL_261 = _EVAL_294[4];
  assign _EVAL_341 = _EVAL_261 & _EVAL_31;
  assign _EVAL_323 = _EVAL_410 ? _EVAL_341 : _EVAL_212;
  assign _EVAL_378 = {_EVAL_58,_EVAL_132,_EVAL_229,_EVAL_46,_EVAL_76,_EVAL_123,_EVAL_1,_EVAL_72};
  assign _EVAL_302 = _EVAL_323 ? _EVAL_378 : 51'h0;
  assign _EVAL_369 = {{1'd0}, _EVAL_11};
  assign _EVAL_195 = 21'h3f << _EVAL_369;
  assign _EVAL_413 = _EVAL_207 ? _EVAL_260 : 6'h0;
  assign _EVAL_145 = _EVAL_102[0];
  assign _EVAL_372 = 21'h3f << _EVAL_364;
  assign _EVAL_411 = _EVAL_372[5:0];
  assign _EVAL_300 = ~ _EVAL_411;
  assign _EVAL_247 = _EVAL_300[5:2];
  assign _EVAL_157 = _EVAL_145 ? _EVAL_247 : 4'h0;
  assign _EVAL_293 = _EVAL_222 ? _EVAL_157 : 4'h0;
  assign _EVAL_330 = {{2'd0}, _EVAL_293};
  assign _EVAL_384 = _EVAL_413 | _EVAL_330;
  assign _EVAL_167 = {{2'd0}, _EVAL_343};
  assign _EVAL_196 = _EVAL_384 | _EVAL_167;
  assign _EVAL_314 = _EVAL_294[3];
  assign _EVAL_270 = _EVAL_314 & _EVAL_101;
  assign _EVAL_388 = _EVAL_107[0];
  assign _EVAL_368 = _EVAL_195[5:0];
  assign _EVAL_209 = ~ _EVAL_368;
  assign _EVAL_316 = _EVAL_209[5:2];
  assign _EVAL_370 = _EVAL_388 ? _EVAL_316 : 4'h0;
  assign _EVAL_178 = _EVAL_270 ? _EVAL_370 : 4'h0;
  assign _EVAL_313 = {{2'd0}, _EVAL_178};
  assign _EVAL_161 = _EVAL_196 | _EVAL_313;
  assign _EVAL_239 = _EVAL_58[0];
  assign _EVAL_180 = _EVAL_170[5:0];
  assign _EVAL_350 = ~ _EVAL_180;
  assign _EVAL_389 = _EVAL_350[5:2];
  assign _EVAL_169 = _EVAL_239 ? _EVAL_389 : 4'h0;
  assign _EVAL_171 = _EVAL_341 ? _EVAL_169 : 4'h0;
  assign _EVAL_228 = {{2'd0}, _EVAL_171};
  assign _EVAL_187 = _EVAL_161 | _EVAL_228;
  assign _EVAL_336 = _EVAL_294[5];
  assign _EVAL_275 = _EVAL_336 & _EVAL_70;
  assign _EVAL_357 = _EVAL_22[0];
  assign _EVAL_308 = {{1'd0}, _EVAL_4};
  assign _EVAL_221 = 21'h3f << _EVAL_308;
  assign _EVAL_398 = _EVAL_221[5:0];
  assign _EVAL_402 = ~ _EVAL_398;
  assign _EVAL_347 = _EVAL_402[5:2];
  assign _EVAL_184 = _EVAL_357 ? _EVAL_347 : 4'h0;
  assign _EVAL_355 = _EVAL_275 ? _EVAL_184 : 4'h0;
  assign _EVAL_367 = {{2'd0}, _EVAL_355};
  assign _EVAL_264 = _EVAL_187 | _EVAL_367;
  assign _EVAL_286 = _EVAL_294[6];
  assign _EVAL_310 = _EVAL_286 & _EVAL_63;
  assign _EVAL_280 = _EVAL_116[0];
  assign _EVAL_278 = {{1'd0}, _EVAL_139};
  assign _EVAL_346 = 21'h3f << _EVAL_278;
  assign _EVAL_219 = _EVAL_346[5:0];
  assign _EVAL_408 = ~ _EVAL_219;
  assign _EVAL_149 = _EVAL_408[5:2];
  assign _EVAL_379 = _EVAL_280 ? _EVAL_149 : 4'h0;
  assign _EVAL_153 = _EVAL_310 ? _EVAL_379 : 4'h0;
  assign _EVAL_183 = {{2'd0}, _EVAL_153};
  assign _EVAL_189 = _EVAL_264 | _EVAL_183;
  assign _EVAL_371 = _EVAL_10 ^ 30'h4000;
  assign _EVAL_220 = {1'b0,$signed(_EVAL_371)};
  assign _EVAL_224 = $signed(_EVAL_220) & $signed(31'sh2b005000);
  assign _EVAL_390 = $signed(_EVAL_224);
  assign _EVAL_337 = _EVAL_410 ? _EVAL_314 : _EVAL_223;
  assign _EVAL_181 = $signed(_EVAL_390) == $signed(31'sh0);
  assign _EVAL_363 = _EVAL_181 ? _EVAL_77 : 1'h0;
  assign _EVAL_186 = _EVAL_206 ? _EVAL_17 : 1'h0;
  assign _EVAL_297 = _EVAL_128 | _EVAL_3;
  assign _EVAL_309 = _EVAL_297 | _EVAL_17;
  assign _EVAL_358 = _EVAL_309 | _EVAL_101;
  assign _EVAL_394 = _EVAL_358 | _EVAL_31;
  assign _EVAL_385 = _EVAL_394 | _EVAL_70;
  assign _EVAL_159 = _EVAL_385 | _EVAL_63;
  assign _EVAL_266 = $signed(_EVAL_396) & $signed(31'sh2b000000);
  assign _EVAL_165 = $signed(_EVAL_266);
  assign _EVAL_298 = $signed(_EVAL_165) == $signed(31'sh0);
  assign _EVAL_267 = _EVAL_298 | _EVAL_301;
  assign _EVAL_254 = _EVAL_267 ? _EVAL_82 : 1'h0;
  assign _EVAL_252 = _EVAL_10 ^ 30'h8000000;
  assign _EVAL_377 = {1'b0,$signed(_EVAL_252)};
  assign _EVAL_375 = $signed(_EVAL_377) & $signed(31'sh28000000);
  assign _EVAL_241 = $signed(_EVAL_375);
  assign _EVAL_194 = {1'b0,$signed(_EVAL_10)};
  assign _EVAL_151 = $signed(_EVAL_194) & $signed(31'sh2b005000);
  assign _EVAL_190 = $signed(_EVAL_151);
  assign _EVAL_318 = _EVAL_410 ? _EVAL_391 : _EVAL_206;
  assign _EVAL_147 = _EVAL_10 ^ 30'h20000000;
  assign _EVAL_202 = _EVAL_410 ? _EVAL_270 : _EVAL_223;
  assign _EVAL_292 = {_EVAL_107,2'h0,_EVAL_369,_EVAL_108,2'h0,_EVAL_106,1'h0};
  assign _EVAL_328 = _EVAL_202 ? _EVAL_292 : 51'h0;
  assign _EVAL_248 = _EVAL_244 | _EVAL_328;
  assign _EVAL_175 = _EVAL_248 | _EVAL_302;
  assign _EVAL_365 = _EVAL_410 ? _EVAL_275 : _EVAL_164;
  assign _EVAL_380 = {_EVAL_22,2'h0,_EVAL_308,_EVAL_75,2'h0,_EVAL_138,1'h0};
  assign _EVAL_409 = _EVAL_365 ? _EVAL_380 : 51'h0;
  assign _EVAL_234 = _EVAL_175 | _EVAL_409;
  assign _EVAL_332 = _EVAL_410 ? _EVAL_310 : _EVAL_255;
  assign _EVAL_290 = {_EVAL_116,2'h0,_EVAL_278,_EVAL_20,1'h0,_EVAL_73,_EVAL_40,_EVAL_24};
  assign _EVAL_179 = _EVAL_332 ? _EVAL_290 : 51'h0;
  assign _EVAL_322 = _EVAL_234 | _EVAL_179;
  assign _EVAL_320 = _EVAL_410 ? _EVAL_329 : _EVAL_397;
  assign _EVAL_353 = _EVAL_10 ^ 30'h1000;
  assign _EVAL_348 = {1'b0,$signed(_EVAL_353)};
  assign _EVAL_163 = $signed(_EVAL_348) & $signed(31'sh2b005000);
  assign _EVAL_374 = $signed(_EVAL_163);
  assign _EVAL_158 = $signed(_EVAL_374) == $signed(31'sh0);
  assign _EVAL_200 = _EVAL_158 ? _EVAL_29 : 1'h0;
  assign _EVAL_284 = $signed(_EVAL_241) == $signed(31'sh0);
  assign _EVAL_257 = _EVAL_284 ? _EVAL_129 : 1'h0;
  assign _EVAL_177 = _EVAL_200 | _EVAL_257;
  assign _EVAL_331 = $signed(_EVAL_356) == $signed(31'sh0);
  assign _EVAL_182 = _EVAL_331 ? _EVAL_45 : 1'h0;
  assign _EVAL_185 = _EVAL_177 | _EVAL_182;
  assign _EVAL_150 = {1'b0,$signed(_EVAL_147)};
  assign _EVAL_245 = $signed(_EVAL_150) & $signed(31'sh2b004000);
  assign _EVAL_152 = $signed(_EVAL_245);
  assign _EVAL_304 = $signed(_EVAL_152) == $signed(31'sh0);
  assign _EVAL_237 = _EVAL_223 ? _EVAL_101 : 1'h0;
  assign _EVAL_412 = _EVAL_410 & _EVAL_25;
  assign _EVAL_249 = _EVAL_412 & _EVAL_225;
  assign _EVAL_173 = _EVAL_410 ? _EVAL_261 : _EVAL_212;
  assign _EVAL_265 = _EVAL_326 | _EVAL_186;
  assign _EVAL_154 = _EVAL_265 | _EVAL_237;
  assign _EVAL_406 = _EVAL_212 ? _EVAL_31 : 1'h0;
  assign _EVAL_230 = _EVAL_154 | _EVAL_406;
  assign _EVAL_263 = _EVAL_164 ? _EVAL_70 : 1'h0;
  assign _EVAL_218 = _EVAL_230 | _EVAL_263;
  assign _EVAL_401 = _EVAL_255 ? _EVAL_63 : 1'h0;
  assign _EVAL_166 = _EVAL_218 | _EVAL_401;
  assign _EVAL_340 = _EVAL_410 ? _EVAL_159 : _EVAL_166;
  assign _EVAL_296 = _EVAL_25 & _EVAL_340;
  assign _EVAL_335 = {{5'd0}, _EVAL_296};
  assign _EVAL_233 = _EVAL_208 - _EVAL_335;
  assign _EVAL_285 = $signed(_EVAL_190) == $signed(31'sh0);
  assign _EVAL_351 = _EVAL_285 ? _EVAL_33 : 1'h0;
  assign _EVAL_203 = _EVAL_185 | _EVAL_351;
  assign _EVAL_226 = _EVAL_203 | _EVAL_254;
  assign _EVAL_283 = _EVAL_410 ? _EVAL_286 : _EVAL_255;
  assign _EVAL_311 = _EVAL_410 ? _EVAL_336 : _EVAL_164;
  assign _EVAL_217 = _EVAL_304 ? _EVAL_92 : 1'h0;
  assign _EVAL_305 = _EVAL_226 | _EVAL_363;
  assign _EVAL_160 = _EVAL_410 ? _EVAL_325 : _EVAL_215;
  assign _EVAL_90 = _EVAL_322[41:35];
  assign _EVAL_97 = _EVAL_25 & _EVAL_311;
  assign _EVAL_131 = _EVAL_64;
  assign _EVAL_86 = _EVAL_53;
  assign _EVAL_13 = _EVAL_305 | _EVAL_217;
  assign _EVAL_12 = _EVAL_127;
  assign _EVAL_8 = _EVAL_113[2:0];
  assign _EVAL_78 = _EVAL_64;
  assign _EVAL_122 = _EVAL_64;
  assign _EVAL_115 = _EVAL_10[11:0];
  assign _EVAL_28 = _EVAL_133;
  assign _EVAL_103 = _EVAL_25 & _EVAL_320;
  assign _EVAL_65 = _EVAL_96;
  assign _EVAL_134 = _EVAL_61 & _EVAL_158;
  assign _EVAL_118 = _EVAL_61 & _EVAL_304;
  assign _EVAL_117 = _EVAL_133;
  assign _EVAL_80 = _EVAL_25 & _EVAL_283;
  assign _EVAL_34 = _EVAL_322[45:42];
  assign _EVAL_125 = _EVAL_133;
  assign _EVAL_42 = _EVAL_133;
  assign _EVAL_83 = _EVAL_10[24:0];
  assign _EVAL_120 = _EVAL_96;
  assign _EVAL_79 = _EVAL_25 & _EVAL_318;
  assign _EVAL_105 = _EVAL_322[50:48];
  assign _EVAL_137 = _EVAL_25 & _EVAL_173;
  assign _EVAL_85 = _EVAL_121;
  assign _EVAL_126 = _EVAL_113[2:0];
  assign _EVAL_14 = _EVAL_410 ? _EVAL_159 : _EVAL_166;
  assign _EVAL_98 = _EVAL_10[25:0];
  assign _EVAL_59 = _EVAL_127;
  assign _EVAL_109 = _EVAL_61 & _EVAL_267;
  assign _EVAL_71 = _EVAL_113;
  assign _EVAL_124 = _EVAL_64;
  assign _EVAL_57 = _EVAL_322[34];
  assign _EVAL = _EVAL_10[27:0];
  assign _EVAL_36 = _EVAL_53;
  assign _EVAL_67 = _EVAL_61 & _EVAL_284;
  assign _EVAL_130 = _EVAL_64;
  assign _EVAL_54 = _EVAL_53;
  assign _EVAL_39 = _EVAL_25 & _EVAL_160;
  assign _EVAL_140 = _EVAL_96;
  assign _EVAL_51 = _EVAL_133;
  assign _EVAL_38 = _EVAL_10;
  assign _EVAL_99 = _EVAL_127;
  assign _EVAL_62 = _EVAL_121;
  assign _EVAL_69 = _EVAL_127;
  assign _EVAL_50 = _EVAL_53;
  assign _EVAL_0 = _EVAL_64;
  assign _EVAL_30 = _EVAL_121;
  assign _EVAL_95 = _EVAL_133;
  assign _EVAL_37 = _EVAL_64;
  assign _EVAL_6 = _EVAL_127;
  assign _EVAL_104 = _EVAL_113[2:0];
  assign _EVAL_100 = _EVAL_322[33];
  assign _EVAL_88 = _EVAL_322[0];
  assign _EVAL_47 = _EVAL_121;
  assign _EVAL_74 = _EVAL_322[32:1];
  assign _EVAL_87 = _EVAL_61 & _EVAL_285;
  assign _EVAL_111 = _EVAL_133;
  assign _EVAL_23 = _EVAL_10[13:0];
  assign _EVAL_35 = _EVAL_53;
  assign _EVAL_43 = _EVAL_113[2:0];
  assign _EVAL_114 = _EVAL_53;
  assign _EVAL_93 = _EVAL_96;
  assign _EVAL_136 = _EVAL_121;
  assign _EVAL_7 = _EVAL_61 & _EVAL_331;
  assign _EVAL_119 = _EVAL_96;
  assign _EVAL_94 = _EVAL_127;
  assign _EVAL_26 = _EVAL_53;
  assign _EVAL_89 = _EVAL_322[47:46];
  assign _EVAL_110 = _EVAL_96;
  assign _EVAL_112 = _EVAL_25 & _EVAL_337;
  assign _EVAL_18 = _EVAL_113[2:0];
  assign _EVAL_21 = _EVAL_121;
  assign _EVAL_41 = _EVAL_61 & _EVAL_181;
  assign _EVAL_55 = _EVAL_10[14:0];
  assign _EVAL_32 = _EVAL_121;
  assign _EVAL_68 = _EVAL_127;
  assign _EVAL_141 = _EVAL_113[2:0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_164 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_206 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_208 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_212 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_215 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_223 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_255 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_393 = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_397 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_49) begin
    if (_EVAL_16) begin
      _EVAL_164 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_164 <= _EVAL_275;
      end
    end
    if (_EVAL_16) begin
      _EVAL_206 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_206 <= _EVAL_148;
      end
    end
    if (_EVAL_16) begin
      _EVAL_208 <= 6'h0;
    end else begin
      if (_EVAL_412) begin
        _EVAL_208 <= _EVAL_189;
      end else begin
        _EVAL_208 <= _EVAL_233;
      end
    end
    if (_EVAL_16) begin
      _EVAL_212 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_212 <= _EVAL_341;
      end
    end
    if (_EVAL_16) begin
      _EVAL_215 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_215 <= _EVAL_207;
      end
    end
    if (_EVAL_16) begin
      _EVAL_223 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_223 <= _EVAL_270;
      end
    end
    if (_EVAL_16) begin
      _EVAL_255 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_255 <= _EVAL_310;
      end
    end
    if (_EVAL_16) begin
      _EVAL_393 <= 7'h7f;
    end else begin
      if (_EVAL_249) begin
        _EVAL_393 <= _EVAL_324;
      end
    end
    if (_EVAL_16) begin
      _EVAL_397 <= 1'h0;
    end else begin
      if (_EVAL_410) begin
        _EVAL_397 <= _EVAL_222;
      end
    end
  end
endmodule
