//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_49(
  output        _EVAL,
  input  [3:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  input  [7:0]  _EVAL_2,
  output [2:0]  _EVAL_3,
  input  [63:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  output [3:0]  _EVAL_8,
  output [63:0] _EVAL_9,
  input  [1:0]  _EVAL_10,
  output [31:0] _EVAL_11,
  output [3:0]  _EVAL_12,
  output [1:0]  _EVAL_13,
  input         _EVAL_14,
  output [7:0]  _EVAL_15,
  input  [31:0] _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  output        _EVAL_19,
  output [2:0]  _EVAL_20,
  input  [1:0]  _EVAL_21,
  output [1:0]  _EVAL_22,
  output [2:0]  _EVAL_23,
  output [1:0]  _EVAL_24,
  output [6:0]  _EVAL_25,
  output [3:0]  _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  output [3:0]  _EVAL_29,
  output [30:0] _EVAL_30,
  input         _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input  [3:0]  _EVAL_34,
  input  [2:0]  _EVAL_35,
  output [3:0]  _EVAL_36,
  input  [2:0]  _EVAL_37,
  output [3:0]  _EVAL_38,
  output [2:0]  _EVAL_39,
  input  [2:0]  _EVAL_40,
  input         _EVAL_41,
  output [2:0]  _EVAL_42,
  input         _EVAL_43,
  input  [5:0]  _EVAL_44,
  input  [1:0]  _EVAL_45,
  input         _EVAL_46,
  input  [3:0]  _EVAL_47,
  input  [31:0] _EVAL_48,
  output [2:0]  _EVAL_49,
  input         _EVAL_50,
  output [1:0]  _EVAL_51,
  output        _EVAL_52,
  output        _EVAL_53,
  input  [1:0]  _EVAL_54,
  output [3:0]  _EVAL_55,
  input         _EVAL_56,
  output        _EVAL_57,
  output        _EVAL_58,
  input  [1:0]  _EVAL_59,
  output [2:0]  _EVAL_60,
  output        _EVAL_61,
  input  [31:0] _EVAL_62,
  output        _EVAL_63,
  output [6:0]  _EVAL_64,
  output [2:0]  _EVAL_65,
  input  [31:0] _EVAL_66,
  input         _EVAL_67,
  output [1:0]  _EVAL_68,
  input         _EVAL_69,
  input  [63:0] _EVAL_70,
  output [63:0] _EVAL_71,
  output [30:0] _EVAL_72,
  output [63:0] _EVAL_73,
  input  [63:0] _EVAL_74,
  output [31:0] _EVAL_75,
  input         _EVAL_76,
  output [1:0]  _EVAL_77,
  output [2:0]  _EVAL_78,
  input  [3:0]  _EVAL_79,
  output [6:0]  _EVAL_80,
  output [3:0]  _EVAL_81,
  output        _EVAL_82,
  output        _EVAL_83,
  output [31:0] _EVAL_84,
  input  [2:0]  _EVAL_85,
  input  [2:0]  _EVAL_86,
  output [1:0]  _EVAL_87,
  input  [6:0]  _EVAL_88,
  input  [31:0] _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  output [31:0] _EVAL_92,
  input  [31:0] _EVAL_93,
  output [1:0]  _EVAL_94,
  input  [2:0]  _EVAL_95,
  output [31:0] _EVAL_96,
  input  [1:0]  _EVAL_97,
  input         _EVAL_98,
  input  [3:0]  _EVAL_99,
  output [1:0]  _EVAL_100,
  input         _EVAL_101,
  output [7:0]  _EVAL_102,
  output        _EVAL_103,
  input         _EVAL_104,
  input  [63:0] _EVAL_105,
  input         _EVAL_106,
  output [3:0]  _EVAL_107,
  input  [1:0]  _EVAL_108,
  output [3:0]  _EVAL_109,
  input         _EVAL_110,
  output [2:0]  _EVAL_111,
  input  [2:0]  _EVAL_112,
  output        _EVAL_113,
  input         _EVAL_114,
  input         _EVAL_115,
  input  [6:0]  _EVAL_116,
  output [3:0]  _EVAL_117,
  input  [3:0]  _EVAL_118,
  output [6:0]  _EVAL_119,
  input  [3:0]  _EVAL_120,
  output        _EVAL_121,
  output        _EVAL_122,
  input  [1:0]  _EVAL_123,
  output        _EVAL_124,
  output [29:0] _EVAL_125,
  input         _EVAL_126,
  input         _EVAL_127,
  input  [6:0]  _EVAL_128,
  output        _EVAL_129,
  input  [2:0]  _EVAL_130,
  input  [3:0]  _EVAL_131,
  output [2:0]  _EVAL_132,
  input         _EVAL_133,
  input         _EVAL_134,
  input         _EVAL_135,
  output        _EVAL_136,
  input         _EVAL_137,
  input  [3:0]  _EVAL_138,
  output        _EVAL_139,
  output [2:0]  _EVAL_140,
  output        _EVAL_141,
  output [7:0]  _EVAL_142,
  input  [63:0] _EVAL_143,
  input         _EVAL_144,
  input  [31:0] _EVAL_145,
  output        _EVAL_146,
  output        _EVAL_147,
  output        _EVAL_148,
  input         _EVAL_149,
  input         _EVAL_150,
  input  [3:0]  _EVAL_151,
  output [6:0]  _EVAL_152,
  input         _EVAL_153,
  output        _EVAL_154,
  output [2:0]  _EVAL_155,
  output        _EVAL_156,
  input  [2:0]  _EVAL_157,
  input  [2:0]  _EVAL_158,
  input         _EVAL_159,
  output        _EVAL_160,
  input  [1:0]  _EVAL_161,
  output [2:0]  _EVAL_162,
  input  [3:0]  _EVAL_163,
  output        _EVAL_164,
  output        _EVAL_165,
  input         _EVAL_166,
  output        _EVAL_167,
  input  [7:0]  _EVAL_168,
  input         _EVAL_169,
  output        _EVAL_170,
  output        _EVAL_171,
  input  [31:0] _EVAL_172,
  input  [3:0]  _EVAL_173,
  output [1:0]  _EVAL_174,
  output [3:0]  _EVAL_175,
  output [3:0]  _EVAL_176,
  output [31:0] _EVAL_177,
  input         _EVAL_178,
  input  [3:0]  _EVAL_179,
  output [31:0] _EVAL_180,
  output [29:0] _EVAL_181,
  input  [3:0]  _EVAL_182,
  output        _EVAL_183,
  output [63:0] _EVAL_184,
  output [7:0]  _EVAL_185,
  input  [2:0]  _EVAL_186,
  input  [31:0] _EVAL_187,
  output [5:0]  _EVAL_188,
  input  [2:0]  _EVAL_189,
  input  [63:0] _EVAL_190,
  input  [2:0]  _EVAL_191,
  input  [6:0]  _EVAL_192,
  output [63:0] _EVAL_193,
  input  [2:0]  _EVAL_194,
  output        _EVAL_195,
  output [3:0]  _EVAL_196,
  input  [63:0] _EVAL_197,
  output [1:0]  _EVAL_198,
  input  [29:0] _EVAL_199,
  output [63:0] _EVAL_200,
  output [3:0]  _EVAL_201,
  output        _EVAL_202,
  input         _EVAL_203,
  input  [1:0]  _EVAL_204,
  output        _EVAL_205,
  output [2:0]  _EVAL_206,
  input         _EVAL_207,
  output [1:0]  _EVAL_208,
  input  [2:0]  _EVAL_209,
  input  [7:0]  _EVAL_210,
  input         _EVAL_211,
  output        _EVAL_212,
  output        _EVAL_213,
  output        _EVAL_214,
  output [1:0]  _EVAL_215,
  output        _EVAL_216,
  output [2:0]  _EVAL_217,
  output        _EVAL_218,
  output        _EVAL_219,
  output        _EVAL_220,
  input  [3:0]  _EVAL_221,
  input         _EVAL_222,
  output [3:0]  _EVAL_223,
  output [2:0]  _EVAL_224
);
  wire [6:0] coupler_to_bus_named_cbus__EVAL;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_0;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_1;
  wire  coupler_to_bus_named_cbus__EVAL_2;
  wire  coupler_to_bus_named_cbus__EVAL_3;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_4;
  wire  coupler_to_bus_named_cbus__EVAL_5;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_6;
  wire  coupler_to_bus_named_cbus__EVAL_7;
  wire [6:0] coupler_to_bus_named_cbus__EVAL_8;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_9;
  wire  coupler_to_bus_named_cbus__EVAL_10;
  wire  coupler_to_bus_named_cbus__EVAL_11;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_12;
  wire  coupler_to_bus_named_cbus__EVAL_13;
  wire  coupler_to_bus_named_cbus__EVAL_14;
  wire  coupler_to_bus_named_cbus__EVAL_15;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_16;
  wire [31:0] coupler_to_bus_named_cbus__EVAL_17;
  wire [63:0] coupler_to_bus_named_cbus__EVAL_18;
  wire [7:0] coupler_to_bus_named_cbus__EVAL_19;
  wire [31:0] coupler_to_bus_named_cbus__EVAL_20;
  wire  coupler_to_bus_named_cbus__EVAL_21;
  wire  coupler_to_bus_named_cbus__EVAL_22;
  wire [6:0] coupler_to_bus_named_cbus__EVAL_23;
  wire [63:0] coupler_to_bus_named_cbus__EVAL_24;
  wire [29:0] coupler_to_bus_named_cbus__EVAL_25;
  wire  coupler_to_bus_named_cbus__EVAL_26;
  wire  coupler_to_bus_named_cbus__EVAL_27;
  wire [29:0] coupler_to_bus_named_cbus__EVAL_28;
  wire [1:0] coupler_to_bus_named_cbus__EVAL_29;
  wire [1:0] coupler_to_bus_named_cbus__EVAL_30;
  wire  coupler_to_bus_named_cbus__EVAL_31;
  wire  coupler_to_bus_named_cbus__EVAL_32;
  wire  coupler_to_bus_named_cbus__EVAL_33;
  wire [6:0] coupler_to_bus_named_cbus__EVAL_34;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_35;
  wire  coupler_to_bus_named_cbus__EVAL_36;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_37;
  wire  coupler_to_bus_named_cbus__EVAL_38;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_39;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_40;
  wire  system_bus_xbar__EVAL;
  wire [2:0] system_bus_xbar__EVAL_0;
  wire  system_bus_xbar__EVAL_1;
  wire [6:0] system_bus_xbar__EVAL_2;
  wire [2:0] system_bus_xbar__EVAL_3;
  wire [6:0] system_bus_xbar__EVAL_4;
  wire [7:0] system_bus_xbar__EVAL_5;
  wire [3:0] system_bus_xbar__EVAL_6;
  wire [2:0] system_bus_xbar__EVAL_7;
  wire [2:0] system_bus_xbar__EVAL_8;
  wire  system_bus_xbar__EVAL_9;
  wire  system_bus_xbar__EVAL_10;
  wire [2:0] system_bus_xbar__EVAL_11;
  wire [31:0] system_bus_xbar__EVAL_12;
  wire [31:0] system_bus_xbar__EVAL_13;
  wire [2:0] system_bus_xbar__EVAL_14;
  wire  system_bus_xbar__EVAL_15;
  wire  system_bus_xbar__EVAL_16;
  wire [2:0] system_bus_xbar__EVAL_17;
  wire [2:0] system_bus_xbar__EVAL_18;
  wire [63:0] system_bus_xbar__EVAL_19;
  wire [6:0] system_bus_xbar__EVAL_20;
  wire [63:0] system_bus_xbar__EVAL_21;
  wire [2:0] system_bus_xbar__EVAL_22;
  wire  system_bus_xbar__EVAL_23;
  wire  system_bus_xbar__EVAL_24;
  wire  system_bus_xbar__EVAL_25;
  wire [6:0] system_bus_xbar__EVAL_26;
  wire [31:0] system_bus_xbar__EVAL_27;
  wire [3:0] system_bus_xbar__EVAL_28;
  wire  system_bus_xbar__EVAL_29;
  wire  system_bus_xbar__EVAL_30;
  wire [1:0] system_bus_xbar__EVAL_31;
  wire [2:0] system_bus_xbar__EVAL_32;
  wire [31:0] system_bus_xbar__EVAL_33;
  wire [6:0] system_bus_xbar__EVAL_34;
  wire [2:0] system_bus_xbar__EVAL_35;
  wire  system_bus_xbar__EVAL_36;
  wire [2:0] system_bus_xbar__EVAL_37;
  wire  system_bus_xbar__EVAL_38;
  wire  system_bus_xbar__EVAL_39;
  wire [3:0] system_bus_xbar__EVAL_40;
  wire [2:0] system_bus_xbar__EVAL_41;
  wire  system_bus_xbar__EVAL_42;
  wire  system_bus_xbar__EVAL_43;
  wire  system_bus_xbar__EVAL_44;
  wire [2:0] system_bus_xbar__EVAL_45;
  wire  system_bus_xbar__EVAL_46;
  wire [63:0] system_bus_xbar__EVAL_47;
  wire [2:0] system_bus_xbar__EVAL_48;
  wire  system_bus_xbar__EVAL_49;
  wire  system_bus_xbar__EVAL_50;
  wire  system_bus_xbar__EVAL_51;
  wire [63:0] system_bus_xbar__EVAL_52;
  wire [31:0] system_bus_xbar__EVAL_53;
  wire  system_bus_xbar__EVAL_54;
  wire [29:0] system_bus_xbar__EVAL_55;
  wire [3:0] system_bus_xbar__EVAL_56;
  wire  system_bus_xbar__EVAL_57;
  wire [2:0] system_bus_xbar__EVAL_58;
  wire [1:0] system_bus_xbar__EVAL_59;
  wire  system_bus_xbar__EVAL_60;
  wire [2:0] system_bus_xbar__EVAL_61;
  wire [2:0] system_bus_xbar__EVAL_62;
  wire  system_bus_xbar__EVAL_63;
  wire  system_bus_xbar__EVAL_64;
  wire  system_bus_xbar__EVAL_65;
  wire  system_bus_xbar__EVAL_66;
  wire [7:0] system_bus_xbar__EVAL_67;
  wire [1:0] system_bus_xbar__EVAL_68;
  wire [31:0] system_bus_xbar__EVAL_69;
  wire [63:0] system_bus_xbar__EVAL_70;
  wire [3:0] system_bus_xbar__EVAL_71;
  wire  system_bus_xbar__EVAL_72;
  wire  system_bus_xbar__EVAL_73;
  wire  system_bus_xbar__EVAL_74;
  wire [2:0] system_bus_xbar__EVAL_75;
  wire [63:0] system_bus_xbar__EVAL_76;
  wire [3:0] system_bus_xbar__EVAL_77;
  wire  system_bus_xbar__EVAL_78;
  wire [63:0] system_bus_xbar__EVAL_79;
  wire [1:0] system_bus_xbar__EVAL_80;
  wire  system_bus_xbar__EVAL_81;
  wire  system_bus_xbar__EVAL_82;
  wire  system_bus_xbar__EVAL_83;
  wire  system_bus_xbar__EVAL_84;
  wire [6:0] system_bus_xbar__EVAL_85;
  wire  system_bus_xbar__EVAL_86;
  wire [63:0] system_bus_xbar__EVAL_87;
  wire [7:0] system_bus_xbar__EVAL_88;
  wire [5:0] system_bus_xbar__EVAL_89;
  wire [2:0] system_bus_xbar__EVAL_90;
  wire  system_bus_xbar__EVAL_91;
  wire  system_bus_xbar__EVAL_92;
  wire [7:0] system_bus_xbar__EVAL_93;
  wire [63:0] system_bus_xbar__EVAL_94;
  wire [3:0] system_bus_xbar__EVAL_95;
  wire  system_bus_xbar__EVAL_96;
  wire  system_bus_xbar__EVAL_97;
  wire [2:0] system_bus_xbar__EVAL_98;
  wire  system_bus_xbar__EVAL_99;
  wire  system_bus_xbar__EVAL_100;
  wire  system_bus_xbar__EVAL_101;
  wire [3:0] system_bus_xbar__EVAL_102;
  wire  system_bus_xbar__EVAL_103;
  wire [3:0] system_bus_xbar__EVAL_104;
  wire  system_bus_xbar__EVAL_105;
  wire  system_bus_xbar__EVAL_106;
  wire  system_bus_xbar__EVAL_107;
  wire [2:0] system_bus_xbar__EVAL_108;
  wire [1:0] system_bus_xbar__EVAL_109;
  wire [1:0] system_bus_xbar__EVAL_110;
  wire [63:0] system_bus_xbar__EVAL_111;
  wire [63:0] system_bus_xbar__EVAL_112;
  wire  system_bus_xbar__EVAL_113;
  wire [31:0] system_bus_xbar__EVAL_114;
  wire  system_bus_xbar__EVAL_115;
  wire [30:0] system_bus_xbar__EVAL_116;
  wire [3:0] system_bus_xbar__EVAL_117;
  wire [2:0] system_bus_xbar__EVAL_118;
  wire [63:0] system_bus_xbar__EVAL_119;
  wire  system_bus_xbar__EVAL_120;
  wire [7:0] system_bus_xbar__EVAL_121;
  wire  system_bus_xbar__EVAL_122;
  wire  system_bus_xbar__EVAL_123;
  wire  system_bus_xbar__EVAL_124;
  wire [6:0] system_bus_xbar__EVAL_125;
  wire  system_bus_xbar__EVAL_126;
  wire [5:0] system_bus_xbar__EVAL_127;
  wire [2:0] system_bus_xbar__EVAL_128;
  wire [3:0] coupler_from_tile_with_no_name__EVAL;
  wire  coupler_from_tile_with_no_name__EVAL_0;
  wire  coupler_from_tile_with_no_name__EVAL_1;
  wire  coupler_from_tile_with_no_name__EVAL_2;
  wire  coupler_from_tile_with_no_name__EVAL_3;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_4;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_5;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_6;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_7;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_8;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_9;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_10;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_11;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_12;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_13;
  wire  coupler_from_tile_with_no_name__EVAL_14;
  wire [7:0] coupler_from_tile_with_no_name__EVAL_15;
  wire  coupler_from_tile_with_no_name__EVAL_16;
  wire  coupler_from_tile_with_no_name__EVAL_17;
  wire  coupler_from_tile_with_no_name__EVAL_18;
  wire  coupler_from_tile_with_no_name__EVAL_19;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_20;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_21;
  wire  coupler_from_tile_with_no_name__EVAL_22;
  wire  coupler_from_tile_with_no_name__EVAL_23;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_24;
  wire  coupler_from_tile_with_no_name__EVAL_25;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_26;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_27;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_28;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_29;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_30;
  wire  coupler_from_tile_with_no_name__EVAL_31;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_32;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_33;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_34;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_35;
  wire  coupler_from_tile_with_no_name__EVAL_36;
  wire  coupler_from_tile_with_no_name__EVAL_37;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_38;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_39;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_40;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_41;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_42;
  wire  coupler_from_tile_with_no_name__EVAL_43;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_44;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_45;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_46;
  wire  coupler_from_tile_with_no_name__EVAL_47;
  wire  coupler_from_tile_with_no_name__EVAL_48;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_49;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_50;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_51;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_52;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_53;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_54;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_55;
  wire  coupler_from_tile_with_no_name__EVAL_56;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_57;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_58;
  wire [7:0] coupler_from_tile_with_no_name__EVAL_59;
  wire  coupler_from_tile_with_no_name__EVAL_60;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_61;
  wire  coupler_from_tile_with_no_name__EVAL_62;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_63;
  wire  coupler_from_tile_with_no_name__EVAL_64;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_65;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_66;
  wire  coupler_from_tile_with_no_name__EVAL_67;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_68;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_69;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_70;
  wire  coupler_from_tile_with_no_name__EVAL_71;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_72;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_73;
  wire  coupler_from_tile_with_no_name__EVAL_74;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_75;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_76;
  wire  coupler_from_tile_with_no_name__EVAL_77;
  wire  coupler_from_tile_with_no_name__EVAL_78;
  wire  coupler_from_tile_with_no_name__EVAL_79;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_80;
  wire  coupler_from_tile_with_no_name__EVAL_81;
  wire  coupler_from_tile_with_no_name__EVAL_82;
  wire  coupler_from_tile_with_no_name__EVAL_83;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_84;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_85;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_86;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_87;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_88;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_89;
  wire  coupler_from_tile_with_no_name__EVAL_90;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_91;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_92;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_93;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_94;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_95;
  wire  coupler_from_tile_with_no_name__EVAL_96;
  wire  coupler_from_tile_with_no_name__EVAL_97;
  wire  coupler_from_tile_with_no_name__EVAL_98;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_99;
  wire  coupler_from_tile_with_no_name__EVAL_100;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_101;
  wire [63:0] coupler_from_tile_with_no_name__EVAL_102;
  wire  coupler_from_tile_with_no_name__EVAL_103;
  wire  coupler_from_tile_with_no_name__EVAL_104;
  wire [7:0] coupler_from_tile_with_no_name__EVAL_105;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_106;
  wire  coupler_from_tile_with_no_name__EVAL_107;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_0;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_1;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_2;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_3;
  wire [1:0] coupler_to_port_named_axi4_sys_port__EVAL_4;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_5;
  wire [63:0] coupler_to_port_named_axi4_sys_port__EVAL_6;
  wire [1:0] coupler_to_port_named_axi4_sys_port__EVAL_7;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_8;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_9;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_10;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_11;
  wire [1:0] coupler_to_port_named_axi4_sys_port__EVAL_12;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_13;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_14;
  wire [1:0] coupler_to_port_named_axi4_sys_port__EVAL_15;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_16;
  wire [30:0] coupler_to_port_named_axi4_sys_port__EVAL_17;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_18;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_19;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_20;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_21;
  wire [63:0] coupler_to_port_named_axi4_sys_port__EVAL_22;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_23;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_24;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_25;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_26;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_27;
  wire [6:0] coupler_to_port_named_axi4_sys_port__EVAL_28;
  wire [30:0] coupler_to_port_named_axi4_sys_port__EVAL_29;
  wire [31:0] coupler_to_port_named_axi4_sys_port__EVAL_30;
  wire [6:0] coupler_to_port_named_axi4_sys_port__EVAL_31;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_32;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_33;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_34;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_35;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_36;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_37;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_38;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_39;
  wire [31:0] coupler_to_port_named_axi4_sys_port__EVAL_40;
  wire [30:0] coupler_to_port_named_axi4_sys_port__EVAL_41;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_42;
  wire [7:0] coupler_to_port_named_axi4_sys_port__EVAL_43;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_44;
  wire [7:0] coupler_to_port_named_axi4_sys_port__EVAL_45;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_46;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_47;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_48;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_49;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_50;
  wire [2:0] coupler_to_port_named_axi4_sys_port__EVAL_51;
  wire [7:0] coupler_to_port_named_axi4_sys_port__EVAL_52;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_53;
  wire  coupler_to_port_named_axi4_sys_port__EVAL_54;
  wire [3:0] coupler_to_port_named_axi4_sys_port__EVAL_55;
  wire  coupler_from_bus_named_front_bus__EVAL;
  wire [5:0] coupler_from_bus_named_front_bus__EVAL_0;
  wire [63:0] coupler_from_bus_named_front_bus__EVAL_1;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_2;
  wire [1:0] coupler_from_bus_named_front_bus__EVAL_3;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_4;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_5;
  wire  coupler_from_bus_named_front_bus__EVAL_6;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_7;
  wire  coupler_from_bus_named_front_bus__EVAL_8;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_9;
  wire [63:0] coupler_from_bus_named_front_bus__EVAL_10;
  wire [1:0] coupler_from_bus_named_front_bus__EVAL_11;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_12;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_13;
  wire  coupler_from_bus_named_front_bus__EVAL_14;
  wire  coupler_from_bus_named_front_bus__EVAL_15;
  wire  coupler_from_bus_named_front_bus__EVAL_16;
  wire  coupler_from_bus_named_front_bus__EVAL_17;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_18;
  wire [5:0] coupler_from_bus_named_front_bus__EVAL_19;
  wire  coupler_from_bus_named_front_bus__EVAL_20;
  wire  coupler_from_bus_named_front_bus__EVAL_21;
  wire  coupler_from_bus_named_front_bus__EVAL_22;
  wire  coupler_from_bus_named_front_bus__EVAL_23;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_24;
  wire  coupler_from_bus_named_front_bus__EVAL_25;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_26;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_27;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_28;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_29;
  wire [7:0] coupler_from_bus_named_front_bus__EVAL_30;
  wire  coupler_from_bus_named_front_bus__EVAL_31;
  wire  coupler_from_bus_named_front_bus__EVAL_32;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_33;
  wire  coupler_from_bus_named_front_bus__EVAL_34;
  wire [5:0] coupler_from_bus_named_front_bus__EVAL_35;
  wire  coupler_from_bus_named_front_bus__EVAL_36;
  wire  coupler_from_bus_named_front_bus__EVAL_37;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_38;
  wire [5:0] coupler_from_bus_named_front_bus__EVAL_39;
  wire  coupler_from_bus_named_front_bus__EVAL_40;
  SiFive__EVAL_44 coupler_to_bus_named_cbus (
    ._EVAL(coupler_to_bus_named_cbus__EVAL),
    ._EVAL_0(coupler_to_bus_named_cbus__EVAL_0),
    ._EVAL_1(coupler_to_bus_named_cbus__EVAL_1),
    ._EVAL_2(coupler_to_bus_named_cbus__EVAL_2),
    ._EVAL_3(coupler_to_bus_named_cbus__EVAL_3),
    ._EVAL_4(coupler_to_bus_named_cbus__EVAL_4),
    ._EVAL_5(coupler_to_bus_named_cbus__EVAL_5),
    ._EVAL_6(coupler_to_bus_named_cbus__EVAL_6),
    ._EVAL_7(coupler_to_bus_named_cbus__EVAL_7),
    ._EVAL_8(coupler_to_bus_named_cbus__EVAL_8),
    ._EVAL_9(coupler_to_bus_named_cbus__EVAL_9),
    ._EVAL_10(coupler_to_bus_named_cbus__EVAL_10),
    ._EVAL_11(coupler_to_bus_named_cbus__EVAL_11),
    ._EVAL_12(coupler_to_bus_named_cbus__EVAL_12),
    ._EVAL_13(coupler_to_bus_named_cbus__EVAL_13),
    ._EVAL_14(coupler_to_bus_named_cbus__EVAL_14),
    ._EVAL_15(coupler_to_bus_named_cbus__EVAL_15),
    ._EVAL_16(coupler_to_bus_named_cbus__EVAL_16),
    ._EVAL_17(coupler_to_bus_named_cbus__EVAL_17),
    ._EVAL_18(coupler_to_bus_named_cbus__EVAL_18),
    ._EVAL_19(coupler_to_bus_named_cbus__EVAL_19),
    ._EVAL_20(coupler_to_bus_named_cbus__EVAL_20),
    ._EVAL_21(coupler_to_bus_named_cbus__EVAL_21),
    ._EVAL_22(coupler_to_bus_named_cbus__EVAL_22),
    ._EVAL_23(coupler_to_bus_named_cbus__EVAL_23),
    ._EVAL_24(coupler_to_bus_named_cbus__EVAL_24),
    ._EVAL_25(coupler_to_bus_named_cbus__EVAL_25),
    ._EVAL_26(coupler_to_bus_named_cbus__EVAL_26),
    ._EVAL_27(coupler_to_bus_named_cbus__EVAL_27),
    ._EVAL_28(coupler_to_bus_named_cbus__EVAL_28),
    ._EVAL_29(coupler_to_bus_named_cbus__EVAL_29),
    ._EVAL_30(coupler_to_bus_named_cbus__EVAL_30),
    ._EVAL_31(coupler_to_bus_named_cbus__EVAL_31),
    ._EVAL_32(coupler_to_bus_named_cbus__EVAL_32),
    ._EVAL_33(coupler_to_bus_named_cbus__EVAL_33),
    ._EVAL_34(coupler_to_bus_named_cbus__EVAL_34),
    ._EVAL_35(coupler_to_bus_named_cbus__EVAL_35),
    ._EVAL_36(coupler_to_bus_named_cbus__EVAL_36),
    ._EVAL_37(coupler_to_bus_named_cbus__EVAL_37),
    ._EVAL_38(coupler_to_bus_named_cbus__EVAL_38),
    ._EVAL_39(coupler_to_bus_named_cbus__EVAL_39),
    ._EVAL_40(coupler_to_bus_named_cbus__EVAL_40)
  );
  SiFive__EVAL_2 system_bus_xbar (
    ._EVAL(system_bus_xbar__EVAL),
    ._EVAL_0(system_bus_xbar__EVAL_0),
    ._EVAL_1(system_bus_xbar__EVAL_1),
    ._EVAL_2(system_bus_xbar__EVAL_2),
    ._EVAL_3(system_bus_xbar__EVAL_3),
    ._EVAL_4(system_bus_xbar__EVAL_4),
    ._EVAL_5(system_bus_xbar__EVAL_5),
    ._EVAL_6(system_bus_xbar__EVAL_6),
    ._EVAL_7(system_bus_xbar__EVAL_7),
    ._EVAL_8(system_bus_xbar__EVAL_8),
    ._EVAL_9(system_bus_xbar__EVAL_9),
    ._EVAL_10(system_bus_xbar__EVAL_10),
    ._EVAL_11(system_bus_xbar__EVAL_11),
    ._EVAL_12(system_bus_xbar__EVAL_12),
    ._EVAL_13(system_bus_xbar__EVAL_13),
    ._EVAL_14(system_bus_xbar__EVAL_14),
    ._EVAL_15(system_bus_xbar__EVAL_15),
    ._EVAL_16(system_bus_xbar__EVAL_16),
    ._EVAL_17(system_bus_xbar__EVAL_17),
    ._EVAL_18(system_bus_xbar__EVAL_18),
    ._EVAL_19(system_bus_xbar__EVAL_19),
    ._EVAL_20(system_bus_xbar__EVAL_20),
    ._EVAL_21(system_bus_xbar__EVAL_21),
    ._EVAL_22(system_bus_xbar__EVAL_22),
    ._EVAL_23(system_bus_xbar__EVAL_23),
    ._EVAL_24(system_bus_xbar__EVAL_24),
    ._EVAL_25(system_bus_xbar__EVAL_25),
    ._EVAL_26(system_bus_xbar__EVAL_26),
    ._EVAL_27(system_bus_xbar__EVAL_27),
    ._EVAL_28(system_bus_xbar__EVAL_28),
    ._EVAL_29(system_bus_xbar__EVAL_29),
    ._EVAL_30(system_bus_xbar__EVAL_30),
    ._EVAL_31(system_bus_xbar__EVAL_31),
    ._EVAL_32(system_bus_xbar__EVAL_32),
    ._EVAL_33(system_bus_xbar__EVAL_33),
    ._EVAL_34(system_bus_xbar__EVAL_34),
    ._EVAL_35(system_bus_xbar__EVAL_35),
    ._EVAL_36(system_bus_xbar__EVAL_36),
    ._EVAL_37(system_bus_xbar__EVAL_37),
    ._EVAL_38(system_bus_xbar__EVAL_38),
    ._EVAL_39(system_bus_xbar__EVAL_39),
    ._EVAL_40(system_bus_xbar__EVAL_40),
    ._EVAL_41(system_bus_xbar__EVAL_41),
    ._EVAL_42(system_bus_xbar__EVAL_42),
    ._EVAL_43(system_bus_xbar__EVAL_43),
    ._EVAL_44(system_bus_xbar__EVAL_44),
    ._EVAL_45(system_bus_xbar__EVAL_45),
    ._EVAL_46(system_bus_xbar__EVAL_46),
    ._EVAL_47(system_bus_xbar__EVAL_47),
    ._EVAL_48(system_bus_xbar__EVAL_48),
    ._EVAL_49(system_bus_xbar__EVAL_49),
    ._EVAL_50(system_bus_xbar__EVAL_50),
    ._EVAL_51(system_bus_xbar__EVAL_51),
    ._EVAL_52(system_bus_xbar__EVAL_52),
    ._EVAL_53(system_bus_xbar__EVAL_53),
    ._EVAL_54(system_bus_xbar__EVAL_54),
    ._EVAL_55(system_bus_xbar__EVAL_55),
    ._EVAL_56(system_bus_xbar__EVAL_56),
    ._EVAL_57(system_bus_xbar__EVAL_57),
    ._EVAL_58(system_bus_xbar__EVAL_58),
    ._EVAL_59(system_bus_xbar__EVAL_59),
    ._EVAL_60(system_bus_xbar__EVAL_60),
    ._EVAL_61(system_bus_xbar__EVAL_61),
    ._EVAL_62(system_bus_xbar__EVAL_62),
    ._EVAL_63(system_bus_xbar__EVAL_63),
    ._EVAL_64(system_bus_xbar__EVAL_64),
    ._EVAL_65(system_bus_xbar__EVAL_65),
    ._EVAL_66(system_bus_xbar__EVAL_66),
    ._EVAL_67(system_bus_xbar__EVAL_67),
    ._EVAL_68(system_bus_xbar__EVAL_68),
    ._EVAL_69(system_bus_xbar__EVAL_69),
    ._EVAL_70(system_bus_xbar__EVAL_70),
    ._EVAL_71(system_bus_xbar__EVAL_71),
    ._EVAL_72(system_bus_xbar__EVAL_72),
    ._EVAL_73(system_bus_xbar__EVAL_73),
    ._EVAL_74(system_bus_xbar__EVAL_74),
    ._EVAL_75(system_bus_xbar__EVAL_75),
    ._EVAL_76(system_bus_xbar__EVAL_76),
    ._EVAL_77(system_bus_xbar__EVAL_77),
    ._EVAL_78(system_bus_xbar__EVAL_78),
    ._EVAL_79(system_bus_xbar__EVAL_79),
    ._EVAL_80(system_bus_xbar__EVAL_80),
    ._EVAL_81(system_bus_xbar__EVAL_81),
    ._EVAL_82(system_bus_xbar__EVAL_82),
    ._EVAL_83(system_bus_xbar__EVAL_83),
    ._EVAL_84(system_bus_xbar__EVAL_84),
    ._EVAL_85(system_bus_xbar__EVAL_85),
    ._EVAL_86(system_bus_xbar__EVAL_86),
    ._EVAL_87(system_bus_xbar__EVAL_87),
    ._EVAL_88(system_bus_xbar__EVAL_88),
    ._EVAL_89(system_bus_xbar__EVAL_89),
    ._EVAL_90(system_bus_xbar__EVAL_90),
    ._EVAL_91(system_bus_xbar__EVAL_91),
    ._EVAL_92(system_bus_xbar__EVAL_92),
    ._EVAL_93(system_bus_xbar__EVAL_93),
    ._EVAL_94(system_bus_xbar__EVAL_94),
    ._EVAL_95(system_bus_xbar__EVAL_95),
    ._EVAL_96(system_bus_xbar__EVAL_96),
    ._EVAL_97(system_bus_xbar__EVAL_97),
    ._EVAL_98(system_bus_xbar__EVAL_98),
    ._EVAL_99(system_bus_xbar__EVAL_99),
    ._EVAL_100(system_bus_xbar__EVAL_100),
    ._EVAL_101(system_bus_xbar__EVAL_101),
    ._EVAL_102(system_bus_xbar__EVAL_102),
    ._EVAL_103(system_bus_xbar__EVAL_103),
    ._EVAL_104(system_bus_xbar__EVAL_104),
    ._EVAL_105(system_bus_xbar__EVAL_105),
    ._EVAL_106(system_bus_xbar__EVAL_106),
    ._EVAL_107(system_bus_xbar__EVAL_107),
    ._EVAL_108(system_bus_xbar__EVAL_108),
    ._EVAL_109(system_bus_xbar__EVAL_109),
    ._EVAL_110(system_bus_xbar__EVAL_110),
    ._EVAL_111(system_bus_xbar__EVAL_111),
    ._EVAL_112(system_bus_xbar__EVAL_112),
    ._EVAL_113(system_bus_xbar__EVAL_113),
    ._EVAL_114(system_bus_xbar__EVAL_114),
    ._EVAL_115(system_bus_xbar__EVAL_115),
    ._EVAL_116(system_bus_xbar__EVAL_116),
    ._EVAL_117(system_bus_xbar__EVAL_117),
    ._EVAL_118(system_bus_xbar__EVAL_118),
    ._EVAL_119(system_bus_xbar__EVAL_119),
    ._EVAL_120(system_bus_xbar__EVAL_120),
    ._EVAL_121(system_bus_xbar__EVAL_121),
    ._EVAL_122(system_bus_xbar__EVAL_122),
    ._EVAL_123(system_bus_xbar__EVAL_123),
    ._EVAL_124(system_bus_xbar__EVAL_124),
    ._EVAL_125(system_bus_xbar__EVAL_125),
    ._EVAL_126(system_bus_xbar__EVAL_126),
    ._EVAL_127(system_bus_xbar__EVAL_127),
    ._EVAL_128(system_bus_xbar__EVAL_128)
  );
  SiFive__EVAL_18 coupler_from_tile_with_no_name (
    ._EVAL(coupler_from_tile_with_no_name__EVAL),
    ._EVAL_0(coupler_from_tile_with_no_name__EVAL_0),
    ._EVAL_1(coupler_from_tile_with_no_name__EVAL_1),
    ._EVAL_2(coupler_from_tile_with_no_name__EVAL_2),
    ._EVAL_3(coupler_from_tile_with_no_name__EVAL_3),
    ._EVAL_4(coupler_from_tile_with_no_name__EVAL_4),
    ._EVAL_5(coupler_from_tile_with_no_name__EVAL_5),
    ._EVAL_6(coupler_from_tile_with_no_name__EVAL_6),
    ._EVAL_7(coupler_from_tile_with_no_name__EVAL_7),
    ._EVAL_8(coupler_from_tile_with_no_name__EVAL_8),
    ._EVAL_9(coupler_from_tile_with_no_name__EVAL_9),
    ._EVAL_10(coupler_from_tile_with_no_name__EVAL_10),
    ._EVAL_11(coupler_from_tile_with_no_name__EVAL_11),
    ._EVAL_12(coupler_from_tile_with_no_name__EVAL_12),
    ._EVAL_13(coupler_from_tile_with_no_name__EVAL_13),
    ._EVAL_14(coupler_from_tile_with_no_name__EVAL_14),
    ._EVAL_15(coupler_from_tile_with_no_name__EVAL_15),
    ._EVAL_16(coupler_from_tile_with_no_name__EVAL_16),
    ._EVAL_17(coupler_from_tile_with_no_name__EVAL_17),
    ._EVAL_18(coupler_from_tile_with_no_name__EVAL_18),
    ._EVAL_19(coupler_from_tile_with_no_name__EVAL_19),
    ._EVAL_20(coupler_from_tile_with_no_name__EVAL_20),
    ._EVAL_21(coupler_from_tile_with_no_name__EVAL_21),
    ._EVAL_22(coupler_from_tile_with_no_name__EVAL_22),
    ._EVAL_23(coupler_from_tile_with_no_name__EVAL_23),
    ._EVAL_24(coupler_from_tile_with_no_name__EVAL_24),
    ._EVAL_25(coupler_from_tile_with_no_name__EVAL_25),
    ._EVAL_26(coupler_from_tile_with_no_name__EVAL_26),
    ._EVAL_27(coupler_from_tile_with_no_name__EVAL_27),
    ._EVAL_28(coupler_from_tile_with_no_name__EVAL_28),
    ._EVAL_29(coupler_from_tile_with_no_name__EVAL_29),
    ._EVAL_30(coupler_from_tile_with_no_name__EVAL_30),
    ._EVAL_31(coupler_from_tile_with_no_name__EVAL_31),
    ._EVAL_32(coupler_from_tile_with_no_name__EVAL_32),
    ._EVAL_33(coupler_from_tile_with_no_name__EVAL_33),
    ._EVAL_34(coupler_from_tile_with_no_name__EVAL_34),
    ._EVAL_35(coupler_from_tile_with_no_name__EVAL_35),
    ._EVAL_36(coupler_from_tile_with_no_name__EVAL_36),
    ._EVAL_37(coupler_from_tile_with_no_name__EVAL_37),
    ._EVAL_38(coupler_from_tile_with_no_name__EVAL_38),
    ._EVAL_39(coupler_from_tile_with_no_name__EVAL_39),
    ._EVAL_40(coupler_from_tile_with_no_name__EVAL_40),
    ._EVAL_41(coupler_from_tile_with_no_name__EVAL_41),
    ._EVAL_42(coupler_from_tile_with_no_name__EVAL_42),
    ._EVAL_43(coupler_from_tile_with_no_name__EVAL_43),
    ._EVAL_44(coupler_from_tile_with_no_name__EVAL_44),
    ._EVAL_45(coupler_from_tile_with_no_name__EVAL_45),
    ._EVAL_46(coupler_from_tile_with_no_name__EVAL_46),
    ._EVAL_47(coupler_from_tile_with_no_name__EVAL_47),
    ._EVAL_48(coupler_from_tile_with_no_name__EVAL_48),
    ._EVAL_49(coupler_from_tile_with_no_name__EVAL_49),
    ._EVAL_50(coupler_from_tile_with_no_name__EVAL_50),
    ._EVAL_51(coupler_from_tile_with_no_name__EVAL_51),
    ._EVAL_52(coupler_from_tile_with_no_name__EVAL_52),
    ._EVAL_53(coupler_from_tile_with_no_name__EVAL_53),
    ._EVAL_54(coupler_from_tile_with_no_name__EVAL_54),
    ._EVAL_55(coupler_from_tile_with_no_name__EVAL_55),
    ._EVAL_56(coupler_from_tile_with_no_name__EVAL_56),
    ._EVAL_57(coupler_from_tile_with_no_name__EVAL_57),
    ._EVAL_58(coupler_from_tile_with_no_name__EVAL_58),
    ._EVAL_59(coupler_from_tile_with_no_name__EVAL_59),
    ._EVAL_60(coupler_from_tile_with_no_name__EVAL_60),
    ._EVAL_61(coupler_from_tile_with_no_name__EVAL_61),
    ._EVAL_62(coupler_from_tile_with_no_name__EVAL_62),
    ._EVAL_63(coupler_from_tile_with_no_name__EVAL_63),
    ._EVAL_64(coupler_from_tile_with_no_name__EVAL_64),
    ._EVAL_65(coupler_from_tile_with_no_name__EVAL_65),
    ._EVAL_66(coupler_from_tile_with_no_name__EVAL_66),
    ._EVAL_67(coupler_from_tile_with_no_name__EVAL_67),
    ._EVAL_68(coupler_from_tile_with_no_name__EVAL_68),
    ._EVAL_69(coupler_from_tile_with_no_name__EVAL_69),
    ._EVAL_70(coupler_from_tile_with_no_name__EVAL_70),
    ._EVAL_71(coupler_from_tile_with_no_name__EVAL_71),
    ._EVAL_72(coupler_from_tile_with_no_name__EVAL_72),
    ._EVAL_73(coupler_from_tile_with_no_name__EVAL_73),
    ._EVAL_74(coupler_from_tile_with_no_name__EVAL_74),
    ._EVAL_75(coupler_from_tile_with_no_name__EVAL_75),
    ._EVAL_76(coupler_from_tile_with_no_name__EVAL_76),
    ._EVAL_77(coupler_from_tile_with_no_name__EVAL_77),
    ._EVAL_78(coupler_from_tile_with_no_name__EVAL_78),
    ._EVAL_79(coupler_from_tile_with_no_name__EVAL_79),
    ._EVAL_80(coupler_from_tile_with_no_name__EVAL_80),
    ._EVAL_81(coupler_from_tile_with_no_name__EVAL_81),
    ._EVAL_82(coupler_from_tile_with_no_name__EVAL_82),
    ._EVAL_83(coupler_from_tile_with_no_name__EVAL_83),
    ._EVAL_84(coupler_from_tile_with_no_name__EVAL_84),
    ._EVAL_85(coupler_from_tile_with_no_name__EVAL_85),
    ._EVAL_86(coupler_from_tile_with_no_name__EVAL_86),
    ._EVAL_87(coupler_from_tile_with_no_name__EVAL_87),
    ._EVAL_88(coupler_from_tile_with_no_name__EVAL_88),
    ._EVAL_89(coupler_from_tile_with_no_name__EVAL_89),
    ._EVAL_90(coupler_from_tile_with_no_name__EVAL_90),
    ._EVAL_91(coupler_from_tile_with_no_name__EVAL_91),
    ._EVAL_92(coupler_from_tile_with_no_name__EVAL_92),
    ._EVAL_93(coupler_from_tile_with_no_name__EVAL_93),
    ._EVAL_94(coupler_from_tile_with_no_name__EVAL_94),
    ._EVAL_95(coupler_from_tile_with_no_name__EVAL_95),
    ._EVAL_96(coupler_from_tile_with_no_name__EVAL_96),
    ._EVAL_97(coupler_from_tile_with_no_name__EVAL_97),
    ._EVAL_98(coupler_from_tile_with_no_name__EVAL_98),
    ._EVAL_99(coupler_from_tile_with_no_name__EVAL_99),
    ._EVAL_100(coupler_from_tile_with_no_name__EVAL_100),
    ._EVAL_101(coupler_from_tile_with_no_name__EVAL_101),
    ._EVAL_102(coupler_from_tile_with_no_name__EVAL_102),
    ._EVAL_103(coupler_from_tile_with_no_name__EVAL_103),
    ._EVAL_104(coupler_from_tile_with_no_name__EVAL_104),
    ._EVAL_105(coupler_from_tile_with_no_name__EVAL_105),
    ._EVAL_106(coupler_from_tile_with_no_name__EVAL_106),
    ._EVAL_107(coupler_from_tile_with_no_name__EVAL_107)
  );
  SiFive__EVAL_40 coupler_to_port_named_axi4_sys_port (
    ._EVAL(coupler_to_port_named_axi4_sys_port__EVAL),
    ._EVAL_0(coupler_to_port_named_axi4_sys_port__EVAL_0),
    ._EVAL_1(coupler_to_port_named_axi4_sys_port__EVAL_1),
    ._EVAL_2(coupler_to_port_named_axi4_sys_port__EVAL_2),
    ._EVAL_3(coupler_to_port_named_axi4_sys_port__EVAL_3),
    ._EVAL_4(coupler_to_port_named_axi4_sys_port__EVAL_4),
    ._EVAL_5(coupler_to_port_named_axi4_sys_port__EVAL_5),
    ._EVAL_6(coupler_to_port_named_axi4_sys_port__EVAL_6),
    ._EVAL_7(coupler_to_port_named_axi4_sys_port__EVAL_7),
    ._EVAL_8(coupler_to_port_named_axi4_sys_port__EVAL_8),
    ._EVAL_9(coupler_to_port_named_axi4_sys_port__EVAL_9),
    ._EVAL_10(coupler_to_port_named_axi4_sys_port__EVAL_10),
    ._EVAL_11(coupler_to_port_named_axi4_sys_port__EVAL_11),
    ._EVAL_12(coupler_to_port_named_axi4_sys_port__EVAL_12),
    ._EVAL_13(coupler_to_port_named_axi4_sys_port__EVAL_13),
    ._EVAL_14(coupler_to_port_named_axi4_sys_port__EVAL_14),
    ._EVAL_15(coupler_to_port_named_axi4_sys_port__EVAL_15),
    ._EVAL_16(coupler_to_port_named_axi4_sys_port__EVAL_16),
    ._EVAL_17(coupler_to_port_named_axi4_sys_port__EVAL_17),
    ._EVAL_18(coupler_to_port_named_axi4_sys_port__EVAL_18),
    ._EVAL_19(coupler_to_port_named_axi4_sys_port__EVAL_19),
    ._EVAL_20(coupler_to_port_named_axi4_sys_port__EVAL_20),
    ._EVAL_21(coupler_to_port_named_axi4_sys_port__EVAL_21),
    ._EVAL_22(coupler_to_port_named_axi4_sys_port__EVAL_22),
    ._EVAL_23(coupler_to_port_named_axi4_sys_port__EVAL_23),
    ._EVAL_24(coupler_to_port_named_axi4_sys_port__EVAL_24),
    ._EVAL_25(coupler_to_port_named_axi4_sys_port__EVAL_25),
    ._EVAL_26(coupler_to_port_named_axi4_sys_port__EVAL_26),
    ._EVAL_27(coupler_to_port_named_axi4_sys_port__EVAL_27),
    ._EVAL_28(coupler_to_port_named_axi4_sys_port__EVAL_28),
    ._EVAL_29(coupler_to_port_named_axi4_sys_port__EVAL_29),
    ._EVAL_30(coupler_to_port_named_axi4_sys_port__EVAL_30),
    ._EVAL_31(coupler_to_port_named_axi4_sys_port__EVAL_31),
    ._EVAL_32(coupler_to_port_named_axi4_sys_port__EVAL_32),
    ._EVAL_33(coupler_to_port_named_axi4_sys_port__EVAL_33),
    ._EVAL_34(coupler_to_port_named_axi4_sys_port__EVAL_34),
    ._EVAL_35(coupler_to_port_named_axi4_sys_port__EVAL_35),
    ._EVAL_36(coupler_to_port_named_axi4_sys_port__EVAL_36),
    ._EVAL_37(coupler_to_port_named_axi4_sys_port__EVAL_37),
    ._EVAL_38(coupler_to_port_named_axi4_sys_port__EVAL_38),
    ._EVAL_39(coupler_to_port_named_axi4_sys_port__EVAL_39),
    ._EVAL_40(coupler_to_port_named_axi4_sys_port__EVAL_40),
    ._EVAL_41(coupler_to_port_named_axi4_sys_port__EVAL_41),
    ._EVAL_42(coupler_to_port_named_axi4_sys_port__EVAL_42),
    ._EVAL_43(coupler_to_port_named_axi4_sys_port__EVAL_43),
    ._EVAL_44(coupler_to_port_named_axi4_sys_port__EVAL_44),
    ._EVAL_45(coupler_to_port_named_axi4_sys_port__EVAL_45),
    ._EVAL_46(coupler_to_port_named_axi4_sys_port__EVAL_46),
    ._EVAL_47(coupler_to_port_named_axi4_sys_port__EVAL_47),
    ._EVAL_48(coupler_to_port_named_axi4_sys_port__EVAL_48),
    ._EVAL_49(coupler_to_port_named_axi4_sys_port__EVAL_49),
    ._EVAL_50(coupler_to_port_named_axi4_sys_port__EVAL_50),
    ._EVAL_51(coupler_to_port_named_axi4_sys_port__EVAL_51),
    ._EVAL_52(coupler_to_port_named_axi4_sys_port__EVAL_52),
    ._EVAL_53(coupler_to_port_named_axi4_sys_port__EVAL_53),
    ._EVAL_54(coupler_to_port_named_axi4_sys_port__EVAL_54),
    ._EVAL_55(coupler_to_port_named_axi4_sys_port__EVAL_55)
  );
  SiFive__EVAL_48 coupler_from_bus_named_front_bus (
    ._EVAL(coupler_from_bus_named_front_bus__EVAL),
    ._EVAL_0(coupler_from_bus_named_front_bus__EVAL_0),
    ._EVAL_1(coupler_from_bus_named_front_bus__EVAL_1),
    ._EVAL_2(coupler_from_bus_named_front_bus__EVAL_2),
    ._EVAL_3(coupler_from_bus_named_front_bus__EVAL_3),
    ._EVAL_4(coupler_from_bus_named_front_bus__EVAL_4),
    ._EVAL_5(coupler_from_bus_named_front_bus__EVAL_5),
    ._EVAL_6(coupler_from_bus_named_front_bus__EVAL_6),
    ._EVAL_7(coupler_from_bus_named_front_bus__EVAL_7),
    ._EVAL_8(coupler_from_bus_named_front_bus__EVAL_8),
    ._EVAL_9(coupler_from_bus_named_front_bus__EVAL_9),
    ._EVAL_10(coupler_from_bus_named_front_bus__EVAL_10),
    ._EVAL_11(coupler_from_bus_named_front_bus__EVAL_11),
    ._EVAL_12(coupler_from_bus_named_front_bus__EVAL_12),
    ._EVAL_13(coupler_from_bus_named_front_bus__EVAL_13),
    ._EVAL_14(coupler_from_bus_named_front_bus__EVAL_14),
    ._EVAL_15(coupler_from_bus_named_front_bus__EVAL_15),
    ._EVAL_16(coupler_from_bus_named_front_bus__EVAL_16),
    ._EVAL_17(coupler_from_bus_named_front_bus__EVAL_17),
    ._EVAL_18(coupler_from_bus_named_front_bus__EVAL_18),
    ._EVAL_19(coupler_from_bus_named_front_bus__EVAL_19),
    ._EVAL_20(coupler_from_bus_named_front_bus__EVAL_20),
    ._EVAL_21(coupler_from_bus_named_front_bus__EVAL_21),
    ._EVAL_22(coupler_from_bus_named_front_bus__EVAL_22),
    ._EVAL_23(coupler_from_bus_named_front_bus__EVAL_23),
    ._EVAL_24(coupler_from_bus_named_front_bus__EVAL_24),
    ._EVAL_25(coupler_from_bus_named_front_bus__EVAL_25),
    ._EVAL_26(coupler_from_bus_named_front_bus__EVAL_26),
    ._EVAL_27(coupler_from_bus_named_front_bus__EVAL_27),
    ._EVAL_28(coupler_from_bus_named_front_bus__EVAL_28),
    ._EVAL_29(coupler_from_bus_named_front_bus__EVAL_29),
    ._EVAL_30(coupler_from_bus_named_front_bus__EVAL_30),
    ._EVAL_31(coupler_from_bus_named_front_bus__EVAL_31),
    ._EVAL_32(coupler_from_bus_named_front_bus__EVAL_32),
    ._EVAL_33(coupler_from_bus_named_front_bus__EVAL_33),
    ._EVAL_34(coupler_from_bus_named_front_bus__EVAL_34),
    ._EVAL_35(coupler_from_bus_named_front_bus__EVAL_35),
    ._EVAL_36(coupler_from_bus_named_front_bus__EVAL_36),
    ._EVAL_37(coupler_from_bus_named_front_bus__EVAL_37),
    ._EVAL_38(coupler_from_bus_named_front_bus__EVAL_38),
    ._EVAL_39(coupler_from_bus_named_front_bus__EVAL_39),
    ._EVAL_40(coupler_from_bus_named_front_bus__EVAL_40)
  );
  assign _EVAL_218 = coupler_to_port_named_axi4_sys_port__EVAL_48;
  assign coupler_to_port_named_axi4_sys_port__EVAL_31 = system_bus_xbar__EVAL_2;
  assign _EVAL_176 = coupler_from_tile_with_no_name__EVAL_61;
  assign _EVAL_177 = coupler_from_tile_with_no_name__EVAL_50;
  assign system_bus_xbar__EVAL_67 = coupler_from_tile_with_no_name__EVAL_59;
  assign _EVAL_96 = coupler_to_bus_named_cbus__EVAL_17;
  assign coupler_to_port_named_axi4_sys_port__EVAL_10 = _EVAL_98;
  assign coupler_from_bus_named_front_bus__EVAL_14 = system_bus_xbar__EVAL_66;
  assign _EVAL_160 = system_bus_xbar__EVAL_25;
  assign coupler_to_bus_named_cbus__EVAL_20 = _EVAL_62;
  assign system_bus_xbar__EVAL_84 = coupler_from_bus_named_front_bus__EVAL_37;
  assign system_bus_xbar__EVAL_101 = _EVAL_137;
  assign system_bus_xbar__EVAL_38 = coupler_from_tile_with_no_name__EVAL_74;
  assign _EVAL_32 = coupler_to_bus_named_cbus__EVAL_32;
  assign system_bus_xbar__EVAL_59 = _EVAL_1;
  assign _EVAL_167 = coupler_to_port_named_axi4_sys_port__EVAL_2;
  assign _EVAL_26 = coupler_to_bus_named_cbus__EVAL_37;
  assign system_bus_xbar__EVAL_99 = coupler_to_port_named_axi4_sys_port__EVAL_33;
  assign _EVAL_124 = coupler_from_tile_with_no_name__EVAL_3;
  assign coupler_from_bus_named_front_bus__EVAL_31 = _EVAL_27;
  assign system_bus_xbar__EVAL_118 = coupler_to_port_named_axi4_sys_port__EVAL_19;
  assign coupler_from_tile_with_no_name__EVAL_24 = _EVAL_40;
  assign coupler_from_tile_with_no_name__EVAL_40 = _EVAL_10;
  assign _EVAL_78 = system_bus_xbar__EVAL_58;
  assign _EVAL_64 = system_bus_xbar__EVAL_26;
  assign system_bus_xbar__EVAL_119 = coupler_from_tile_with_no_name__EVAL_51;
  assign coupler_to_bus_named_cbus__EVAL_21 = _EVAL_169;
  assign coupler_from_tile_with_no_name__EVAL_34 = _EVAL_191;
  assign coupler_from_tile_with_no_name__EVAL_0 = system_bus_xbar__EVAL_72;
  assign coupler_from_tile_with_no_name__EVAL_82 = _EVAL_144;
  assign _EVAL_33 = coupler_to_bus_named_cbus__EVAL_3;
  assign system_bus_xbar__EVAL_1 = coupler_from_tile_with_no_name__EVAL_67;
  assign _EVAL_61 = coupler_to_port_named_axi4_sys_port__EVAL_53;
  assign coupler_to_port_named_axi4_sys_port__EVAL_16 = _EVAL_31;
  assign system_bus_xbar__EVAL_77 = coupler_from_tile_with_no_name__EVAL_38;
  assign system_bus_xbar__EVAL_68 = _EVAL_45;
  assign system_bus_xbar__EVAL_56 = coupler_from_tile_with_no_name__EVAL_86;
  assign coupler_to_port_named_axi4_sys_port__EVAL_3 = _EVAL_149;
  assign system_bus_xbar__EVAL_122 = coupler_from_tile_with_no_name__EVAL_43;
  assign _EVAL_109 = coupler_to_port_named_axi4_sys_port__EVAL_49;
  assign _EVAL_216 = coupler_to_port_named_axi4_sys_port__EVAL_46;
  assign _EVAL_205 = coupler_from_bus_named_front_bus__EVAL_34;
  assign _EVAL_42 = coupler_to_port_named_axi4_sys_port__EVAL_36;
  assign coupler_from_tile_with_no_name__EVAL_25 = system_bus_xbar__EVAL_16;
  assign coupler_from_bus_named_front_bus__EVAL_23 = _EVAL_137;
  assign system_bus_xbar__EVAL_123 = coupler_to_port_named_axi4_sys_port__EVAL_32;
  assign coupler_from_tile_with_no_name__EVAL_55 = system_bus_xbar__EVAL_104;
  assign system_bus_xbar__EVAL_51 = _EVAL_159;
  assign coupler_from_bus_named_front_bus__EVAL_16 = system_bus_xbar__EVAL_65;
  assign _EVAL_152 = coupler_to_bus_named_cbus__EVAL_23;
  assign _EVAL_220 = coupler_from_tile_with_no_name__EVAL_96;
  assign _EVAL_217 = coupler_to_bus_named_cbus__EVAL_39;
  assign coupler_from_bus_named_front_bus__EVAL_35 = system_bus_xbar__EVAL_89;
  assign system_bus_xbar__EVAL_76 = coupler_from_tile_with_no_name__EVAL_89;
  assign system_bus_xbar__EVAL_127 = coupler_from_bus_named_front_bus__EVAL_0;
  assign _EVAL_215 = coupler_to_port_named_axi4_sys_port__EVAL_15;
  assign coupler_to_bus_named_cbus__EVAL_10 = _EVAL_90;
  assign _EVAL_81 = coupler_to_bus_named_cbus__EVAL_9;
  assign coupler_to_port_named_axi4_sys_port__EVAL_1 = system_bus_xbar__EVAL_105;
  assign coupler_from_tile_with_no_name__EVAL = _EVAL_120;
  assign coupler_to_port_named_axi4_sys_port__EVAL_50 = _EVAL_159;
  assign _EVAL_213 = coupler_from_tile_with_no_name__EVAL_48;
  assign coupler_from_tile_with_no_name__EVAL_95 = _EVAL_179;
  assign system_bus_xbar__EVAL_69 = coupler_from_tile_with_no_name__EVAL_6;
  assign coupler_from_tile_with_no_name__EVAL_23 = _EVAL_222;
  assign _EVAL_82 = coupler_to_port_named_axi4_sys_port__EVAL_54;
  assign _EVAL_58 = coupler_to_bus_named_cbus__EVAL_5;
  assign _EVAL_140 = system_bus_xbar__EVAL_37;
  assign _EVAL_181 = coupler_to_bus_named_cbus__EVAL_28;
  assign coupler_to_port_named_axi4_sys_port__EVAL_6 = system_bus_xbar__EVAL_87;
  assign coupler_from_bus_named_front_bus__EVAL_8 = _EVAL_76;
  assign system_bus_xbar__EVAL_42 = coupler_from_tile_with_no_name__EVAL_81;
  assign _EVAL_100 = coupler_from_tile_with_no_name__EVAL_80;
  assign _EVAL_121 = system_bus_xbar__EVAL_115;
  assign _EVAL_53 = coupler_from_bus_named_front_bus__EVAL_40;
  assign _EVAL_24 = coupler_from_tile_with_no_name__EVAL_28;
  assign coupler_to_bus_named_cbus__EVAL_8 = _EVAL_88;
  assign _EVAL_188 = coupler_from_bus_named_front_bus__EVAL_19;
  assign coupler_to_bus_named_cbus__EVAL_6 = _EVAL_186;
  assign _EVAL_156 = coupler_to_bus_named_cbus__EVAL_2;
  assign coupler_from_tile_with_no_name__EVAL_107 = system_bus_xbar__EVAL_81;
  assign _EVAL_129 = system_bus_xbar__EVAL_73;
  assign _EVAL_51 = coupler_from_tile_with_no_name__EVAL_58;
  assign _EVAL_141 = coupler_from_bus_named_front_bus__EVAL_21;
  assign system_bus_xbar__EVAL_45 = coupler_from_bus_named_front_bus__EVAL_26;
  assign coupler_from_tile_with_no_name__EVAL_98 = _EVAL_17;
  assign coupler_from_tile_with_no_name__EVAL_92 = _EVAL_70;
  assign system_bus_xbar__EVAL_20 = _EVAL_192;
  assign _EVAL_148 = system_bus_xbar__EVAL_10;
  assign _EVAL_171 = system_bus_xbar__EVAL_86;
  assign _EVAL_174 = coupler_from_tile_with_no_name__EVAL_66;
  assign coupler_from_tile_with_no_name__EVAL_12 = _EVAL_131;
  assign coupler_from_tile_with_no_name__EVAL_46 = _EVAL_189;
  assign system_bus_xbar__EVAL_100 = coupler_to_port_named_axi4_sys_port__EVAL_24;
  assign system_bus_xbar__EVAL_34 = coupler_to_port_named_axi4_sys_port__EVAL_28;
  assign coupler_to_port_named_axi4_sys_port__EVAL_14 = system_bus_xbar__EVAL_78;
  assign _EVAL_84 = coupler_from_bus_named_front_bus__EVAL_29;
  assign coupler_from_tile_with_no_name__EVAL_99 = _EVAL_21;
  assign system_bus_xbar__EVAL_47 = _EVAL_4;
  assign coupler_from_tile_with_no_name__EVAL_83 = system_bus_xbar__EVAL_64;
  assign _EVAL_200 = system_bus_xbar__EVAL_19;
  assign coupler_to_port_named_axi4_sys_port__EVAL_27 = system_bus_xbar__EVAL_0;
  assign _EVAL_193 = coupler_to_bus_named_cbus__EVAL_24;
  assign _EVAL_170 = coupler_to_bus_named_cbus__EVAL_7;
  assign coupler_to_port_named_axi4_sys_port__EVAL_12 = _EVAL_59;
  assign system_bus_xbar__EVAL_113 = _EVAL_126;
  assign _EVAL_68 = coupler_from_tile_with_no_name__EVAL_7;
  assign coupler_from_tile_with_no_name__EVAL_90 = _EVAL_110;
  assign coupler_from_tile_with_no_name__EVAL_65 = _EVAL_79;
  assign coupler_from_tile_with_no_name__EVAL_9 = system_bus_xbar__EVAL_28;
  assign coupler_from_tile_with_no_name__EVAL_19 = system_bus_xbar__EVAL_107;
  assign coupler_from_bus_named_front_bus__EVAL_17 = _EVAL_104;
  assign coupler_from_tile_with_no_name__EVAL_104 = _EVAL_41;
  assign system_bus_xbar__EVAL_60 = coupler_from_bus_named_front_bus__EVAL_25;
  assign coupler_to_bus_named_cbus__EVAL_29 = _EVAL_108;
  assign coupler_from_tile_with_no_name__EVAL_42 = _EVAL_85;
  assign coupler_from_tile_with_no_name__EVAL_4 = _EVAL_204;
  assign coupler_from_tile_with_no_name__EVAL_53 = _EVAL_97;
  assign system_bus_xbar__EVAL_61 = coupler_from_tile_with_no_name__EVAL_76;
  assign system_bus_xbar__EVAL_74 = _EVAL_114;
  assign _EVAL_92 = system_bus_xbar__EVAL_12;
  assign system_bus_xbar__EVAL_40 = coupler_from_tile_with_no_name__EVAL_39;
  assign coupler_from_bus_named_front_bus__EVAL_11 = system_bus_xbar__EVAL_109;
  assign system_bus_xbar__EVAL_117 = coupler_from_bus_named_front_bus__EVAL_27;
  assign system_bus_xbar__EVAL_32 = coupler_from_tile_with_no_name__EVAL_21;
  assign _EVAL_154 = system_bus_xbar__EVAL_120;
  assign _EVAL_22 = coupler_to_port_named_axi4_sys_port__EVAL_4;
  assign coupler_to_bus_named_cbus__EVAL_31 = _EVAL_153;
  assign coupler_from_tile_with_no_name__EVAL_97 = _EVAL_137;
  assign system_bus_xbar__EVAL_24 = _EVAL_178;
  assign _EVAL_111 = system_bus_xbar__EVAL_75;
  assign system_bus_xbar__EVAL_85 = _EVAL_116;
  assign system_bus_xbar__EVAL_71 = coupler_from_tile_with_no_name__EVAL_11;
  assign coupler_from_tile_with_no_name__EVAL_15 = _EVAL_168;
  assign coupler_from_tile_with_no_name__EVAL_106 = system_bus_xbar__EVAL_80;
  assign coupler_to_port_named_axi4_sys_port__EVAL_35 = system_bus_xbar__EVAL_46;
  assign _EVAL_9 = system_bus_xbar__EVAL_70;
  assign _EVAL_184 = coupler_from_tile_with_no_name__EVAL_72;
  assign _EVAL_71 = coupler_from_tile_with_no_name__EVAL_33;
  assign coupler_to_bus_named_cbus__EVAL_18 = _EVAL_190;
  assign coupler_from_tile_with_no_name__EVAL_2 = _EVAL_159;
  assign coupler_from_bus_named_front_bus__EVAL_5 = _EVAL_118;
  assign coupler_from_tile_with_no_name__EVAL_105 = _EVAL_210;
  assign _EVAL_12 = coupler_from_bus_named_front_bus__EVAL_4;
  assign _EVAL_223 = coupler_from_tile_with_no_name__EVAL_54;
  assign coupler_from_bus_named_front_bus__EVAL_13 = system_bus_xbar__EVAL_6;
  assign system_bus_xbar__EVAL_48 = coupler_to_port_named_axi4_sys_port__EVAL_8;
  assign coupler_to_bus_named_cbus__EVAL_19 = _EVAL_2;
  assign _EVAL = coupler_from_tile_with_no_name__EVAL_1;
  assign _EVAL_139 = coupler_to_bus_named_cbus__EVAL_33;
  assign coupler_from_bus_named_front_bus__EVAL_39 = _EVAL_44;
  assign coupler_from_bus_named_front_bus__EVAL_18 = _EVAL_173;
  assign _EVAL_219 = coupler_to_port_named_axi4_sys_port__EVAL_47;
  assign _EVAL_60 = coupler_to_bus_named_cbus__EVAL_12;
  assign system_bus_xbar__EVAL_13 = coupler_from_bus_named_front_bus__EVAL_33;
  assign coupler_from_bus_named_front_bus__EVAL = _EVAL_159;
  assign _EVAL_36 = coupler_to_port_named_axi4_sys_port__EVAL_20;
  assign _EVAL_18 = system_bus_xbar__EVAL_41;
  assign _EVAL_52 = coupler_to_port_named_axi4_sys_port__EVAL_0;
  assign coupler_to_bus_named_cbus__EVAL_0 = _EVAL_157;
  assign coupler_from_tile_with_no_name__EVAL_26 = system_bus_xbar__EVAL_111;
  assign coupler_from_tile_with_no_name__EVAL_45 = _EVAL_112;
  assign system_bus_xbar__EVAL_23 = _EVAL_101;
  assign system_bus_xbar__EVAL_39 = _EVAL_166;
  assign _EVAL_224 = coupler_to_port_named_axi4_sys_port__EVAL_42;
  assign coupler_from_bus_named_front_bus__EVAL_7 = _EVAL_194;
  assign _EVAL_208 = coupler_from_bus_named_front_bus__EVAL_3;
  assign coupler_from_tile_with_no_name__EVAL_71 = system_bus_xbar__EVAL_96;
  assign coupler_to_bus_named_cbus__EVAL_38 = _EVAL_137;
  assign system_bus_xbar__EVAL_49 = _EVAL_6;
  assign coupler_from_tile_with_no_name__EVAL_29 = system_bus_xbar__EVAL_128;
  assign _EVAL_155 = system_bus_xbar__EVAL_8;
  assign coupler_to_bus_named_cbus__EVAL_13 = _EVAL_69;
  assign coupler_from_tile_with_no_name__EVAL_75 = _EVAL_105;
  assign _EVAL_3 = system_bus_xbar__EVAL_18;
  assign _EVAL_180 = coupler_from_tile_with_no_name__EVAL_91;
  assign coupler_from_bus_named_front_bus__EVAL_15 = system_bus_xbar__EVAL_97;
  assign coupler_from_bus_named_front_bus__EVAL_38 = _EVAL_158;
  assign coupler_to_port_named_axi4_sys_port__EVAL_30 = _EVAL_66;
  assign _EVAL_201 = coupler_to_port_named_axi4_sys_port__EVAL_55;
  assign _EVAL_8 = coupler_to_port_named_axi4_sys_port__EVAL;
  assign _EVAL_94 = coupler_from_tile_with_no_name__EVAL_57;
  assign coupler_from_bus_named_front_bus__EVAL_28 = _EVAL_93;
  assign _EVAL_20 = coupler_to_bus_named_cbus__EVAL_35;
  assign _EVAL_55 = coupler_from_tile_with_no_name__EVAL_88;
  assign _EVAL_80 = system_bus_xbar__EVAL_4;
  assign coupler_from_tile_with_no_name__EVAL_13 = _EVAL_16;
  assign coupler_from_tile_with_no_name__EVAL_31 = _EVAL_127;
  assign coupler_to_port_named_axi4_sys_port__EVAL_25 = _EVAL_47;
  assign _EVAL_132 = coupler_from_bus_named_front_bus__EVAL_2;
  assign _EVAL_83 = coupler_from_tile_with_no_name__EVAL_56;
  assign coupler_from_tile_with_no_name__EVAL_18 = _EVAL_91;
  assign system_bus_xbar__EVAL_82 = coupler_from_tile_with_no_name__EVAL_22;
  assign coupler_from_tile_with_no_name__EVAL_32 = system_bus_xbar__EVAL_110;
  assign coupler_from_tile_with_no_name__EVAL_101 = system_bus_xbar__EVAL_27;
  assign coupler_from_tile_with_no_name__EVAL_36 = _EVAL_115;
  assign coupler_from_bus_named_front_bus__EVAL_10 = system_bus_xbar__EVAL_52;
  assign coupler_from_tile_with_no_name__EVAL_102 = _EVAL_197;
  assign system_bus_xbar__EVAL = coupler_to_port_named_axi4_sys_port__EVAL_9;
  assign _EVAL_214 = coupler_from_tile_with_no_name__EVAL_60;
  assign _EVAL_75 = coupler_to_port_named_axi4_sys_port__EVAL_40;
  assign system_bus_xbar__EVAL_36 = _EVAL_207;
  assign coupler_from_tile_with_no_name__EVAL_100 = system_bus_xbar__EVAL_63;
  assign _EVAL_77 = coupler_from_tile_with_no_name__EVAL_94;
  assign _EVAL_125 = system_bus_xbar__EVAL_55;
  assign _EVAL_65 = system_bus_xbar__EVAL_108;
  assign _EVAL_198 = coupler_from_tile_with_no_name__EVAL_52;
  assign coupler_from_tile_with_no_name__EVAL_8 = _EVAL_89;
  assign system_bus_xbar__EVAL_95 = _EVAL_182;
  assign _EVAL_49 = coupler_to_port_named_axi4_sys_port__EVAL_51;
  assign system_bus_xbar__EVAL_22 = _EVAL_130;
  assign coupler_from_bus_named_front_bus__EVAL_12 = system_bus_xbar__EVAL_7;
  assign _EVAL_107 = coupler_from_tile_with_no_name__EVAL_87;
  assign coupler_to_port_named_axi4_sys_port__EVAL_11 = _EVAL_134;
  assign coupler_to_port_named_axi4_sys_port__EVAL_34 = _EVAL_46;
  assign coupler_to_port_named_axi4_sys_port__EVAL_45 = system_bus_xbar__EVAL_93;
  assign system_bus_xbar__EVAL_112 = _EVAL_74;
  assign coupler_to_bus_named_cbus__EVAL_40 = _EVAL_37;
  assign system_bus_xbar__EVAL_33 = coupler_from_tile_with_no_name__EVAL_85;
  assign system_bus_xbar__EVAL_21 = coupler_to_port_named_axi4_sys_port__EVAL_22;
  assign system_bus_xbar__EVAL_43 = _EVAL_211;
  assign system_bus_xbar__EVAL_121 = coupler_from_bus_named_front_bus__EVAL_30;
  assign _EVAL_212 = system_bus_xbar__EVAL_29;
  assign coupler_from_tile_with_no_name__EVAL_68 = _EVAL_123;
  assign _EVAL_57 = coupler_to_bus_named_cbus__EVAL_11;
  assign coupler_from_tile_with_no_name__EVAL_35 = _EVAL_34;
  assign _EVAL_13 = coupler_from_tile_with_no_name__EVAL_73;
  assign coupler_from_tile_with_no_name__EVAL_5 = _EVAL_143;
  assign _EVAL_142 = coupler_to_port_named_axi4_sys_port__EVAL_43;
  assign coupler_to_port_named_axi4_sys_port__EVAL_39 = _EVAL_150;
  assign _EVAL_73 = system_bus_xbar__EVAL_94;
  assign system_bus_xbar__EVAL_83 = _EVAL_56;
  assign coupler_to_bus_named_cbus__EVAL_26 = _EVAL_67;
  assign coupler_to_bus_named_cbus__EVAL_25 = _EVAL_199;
  assign system_bus_xbar__EVAL_15 = coupler_from_bus_named_front_bus__EVAL_36;
  assign _EVAL_19 = coupler_from_tile_with_no_name__EVAL_37;
  assign _EVAL_195 = coupler_from_bus_named_front_bus__EVAL_32;
  assign system_bus_xbar__EVAL_31 = _EVAL_161;
  assign _EVAL_206 = coupler_from_tile_with_no_name__EVAL_93;
  assign system_bus_xbar__EVAL_62 = coupler_from_tile_with_no_name__EVAL_49;
  assign coupler_to_bus_named_cbus__EVAL_34 = _EVAL_128;
  assign system_bus_xbar__EVAL_54 = coupler_from_tile_with_no_name__EVAL_103;
  assign _EVAL_119 = coupler_to_bus_named_cbus__EVAL;
  assign _EVAL_146 = coupler_from_tile_with_no_name__EVAL_78;
  assign _EVAL_183 = coupler_to_bus_named_cbus__EVAL_36;
  assign coupler_to_port_named_axi4_sys_port__EVAL_21 = _EVAL_137;
  assign coupler_from_tile_with_no_name__EVAL_10 = _EVAL_0;
  assign coupler_from_tile_with_no_name__EVAL_14 = _EVAL_133;
  assign coupler_from_tile_with_no_name__EVAL_41 = _EVAL_145;
  assign coupler_from_tile_with_no_name__EVAL_63 = _EVAL_35;
  assign system_bus_xbar__EVAL_3 = coupler_from_bus_named_front_bus__EVAL_9;
  assign system_bus_xbar__EVAL_126 = _EVAL_5;
  assign system_bus_xbar__EVAL_90 = coupler_from_tile_with_no_name__EVAL_20;
  assign _EVAL_175 = coupler_to_port_named_axi4_sys_port__EVAL_18;
  assign _EVAL_23 = coupler_to_port_named_axi4_sys_port__EVAL_37;
  assign _EVAL_39 = system_bus_xbar__EVAL_17;
  assign system_bus_xbar__EVAL_11 = _EVAL_86;
  assign coupler_to_bus_named_cbus__EVAL_14 = _EVAL_135;
  assign _EVAL_87 = coupler_to_bus_named_cbus__EVAL_30;
  assign _EVAL_164 = coupler_from_tile_with_no_name__EVAL_17;
  assign _EVAL_117 = coupler_to_port_named_axi4_sys_port__EVAL_23;
  assign coupler_to_bus_named_cbus__EVAL_15 = _EVAL_203;
  assign _EVAL_63 = system_bus_xbar__EVAL_30;
  assign coupler_to_port_named_axi4_sys_port__EVAL_5 = system_bus_xbar__EVAL_14;
  assign coupler_to_port_named_axi4_sys_port__EVAL_7 = _EVAL_54;
  assign coupler_to_bus_named_cbus__EVAL_27 = _EVAL_159;
  assign _EVAL_15 = coupler_to_port_named_axi4_sys_port__EVAL_52;
  assign system_bus_xbar__EVAL_98 = _EVAL_28;
  assign coupler_to_port_named_axi4_sys_port__EVAL_44 = system_bus_xbar__EVAL_35;
  assign coupler_from_bus_named_front_bus__EVAL_24 = _EVAL_48;
  assign coupler_to_port_named_axi4_sys_port__EVAL_13 = _EVAL_138;
  assign _EVAL_38 = coupler_to_bus_named_cbus__EVAL_4;
  assign _EVAL_122 = coupler_to_port_named_axi4_sys_port__EVAL_26;
  assign coupler_to_bus_named_cbus__EVAL_16 = _EVAL_163;
  assign _EVAL_29 = system_bus_xbar__EVAL_102;
  assign coupler_to_bus_named_cbus__EVAL_1 = _EVAL_99;
  assign coupler_to_port_named_axi4_sys_port__EVAL_41 = system_bus_xbar__EVAL_116;
  assign coupler_from_tile_with_no_name__EVAL_84 = _EVAL_151;
  assign _EVAL_103 = system_bus_xbar__EVAL_106;
  assign coupler_from_tile_with_no_name__EVAL_70 = _EVAL_221;
  assign _EVAL_113 = coupler_from_tile_with_no_name__EVAL_16;
  assign _EVAL_25 = system_bus_xbar__EVAL_125;
  assign _EVAL_11 = system_bus_xbar__EVAL_53;
  assign coupler_from_tile_with_no_name__EVAL_44 = _EVAL_187;
  assign coupler_to_bus_named_cbus__EVAL_22 = _EVAL_50;
  assign coupler_from_bus_named_front_bus__EVAL_6 = system_bus_xbar__EVAL_44;
  assign _EVAL_162 = coupler_from_tile_with_no_name__EVAL_27;
  assign coupler_from_tile_with_no_name__EVAL_64 = _EVAL_7;
  assign _EVAL_147 = coupler_from_tile_with_no_name__EVAL_77;
  assign system_bus_xbar__EVAL_9 = coupler_from_tile_with_no_name__EVAL_79;
  assign _EVAL_165 = coupler_from_bus_named_front_bus__EVAL_20;
  assign _EVAL_136 = system_bus_xbar__EVAL_50;
  assign _EVAL_202 = system_bus_xbar__EVAL_92;
  assign _EVAL_30 = coupler_to_port_named_axi4_sys_port__EVAL_17;
  assign _EVAL_196 = coupler_to_port_named_axi4_sys_port__EVAL_38;
  assign _EVAL_185 = system_bus_xbar__EVAL_5;
  assign _EVAL_72 = coupler_to_port_named_axi4_sys_port__EVAL_29;
  assign system_bus_xbar__EVAL_124 = _EVAL_43;
  assign coupler_from_bus_named_front_bus__EVAL_22 = system_bus_xbar__EVAL_57;
  assign _EVAL_102 = system_bus_xbar__EVAL_88;
  assign coupler_from_tile_with_no_name__EVAL_69 = _EVAL_209;
  assign system_bus_xbar__EVAL_103 = coupler_from_tile_with_no_name__EVAL_47;
  assign system_bus_xbar__EVAL_91 = _EVAL_14;
  assign system_bus_xbar__EVAL_114 = _EVAL_172;
  assign coupler_from_tile_with_no_name__EVAL_30 = _EVAL_95;
  assign coupler_from_tile_with_no_name__EVAL_62 = _EVAL_106;
  assign system_bus_xbar__EVAL_79 = coupler_from_bus_named_front_bus__EVAL_1;
endmodule
