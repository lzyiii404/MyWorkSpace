//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_257(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  input  [29:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input  [29:0] _EVAL_15,
  input         _EVAL_16,
  input  [29:0] _EVAL_17,
  output        _EVAL_18,
  input  [29:0] _EVAL_19,
  input  [1:0]  _EVAL_20,
  input  [31:0] _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [31:0] _EVAL_24,
  input  [1:0]  _EVAL_25,
  input         _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [29:0] _EVAL_28,
  input  [31:0] _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [1:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input         _EVAL_34,
  input  [29:0] _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [31:0] _EVAL_38,
  input         _EVAL_39,
  input  [1:0]  _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  input  [4:0]  _EVAL_49,
  input  [29:0] _EVAL_50,
  input         _EVAL_51,
  output        _EVAL_52,
  input  [1:0]  _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input  [1:0]  _EVAL_56,
  input         _EVAL_57,
  output        _EVAL_58,
  input  [31:0] _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  input         _EVAL_62,
  input  [1:0]  _EVAL_63,
  output        _EVAL_64,
  input  [29:0] _EVAL_65,
  input  [31:0] _EVAL_66,
  input         _EVAL_67,
  output        _EVAL_68,
  output        _EVAL_69,
  input         _EVAL_70,
  input  [1:0]  _EVAL_71
);
  wire  pmp__EVAL;
  wire [31:0] pmp__EVAL_0;
  wire [29:0] pmp__EVAL_1;
  wire  pmp__EVAL_2;
  wire [31:0] pmp__EVAL_3;
  wire  pmp__EVAL_4;
  wire  pmp__EVAL_5;
  wire  pmp__EVAL_6;
  wire  pmp__EVAL_7;
  wire  pmp__EVAL_8;
  wire [1:0] pmp__EVAL_9;
  wire  pmp__EVAL_10;
  wire  pmp__EVAL_11;
  wire [31:0] pmp__EVAL_12;
  wire [29:0] pmp__EVAL_13;
  wire  pmp__EVAL_14;
  wire [31:0] pmp__EVAL_15;
  wire [31:0] pmp__EVAL_16;
  wire  pmp__EVAL_17;
  wire  pmp__EVAL_18;
  wire [31:0] pmp__EVAL_19;
  wire [29:0] pmp__EVAL_20;
  wire [1:0] pmp__EVAL_21;
  wire [29:0] pmp__EVAL_22;
  wire  pmp__EVAL_23;
  wire [1:0] pmp__EVAL_24;
  wire  pmp__EVAL_25;
  wire  pmp__EVAL_26;
  wire [29:0] pmp__EVAL_27;
  wire  pmp__EVAL_28;
  wire  pmp__EVAL_29;
  wire  pmp__EVAL_30;
  wire  pmp__EVAL_31;
  wire  pmp__EVAL_32;
  wire [1:0] pmp__EVAL_33;
  wire [1:0] pmp__EVAL_34;
  wire  pmp__EVAL_35;
  wire  pmp__EVAL_36;
  wire [31:0] pmp__EVAL_37;
  wire  pmp__EVAL_38;
  wire [1:0] pmp__EVAL_39;
  wire  pmp__EVAL_40;
  wire [1:0] pmp__EVAL_41;
  wire  pmp__EVAL_42;
  wire [29:0] pmp__EVAL_43;
  wire [1:0] pmp__EVAL_44;
  wire  pmp__EVAL_45;
  wire  pmp__EVAL_46;
  wire  pmp__EVAL_47;
  wire [29:0] pmp__EVAL_48;
  wire [31:0] pmp__EVAL_49;
  wire  pmp__EVAL_50;
  wire  pmp__EVAL_51;
  wire  pmp__EVAL_52;
  wire  pmp__EVAL_53;
  wire [1:0] pmp__EVAL_54;
  wire  pmp__EVAL_55;
  wire [31:0] pmp__EVAL_56;
  wire [29:0] pmp__EVAL_57;
  wire  pmp__EVAL_58;
  wire  pmp__EVAL_59;
  wire  pmp__EVAL_60;
  wire [19:0] _EVAL_78;
  wire [11:0] _EVAL_184;
  wire [31:0] _EVAL_153;
  wire [31:0] _EVAL_90;
  wire [31:0] _EVAL_257;
  wire  _EVAL_116;
  wire  _EVAL_178;
  wire  _EVAL_234;
  wire  _EVAL_92;
  wire  _EVAL_204;
  wire  _EVAL_243;
  wire  _EVAL_113;
  wire [31:0] _EVAL_223;
  wire [32:0] _EVAL_121;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_132;
  wire [32:0] _EVAL_226;
  wire [32:0] _EVAL_103;
  wire [32:0] _EVAL_161;
  wire  _EVAL_154;
  wire [31:0] _EVAL_254;
  wire [32:0] _EVAL_207;
  wire [32:0] _EVAL_114;
  wire [32:0] _EVAL_141;
  wire  _EVAL_152;
  wire  _EVAL_244;
  wire [31:0] _EVAL_227;
  wire [32:0] _EVAL_145;
  wire [32:0] _EVAL_239;
  wire [32:0] _EVAL_206;
  wire  _EVAL_238;
  wire  _EVAL_188;
  wire [32:0] _EVAL_137;
  wire [32:0] _EVAL_196;
  wire [32:0] _EVAL_255;
  wire  _EVAL_199;
  wire  _EVAL_105;
  wire [31:0] _EVAL_185;
  wire [32:0] _EVAL_86;
  wire [32:0] _EVAL_248;
  wire [32:0] _EVAL_171;
  wire  _EVAL_100;
  wire  _EVAL_148;
  wire [32:0] _EVAL_82;
  wire [32:0] _EVAL_117;
  wire  _EVAL_216;
  wire  _EVAL_225;
  wire [32:0] _EVAL_193;
  wire [32:0] _EVAL_101;
  wire [32:0] _EVAL_191;
  wire  _EVAL_176;
  wire  _EVAL_230;
  wire [31:0] _EVAL_218;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_129;
  wire  _EVAL_83;
  wire  _EVAL_98;
  wire [31:0] _EVAL_173;
  wire [32:0] _EVAL_135;
  wire [32:0] _EVAL_236;
  wire [32:0] _EVAL_138;
  wire  _EVAL_195;
  wire  _EVAL_157;
  wire [31:0] _EVAL_233;
  wire [32:0] _EVAL_134;
  wire [32:0] _EVAL_232;
  wire [32:0] _EVAL_237;
  wire  _EVAL_74;
  wire  _EVAL_253;
  wire [32:0] _EVAL_147;
  wire [32:0] _EVAL_136;
  wire  _EVAL_215;
  wire [31:0] _EVAL_213;
  wire [32:0] _EVAL_77;
  wire [32:0] _EVAL_242;
  wire [32:0] _EVAL_120;
  wire  _EVAL_179;
  wire  _EVAL_219;
  wire  _EVAL_130;
  wire  _EVAL_122;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_201;
  wire  _EVAL_115;
  wire  _EVAL_89;
  wire  _EVAL_142;
  wire [1:0] _EVAL_240;
  wire [15:0] _EVAL_210;
  wire [32:0] _EVAL_144;
  wire [32:0] _EVAL_107;
  wire  _EVAL_118;
  wire  _EVAL_169;
  wire [1:0] _EVAL_246;
  wire [15:0] _EVAL_84;
  wire [15:0] _EVAL_256;
  wire [15:0] _EVAL_245;
  wire [15:0] _EVAL_250;
  wire  _EVAL_94;
  wire  _EVAL_126;
  wire  _EVAL_241;
  wire  _EVAL_181;
  wire  _EVAL_192;
  wire  _EVAL_175;
  wire  _EVAL_251;
  wire  _EVAL_127;
  wire  _EVAL_231;
  wire  _EVAL_87;
  wire  _EVAL_96;
  wire  _EVAL_79;
  wire  _EVAL_158;
  wire  _EVAL_109;
  wire  _EVAL_91;
  wire  _EVAL_212;
  wire  _EVAL_221;
  wire  _EVAL_123;
  wire [3:0] _EVAL_177;
  wire [3:0] _EVAL_155;
  wire [31:0] _EVAL_143;
  wire [31:0] _EVAL_162;
  wire  _EVAL_76;
  wire [32:0] _EVAL_146;
  wire [32:0] _EVAL_72;
  wire  _EVAL_205;
  wire  _EVAL_228;
  wire  _EVAL_187;
  wire [32:0] _EVAL_108;
  wire [32:0] _EVAL_110;
  wire  _EVAL_168;
  wire  _EVAL_81;
  wire  _EVAL_220;
  wire  _EVAL_133;
  wire [1:0] _EVAL_166;
  wire [15:0] _EVAL_189;
  wire [15:0] _EVAL_249;
  wire  _EVAL_235;
  wire  _EVAL_252;
  wire [15:0] _EVAL_167;
  wire [15:0] _EVAL_131;
  wire [15:0] _EVAL_214;
  wire [2:0] _EVAL_73;
  wire  _EVAL_183;
  wire  _EVAL_222;
  wire  _EVAL_128;
  wire  _EVAL_97;
  wire  _EVAL_180;
  wire [1:0] _EVAL_202;
  wire [15:0] _EVAL_88;
  wire [15:0] _EVAL_174;
  wire [15:0] _EVAL_190;
  wire [15:0] _EVAL_165;
  wire [15:0] _EVAL_95;
  wire [15:0] _EVAL_217;
  wire [15:0] _EVAL_200;
  wire [15:0] _EVAL_198;
  wire [15:0] _EVAL_229;
  wire  _EVAL_194;
  wire [15:0] _EVAL_164;
  wire [15:0] _EVAL_182;
  wire  _EVAL_160;
  wire [1:0] _EVAL_112;
  wire [15:0] _EVAL_247;
  wire [15:0] _EVAL_125;
  wire [15:0] _EVAL_102;
  wire [15:0] _EVAL_203;
  wire [15:0] _EVAL_208;
  wire [15:0] _EVAL_106;
  wire [15:0] _EVAL_75;
  wire  _EVAL_211;
  wire  _EVAL_224;
  wire  _EVAL_80;
  wire  _EVAL_209;
  wire [15:0] _EVAL_139;
  wire [15:0] _EVAL_151;
  wire [15:0] _EVAL_140;
  wire [15:0] _EVAL_156;
  wire [15:0] _EVAL_197;
  wire [15:0] _EVAL_93;
  wire [15:0] _EVAL_170;
  wire [19:0] _EVAL_111;
  wire  _EVAL_149;
  wire [15:0] _EVAL_186;
  wire [15:0] _EVAL_159;
  wire [15:0] _EVAL_85;
  wire [15:0] _EVAL_119;
  wire [15:0] _EVAL_99;
  SiFive__EVAL_256 pmp (
    ._EVAL(pmp__EVAL),
    ._EVAL_0(pmp__EVAL_0),
    ._EVAL_1(pmp__EVAL_1),
    ._EVAL_2(pmp__EVAL_2),
    ._EVAL_3(pmp__EVAL_3),
    ._EVAL_4(pmp__EVAL_4),
    ._EVAL_5(pmp__EVAL_5),
    ._EVAL_6(pmp__EVAL_6),
    ._EVAL_7(pmp__EVAL_7),
    ._EVAL_8(pmp__EVAL_8),
    ._EVAL_9(pmp__EVAL_9),
    ._EVAL_10(pmp__EVAL_10),
    ._EVAL_11(pmp__EVAL_11),
    ._EVAL_12(pmp__EVAL_12),
    ._EVAL_13(pmp__EVAL_13),
    ._EVAL_14(pmp__EVAL_14),
    ._EVAL_15(pmp__EVAL_15),
    ._EVAL_16(pmp__EVAL_16),
    ._EVAL_17(pmp__EVAL_17),
    ._EVAL_18(pmp__EVAL_18),
    ._EVAL_19(pmp__EVAL_19),
    ._EVAL_20(pmp__EVAL_20),
    ._EVAL_21(pmp__EVAL_21),
    ._EVAL_22(pmp__EVAL_22),
    ._EVAL_23(pmp__EVAL_23),
    ._EVAL_24(pmp__EVAL_24),
    ._EVAL_25(pmp__EVAL_25),
    ._EVAL_26(pmp__EVAL_26),
    ._EVAL_27(pmp__EVAL_27),
    ._EVAL_28(pmp__EVAL_28),
    ._EVAL_29(pmp__EVAL_29),
    ._EVAL_30(pmp__EVAL_30),
    ._EVAL_31(pmp__EVAL_31),
    ._EVAL_32(pmp__EVAL_32),
    ._EVAL_33(pmp__EVAL_33),
    ._EVAL_34(pmp__EVAL_34),
    ._EVAL_35(pmp__EVAL_35),
    ._EVAL_36(pmp__EVAL_36),
    ._EVAL_37(pmp__EVAL_37),
    ._EVAL_38(pmp__EVAL_38),
    ._EVAL_39(pmp__EVAL_39),
    ._EVAL_40(pmp__EVAL_40),
    ._EVAL_41(pmp__EVAL_41),
    ._EVAL_42(pmp__EVAL_42),
    ._EVAL_43(pmp__EVAL_43),
    ._EVAL_44(pmp__EVAL_44),
    ._EVAL_45(pmp__EVAL_45),
    ._EVAL_46(pmp__EVAL_46),
    ._EVAL_47(pmp__EVAL_47),
    ._EVAL_48(pmp__EVAL_48),
    ._EVAL_49(pmp__EVAL_49),
    ._EVAL_50(pmp__EVAL_50),
    ._EVAL_51(pmp__EVAL_51),
    ._EVAL_52(pmp__EVAL_52),
    ._EVAL_53(pmp__EVAL_53),
    ._EVAL_54(pmp__EVAL_54),
    ._EVAL_55(pmp__EVAL_55),
    ._EVAL_56(pmp__EVAL_56),
    ._EVAL_57(pmp__EVAL_57),
    ._EVAL_58(pmp__EVAL_58),
    ._EVAL_59(pmp__EVAL_59),
    ._EVAL_60(pmp__EVAL_60)
  );
  assign _EVAL_78 = _EVAL_29[31:12];
  assign _EVAL_184 = _EVAL_29[11:0];
  assign _EVAL_153 = {_EVAL_78,_EVAL_184};
  assign _EVAL_90 = _EVAL_153 ^ 32'h3000;
  assign _EVAL_257 = _EVAL_153 ^ 32'h1900000;
  assign _EVAL_116 = _EVAL_49 == 5'h4;
  assign _EVAL_178 = _EVAL_49 == 5'h9;
  assign _EVAL_234 = _EVAL_116 | _EVAL_178;
  assign _EVAL_92 = _EVAL_49 == 5'ha;
  assign _EVAL_204 = _EVAL_234 | _EVAL_92;
  assign _EVAL_243 = _EVAL_49 == 5'hb;
  assign _EVAL_113 = _EVAL_204 | _EVAL_243;
  assign _EVAL_223 = _EVAL_153 ^ 32'h2000000;
  assign _EVAL_121 = {1'b0,$signed(_EVAL_223)};
  assign _EVAL_163 = $signed(_EVAL_121) & $signed(33'sheb000000);
  assign _EVAL_132 = $signed(_EVAL_163);
  assign _EVAL_226 = {1'b0,$signed(_EVAL_257)};
  assign _EVAL_103 = $signed(_EVAL_226) & $signed(-33'sh2000);
  assign _EVAL_161 = $signed(_EVAL_103);
  assign _EVAL_154 = $signed(_EVAL_161) == $signed(33'sh0);
  assign _EVAL_254 = _EVAL_153 ^ 32'h40000000;
  assign _EVAL_207 = {1'b0,$signed(_EVAL_254)};
  assign _EVAL_114 = $signed(_EVAL_207) & $signed(-33'sh2000);
  assign _EVAL_141 = $signed(_EVAL_114);
  assign _EVAL_152 = $signed(_EVAL_141) == $signed(33'sh0);
  assign _EVAL_244 = _EVAL_154 | _EVAL_152;
  assign _EVAL_227 = _EVAL_153 ^ 32'h80000000;
  assign _EVAL_145 = {1'b0,$signed(_EVAL_227)};
  assign _EVAL_239 = $signed(_EVAL_145) & $signed(-33'sh20000);
  assign _EVAL_206 = $signed(_EVAL_239);
  assign _EVAL_238 = $signed(_EVAL_206) == $signed(33'sh0);
  assign _EVAL_188 = _EVAL_244 | _EVAL_238;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_90)};
  assign _EVAL_196 = $signed(_EVAL_137) & $signed(-33'sh1000);
  assign _EVAL_255 = $signed(_EVAL_196);
  assign _EVAL_199 = $signed(_EVAL_255) == $signed(33'sh0);
  assign _EVAL_105 = _EVAL_188 | _EVAL_199;
  assign _EVAL_185 = _EVAL_153 ^ 32'hc000000;
  assign _EVAL_86 = {1'b0,$signed(_EVAL_185)};
  assign _EVAL_248 = $signed(_EVAL_86) & $signed(-33'sh4000000);
  assign _EVAL_171 = $signed(_EVAL_248);
  assign _EVAL_100 = $signed(_EVAL_171) == $signed(33'sh0);
  assign _EVAL_148 = _EVAL_105 | _EVAL_100;
  assign _EVAL_82 = $signed(_EVAL_121) & $signed(-33'sh10000);
  assign _EVAL_117 = $signed(_EVAL_82);
  assign _EVAL_216 = $signed(_EVAL_117) == $signed(33'sh0);
  assign _EVAL_225 = _EVAL_148 | _EVAL_216;
  assign _EVAL_193 = {1'b0,$signed(_EVAL_153)};
  assign _EVAL_101 = $signed(_EVAL_193) & $signed(-33'sh1000);
  assign _EVAL_191 = $signed(_EVAL_101);
  assign _EVAL_176 = $signed(_EVAL_191) == $signed(33'sh0);
  assign _EVAL_230 = _EVAL_225 | _EVAL_176;
  assign _EVAL_218 = _EVAL_153 ^ 32'h1800000;
  assign _EVAL_104 = {1'b0,$signed(_EVAL_218)};
  assign _EVAL_172 = $signed(_EVAL_104) & $signed(-33'sh8000);
  assign _EVAL_129 = $signed(_EVAL_172);
  assign _EVAL_83 = $signed(_EVAL_129) == $signed(33'sh0);
  assign _EVAL_98 = _EVAL_230 | _EVAL_83;
  assign _EVAL_173 = _EVAL_153 ^ 32'h4000;
  assign _EVAL_135 = {1'b0,$signed(_EVAL_173)};
  assign _EVAL_236 = $signed(_EVAL_135) & $signed(-33'sh1000);
  assign _EVAL_138 = $signed(_EVAL_236);
  assign _EVAL_195 = $signed(_EVAL_138) == $signed(33'sh0);
  assign _EVAL_157 = _EVAL_98 | _EVAL_195;
  assign _EVAL_233 = _EVAL_153 ^ 32'h20000000;
  assign _EVAL_134 = {1'b0,$signed(_EVAL_233)};
  assign _EVAL_232 = $signed(_EVAL_134) & $signed(-33'sh2000);
  assign _EVAL_237 = $signed(_EVAL_232);
  assign _EVAL_74 = $signed(_EVAL_237) == $signed(33'sh0);
  assign _EVAL_253 = _EVAL_157 | _EVAL_74;
  assign _EVAL_147 = $signed(_EVAL_193) & $signed(33'shea000000);
  assign _EVAL_136 = $signed(_EVAL_147);
  assign _EVAL_215 = $signed(_EVAL_136) == $signed(33'sh0);
  assign _EVAL_213 = _EVAL_153 ^ 32'h8000000;
  assign _EVAL_77 = {1'b0,$signed(_EVAL_213)};
  assign _EVAL_242 = $signed(_EVAL_77) & $signed(33'she8000000);
  assign _EVAL_120 = $signed(_EVAL_242);
  assign _EVAL_179 = $signed(_EVAL_120) == $signed(33'sh0);
  assign _EVAL_219 = _EVAL_215 | _EVAL_179;
  assign _EVAL_130 = $signed(_EVAL_132) == $signed(33'sh0);
  assign _EVAL_122 = _EVAL_219 | _EVAL_130;
  assign _EVAL_150 = $signed(_EVAL_134) & $signed(33'sheb000000);
  assign _EVAL_201 = $signed(_EVAL_150);
  assign _EVAL_115 = $signed(_EVAL_201) == $signed(33'sh0);
  assign _EVAL_89 = _EVAL_122 | _EVAL_115;
  assign _EVAL_142 = _EVAL_253 & _EVAL_89;
  assign _EVAL_240 = _EVAL_142 ? 2'h3 : 2'h0;
  assign _EVAL_210 = {_EVAL_240,14'h0};
  assign _EVAL_144 = $signed(_EVAL_145) & $signed(33'sh80000000);
  assign _EVAL_107 = $signed(_EVAL_144);
  assign _EVAL_118 = $signed(_EVAL_107) == $signed(33'sh0);
  assign _EVAL_169 = _EVAL_253 & _EVAL_118;
  assign _EVAL_246 = _EVAL_169 ? 2'h3 : 2'h0;
  assign _EVAL_84 = {_EVAL_246,14'h0};
  assign _EVAL_256 = _EVAL_210 | _EVAL_84;
  assign _EVAL_245 = ~ _EVAL_256;
  assign _EVAL_250 = _EVAL_113 ? _EVAL_245 : 16'h0;
  assign _EVAL_94 = _EVAL_49 == 5'he;
  assign _EVAL_126 = _EVAL_49 == 5'h1;
  assign _EVAL_241 = _EVAL_49 == 5'h11;
  assign _EVAL_181 = _EVAL_126 | _EVAL_241;
  assign _EVAL_192 = _EVAL_49 == 5'h7;
  assign _EVAL_175 = _EVAL_181 | _EVAL_192;
  assign _EVAL_251 = _EVAL_49 == 5'h8;
  assign _EVAL_127 = _EVAL_49 == 5'hc;
  assign _EVAL_231 = _EVAL_251 | _EVAL_127;
  assign _EVAL_87 = _EVAL_49 == 5'hd;
  assign _EVAL_96 = _EVAL_231 | _EVAL_87;
  assign _EVAL_79 = _EVAL_96 | _EVAL_94;
  assign _EVAL_158 = _EVAL_49 == 5'hf;
  assign _EVAL_109 = _EVAL_79 | _EVAL_158;
  assign _EVAL_91 = _EVAL_113 | _EVAL_109;
  assign _EVAL_212 = _EVAL_175 | _EVAL_91;
  assign _EVAL_221 = _EVAL_49 == 5'h5;
  assign _EVAL_123 = _EVAL_212 | _EVAL_221;
  assign _EVAL_177 = 4'h1 << _EVAL_2;
  assign _EVAL_155 = _EVAL_177 - 4'h1;
  assign _EVAL_143 = {{28'd0}, _EVAL_155};
  assign _EVAL_162 = _EVAL_29 & _EVAL_143;
  assign _EVAL_76 = _EVAL_162 != 32'h0;
  assign _EVAL_146 = $signed(_EVAL_207) & $signed(33'sheb000000);
  assign _EVAL_72 = $signed(_EVAL_146);
  assign _EVAL_205 = $signed(_EVAL_72) == $signed(33'sh0);
  assign _EVAL_228 = _EVAL_205 | _EVAL_179;
  assign _EVAL_187 = _EVAL_228 | _EVAL_130;
  assign _EVAL_108 = $signed(_EVAL_193) & $signed(33'sheb001000);
  assign _EVAL_110 = $signed(_EVAL_108);
  assign _EVAL_168 = $signed(_EVAL_110) == $signed(33'sh0);
  assign _EVAL_81 = _EVAL_187 | _EVAL_168;
  assign _EVAL_220 = _EVAL_81 | _EVAL_115;
  assign _EVAL_133 = _EVAL_253 & _EVAL_220;
  assign _EVAL_166 = _EVAL_133 ? 2'h3 : 2'h0;
  assign _EVAL_189 = {_EVAL_166,14'h0};
  assign _EVAL_249 = _EVAL_76 ? _EVAL_189 : 16'h0;
  assign _EVAL_235 = _EVAL_49 == 5'h6;
  assign _EVAL_252 = _EVAL_235 | _EVAL_192;
  assign _EVAL_167 = ~ _EVAL_84;
  assign _EVAL_131 = _EVAL_252 ? _EVAL_167 : 16'h0;
  assign _EVAL_214 = _EVAL_249 | _EVAL_131;
  assign _EVAL_73 = {_EVAL_39,_EVAL_32};
  assign _EVAL_183 = _EVAL_73 <= 3'h3;
  assign _EVAL_222 = _EVAL_183 & _EVAL_176;
  assign _EVAL_128 = _EVAL_222 == 1'h0;
  assign _EVAL_97 = _EVAL_253 & _EVAL_128;
  assign _EVAL_180 = _EVAL_97 & pmp__EVAL_42;
  assign _EVAL_202 = _EVAL_180 ? 2'h3 : 2'h0;
  assign _EVAL_88 = {_EVAL_202,14'h0};
  assign _EVAL_174 = ~ _EVAL_88;
  assign _EVAL_190 = _EVAL_214 | _EVAL_174;
  assign _EVAL_165 = _EVAL_123 ? _EVAL_190 : 16'h0;
  assign _EVAL_95 = _EVAL_165 | _EVAL_250;
  assign _EVAL_217 = ~ _EVAL_210;
  assign _EVAL_200 = _EVAL_113 ? _EVAL_217 : 16'h0;
  assign _EVAL_198 = _EVAL_109 ? _EVAL_217 : 16'h0;
  assign _EVAL_229 = _EVAL_200 | _EVAL_198;
  assign _EVAL_194 = _EVAL_76 & _EVAL_212;
  assign _EVAL_164 = ~ _EVAL_189;
  assign _EVAL_182 = _EVAL_194 ? _EVAL_164 : 16'h0;
  assign _EVAL_160 = _EVAL_97 & pmp__EVAL_6;
  assign _EVAL_112 = _EVAL_160 ? 2'h3 : 2'h0;
  assign _EVAL_247 = {_EVAL_112,14'h0};
  assign _EVAL_125 = _EVAL_84 & 16'h8000;
  assign _EVAL_102 = _EVAL_109 ? _EVAL_245 : 16'h0;
  assign _EVAL_203 = _EVAL_95 | _EVAL_102;
  assign _EVAL_208 = _EVAL_252 ? 16'hffff : 16'h0;
  assign _EVAL_106 = _EVAL_229 | _EVAL_208;
  assign _EVAL_75 = ~ _EVAL_247;
  assign _EVAL_211 = _EVAL_49 == 5'h0;
  assign _EVAL_224 = _EVAL_211 | _EVAL_235;
  assign _EVAL_80 = _EVAL_224 | _EVAL_192;
  assign _EVAL_209 = _EVAL_80 | _EVAL_91;
  assign _EVAL_139 = _EVAL_214 | _EVAL_75;
  assign _EVAL_151 = _EVAL_209 ? _EVAL_139 : 16'h0;
  assign _EVAL_140 = _EVAL_151 & 16'h8000;
  assign _EVAL_156 = _EVAL_123 ? 16'h7fff : 16'h0;
  assign _EVAL_197 = _EVAL_156 & 16'h8000;
  assign _EVAL_93 = _EVAL_209 ? 16'h7fff : 16'h0;
  assign _EVAL_170 = _EVAL_93 & 16'h8000;
  assign _EVAL_111 = _EVAL_29[31:12];
  assign _EVAL_149 = _EVAL_76 & _EVAL_209;
  assign _EVAL_186 = _EVAL_149 ? _EVAL_164 : 16'h0;
  assign _EVAL_159 = _EVAL_203 & 16'h8000;
  assign _EVAL_85 = _EVAL_182 & 16'h8000;
  assign _EVAL_119 = _EVAL_106 & 16'h8000;
  assign _EVAL_99 = _EVAL_186 & 16'h8000;
  assign pmp__EVAL_50 = _EVAL_46;
  assign pmp__EVAL_45 = _EVAL_67;
  assign pmp__EVAL_11 = _EVAL_55;
  assign pmp__EVAL_12 = _EVAL_33;
  assign pmp__EVAL_21 = _EVAL_53;
  assign pmp__EVAL_0 = _EVAL_24;
  assign pmp__EVAL_1 = _EVAL_28;
  assign pmp__EVAL_9 = _EVAL_20;
  assign pmp__EVAL_41 = _EVAL_40;
  assign pmp__EVAL_56 = {_EVAL_78,_EVAL_184};
  assign pmp__EVAL_26 = _EVAL_43;
  assign pmp__EVAL_7 = _EVAL_57;
  assign _EVAL_58 = _EVAL_197 != 16'h0;
  assign pmp__EVAL = _EVAL_1;
  assign pmp__EVAL_33 = _EVAL_73[1:0];
  assign pmp__EVAL_49 = _EVAL_3;
  assign pmp__EVAL_10 = _EVAL_45;
  assign pmp__EVAL_27 = _EVAL_35;
  assign pmp__EVAL_19 = _EVAL_27;
  assign pmp__EVAL_28 = _EVAL_10;
  assign pmp__EVAL_48 = _EVAL_17;
  assign pmp__EVAL_14 = _EVAL_48;
  assign pmp__EVAL_37 = _EVAL_66;
  assign pmp__EVAL_13 = _EVAL_19;
  assign pmp__EVAL_51 = _EVAL_44;
  assign pmp__EVAL_39 = _EVAL_63;
  assign pmp__EVAL_4 = _EVAL_31;
  assign pmp__EVAL_38 = _EVAL_8;
  assign pmp__EVAL_23 = _EVAL_62;
  assign pmp__EVAL_20 = _EVAL_65;
  assign pmp__EVAL_57 = _EVAL_50;
  assign pmp__EVAL_16 = _EVAL_13;
  assign pmp__EVAL_53 = _EVAL_47;
  assign pmp__EVAL_59 = _EVAL_14;
  assign _EVAL_68 = _EVAL_125 != 16'h0;
  assign pmp__EVAL_32 = _EVAL_30;
  assign _EVAL_9 = _EVAL_99 != 16'h0;
  assign pmp__EVAL_25 = _EVAL_70;
  assign pmp__EVAL_55 = _EVAL;
  assign _EVAL_18 = _EVAL_159 != 16'h0;
  assign pmp__EVAL_47 = _EVAL_16;
  assign pmp__EVAL_46 = _EVAL_42;
  assign pmp__EVAL_30 = _EVAL_37;
  assign pmp__EVAL_31 = _EVAL_11;
  assign pmp__EVAL_22 = _EVAL_4;
  assign pmp__EVAL_3 = _EVAL_59;
  assign pmp__EVAL_2 = _EVAL_61;
  assign pmp__EVAL_15 = _EVAL_21;
  assign _EVAL_52 = _EVAL_170 != 16'h0;
  assign pmp__EVAL_60 = _EVAL_54;
  assign pmp__EVAL_43 = _EVAL_15;
  assign pmp__EVAL_44 = _EVAL_25;
  assign pmp__EVAL_40 = _EVAL_6;
  assign _EVAL_38 = {_EVAL_111,_EVAL_184};
  assign pmp__EVAL_29 = _EVAL_26;
  assign pmp__EVAL_8 = _EVAL_7;
  assign pmp__EVAL_17 = _EVAL_34;
  assign pmp__EVAL_5 = _EVAL_0;
  assign pmp__EVAL_58 = _EVAL_36;
  assign _EVAL_23 = _EVAL_119 != 16'h0;
  assign pmp__EVAL_52 = _EVAL_22;
  assign pmp__EVAL_35 = _EVAL_51;
  assign _EVAL_64 = _EVAL_85 != 16'h0;
  assign pmp__EVAL_54 = _EVAL_12;
  assign pmp__EVAL_36 = _EVAL_5;
  assign pmp__EVAL_18 = _EVAL_60;
  assign pmp__EVAL_34 = _EVAL_56;
  assign pmp__EVAL_24 = _EVAL_71;
  assign _EVAL_69 = _EVAL_140 != 16'h0;
endmodule
