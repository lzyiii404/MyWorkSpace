//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_254(
  output [63:0] _EVAL,
  input         _EVAL_0,
  output [63:0] _EVAL_1,
  input  [3:0]  _EVAL_2,
  input         _EVAL_3,
  input  [11:0] _EVAL_4,
  output [63:0] _EVAL_5,
  input  [3:0]  _EVAL_6,
  output [63:0] _EVAL_7,
  input  [63:0] _EVAL_8,
  input  [1:0]  _EVAL_9,
  input         _EVAL_10
);
  wire [7:0] data_arrays_0__EVAL;
  wire [7:0] data_arrays_0__EVAL_0;
  wire [7:0] data_arrays_0__EVAL_1;
  wire  data_arrays_0__EVAL_2;
  wire [7:0] data_arrays_0__EVAL_3;
  wire  data_arrays_0__EVAL_4;
  wire  data_arrays_0__EVAL_5;
  wire [7:0] data_arrays_0__EVAL_6;
  wire  data_arrays_0__EVAL_7;
  wire [7:0] data_arrays_0__EVAL_8;
  wire  data_arrays_0__EVAL_9;
  wire [7:0] data_arrays_0__EVAL_10;
  wire [8:0] data_arrays_0__EVAL_11;
  wire [7:0] data_arrays_0__EVAL_12;
  wire  data_arrays_0__EVAL_13;
  wire [7:0] data_arrays_0__EVAL_14;
  wire [7:0] data_arrays_0__EVAL_15;
  wire  data_arrays_0__EVAL_16;
  wire [7:0] data_arrays_0__EVAL_17;
  wire  data_arrays_0__EVAL_18;
  wire [7:0] data_arrays_0__EVAL_19;
  wire [7:0] data_arrays_0__EVAL_20;
  wire [7:0] data_arrays_0__EVAL_21;
  wire  data_arrays_0__EVAL_22;
  wire  data_arrays_0__EVAL_23;
  wire [7:0] data_arrays_0__EVAL_24;
  wire  data_arrays_0__EVAL_25;
  wire [7:0] data_arrays_0__EVAL_26;
  wire [7:0] data_arrays_0__EVAL_27;
  wire [7:0] data_arrays_0__EVAL_28;
  wire [7:0] data_arrays_0__EVAL_29;
  wire  data_arrays_0__EVAL_30;
  wire [7:0] data_arrays_0__EVAL_31;
  wire [7:0] data_arrays_0__EVAL_32;
  wire [7:0] data_arrays_0__EVAL_33;
  wire [7:0] data_arrays_0__EVAL_34;
  wire [7:0] data_arrays_0__EVAL_35;
  wire  data_arrays_0__EVAL_36;
  wire [7:0] data_arrays_0__EVAL_37;
  wire [7:0] data_arrays_0__EVAL_38;
  wire [7:0] data_arrays_0__EVAL_39;
  wire [7:0] data_arrays_0__EVAL_40;
  wire  data_arrays_0__EVAL_41;
  wire [7:0] data_arrays_0__EVAL_42;
  wire  data_arrays_0__EVAL_43;
  wire [7:0] data_arrays_0__EVAL_44;
  wire  data_arrays_0__EVAL_45;
  wire  data_arrays_0__EVAL_46;
  wire [7:0] data_arrays_0__EVAL_47;
  wire [7:0] data_arrays_0__EVAL_48;
  wire  data_arrays_0__EVAL_49;
  wire  data_arrays_0__EVAL_50;
  wire [7:0] data_arrays_1__EVAL;
  wire [7:0] data_arrays_1__EVAL_0;
  wire [7:0] data_arrays_1__EVAL_1;
  wire  data_arrays_1__EVAL_2;
  wire [7:0] data_arrays_1__EVAL_3;
  wire  data_arrays_1__EVAL_4;
  wire  data_arrays_1__EVAL_5;
  wire [7:0] data_arrays_1__EVAL_6;
  wire  data_arrays_1__EVAL_7;
  wire [7:0] data_arrays_1__EVAL_8;
  wire  data_arrays_1__EVAL_9;
  wire [7:0] data_arrays_1__EVAL_10;
  wire [8:0] data_arrays_1__EVAL_11;
  wire [7:0] data_arrays_1__EVAL_12;
  wire  data_arrays_1__EVAL_13;
  wire [7:0] data_arrays_1__EVAL_14;
  wire [7:0] data_arrays_1__EVAL_15;
  wire  data_arrays_1__EVAL_16;
  wire [7:0] data_arrays_1__EVAL_17;
  wire  data_arrays_1__EVAL_18;
  wire [7:0] data_arrays_1__EVAL_19;
  wire [7:0] data_arrays_1__EVAL_20;
  wire [7:0] data_arrays_1__EVAL_21;
  wire  data_arrays_1__EVAL_22;
  wire  data_arrays_1__EVAL_23;
  wire [7:0] data_arrays_1__EVAL_24;
  wire  data_arrays_1__EVAL_25;
  wire [7:0] data_arrays_1__EVAL_26;
  wire [7:0] data_arrays_1__EVAL_27;
  wire [7:0] data_arrays_1__EVAL_28;
  wire [7:0] data_arrays_1__EVAL_29;
  wire  data_arrays_1__EVAL_30;
  wire [7:0] data_arrays_1__EVAL_31;
  wire [7:0] data_arrays_1__EVAL_32;
  wire [7:0] data_arrays_1__EVAL_33;
  wire [7:0] data_arrays_1__EVAL_34;
  wire [7:0] data_arrays_1__EVAL_35;
  wire  data_arrays_1__EVAL_36;
  wire [7:0] data_arrays_1__EVAL_37;
  wire [7:0] data_arrays_1__EVAL_38;
  wire [7:0] data_arrays_1__EVAL_39;
  wire [7:0] data_arrays_1__EVAL_40;
  wire  data_arrays_1__EVAL_41;
  wire [7:0] data_arrays_1__EVAL_42;
  wire  data_arrays_1__EVAL_43;
  wire [7:0] data_arrays_1__EVAL_44;
  wire  data_arrays_1__EVAL_45;
  wire  data_arrays_1__EVAL_46;
  wire [7:0] data_arrays_1__EVAL_47;
  wire [7:0] data_arrays_1__EVAL_48;
  wire  data_arrays_1__EVAL_49;
  wire  data_arrays_1__EVAL_50;
  wire  _EVAL_35;
  wire [31:0] _EVAL_22;
  wire  _EVAL_24;
  wire  _EVAL_11;
  wire [31:0] _EVAL_36;
  wire [31:0] _EVAL_30;
  wire [31:0] _EVAL_12;
  wire  _EVAL_18;
  wire  _EVAL_29;
  wire  _EVAL_25;
  wire  _EVAL_27;
  wire [31:0] _EVAL_23;
  wire  _EVAL_26;
  wire  _EVAL_28;
  wire  _EVAL_34;
  wire  _EVAL_17;
  wire  _EVAL_31;
  wire  _EVAL_15;
  wire  _EVAL_32;
  wire [31:0] _EVAL_33;
  wire  _EVAL_37;
  wire [31:0] _EVAL_14;
  wire [31:0] _EVAL_19;
  wire [31:0] _EVAL_20;
  wire  _EVAL_16;
  wire [31:0] _EVAL_21;
  wire  _EVAL_13;
  SiFive__EVAL_343 data_arrays_0 (
    ._EVAL(data_arrays_0__EVAL),
    ._EVAL_0(data_arrays_0__EVAL_0),
    ._EVAL_1(data_arrays_0__EVAL_1),
    ._EVAL_2(data_arrays_0__EVAL_2),
    ._EVAL_3(data_arrays_0__EVAL_3),
    ._EVAL_4(data_arrays_0__EVAL_4),
    ._EVAL_5(data_arrays_0__EVAL_5),
    ._EVAL_6(data_arrays_0__EVAL_6),
    ._EVAL_7(data_arrays_0__EVAL_7),
    ._EVAL_8(data_arrays_0__EVAL_8),
    ._EVAL_9(data_arrays_0__EVAL_9),
    ._EVAL_10(data_arrays_0__EVAL_10),
    ._EVAL_11(data_arrays_0__EVAL_11),
    ._EVAL_12(data_arrays_0__EVAL_12),
    ._EVAL_13(data_arrays_0__EVAL_13),
    ._EVAL_14(data_arrays_0__EVAL_14),
    ._EVAL_15(data_arrays_0__EVAL_15),
    ._EVAL_16(data_arrays_0__EVAL_16),
    ._EVAL_17(data_arrays_0__EVAL_17),
    ._EVAL_18(data_arrays_0__EVAL_18),
    ._EVAL_19(data_arrays_0__EVAL_19),
    ._EVAL_20(data_arrays_0__EVAL_20),
    ._EVAL_21(data_arrays_0__EVAL_21),
    ._EVAL_22(data_arrays_0__EVAL_22),
    ._EVAL_23(data_arrays_0__EVAL_23),
    ._EVAL_24(data_arrays_0__EVAL_24),
    ._EVAL_25(data_arrays_0__EVAL_25),
    ._EVAL_26(data_arrays_0__EVAL_26),
    ._EVAL_27(data_arrays_0__EVAL_27),
    ._EVAL_28(data_arrays_0__EVAL_28),
    ._EVAL_29(data_arrays_0__EVAL_29),
    ._EVAL_30(data_arrays_0__EVAL_30),
    ._EVAL_31(data_arrays_0__EVAL_31),
    ._EVAL_32(data_arrays_0__EVAL_32),
    ._EVAL_33(data_arrays_0__EVAL_33),
    ._EVAL_34(data_arrays_0__EVAL_34),
    ._EVAL_35(data_arrays_0__EVAL_35),
    ._EVAL_36(data_arrays_0__EVAL_36),
    ._EVAL_37(data_arrays_0__EVAL_37),
    ._EVAL_38(data_arrays_0__EVAL_38),
    ._EVAL_39(data_arrays_0__EVAL_39),
    ._EVAL_40(data_arrays_0__EVAL_40),
    ._EVAL_41(data_arrays_0__EVAL_41),
    ._EVAL_42(data_arrays_0__EVAL_42),
    ._EVAL_43(data_arrays_0__EVAL_43),
    ._EVAL_44(data_arrays_0__EVAL_44),
    ._EVAL_45(data_arrays_0__EVAL_45),
    ._EVAL_46(data_arrays_0__EVAL_46),
    ._EVAL_47(data_arrays_0__EVAL_47),
    ._EVAL_48(data_arrays_0__EVAL_48),
    ._EVAL_49(data_arrays_0__EVAL_49),
    ._EVAL_50(data_arrays_0__EVAL_50)
  );
  SiFive__EVAL_343 data_arrays_1 (
    ._EVAL(data_arrays_1__EVAL),
    ._EVAL_0(data_arrays_1__EVAL_0),
    ._EVAL_1(data_arrays_1__EVAL_1),
    ._EVAL_2(data_arrays_1__EVAL_2),
    ._EVAL_3(data_arrays_1__EVAL_3),
    ._EVAL_4(data_arrays_1__EVAL_4),
    ._EVAL_5(data_arrays_1__EVAL_5),
    ._EVAL_6(data_arrays_1__EVAL_6),
    ._EVAL_7(data_arrays_1__EVAL_7),
    ._EVAL_8(data_arrays_1__EVAL_8),
    ._EVAL_9(data_arrays_1__EVAL_9),
    ._EVAL_10(data_arrays_1__EVAL_10),
    ._EVAL_11(data_arrays_1__EVAL_11),
    ._EVAL_12(data_arrays_1__EVAL_12),
    ._EVAL_13(data_arrays_1__EVAL_13),
    ._EVAL_14(data_arrays_1__EVAL_14),
    ._EVAL_15(data_arrays_1__EVAL_15),
    ._EVAL_16(data_arrays_1__EVAL_16),
    ._EVAL_17(data_arrays_1__EVAL_17),
    ._EVAL_18(data_arrays_1__EVAL_18),
    ._EVAL_19(data_arrays_1__EVAL_19),
    ._EVAL_20(data_arrays_1__EVAL_20),
    ._EVAL_21(data_arrays_1__EVAL_21),
    ._EVAL_22(data_arrays_1__EVAL_22),
    ._EVAL_23(data_arrays_1__EVAL_23),
    ._EVAL_24(data_arrays_1__EVAL_24),
    ._EVAL_25(data_arrays_1__EVAL_25),
    ._EVAL_26(data_arrays_1__EVAL_26),
    ._EVAL_27(data_arrays_1__EVAL_27),
    ._EVAL_28(data_arrays_1__EVAL_28),
    ._EVAL_29(data_arrays_1__EVAL_29),
    ._EVAL_30(data_arrays_1__EVAL_30),
    ._EVAL_31(data_arrays_1__EVAL_31),
    ._EVAL_32(data_arrays_1__EVAL_32),
    ._EVAL_33(data_arrays_1__EVAL_33),
    ._EVAL_34(data_arrays_1__EVAL_34),
    ._EVAL_35(data_arrays_1__EVAL_35),
    ._EVAL_36(data_arrays_1__EVAL_36),
    ._EVAL_37(data_arrays_1__EVAL_37),
    ._EVAL_38(data_arrays_1__EVAL_38),
    ._EVAL_39(data_arrays_1__EVAL_39),
    ._EVAL_40(data_arrays_1__EVAL_40),
    ._EVAL_41(data_arrays_1__EVAL_41),
    ._EVAL_42(data_arrays_1__EVAL_42),
    ._EVAL_43(data_arrays_1__EVAL_43),
    ._EVAL_44(data_arrays_1__EVAL_44),
    ._EVAL_45(data_arrays_1__EVAL_45),
    ._EVAL_46(data_arrays_1__EVAL_46),
    ._EVAL_47(data_arrays_1__EVAL_47),
    ._EVAL_48(data_arrays_1__EVAL_48),
    ._EVAL_49(data_arrays_1__EVAL_49),
    ._EVAL_50(data_arrays_1__EVAL_50)
  );
  assign _EVAL_35 = _EVAL_6[3];
  assign _EVAL_22 = _EVAL_8[63:32];
  assign _EVAL_24 = _EVAL_2[0];
  assign _EVAL_11 = _EVAL_6[1];
  assign _EVAL_36 = {data_arrays_1__EVAL_21,data_arrays_1__EVAL_39,data_arrays_1__EVAL_35,data_arrays_1__EVAL_14};
  assign _EVAL_30 = {data_arrays_0__EVAL_1,data_arrays_0__EVAL_37,data_arrays_0__EVAL_48,data_arrays_0__EVAL_33};
  assign _EVAL_12 = {data_arrays_1__EVAL_26,data_arrays_1__EVAL_17,data_arrays_1__EVAL_42,data_arrays_1__EVAL_15};
  assign _EVAL_18 = _EVAL_9[1];
  assign _EVAL_29 = _EVAL_9[0];
  assign _EVAL_25 = _EVAL_3 & _EVAL_29;
  assign _EVAL_27 = _EVAL_25 & _EVAL_10;
  assign _EVAL_23 = {data_arrays_0__EVAL_38,data_arrays_0__EVAL_0,data_arrays_0__EVAL_20,data_arrays_0__EVAL};
  assign _EVAL_26 = _EVAL_10 == 1'h0;
  assign _EVAL_28 = _EVAL_25 & _EVAL_26;
  assign _EVAL_34 = _EVAL_3 & _EVAL_18;
  assign _EVAL_17 = _EVAL_34 & _EVAL_26;
  assign _EVAL_31 = _EVAL_34 & _EVAL_10;
  assign _EVAL_15 = _EVAL_2[1];
  assign _EVAL_32 = _EVAL_6[0];
  assign _EVAL_33 = {data_arrays_0__EVAL_26,data_arrays_0__EVAL_17,data_arrays_0__EVAL_42,data_arrays_0__EVAL_15};
  assign _EVAL_37 = _EVAL_6[2];
  assign _EVAL_14 = {data_arrays_1__EVAL_38,data_arrays_1__EVAL_0,data_arrays_1__EVAL_20,data_arrays_1__EVAL};
  assign _EVAL_19 = _EVAL_8[31:0];
  assign _EVAL_20 = {data_arrays_1__EVAL_1,data_arrays_1__EVAL_37,data_arrays_1__EVAL_48,data_arrays_1__EVAL_33};
  assign _EVAL_16 = _EVAL_2[2];
  assign _EVAL_21 = {data_arrays_0__EVAL_21,data_arrays_0__EVAL_39,data_arrays_0__EVAL_35,data_arrays_0__EVAL_14};
  assign _EVAL_13 = _EVAL_2[3];
  assign data_arrays_1__EVAL_5 = _EVAL_24 & _EVAL_11;
  assign data_arrays_0__EVAL_18 = _EVAL_0;
  assign data_arrays_1__EVAL_41 = _EVAL_24 & _EVAL_35;
  assign data_arrays_0__EVAL_46 = _EVAL_28 | _EVAL_27;
  assign data_arrays_0__EVAL_9 = _EVAL_16 & _EVAL_37;
  assign data_arrays_1__EVAL_7 = _EVAL_10;
  assign data_arrays_0__EVAL_5 = _EVAL_24 & _EVAL_11;
  assign data_arrays_0__EVAL_27 = _EVAL_19[7:0];
  assign data_arrays_1__EVAL_43 = _EVAL_13 & _EVAL_35;
  assign data_arrays_1__EVAL_10 = _EVAL_22[7:0];
  assign data_arrays_1__EVAL_47 = _EVAL_22[31:24];
  assign data_arrays_1__EVAL_50 = _EVAL_15 & _EVAL_37;
  assign data_arrays_0__EVAL_12 = _EVAL_19[23:16];
  assign data_arrays_0__EVAL_10 = _EVAL_19[7:0];
  assign data_arrays_0__EVAL_50 = _EVAL_15 & _EVAL_37;
  assign data_arrays_1__EVAL_29 = _EVAL_22[31:24];
  assign data_arrays_1__EVAL_22 = _EVAL_24 & _EVAL_32;
  assign data_arrays_0__EVAL_32 = _EVAL_19[23:16];
  assign data_arrays_0__EVAL_31 = _EVAL_19[31:24];
  assign data_arrays_1__EVAL_40 = _EVAL_22[23:16];
  assign data_arrays_0__EVAL_44 = _EVAL_19[15:8];
  assign data_arrays_1__EVAL_45 = _EVAL_13 & _EVAL_37;
  assign data_arrays_1__EVAL_46 = _EVAL_17 | _EVAL_31;
  assign data_arrays_1__EVAL_18 = _EVAL_0;
  assign data_arrays_0__EVAL_19 = _EVAL_19[15:8];
  assign data_arrays_0__EVAL_24 = _EVAL_19[15:8];
  assign data_arrays_0__EVAL_3 = _EVAL_19[7:0];
  assign data_arrays_0__EVAL_4 = _EVAL_16 & _EVAL_35;
  assign data_arrays_1__EVAL_44 = _EVAL_22[15:8];
  assign data_arrays_1__EVAL_11 = _EVAL_4[11:3];
  assign data_arrays_1__EVAL_31 = _EVAL_22[31:24];
  assign data_arrays_0__EVAL_6 = _EVAL_19[23:16];
  assign data_arrays_0__EVAL_34 = _EVAL_19[7:0];
  assign data_arrays_0__EVAL_36 = _EVAL_16 & _EVAL_11;
  assign data_arrays_0__EVAL_41 = _EVAL_24 & _EVAL_35;
  assign data_arrays_0__EVAL_13 = _EVAL_24 & _EVAL_37;
  assign data_arrays_0__EVAL_16 = _EVAL_13 & _EVAL_32;
  assign data_arrays_1__EVAL_49 = _EVAL_16 & _EVAL_32;
  assign data_arrays_0__EVAL_43 = _EVAL_13 & _EVAL_35;
  assign data_arrays_0__EVAL_29 = _EVAL_19[31:24];
  assign _EVAL_5 = {_EVAL_36,_EVAL_21};
  assign data_arrays_1__EVAL_30 = _EVAL_13 & _EVAL_11;
  assign data_arrays_1__EVAL_32 = _EVAL_22[23:16];
  assign data_arrays_0__EVAL_23 = _EVAL_15 & _EVAL_11;
  assign _EVAL_1 = {_EVAL_20,_EVAL_30};
  assign data_arrays_1__EVAL_23 = _EVAL_15 & _EVAL_11;
  assign data_arrays_0__EVAL_30 = _EVAL_13 & _EVAL_11;
  assign data_arrays_0__EVAL_25 = _EVAL_15 & _EVAL_35;
  assign data_arrays_1__EVAL_4 = _EVAL_16 & _EVAL_35;
  assign data_arrays_1__EVAL_16 = _EVAL_13 & _EVAL_32;
  assign data_arrays_1__EVAL_24 = _EVAL_22[15:8];
  assign data_arrays_1__EVAL_13 = _EVAL_24 & _EVAL_37;
  assign data_arrays_1__EVAL_9 = _EVAL_16 & _EVAL_37;
  assign data_arrays_0__EVAL_40 = _EVAL_19[23:16];
  assign data_arrays_1__EVAL_19 = _EVAL_22[15:8];
  assign data_arrays_0__EVAL_11 = _EVAL_4[11:3];
  assign data_arrays_1__EVAL_36 = _EVAL_16 & _EVAL_11;
  assign _EVAL_7 = {_EVAL_14,_EVAL_23};
  assign data_arrays_0__EVAL_28 = _EVAL_19[31:24];
  assign data_arrays_1__EVAL_25 = _EVAL_15 & _EVAL_35;
  assign data_arrays_1__EVAL_3 = _EVAL_22[7:0];
  assign data_arrays_1__EVAL_28 = _EVAL_22[31:24];
  assign data_arrays_0__EVAL_22 = _EVAL_24 & _EVAL_32;
  assign data_arrays_0__EVAL_7 = _EVAL_10;
  assign data_arrays_0__EVAL_8 = _EVAL_19[15:8];
  assign data_arrays_1__EVAL_34 = _EVAL_22[7:0];
  assign data_arrays_0__EVAL_47 = _EVAL_19[31:24];
  assign data_arrays_1__EVAL_6 = _EVAL_22[23:16];
  assign _EVAL = {_EVAL_12,_EVAL_33};
  assign data_arrays_1__EVAL_27 = _EVAL_22[7:0];
  assign data_arrays_0__EVAL_2 = _EVAL_15 & _EVAL_32;
  assign data_arrays_0__EVAL_49 = _EVAL_16 & _EVAL_32;
  assign data_arrays_1__EVAL_2 = _EVAL_15 & _EVAL_32;
  assign data_arrays_1__EVAL_8 = _EVAL_22[15:8];
  assign data_arrays_1__EVAL_12 = _EVAL_22[23:16];
  assign data_arrays_0__EVAL_45 = _EVAL_13 & _EVAL_37;
endmodule
