//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_95(
  output [3:0]  _EVAL,
  output        _EVAL_0,
  input  [1:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  output [2:0]  _EVAL_3,
  output [1:0]  _EVAL_4,
  output [4:0]  _EVAL_5,
  output        _EVAL_6,
  input  [4:0]  _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input  [4:0]  _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output [3:0]  _EVAL_13,
  input         _EVAL_14,
  output [1:0]  _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output [2:0]  _EVAL_18,
  output [3:0]  _EVAL_19,
  input         _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [4:0]  _EVAL_22,
  output [3:0]  _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output [3:0]  _EVAL_26,
  input         _EVAL_27,
  input  [7:0]  _EVAL_28,
  input  [7:0]  _EVAL_29,
  output [7:0]  _EVAL_30,
  output [63:0] _EVAL_31,
  input         _EVAL_32,
  output [7:0]  _EVAL_33,
  input  [3:0]  _EVAL_34,
  output        _EVAL_35,
  output        _EVAL_36,
  input  [1:0]  _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  output [3:0]  _EVAL_40,
  input  [7:0]  _EVAL_41,
  output [31:0] _EVAL_42,
  output        _EVAL_43,
  input  [3:0]  _EVAL_44,
  input  [3:0]  _EVAL_45,
  input         _EVAL_46,
  input  [31:0] _EVAL_47,
  output [1:0]  _EVAL_48,
  input  [1:0]  _EVAL_49,
  input  [3:0]  _EVAL_50,
  input         _EVAL_51,
  input  [3:0]  _EVAL_52,
  output        _EVAL_53,
  input  [2:0]  _EVAL_54,
  input  [31:0] _EVAL_55,
  input         _EVAL_56,
  input  [63:0] _EVAL_57,
  input  [3:0]  _EVAL_58,
  output [2:0]  _EVAL_59,
  input  [63:0] _EVAL_60,
  input  [1:0]  _EVAL_61,
  output [31:0] _EVAL_62,
  output [63:0] _EVAL_63,
  input         _EVAL_64,
  output [7:0]  _EVAL_65,
  input  [4:0]  _EVAL_66,
  input         _EVAL_67,
  output        _EVAL_68,
  output        _EVAL_69,
  output [1:0]  _EVAL_70,
  output [2:0]  _EVAL_71,
  input  [2:0]  _EVAL_72,
  input         _EVAL_73,
  output [4:0]  _EVAL_74,
  input  [4:0]  _EVAL_75,
  input         _EVAL_76,
  output [4:0]  _EVAL_77,
  input         _EVAL_78,
  output        _EVAL_79,
  output        _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82
);
  assign _EVAL_71 = _EVAL_21;
  assign _EVAL_26 = _EVAL_34;
  assign _EVAL_5 = _EVAL_7;
  assign _EVAL_74 = _EVAL_10;
  assign _EVAL_53 = _EVAL_64;
  assign _EVAL_35 = _EVAL_8;
  assign _EVAL_33 = _EVAL_28;
  assign _EVAL_70 = _EVAL_61;
  assign _EVAL_62 = _EVAL_47;
  assign _EVAL_48 = _EVAL_37;
  assign _EVAL_15 = _EVAL_1;
  assign _EVAL_23 = _EVAL_45;
  assign _EVAL_18 = _EVAL_2;
  assign _EVAL_11 = _EVAL_46;
  assign _EVAL_6 = _EVAL_76;
  assign _EVAL_39 = _EVAL_14;
  assign _EVAL_3 = _EVAL_72;
  assign _EVAL_30 = _EVAL_41;
  assign _EVAL_77 = _EVAL_75;
  assign _EVAL_4 = _EVAL_49;
  assign _EVAL_59 = _EVAL_54;
  assign _EVAL_16 = _EVAL_38;
  assign _EVAL_0 = _EVAL_82;
  assign _EVAL_31 = _EVAL_57;
  assign _EVAL_69 = _EVAL_27;
  assign _EVAL_36 = _EVAL_78;
  assign _EVAL_65 = _EVAL_29;
  assign _EVAL_79 = _EVAL_44[0];
  assign _EVAL_19 = _EVAL_50;
  assign _EVAL_9 = _EVAL_73;
  assign _EVAL = _EVAL_58;
  assign _EVAL_22 = _EVAL_66;
  assign _EVAL_42 = _EVAL_55;
  assign _EVAL_17 = _EVAL_32;
  assign _EVAL_43 = _EVAL_20;
  assign _EVAL_13 = {{3'd0}, _EVAL_56};
  assign _EVAL_40 = {{3'd0}, _EVAL_81};
  assign _EVAL_12 = _EVAL_52[0];
  assign _EVAL_25 = _EVAL_51;
  assign _EVAL_63 = _EVAL_60;
  assign _EVAL_68 = _EVAL_67;
  assign _EVAL_80 = _EVAL_24;
endmodule
