//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_21(
  input         _EVAL,
  output [1:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [3:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output [7:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  input         _EVAL_8,
  output [30:0] _EVAL_9,
  output [2:0]  _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  output [3:0]  _EVAL_14,
  output [2:0]  _EVAL_15,
  output        _EVAL_16,
  input  [3:0]  _EVAL_17,
  input  [7:0]  _EVAL_18,
  input  [30:0] _EVAL_19,
  output        _EVAL_20,
  input  [1:0]  _EVAL_21,
  output [3:0]  _EVAL_22
);
  reg [30:0] _EVAL_23 [0:1];
  reg [31:0] _RAND_0;
  wire [30:0] _EVAL_23__EVAL_24_data;
  wire  _EVAL_23__EVAL_24_addr;
  wire [30:0] _EVAL_23__EVAL_25_data;
  wire  _EVAL_23__EVAL_25_addr;
  wire  _EVAL_23__EVAL_25_mask;
  wire  _EVAL_23__EVAL_25_en;
  reg  _EVAL_26 [0:1];
  reg [31:0] _RAND_1;
  wire  _EVAL_26__EVAL_27_data;
  wire  _EVAL_26__EVAL_27_addr;
  wire  _EVAL_26__EVAL_28_data;
  wire  _EVAL_26__EVAL_28_addr;
  wire  _EVAL_26__EVAL_28_mask;
  wire  _EVAL_26__EVAL_28_en;
  reg [2:0] _EVAL_30 [0:1];
  reg [31:0] _RAND_2;
  wire [2:0] _EVAL_30__EVAL_31_data;
  wire  _EVAL_30__EVAL_31_addr;
  wire [2:0] _EVAL_30__EVAL_32_data;
  wire  _EVAL_30__EVAL_32_addr;
  wire  _EVAL_30__EVAL_32_mask;
  wire  _EVAL_30__EVAL_32_en;
  reg [3:0] _EVAL_34 [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] _EVAL_34__EVAL_35_data;
  wire  _EVAL_34__EVAL_35_addr;
  wire [3:0] _EVAL_34__EVAL_36_data;
  wire  _EVAL_34__EVAL_36_addr;
  wire  _EVAL_34__EVAL_36_mask;
  wire  _EVAL_34__EVAL_36_en;
  reg [7:0] _EVAL_46 [0:1];
  reg [31:0] _RAND_4;
  wire [7:0] _EVAL_46__EVAL_47_data;
  wire  _EVAL_46__EVAL_47_addr;
  wire [7:0] _EVAL_46__EVAL_48_data;
  wire  _EVAL_46__EVAL_48_addr;
  wire  _EVAL_46__EVAL_48_mask;
  wire  _EVAL_46__EVAL_48_en;
  reg [1:0] _EVAL_51 [0:1];
  reg [31:0] _RAND_5;
  wire [1:0] _EVAL_51__EVAL_52_data;
  wire  _EVAL_51__EVAL_52_addr;
  wire [1:0] _EVAL_51__EVAL_53_data;
  wire  _EVAL_51__EVAL_53_addr;
  wire  _EVAL_51__EVAL_53_mask;
  wire  _EVAL_51__EVAL_53_en;
  reg [2:0] _EVAL_56 [0:1];
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_56__EVAL_57_data;
  wire  _EVAL_56__EVAL_57_addr;
  wire [2:0] _EVAL_56__EVAL_58_data;
  wire  _EVAL_56__EVAL_58_addr;
  wire  _EVAL_56__EVAL_58_mask;
  wire  _EVAL_56__EVAL_58_en;
  reg [3:0] _EVAL_59 [0:1];
  reg [31:0] _RAND_7;
  wire [3:0] _EVAL_59__EVAL_60_data;
  wire  _EVAL_59__EVAL_60_addr;
  wire [3:0] _EVAL_59__EVAL_61_data;
  wire  _EVAL_59__EVAL_61_addr;
  wire  _EVAL_59__EVAL_61_mask;
  wire  _EVAL_59__EVAL_61_en;
  reg [3:0] _EVAL_62 [0:1];
  reg [31:0] _RAND_8;
  wire [3:0] _EVAL_62__EVAL_63_data;
  wire  _EVAL_62__EVAL_63_addr;
  wire [3:0] _EVAL_62__EVAL_64_data;
  wire  _EVAL_62__EVAL_64_addr;
  wire  _EVAL_62__EVAL_64_mask;
  wire  _EVAL_62__EVAL_64_en;
  reg  _EVAL_33;
  reg [31:0] _RAND_9;
  reg  _EVAL_37;
  reg [31:0] _RAND_10;
  reg  _EVAL_42;
  reg [31:0] _RAND_11;
  wire  _EVAL_38;
  wire  _EVAL_65;
  wire  _EVAL_44;
  wire  _EVAL_39;
  wire  _EVAL_66;
  wire  _EVAL_41;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_40;
  assign _EVAL_23__EVAL_24_addr = _EVAL_33;
  assign _EVAL_23__EVAL_24_data = _EVAL_23[_EVAL_23__EVAL_24_addr];
  assign _EVAL_23__EVAL_25_data = _EVAL_19;
  assign _EVAL_23__EVAL_25_addr = _EVAL_42;
  assign _EVAL_23__EVAL_25_mask = 1'h1;
  assign _EVAL_23__EVAL_25_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_26__EVAL_27_addr = _EVAL_33;
  assign _EVAL_26__EVAL_27_data = _EVAL_26[_EVAL_26__EVAL_27_addr];
  assign _EVAL_26__EVAL_28_data = _EVAL_12;
  assign _EVAL_26__EVAL_28_addr = _EVAL_42;
  assign _EVAL_26__EVAL_28_mask = 1'h1;
  assign _EVAL_26__EVAL_28_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_30__EVAL_31_addr = _EVAL_33;
  assign _EVAL_30__EVAL_31_data = _EVAL_30[_EVAL_30__EVAL_31_addr];
  assign _EVAL_30__EVAL_32_data = _EVAL_13;
  assign _EVAL_30__EVAL_32_addr = _EVAL_42;
  assign _EVAL_30__EVAL_32_mask = 1'h1;
  assign _EVAL_30__EVAL_32_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_34__EVAL_35_addr = _EVAL_33;
  assign _EVAL_34__EVAL_35_data = _EVAL_34[_EVAL_34__EVAL_35_addr];
  assign _EVAL_34__EVAL_36_data = _EVAL_17;
  assign _EVAL_34__EVAL_36_addr = _EVAL_42;
  assign _EVAL_34__EVAL_36_mask = 1'h1;
  assign _EVAL_34__EVAL_36_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_46__EVAL_47_addr = _EVAL_33;
  assign _EVAL_46__EVAL_47_data = _EVAL_46[_EVAL_46__EVAL_47_addr];
  assign _EVAL_46__EVAL_48_data = _EVAL_18;
  assign _EVAL_46__EVAL_48_addr = _EVAL_42;
  assign _EVAL_46__EVAL_48_mask = 1'h1;
  assign _EVAL_46__EVAL_48_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_51__EVAL_52_addr = _EVAL_33;
  assign _EVAL_51__EVAL_52_data = _EVAL_51[_EVAL_51__EVAL_52_addr];
  assign _EVAL_51__EVAL_53_data = _EVAL_21;
  assign _EVAL_51__EVAL_53_addr = _EVAL_42;
  assign _EVAL_51__EVAL_53_mask = 1'h1;
  assign _EVAL_51__EVAL_53_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_56__EVAL_57_addr = _EVAL_33;
  assign _EVAL_56__EVAL_57_data = _EVAL_56[_EVAL_56__EVAL_57_addr];
  assign _EVAL_56__EVAL_58_data = _EVAL_1;
  assign _EVAL_56__EVAL_58_addr = _EVAL_42;
  assign _EVAL_56__EVAL_58_mask = 1'h1;
  assign _EVAL_56__EVAL_58_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_59__EVAL_60_addr = _EVAL_33;
  assign _EVAL_59__EVAL_60_data = _EVAL_59[_EVAL_59__EVAL_60_addr];
  assign _EVAL_59__EVAL_61_data = _EVAL_2;
  assign _EVAL_59__EVAL_61_addr = _EVAL_42;
  assign _EVAL_59__EVAL_61_mask = 1'h1;
  assign _EVAL_59__EVAL_61_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_62__EVAL_63_addr = _EVAL_33;
  assign _EVAL_62__EVAL_63_data = _EVAL_62[_EVAL_62__EVAL_63_addr];
  assign _EVAL_62__EVAL_64_data = _EVAL_6;
  assign _EVAL_62__EVAL_64_addr = _EVAL_42;
  assign _EVAL_62__EVAL_64_mask = 1'h1;
  assign _EVAL_62__EVAL_64_en = _EVAL_16 & _EVAL_3;
  assign _EVAL_38 = _EVAL_16 & _EVAL_3;
  assign _EVAL_65 = _EVAL & _EVAL_20;
  assign _EVAL_44 = _EVAL_38 != _EVAL_65;
  assign _EVAL_39 = _EVAL_37 == 1'h0;
  assign _EVAL_66 = _EVAL_42 == _EVAL_33;
  assign _EVAL_41 = _EVAL_42 + 1'h1;
  assign _EVAL_49 = _EVAL_33 + 1'h1;
  assign _EVAL_50 = _EVAL_66 & _EVAL_39;
  assign _EVAL_40 = _EVAL_66 & _EVAL_37;
  assign _EVAL_20 = _EVAL_50 == 1'h0;
  assign _EVAL_22 = _EVAL_62__EVAL_63_data;
  assign _EVAL_10 = _EVAL_56__EVAL_57_data;
  assign _EVAL_15 = _EVAL_30__EVAL_31_data;
  assign _EVAL_16 = _EVAL_40 == 1'h0;
  assign _EVAL_0 = _EVAL_51__EVAL_52_data;
  assign _EVAL_11 = _EVAL_26__EVAL_27_data;
  assign _EVAL_14 = _EVAL_59__EVAL_60_data;
  assign _EVAL_5 = _EVAL_46__EVAL_47_data;
  assign _EVAL_7 = _EVAL_34__EVAL_35_data;
  assign _EVAL_9 = _EVAL_23__EVAL_24_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_23[initvar] = _RAND_0[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_26[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_30[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_34[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_46[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_51[initvar] = _RAND_5[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_56[initvar] = _RAND_6[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_59[initvar] = _RAND_7[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_62[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_33 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_37 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_42 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_8) begin
    if(_EVAL_23__EVAL_25_en & _EVAL_23__EVAL_25_mask) begin
      _EVAL_23[_EVAL_23__EVAL_25_addr] <= _EVAL_23__EVAL_25_data;
    end
    if(_EVAL_26__EVAL_28_en & _EVAL_26__EVAL_28_mask) begin
      _EVAL_26[_EVAL_26__EVAL_28_addr] <= _EVAL_26__EVAL_28_data;
    end
    if(_EVAL_30__EVAL_32_en & _EVAL_30__EVAL_32_mask) begin
      _EVAL_30[_EVAL_30__EVAL_32_addr] <= _EVAL_30__EVAL_32_data;
    end
    if(_EVAL_34__EVAL_36_en & _EVAL_34__EVAL_36_mask) begin
      _EVAL_34[_EVAL_34__EVAL_36_addr] <= _EVAL_34__EVAL_36_data;
    end
    if(_EVAL_46__EVAL_48_en & _EVAL_46__EVAL_48_mask) begin
      _EVAL_46[_EVAL_46__EVAL_48_addr] <= _EVAL_46__EVAL_48_data;
    end
    if(_EVAL_51__EVAL_53_en & _EVAL_51__EVAL_53_mask) begin
      _EVAL_51[_EVAL_51__EVAL_53_addr] <= _EVAL_51__EVAL_53_data;
    end
    if(_EVAL_56__EVAL_58_en & _EVAL_56__EVAL_58_mask) begin
      _EVAL_56[_EVAL_56__EVAL_58_addr] <= _EVAL_56__EVAL_58_data;
    end
    if(_EVAL_59__EVAL_61_en & _EVAL_59__EVAL_61_mask) begin
      _EVAL_59[_EVAL_59__EVAL_61_addr] <= _EVAL_59__EVAL_61_data;
    end
    if(_EVAL_62__EVAL_64_en & _EVAL_62__EVAL_64_mask) begin
      _EVAL_62[_EVAL_62__EVAL_64_addr] <= _EVAL_62__EVAL_64_data;
    end
    if (_EVAL_4) begin
      _EVAL_33 <= 1'h0;
    end else begin
      if (_EVAL_65) begin
        _EVAL_33 <= _EVAL_49;
      end
    end
    if (_EVAL_4) begin
      _EVAL_37 <= 1'h0;
    end else begin
      if (_EVAL_44) begin
        _EVAL_37 <= _EVAL_38;
      end
    end
    if (_EVAL_4) begin
      _EVAL_42 <= 1'h0;
    end else begin
      if (_EVAL_38) begin
        _EVAL_42 <= _EVAL_41;
      end
    end
  end
endmodule
