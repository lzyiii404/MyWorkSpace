//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_40(
  output [3:0]  _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  output [1:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [63:0] _EVAL_6,
  input  [1:0]  _EVAL_7,
  output [2:0]  _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  output [1:0]  _EVAL_15,
  input         _EVAL_16,
  output [30:0] _EVAL_17,
  output [3:0]  _EVAL_18,
  output [2:0]  _EVAL_19,
  output [3:0]  _EVAL_20,
  input         _EVAL_21,
  output [63:0] _EVAL_22,
  output [3:0]  _EVAL_23,
  output        _EVAL_24,
  input  [3:0]  _EVAL_25,
  output        _EVAL_26,
  input  [2:0]  _EVAL_27,
  output [6:0]  _EVAL_28,
  output [30:0] _EVAL_29,
  input  [31:0] _EVAL_30,
  input  [6:0]  _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  output [2:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  output [3:0]  _EVAL_38,
  input         _EVAL_39,
  output [31:0] _EVAL_40,
  input  [30:0] _EVAL_41,
  output [2:0]  _EVAL_42,
  output [7:0]  _EVAL_43,
  input  [2:0]  _EVAL_44,
  input  [7:0]  _EVAL_45,
  output        _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  output [3:0]  _EVAL_49,
  input         _EVAL_50,
  output [2:0]  _EVAL_51,
  output [7:0]  _EVAL_52,
  output        _EVAL_53,
  output        _EVAL_54,
  output [3:0]  _EVAL_55
);
  wire  bridge_for_axi4_sys_port__EVAL;
  wire  bridge_for_axi4_sys_port__EVAL_0;
  wire [30:0] bridge_for_axi4_sys_port__EVAL_1;
  wire  bridge_for_axi4_sys_port__EVAL_2;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_3;
  wire  bridge_for_axi4_sys_port__EVAL_4;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_5;
  wire  bridge_for_axi4_sys_port__EVAL_6;
  wire  bridge_for_axi4_sys_port__EVAL_7;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_8;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_9;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_10;
  wire [31:0] bridge_for_axi4_sys_port__EVAL_11;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_12;
  wire [1:0] bridge_for_axi4_sys_port__EVAL_13;
  wire [30:0] bridge_for_axi4_sys_port__EVAL_14;
  wire [1:0] bridge_for_axi4_sys_port__EVAL_15;
  wire  bridge_for_axi4_sys_port__EVAL_16;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_17;
  wire  bridge_for_axi4_sys_port__EVAL_18;
  wire  bridge_for_axi4_sys_port__EVAL_19;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_20;
  wire  bridge_for_axi4_sys_port__EVAL_21;
  wire  bridge_for_axi4_sys_port__EVAL_22;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_23;
  wire [6:0] bridge_for_axi4_sys_port__EVAL_24;
  wire  bridge_for_axi4_sys_port__EVAL_25;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_26;
  wire  bridge_for_axi4_sys_port__EVAL_27;
  wire  bridge_for_axi4_sys_port__EVAL_28;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_29;
  wire  bridge_for_axi4_sys_port__EVAL_30;
  wire  bridge_for_axi4_sys_port__EVAL_31;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_32;
  wire  bridge_for_axi4_sys_port__EVAL_33;
  wire [7:0] bridge_for_axi4_sys_port__EVAL_34;
  wire  bridge_for_axi4_sys_port__EVAL_35;
  wire  bridge_for_axi4_sys_port__EVAL_36;
  wire  bridge_for_axi4_sys_port__EVAL_37;
  wire [1:0] bridge_for_axi4_sys_port__EVAL_38;
  wire [6:0] bridge_for_axi4_sys_port__EVAL_39;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_40;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_41;
  wire  bridge_for_axi4_sys_port__EVAL_42;
  wire [1:0] bridge_for_axi4_sys_port__EVAL_43;
  wire [31:0] bridge_for_axi4_sys_port__EVAL_44;
  wire [30:0] bridge_for_axi4_sys_port__EVAL_45;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_46;
  wire [3:0] bridge_for_axi4_sys_port__EVAL_47;
  wire [7:0] bridge_for_axi4_sys_port__EVAL_48;
  wire  bridge_for_axi4_sys_port__EVAL_49;
  wire  bridge_for_axi4_sys_port__EVAL_50;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_51;
  wire [63:0] bridge_for_axi4_sys_port__EVAL_52;
  wire [63:0] bridge_for_axi4_sys_port__EVAL_53;
  wire [7:0] bridge_for_axi4_sys_port__EVAL_54;
  wire [2:0] bridge_for_axi4_sys_port__EVAL_55;
  SiFive__EVAL_39 bridge_for_axi4_sys_port (
    ._EVAL(bridge_for_axi4_sys_port__EVAL),
    ._EVAL_0(bridge_for_axi4_sys_port__EVAL_0),
    ._EVAL_1(bridge_for_axi4_sys_port__EVAL_1),
    ._EVAL_2(bridge_for_axi4_sys_port__EVAL_2),
    ._EVAL_3(bridge_for_axi4_sys_port__EVAL_3),
    ._EVAL_4(bridge_for_axi4_sys_port__EVAL_4),
    ._EVAL_5(bridge_for_axi4_sys_port__EVAL_5),
    ._EVAL_6(bridge_for_axi4_sys_port__EVAL_6),
    ._EVAL_7(bridge_for_axi4_sys_port__EVAL_7),
    ._EVAL_8(bridge_for_axi4_sys_port__EVAL_8),
    ._EVAL_9(bridge_for_axi4_sys_port__EVAL_9),
    ._EVAL_10(bridge_for_axi4_sys_port__EVAL_10),
    ._EVAL_11(bridge_for_axi4_sys_port__EVAL_11),
    ._EVAL_12(bridge_for_axi4_sys_port__EVAL_12),
    ._EVAL_13(bridge_for_axi4_sys_port__EVAL_13),
    ._EVAL_14(bridge_for_axi4_sys_port__EVAL_14),
    ._EVAL_15(bridge_for_axi4_sys_port__EVAL_15),
    ._EVAL_16(bridge_for_axi4_sys_port__EVAL_16),
    ._EVAL_17(bridge_for_axi4_sys_port__EVAL_17),
    ._EVAL_18(bridge_for_axi4_sys_port__EVAL_18),
    ._EVAL_19(bridge_for_axi4_sys_port__EVAL_19),
    ._EVAL_20(bridge_for_axi4_sys_port__EVAL_20),
    ._EVAL_21(bridge_for_axi4_sys_port__EVAL_21),
    ._EVAL_22(bridge_for_axi4_sys_port__EVAL_22),
    ._EVAL_23(bridge_for_axi4_sys_port__EVAL_23),
    ._EVAL_24(bridge_for_axi4_sys_port__EVAL_24),
    ._EVAL_25(bridge_for_axi4_sys_port__EVAL_25),
    ._EVAL_26(bridge_for_axi4_sys_port__EVAL_26),
    ._EVAL_27(bridge_for_axi4_sys_port__EVAL_27),
    ._EVAL_28(bridge_for_axi4_sys_port__EVAL_28),
    ._EVAL_29(bridge_for_axi4_sys_port__EVAL_29),
    ._EVAL_30(bridge_for_axi4_sys_port__EVAL_30),
    ._EVAL_31(bridge_for_axi4_sys_port__EVAL_31),
    ._EVAL_32(bridge_for_axi4_sys_port__EVAL_32),
    ._EVAL_33(bridge_for_axi4_sys_port__EVAL_33),
    ._EVAL_34(bridge_for_axi4_sys_port__EVAL_34),
    ._EVAL_35(bridge_for_axi4_sys_port__EVAL_35),
    ._EVAL_36(bridge_for_axi4_sys_port__EVAL_36),
    ._EVAL_37(bridge_for_axi4_sys_port__EVAL_37),
    ._EVAL_38(bridge_for_axi4_sys_port__EVAL_38),
    ._EVAL_39(bridge_for_axi4_sys_port__EVAL_39),
    ._EVAL_40(bridge_for_axi4_sys_port__EVAL_40),
    ._EVAL_41(bridge_for_axi4_sys_port__EVAL_41),
    ._EVAL_42(bridge_for_axi4_sys_port__EVAL_42),
    ._EVAL_43(bridge_for_axi4_sys_port__EVAL_43),
    ._EVAL_44(bridge_for_axi4_sys_port__EVAL_44),
    ._EVAL_45(bridge_for_axi4_sys_port__EVAL_45),
    ._EVAL_46(bridge_for_axi4_sys_port__EVAL_46),
    ._EVAL_47(bridge_for_axi4_sys_port__EVAL_47),
    ._EVAL_48(bridge_for_axi4_sys_port__EVAL_48),
    ._EVAL_49(bridge_for_axi4_sys_port__EVAL_49),
    ._EVAL_50(bridge_for_axi4_sys_port__EVAL_50),
    ._EVAL_51(bridge_for_axi4_sys_port__EVAL_51),
    ._EVAL_52(bridge_for_axi4_sys_port__EVAL_52),
    ._EVAL_53(bridge_for_axi4_sys_port__EVAL_53),
    ._EVAL_54(bridge_for_axi4_sys_port__EVAL_54),
    ._EVAL_55(bridge_for_axi4_sys_port__EVAL_55)
  );
  assign bridge_for_axi4_sys_port__EVAL_4 = _EVAL_39;
  assign bridge_for_axi4_sys_port__EVAL_39 = _EVAL_31;
  assign _EVAL_43 = bridge_for_axi4_sys_port__EVAL_34;
  assign _EVAL_51 = bridge_for_axi4_sys_port__EVAL_41;
  assign bridge_for_axi4_sys_port__EVAL_5 = _EVAL_44;
  assign bridge_for_axi4_sys_port__EVAL_28 = _EVAL_10;
  assign _EVAL_24 = bridge_for_axi4_sys_port__EVAL_7;
  assign _EVAL_55 = bridge_for_axi4_sys_port__EVAL_29;
  assign _EVAL_40 = bridge_for_axi4_sys_port__EVAL_44;
  assign _EVAL_32 = bridge_for_axi4_sys_port__EVAL_36;
  assign bridge_for_axi4_sys_port__EVAL_35 = _EVAL_34;
  assign bridge_for_axi4_sys_port__EVAL_15 = _EVAL_7;
  assign _EVAL_23 = bridge_for_axi4_sys_port__EVAL_46;
  assign bridge_for_axi4_sys_port__EVAL_11 = _EVAL_30;
  assign _EVAL_53 = bridge_for_axi4_sys_port__EVAL_18;
  assign _EVAL_26 = bridge_for_axi4_sys_port__EVAL_21;
  assign bridge_for_axi4_sys_port__EVAL_37 = _EVAL_50;
  assign bridge_for_axi4_sys_port__EVAL = _EVAL_14;
  assign _EVAL_28 = bridge_for_axi4_sys_port__EVAL_24;
  assign _EVAL_36 = bridge_for_axi4_sys_port__EVAL_23;
  assign _EVAL_15 = bridge_for_axi4_sys_port__EVAL_38;
  assign _EVAL_8 = bridge_for_axi4_sys_port__EVAL_40;
  assign bridge_for_axi4_sys_port__EVAL_51 = _EVAL_27;
  assign _EVAL_4 = bridge_for_axi4_sys_port__EVAL_13;
  assign _EVAL_42 = bridge_for_axi4_sys_port__EVAL_9;
  assign bridge_for_axi4_sys_port__EVAL_45 = _EVAL_41;
  assign _EVAL_0 = bridge_for_axi4_sys_port__EVAL_31;
  assign bridge_for_axi4_sys_port__EVAL_48 = _EVAL_45;
  assign _EVAL = bridge_for_axi4_sys_port__EVAL_17;
  assign _EVAL_47 = bridge_for_axi4_sys_port__EVAL_30;
  assign bridge_for_axi4_sys_port__EVAL_42 = _EVAL_3;
  assign _EVAL_52 = bridge_for_axi4_sys_port__EVAL_54;
  assign _EVAL_38 = bridge_for_axi4_sys_port__EVAL_20;
  assign bridge_for_axi4_sys_port__EVAL_50 = _EVAL_16;
  assign _EVAL_18 = bridge_for_axi4_sys_port__EVAL_26;
  assign bridge_for_axi4_sys_port__EVAL_0 = _EVAL_11;
  assign _EVAL_33 = bridge_for_axi4_sys_port__EVAL_2;
  assign bridge_for_axi4_sys_port__EVAL_53 = _EVAL_6;
  assign _EVAL_17 = bridge_for_axi4_sys_port__EVAL_14;
  assign _EVAL_49 = bridge_for_axi4_sys_port__EVAL_32;
  assign _EVAL_54 = bridge_for_axi4_sys_port__EVAL_33;
  assign bridge_for_axi4_sys_port__EVAL_3 = _EVAL_5;
  assign bridge_for_axi4_sys_port__EVAL_49 = _EVAL_1;
  assign bridge_for_axi4_sys_port__EVAL_8 = _EVAL_13;
  assign _EVAL_9 = bridge_for_axi4_sys_port__EVAL_19;
  assign bridge_for_axi4_sys_port__EVAL_43 = _EVAL_12;
  assign bridge_for_axi4_sys_port__EVAL_16 = _EVAL_35;
  assign _EVAL_19 = bridge_for_axi4_sys_port__EVAL_12;
  assign _EVAL_20 = bridge_for_axi4_sys_port__EVAL_10;
  assign bridge_for_axi4_sys_port__EVAL_25 = _EVAL_21;
  assign _EVAL_2 = bridge_for_axi4_sys_port__EVAL_6;
  assign _EVAL_22 = bridge_for_axi4_sys_port__EVAL_52;
  assign _EVAL_29 = bridge_for_axi4_sys_port__EVAL_1;
  assign _EVAL_48 = bridge_for_axi4_sys_port__EVAL_27;
  assign _EVAL_46 = bridge_for_axi4_sys_port__EVAL_22;
  assign _EVAL_37 = bridge_for_axi4_sys_port__EVAL_55;
  assign bridge_for_axi4_sys_port__EVAL_47 = _EVAL_25;
endmodule
