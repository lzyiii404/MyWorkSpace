//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_156_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [6:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [14:0] _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [6:0]  _EVAL_13,
  input  [2:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_36;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_70;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_89;
  reg [31:0] _RAND_2;
  reg [14:0] _EVAL_118;
  reg [31:0] _RAND_3;
  reg [72:0] _EVAL_122;
  reg [95:0] _RAND_4;
  reg [3:0] _EVAL_126;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_130;
  reg [31:0] _RAND_6;
  reg [6:0] _EVAL_155;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_184;
  reg [31:0] _RAND_8;
  reg [6:0] _EVAL_195;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_206;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_236;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_237;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_279;
  reg [31:0] _RAND_13;
  wire  _EVAL_207;
  wire  _EVAL_85;
  wire  _EVAL_268;
  wire [3:0] _EVAL_29;
  wire  _EVAL_283;
  wire  _EVAL_78;
  wire  _EVAL_249;
  wire  _EVAL_246;
  wire  _EVAL_116;
  wire [12:0] _EVAL_39;
  wire [5:0] _EVAL_240;
  wire [5:0] _EVAL_103;
  wire  _EVAL_60;
  wire  _EVAL_201;
  wire  _EVAL_275;
  wire  _EVAL_219;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_101;
  wire  _EVAL_129;
  wire  _EVAL_262;
  wire  _EVAL_62;
  wire [127:0] _EVAL_228;
  wire [127:0] _EVAL_188;
  wire [72:0] _EVAL_99;
  wire  _EVAL_133;
  wire  _EVAL_91;
  wire [3:0] _EVAL_88;
  wire  _EVAL_254;
  wire [14:0] _EVAL_185;
  wire [15:0] _EVAL_239;
  wire [15:0] _EVAL_233;
  wire [15:0] _EVAL_145;
  wire  _EVAL_248;
  wire  _EVAL_193;
  wire  _EVAL_108;
  wire  _EVAL_286;
  wire  _EVAL_19;
  wire  _EVAL_111;
  wire  _EVAL_71;
  wire  _EVAL_163;
  wire  _EVAL_176;
  wire  _EVAL_117;
  wire [3:0] _EVAL_181;
  wire  _EVAL_199;
  wire  _EVAL_269;
  wire  _EVAL_49;
  wire  _EVAL_76;
  wire [72:0] _EVAL_146;
  wire  _EVAL_231;
  wire  _EVAL_45;
  wire  _EVAL_153;
  wire  _EVAL_52;
  wire  _EVAL_73;
  wire  _EVAL_79;
  wire [127:0] _EVAL_278;
  wire [127:0] _EVAL_144;
  wire [72:0] _EVAL_205;
  wire [72:0] _EVAL_157;
  wire [72:0] _EVAL_128;
  wire [14:0] _EVAL_244;
  wire [14:0] _EVAL_208;
  wire  _EVAL_243;
  wire  _EVAL_149;
  wire  _EVAL_43;
  wire  _EVAL_277;
  wire  _EVAL_284;
  wire [1:0] _EVAL_66;
  wire [1:0] _EVAL_216;
  wire  _EVAL_226;
  wire  _EVAL_222;
  wire  _EVAL_141;
  wire  _EVAL_274;
  wire  _EVAL_192;
  wire  _EVAL_93;
  wire  _EVAL_202;
  wire  _EVAL_166;
  wire  _EVAL_33;
  wire  _EVAL_267;
  wire  _EVAL_28;
  wire  _EVAL_104;
  wire  _EVAL_34;
  wire  _EVAL_161;
  wire  _EVAL_109;
  wire  _EVAL_63;
  wire  _EVAL_56;
  wire  _EVAL_179;
  wire  _EVAL_114;
  wire  _EVAL_217;
  wire  _EVAL_18;
  wire  _EVAL_288;
  wire [3:0] _EVAL_25;
  wire  _EVAL_259;
  wire  _EVAL_112;
  wire  _EVAL_255;
  wire  _EVAL_27;
  wire  _EVAL_137;
  wire  _EVAL_251;
  wire  _EVAL_53;
  wire [3:0] _EVAL_173;
  wire  _EVAL_32;
  wire [3:0] _EVAL_127;
  wire [72:0] _EVAL_272;
  wire  _EVAL_191;
  wire  _EVAL_265;
  wire  _EVAL_230;
  wire  _EVAL_223;
  wire  _EVAL_134;
  wire  _EVAL_225;
  wire  _EVAL_140;
  wire [3:0] _EVAL_110;
  wire  _EVAL_44;
  wire [2:0] _EVAL_35;
  wire  _EVAL_154;
  wire  _EVAL_41;
  wire  _EVAL_263;
  wire  _EVAL_287;
  wire  _EVAL_227;
  wire  _EVAL_106;
  wire  _EVAL_197;
  wire  _EVAL_69;
  wire  _EVAL_143;
  wire  _EVAL_50;
  wire  _EVAL_15;
  wire  _EVAL_31;
  wire  _EVAL_48;
  wire  _EVAL_83;
  wire  _EVAL_105;
  wire  _EVAL_121;
  wire  _EVAL_182;
  wire  _EVAL_187;
  wire [72:0] _EVAL_51;
  wire [72:0] _EVAL_224;
  wire  _EVAL_57;
  wire  _EVAL_22;
  wire  _EVAL_96;
  wire  _EVAL_172;
  wire  _EVAL_242;
  wire  _EVAL_21;
  wire  _EVAL_77;
  wire  _EVAL_194;
  wire  _EVAL_24;
  wire  _EVAL_160;
  wire  _EVAL_98;
  wire [31:0] _EVAL_260;
  wire  _EVAL_189;
  wire  _EVAL_264;
  wire  _EVAL_150;
  wire  _EVAL_253;
  wire  _EVAL_58;
  wire  _EVAL_273;
  wire  _EVAL_186;
  wire  _EVAL_81;
  wire  _EVAL_55;
  wire  _EVAL_280;
  wire  _EVAL_90;
  wire  _EVAL_158;
  wire  _EVAL_229;
  wire  _EVAL_61;
  wire [2:0] _EVAL_271;
  wire  _EVAL_282;
  wire  _EVAL_213;
  wire  _EVAL_221;
  wire  _EVAL_169;
  wire  _EVAL_204;
  wire  _EVAL_148;
  wire  _EVAL_59;
  wire  _EVAL_165;
  wire  _EVAL_198;
  wire  _EVAL_86;
  wire  _EVAL_147;
  wire  _EVAL_218;
  wire [12:0] _EVAL_209;
  wire [5:0] _EVAL_38;
  wire [5:0] _EVAL_132;
  wire [3:0] _EVAL_26;
  wire [3:0] _EVAL_256;
  wire  _EVAL_167;
  wire  _EVAL_84;
  wire  _EVAL_80;
  wire  _EVAL_87;
  wire  _EVAL_238;
  wire  _EVAL_92;
  wire  _EVAL_152;
  wire  _EVAL_136;
  wire  _EVAL_281;
  wire  _EVAL_252;
  wire  _EVAL_95;
  wire [3:0] _EVAL_113;
  wire  _EVAL_23;
  wire  _EVAL_151;
  wire  _EVAL_178;
  wire  _EVAL_177;
  wire  _EVAL_266;
  wire  _EVAL_82;
  wire  _EVAL_17;
  wire  _EVAL_241;
  wire  _EVAL_215;
  wire  _EVAL_54;
  wire  _EVAL_40;
  wire  _EVAL_214;
  wire  _EVAL_171;
  wire  _EVAL_72;
  wire  _EVAL_170;
  wire  _EVAL_100;
  wire  _EVAL_47;
  wire  _EVAL_285;
  wire  _EVAL_175;
  wire  _EVAL_46;
  wire  _EVAL_97;
  wire [3:0] _EVAL_120;
  wire  _EVAL_190;
  wire  _EVAL_220;
  wire  _EVAL_261;
  wire  _EVAL_139;
  wire  _EVAL_212;
  wire  _EVAL_37;
  wire  _EVAL_200;
  wire  _EVAL_16;
  wire  _EVAL_258;
  wire  _EVAL_64;
  wire [3:0] _EVAL_135;
  wire  _EVAL_174;
  wire  _EVAL_211;
  wire  _EVAL_196;
  wire  _EVAL_142;
  wire  _EVAL_20;
  wire  _EVAL_168;
  wire  _EVAL_180;
  wire  _EVAL_42;
  wire  _EVAL_232;
  wire  _EVAL_210;
  wire  _EVAL_164;
  wire  _EVAL_65;
  wire  _EVAL_245;
  wire  _EVAL_235;
  wire  _EVAL_250;
  wire  _EVAL_247;
  wire  _EVAL_125;
  wire  _EVAL_234;
  wire  _EVAL_67;
  wire  _EVAL_203;
  wire  _EVAL_115;
  wire  _EVAL_107;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_207 = _EVAL_13 == _EVAL_155;
  assign _EVAL_85 = _EVAL_207 | _EVAL_12;
  assign _EVAL_268 = _EVAL_85 == 1'h0;
  assign _EVAL_29 = ~ _EVAL_6;
  assign _EVAL_283 = _EVAL_29 == 4'h0;
  assign _EVAL_78 = _EVAL_283 | _EVAL_12;
  assign _EVAL_249 = _EVAL_78 == 1'h0;
  assign _EVAL_246 = _EVAL_5 == 3'h4;
  assign _EVAL_116 = _EVAL_8 & _EVAL_246;
  assign _EVAL_39 = 13'h3f << _EVAL_14;
  assign _EVAL_240 = _EVAL_39[5:0];
  assign _EVAL_103 = ~ _EVAL_240;
  assign _EVAL_60 = _EVAL_122 != 73'h0;
  assign _EVAL_201 = _EVAL_60 == 1'h0;
  assign _EVAL_275 = plusarg_reader_out == 32'h0;
  assign _EVAL_219 = _EVAL_201 | _EVAL_275;
  assign _EVAL_123 = _EVAL_36 < plusarg_reader_out;
  assign _EVAL_124 = _EVAL_219 | _EVAL_123;
  assign _EVAL_101 = _EVAL_124 | _EVAL_12;
  assign _EVAL_129 = _EVAL_4 & _EVAL_8;
  assign _EVAL_262 = _EVAL_126 == 4'h0;
  assign _EVAL_62 = _EVAL_129 & _EVAL_262;
  assign _EVAL_228 = 128'h1 << _EVAL_3;
  assign _EVAL_188 = _EVAL_62 ? _EVAL_228 : 128'h0;
  assign _EVAL_99 = _EVAL_188[72:0];
  assign _EVAL_133 = _EVAL_99 != 73'h0;
  assign _EVAL_91 = _EVAL_133 == 1'h0;
  assign _EVAL_88 = _EVAL_206 - 4'h1;
  assign _EVAL_254 = _EVAL_14 <= 3'h6;
  assign _EVAL_185 = _EVAL_7 ^ 15'h4000;
  assign _EVAL_239 = {1'b0,$signed(_EVAL_185)};
  assign _EVAL_233 = $signed(_EVAL_239) & $signed(-16'sh1000);
  assign _EVAL_145 = $signed(_EVAL_233);
  assign _EVAL_248 = $signed(_EVAL_145) == $signed(16'sh0);
  assign _EVAL_193 = _EVAL_254 & _EVAL_248;
  assign _EVAL_108 = _EVAL_193 | _EVAL_12;
  assign _EVAL_286 = _EVAL_11 == _EVAL_130;
  assign _EVAL_19 = _EVAL_286 | _EVAL_12;
  assign _EVAL_111 = _EVAL_19 == 1'h0;
  assign _EVAL_71 = _EVAL_11 == 3'h4;
  assign _EVAL_163 = _EVAL_0 & _EVAL_71;
  assign _EVAL_176 = _EVAL_5[2];
  assign _EVAL_117 = _EVAL_176 == 1'h0;
  assign _EVAL_181 = _EVAL_103[5:2];
  assign _EVAL_199 = _EVAL_5 == 3'h3;
  assign _EVAL_269 = _EVAL_8 & _EVAL_199;
  assign _EVAL_49 = _EVAL_13 == 7'h40;
  assign _EVAL_76 = _EVAL_1 != 3'h0;
  assign _EVAL_146 = _EVAL_122 | _EVAL_99;
  assign _EVAL_231 = _EVAL_9 & _EVAL_0;
  assign _EVAL_45 = _EVAL_236 == 4'h0;
  assign _EVAL_153 = _EVAL_231 & _EVAL_45;
  assign _EVAL_52 = _EVAL_11 == 3'h6;
  assign _EVAL_73 = _EVAL_52 == 1'h0;
  assign _EVAL_79 = _EVAL_153 & _EVAL_73;
  assign _EVAL_278 = 128'h1 << _EVAL_13;
  assign _EVAL_144 = _EVAL_79 ? _EVAL_278 : 128'h0;
  assign _EVAL_205 = _EVAL_144[72:0];
  assign _EVAL_157 = ~ _EVAL_205;
  assign _EVAL_128 = _EVAL_146 & _EVAL_157;
  assign _EVAL_244 = {{9'd0}, _EVAL_103};
  assign _EVAL_208 = _EVAL_7 & _EVAL_244;
  assign _EVAL_243 = _EVAL_208 == 15'h0;
  assign _EVAL_149 = _EVAL_5 == 3'h5;
  assign _EVAL_43 = _EVAL_8 & _EVAL_149;
  assign _EVAL_277 = _EVAL_14 >= 3'h2;
  assign _EVAL_284 = _EVAL_14[0];
  assign _EVAL_66 = 2'h1 << _EVAL_284;
  assign _EVAL_216 = _EVAL_66 | 2'h1;
  assign _EVAL_226 = _EVAL_216[1];
  assign _EVAL_222 = _EVAL_7[1];
  assign _EVAL_141 = _EVAL_226 & _EVAL_222;
  assign _EVAL_274 = _EVAL_277 | _EVAL_141;
  assign _EVAL_192 = _EVAL_216[0];
  assign _EVAL_93 = _EVAL_7[0];
  assign _EVAL_202 = _EVAL_222 & _EVAL_93;
  assign _EVAL_166 = _EVAL_192 & _EVAL_202;
  assign _EVAL_33 = _EVAL_274 | _EVAL_166;
  assign _EVAL_267 = _EVAL_93 == 1'h0;
  assign _EVAL_28 = _EVAL_222 & _EVAL_267;
  assign _EVAL_104 = _EVAL_192 & _EVAL_28;
  assign _EVAL_34 = _EVAL_274 | _EVAL_104;
  assign _EVAL_161 = _EVAL_222 == 1'h0;
  assign _EVAL_109 = _EVAL_226 & _EVAL_161;
  assign _EVAL_63 = _EVAL_277 | _EVAL_109;
  assign _EVAL_56 = _EVAL_161 & _EVAL_93;
  assign _EVAL_179 = _EVAL_192 & _EVAL_56;
  assign _EVAL_114 = _EVAL_63 | _EVAL_179;
  assign _EVAL_217 = _EVAL_161 & _EVAL_267;
  assign _EVAL_18 = _EVAL_192 & _EVAL_217;
  assign _EVAL_288 = _EVAL_63 | _EVAL_18;
  assign _EVAL_25 = {_EVAL_33,_EVAL_34,_EVAL_114,_EVAL_288};
  assign _EVAL_259 = _EVAL_6 == _EVAL_25;
  assign _EVAL_112 = _EVAL_259 | _EVAL_12;
  assign _EVAL_255 = _EVAL_5 == 3'h6;
  assign _EVAL_27 = _EVAL_3 == 7'h40;
  assign _EVAL_137 = _EVAL_11[0];
  assign _EVAL_251 = _EVAL_5 == _EVAL_184;
  assign _EVAL_53 = _EVAL_251 | _EVAL_12;
  assign _EVAL_173 = _EVAL_13[6:3];
  assign _EVAL_32 = _EVAL_173 == 4'h1;
  assign _EVAL_127 = _EVAL_126 - 4'h1;
  assign _EVAL_272 = _EVAL_122 >> _EVAL_3;
  assign _EVAL_191 = _EVAL_272[0];
  assign _EVAL_265 = _EVAL_191 == 1'h0;
  assign _EVAL_230 = _EVAL_265 | _EVAL_12;
  assign _EVAL_223 = _EVAL_230 == 1'h0;
  assign _EVAL_134 = _EVAL_112 == 1'h0;
  assign _EVAL_225 = _EVAL_3 == 7'h48;
  assign _EVAL_140 = _EVAL_225 | _EVAL_27;
  assign _EVAL_110 = _EVAL_3[6:3];
  assign _EVAL_44 = _EVAL_110 == 4'h8;
  assign _EVAL_35 = _EVAL_3[2:0];
  assign _EVAL_154 = 3'h1 <= _EVAL_35;
  assign _EVAL_41 = _EVAL_44 & _EVAL_154;
  assign _EVAL_263 = _EVAL_140 | _EVAL_41;
  assign _EVAL_287 = _EVAL_3 == 7'h20;
  assign _EVAL_227 = _EVAL_263 | _EVAL_287;
  assign _EVAL_106 = _EVAL_110 == 4'h0;
  assign _EVAL_197 = _EVAL_227 | _EVAL_106;
  assign _EVAL_69 = _EVAL_5 == 3'h0;
  assign _EVAL_143 = _EVAL_10 == 1'h0;
  assign _EVAL_50 = _EVAL_143 | _EVAL_12;
  assign _EVAL_15 = _EVAL_50 == 1'h0;
  assign _EVAL_31 = 3'h6 == _EVAL_14;
  assign _EVAL_48 = _EVAL_27 ? _EVAL_31 : 1'h0;
  assign _EVAL_83 = _EVAL_11 == 3'h5;
  assign _EVAL_105 = _EVAL_99 != _EVAL_205;
  assign _EVAL_121 = _EVAL_105 | _EVAL_91;
  assign _EVAL_182 = _EVAL_121 | _EVAL_12;
  assign _EVAL_187 = _EVAL_11 == 3'h1;
  assign _EVAL_51 = _EVAL_99 | _EVAL_122;
  assign _EVAL_224 = _EVAL_51 >> _EVAL_13;
  assign _EVAL_57 = _EVAL_1 == _EVAL_70;
  assign _EVAL_22 = _EVAL_57 | _EVAL_12;
  assign _EVAL_96 = _EVAL_22 == 1'h0;
  assign _EVAL_172 = _EVAL_89 == 4'h0;
  assign _EVAL_242 = _EVAL_12 == 1'h0;
  assign _EVAL_21 = _EVAL_8 & _EVAL_69;
  assign _EVAL_77 = _EVAL_173 == 4'h0;
  assign _EVAL_194 = _EVAL_108 == 1'h0;
  assign _EVAL_24 = _EVAL_76 | _EVAL_12;
  assign _EVAL_160 = _EVAL_24 == 1'h0;
  assign _EVAL_98 = _EVAL_173 == 4'h2;
  assign _EVAL_260 = _EVAL_36 + 32'h1;
  assign _EVAL_189 = _EVAL_206 == 4'h0;
  assign _EVAL_264 = _EVAL_189 == 1'h0;
  assign _EVAL_150 = _EVAL_8 & _EVAL_264;
  assign _EVAL_253 = _EVAL_5 == 3'h7;
  assign _EVAL_58 = _EVAL_13 == 7'h48;
  assign _EVAL_273 = _EVAL_110 == 4'h2;
  assign _EVAL_186 = _EVAL_224[0];
  assign _EVAL_81 = _EVAL_1 <= 3'h3;
  assign _EVAL_55 = _EVAL_81 | _EVAL_12;
  assign _EVAL_280 = _EVAL >= 3'h2;
  assign _EVAL_90 = _EVAL_280 | _EVAL_12;
  assign _EVAL_158 = _EVAL_90 == 1'h0;
  assign _EVAL_229 = _EVAL_58 | _EVAL_49;
  assign _EVAL_61 = _EVAL_173 == 4'h8;
  assign _EVAL_271 = _EVAL_13[2:0];
  assign _EVAL_282 = 3'h1 <= _EVAL_271;
  assign _EVAL_213 = _EVAL_61 & _EVAL_282;
  assign _EVAL_221 = _EVAL_229 | _EVAL_213;
  assign _EVAL_169 = _EVAL_13 == 7'h20;
  assign _EVAL_204 = _EVAL_221 | _EVAL_169;
  assign _EVAL_148 = _EVAL_204 | _EVAL_77;
  assign _EVAL_59 = _EVAL_148 | _EVAL_32;
  assign _EVAL_165 = _EVAL_186 | _EVAL_12;
  assign _EVAL_198 = _EVAL_165 == 1'h0;
  assign _EVAL_86 = _EVAL_59 | _EVAL_98;
  assign _EVAL_147 = _EVAL_173 == 4'h3;
  assign _EVAL_218 = _EVAL_86 | _EVAL_147;
  assign _EVAL_209 = 13'h3f << _EVAL;
  assign _EVAL_38 = _EVAL_209[5:0];
  assign _EVAL_132 = ~ _EVAL_38;
  assign _EVAL_26 = _EVAL_132[5:2];
  assign _EVAL_256 = ~ _EVAL_25;
  assign _EVAL_167 = _EVAL_11 == 3'h2;
  assign _EVAL_84 = _EVAL_110 == 4'h1;
  assign _EVAL_80 = _EVAL_197 | _EVAL_84;
  assign _EVAL_87 = _EVAL_80 | _EVAL_273;
  assign _EVAL_238 = _EVAL_110 == 4'h3;
  assign _EVAL_92 = _EVAL_87 | _EVAL_238;
  assign _EVAL_152 = _EVAL_92 | _EVAL_12;
  assign _EVAL_136 = _EVAL_152 == 1'h0;
  assign _EVAL_281 = _EVAL_48 | _EVAL_12;
  assign _EVAL_252 = _EVAL_14 == _EVAL_237;
  assign _EVAL_95 = _EVAL_252 | _EVAL_12;
  assign _EVAL_113 = _EVAL_89 - 4'h1;
  assign _EVAL_23 = _EVAL == _EVAL_279;
  assign _EVAL_151 = _EVAL_172 == 1'h0;
  assign _EVAL_178 = _EVAL_11 <= 3'h6;
  assign _EVAL_177 = _EVAL_0 & _EVAL_187;
  assign _EVAL_266 = _EVAL_1 == 3'h0;
  assign _EVAL_82 = _EVAL_3 == _EVAL_195;
  assign _EVAL_17 = _EVAL_82 | _EVAL_12;
  assign _EVAL_241 = _EVAL_178 | _EVAL_12;
  assign _EVAL_215 = _EVAL_241 == 1'h0;
  assign _EVAL_54 = _EVAL_1 <= 3'h2;
  assign _EVAL_40 = _EVAL_54 | _EVAL_12;
  assign _EVAL_214 = _EVAL_40 == 1'h0;
  assign _EVAL_171 = _EVAL_1 <= 3'h4;
  assign _EVAL_72 = _EVAL_171 | _EVAL_12;
  assign _EVAL_170 = _EVAL_72 == 1'h0;
  assign _EVAL_100 = _EVAL_0 & _EVAL_151;
  assign _EVAL_47 = _EVAL_129 | _EVAL_231;
  assign _EVAL_285 = _EVAL_277 | _EVAL_12;
  assign _EVAL_175 = _EVAL_5 == 3'h2;
  assign _EVAL_46 = _EVAL_8 & _EVAL_175;
  assign _EVAL_97 = _EVAL_266 | _EVAL_12;
  assign _EVAL_120 = _EVAL_236 - 4'h1;
  assign _EVAL_190 = _EVAL_8 & _EVAL_253;
  assign _EVAL_220 = _EVAL_0 & _EVAL_167;
  assign _EVAL_261 = _EVAL_285 == 1'h0;
  assign _EVAL_139 = _EVAL_218 | _EVAL_12;
  assign _EVAL_212 = _EVAL_139 == 1'h0;
  assign _EVAL_37 = _EVAL_7 == _EVAL_118;
  assign _EVAL_200 = _EVAL_37 | _EVAL_12;
  assign _EVAL_16 = _EVAL_243 | _EVAL_12;
  assign _EVAL_258 = _EVAL_97 == 1'h0;
  assign _EVAL_64 = _EVAL_8 & _EVAL_255;
  assign _EVAL_135 = _EVAL_6 & _EVAL_256;
  assign _EVAL_174 = _EVAL_135 == 4'h0;
  assign _EVAL_211 = _EVAL_174 | _EVAL_12;
  assign _EVAL_196 = _EVAL_211 == 1'h0;
  assign _EVAL_142 = _EVAL_53 == 1'h0;
  assign _EVAL_20 = _EVAL_17 == 1'h0;
  assign _EVAL_168 = _EVAL_231 & _EVAL_172;
  assign _EVAL_180 = _EVAL_182 == 1'h0;
  assign _EVAL_42 = _EVAL_11 == 3'h0;
  assign _EVAL_232 = _EVAL_0 & _EVAL_42;
  assign _EVAL_210 = _EVAL_129 & _EVAL_189;
  assign _EVAL_164 = _EVAL_16 == 1'h0;
  assign _EVAL_65 = _EVAL_0 & _EVAL_83;
  assign _EVAL_245 = _EVAL_281 == 1'h0;
  assign _EVAL_235 = _EVAL_5 == 3'h1;
  assign _EVAL_250 = _EVAL_8 & _EVAL_235;
  assign _EVAL_247 = _EVAL_55 == 1'h0;
  assign _EVAL_125 = _EVAL_0 & _EVAL_52;
  assign _EVAL_234 = _EVAL_23 | _EVAL_12;
  assign _EVAL_67 = _EVAL_234 == 1'h0;
  assign _EVAL_203 = _EVAL_101 == 1'h0;
  assign _EVAL_115 = _EVAL_200 == 1'h0;
  assign _EVAL_107 = _EVAL_95 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_36 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_70 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_89 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_118 = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  _EVAL_122 = _RAND_4[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_126 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_130 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_155 = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_184 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_195 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_206 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_236 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_237 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_279 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_12) begin
      _EVAL_36 <= 32'h0;
    end else begin
      if (_EVAL_47) begin
        _EVAL_36 <= 32'h0;
      end else begin
        _EVAL_36 <= _EVAL_260;
      end
    end
    if (_EVAL_210) begin
      _EVAL_70 <= _EVAL_1;
    end
    if (_EVAL_12) begin
      _EVAL_89 <= 4'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_172) begin
          if (_EVAL_137) begin
            _EVAL_89 <= _EVAL_26;
          end else begin
            _EVAL_89 <= 4'h0;
          end
        end else begin
          _EVAL_89 <= _EVAL_113;
        end
      end
    end
    if (_EVAL_210) begin
      _EVAL_118 <= _EVAL_7;
    end
    if (_EVAL_12) begin
      _EVAL_122 <= 73'h0;
    end else begin
      _EVAL_122 <= _EVAL_128;
    end
    if (_EVAL_12) begin
      _EVAL_126 <= 4'h0;
    end else begin
      if (_EVAL_129) begin
        if (_EVAL_262) begin
          if (_EVAL_117) begin
            _EVAL_126 <= _EVAL_181;
          end else begin
            _EVAL_126 <= 4'h0;
          end
        end else begin
          _EVAL_126 <= _EVAL_127;
        end
      end
    end
    if (_EVAL_168) begin
      _EVAL_130 <= _EVAL_11;
    end
    if (_EVAL_168) begin
      _EVAL_155 <= _EVAL_13;
    end
    if (_EVAL_210) begin
      _EVAL_184 <= _EVAL_5;
    end
    if (_EVAL_210) begin
      _EVAL_195 <= _EVAL_3;
    end
    if (_EVAL_12) begin
      _EVAL_206 <= 4'h0;
    end else begin
      if (_EVAL_129) begin
        if (_EVAL_189) begin
          if (_EVAL_117) begin
            _EVAL_206 <= _EVAL_181;
          end else begin
            _EVAL_206 <= 4'h0;
          end
        end else begin
          _EVAL_206 <= _EVAL_88;
        end
      end
    end
    if (_EVAL_12) begin
      _EVAL_236 <= 4'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_45) begin
          if (_EVAL_137) begin
            _EVAL_236 <= _EVAL_26;
          end else begin
            _EVAL_236 <= 4'h0;
          end
        end else begin
          _EVAL_236 <= _EVAL_120;
        end
      end
    end
    if (_EVAL_210) begin
      _EVAL_237 <= _EVAL_14;
    end
    if (_EVAL_168) begin
      _EVAL_279 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7746a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3868b797)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b3716a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc08a8f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a22f86f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33d2784)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8206ade2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a084b9a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3090fb8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee5d04b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(172563cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6702cdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c766df9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b53d05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c11b907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aee51283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f51e1c7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9ab6ae1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c5604d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14a37d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(537647f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b8c2ad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(282edf26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac90d79f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35ab4ef6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f469f986)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7df1ae5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e35061c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d130f65e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(893ae7eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bad02596)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98023c7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6249fcd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0a144a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72747584)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4ef97b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab946d38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bd94afc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65db6011)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28283f77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e43dcff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae92ec75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f2f28fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(926209c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49eea6b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1be551ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(456de75a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c417d4a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcdc7dbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30ec002)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1e9cd25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(858f0273)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c454850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3028f83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43b5b74d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edc07cdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ca7322c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10d0945c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccd6b1c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fcae01d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68a7eaf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be8fc856)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba5be1a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c832b31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4cae8e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d778643e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2dd7cbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f8dbb24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cf48ef6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7b578b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c18cd4a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1f72d1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
