//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_208(
  input         _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input  [1:0]  _EVAL_4,
  output [31:0] _EVAL_5,
  output [3:0]  _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [31:0] _EVAL_12,
  output [31:0] _EVAL_13,
  input  [1:0]  _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  output        _EVAL_21,
  output        _EVAL_22,
  output [8:0]  _EVAL_23,
  input         _EVAL_24,
  output [2:0]  _EVAL_25,
  output        _EVAL_26,
  input  [2:0]  _EVAL_27,
  output        _EVAL_28,
  input  [31:0] _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  output [1:0]  _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  output        _EVAL_37,
  output [9:0]  _EVAL_38,
  input         _EVAL_39,
  output        _EVAL_40,
  input  [6:0]  _EVAL_41
);
  wire  dmiXbar__EVAL;
  wire [31:0] dmiXbar__EVAL_0;
  wire  dmiXbar__EVAL_1;
  wire  dmiXbar__EVAL_2;
  wire  dmiXbar__EVAL_3;
  wire [2:0] dmiXbar__EVAL_4;
  wire  dmiXbar__EVAL_5;
  wire [31:0] dmiXbar__EVAL_6;
  wire  dmiXbar__EVAL_7;
  wire [2:0] dmiXbar__EVAL_8;
  wire [1:0] dmiXbar__EVAL_9;
  wire  dmiXbar__EVAL_10;
  wire [31:0] dmiXbar__EVAL_11;
  wire  dmiXbar__EVAL_12;
  wire  dmiXbar__EVAL_13;
  wire [1:0] dmiXbar__EVAL_14;
  wire  dmiXbar__EVAL_15;
  wire  dmiXbar__EVAL_16;
  wire  dmiXbar__EVAL_17;
  wire [3:0] dmiXbar__EVAL_18;
  wire  dmiXbar__EVAL_19;
  wire [31:0] dmiXbar__EVAL_20;
  wire  dmiXbar__EVAL_21;
  wire [2:0] dmiXbar__EVAL_22;
  wire  dmiXbar__EVAL_23;
  wire [8:0] dmiXbar__EVAL_24;
  wire  dmiXbar__EVAL_25;
  wire [2:0] dmiXbar__EVAL_26;
  wire  dmiXbar__EVAL_27;
  wire [3:0] dmiXbar__EVAL_28;
  wire [2:0] dmiXbar__EVAL_29;
  wire [3:0] dmiXbar__EVAL_30;
  wire [31:0] dmiXbar__EVAL_31;
  wire  dmiXbar__EVAL_32;
  wire [31:0] dmiXbar__EVAL_33;
  wire  dmiXbar__EVAL_34;
  wire [6:0] dmiXbar__EVAL_35;
  wire  dmiXbar__EVAL_36;
  wire [8:0] dmiXbar__EVAL_37;
  wire  asource__EVAL;
  wire [2:0] asource__EVAL_0;
  wire  asource__EVAL_1;
  wire  asource__EVAL_2;
  wire  asource__EVAL_3;
  wire [31:0] asource__EVAL_4;
  wire  asource__EVAL_5;
  wire  asource__EVAL_6;
  wire [2:0] asource__EVAL_7;
  wire  asource__EVAL_8;
  wire [31:0] asource__EVAL_9;
  wire [1:0] asource__EVAL_10;
  wire  asource__EVAL_11;
  wire  asource__EVAL_12;
  wire  asource__EVAL_13;
  wire [2:0] asource__EVAL_14;
  wire  asource__EVAL_15;
  wire [3:0] asource__EVAL_16;
  wire [2:0] asource__EVAL_17;
  wire [1:0] asource__EVAL_18;
  wire  asource__EVAL_19;
  wire  asource__EVAL_20;
  wire  asource__EVAL_21;
  wire [1:0] asource__EVAL_22;
  wire [31:0] asource__EVAL_23;
  wire  asource__EVAL_24;
  wire [3:0] asource__EVAL_25;
  wire [8:0] asource__EVAL_26;
  wire  asource__EVAL_27;
  wire  asource__EVAL_28;
  wire  asource__EVAL_29;
  wire [31:0] asource__EVAL_30;
  wire [8:0] asource__EVAL_31;
  wire  asource__EVAL_32;
  wire  asource__EVAL_33;
  wire  asource__EVAL_34;
  wire [9:0] AsyncQueueSource__EVAL;
  wire  AsyncQueueSource__EVAL_0;
  wire  AsyncQueueSource__EVAL_1;
  wire  AsyncQueueSource__EVAL_2;
  wire  AsyncQueueSource__EVAL_3;
  wire  AsyncQueueSource__EVAL_4;
  wire  AsyncQueueSource__EVAL_5;
  wire  AsyncQueueSource__EVAL_6;
  wire  AsyncQueueSource__EVAL_7;
  wire  AsyncQueueSource__EVAL_8;
  wire  AsyncQueueSource__EVAL_9;
  wire  AsyncQueueSource__EVAL_10;
  wire [9:0] AsyncQueueSource__EVAL_11;
  wire  AsyncQueueSource__EVAL_12;
  wire  AsyncQueueSource__EVAL_13;
  wire  AsyncQueueSource__EVAL_14;
  wire  AsyncQueueSource__EVAL_15;
  wire  AsyncQueueSource__EVAL_16;
  wire  intsource__EVAL;
  wire  intsource__EVAL_0;
  wire  dmOuter__EVAL;
  wire  dmOuter__EVAL_0;
  wire [3:0] dmOuter__EVAL_1;
  wire  dmOuter__EVAL_2;
  wire  dmOuter__EVAL_3;
  wire  dmOuter__EVAL_4;
  wire [9:0] dmOuter__EVAL_5;
  wire  dmOuter__EVAL_6;
  wire  dmOuter__EVAL_7;
  wire [6:0] dmOuter__EVAL_8;
  wire  dmOuter__EVAL_9;
  wire  dmOuter__EVAL_10;
  wire [2:0] dmOuter__EVAL_11;
  wire [31:0] dmOuter__EVAL_12;
  wire  dmOuter__EVAL_13;
  wire  dmOuter__EVAL_14;
  wire [2:0] dmOuter__EVAL_15;
  wire [31:0] dmOuter__EVAL_16;
  wire  dmOuter__EVAL_17;
  wire  dmOuter__EVAL_18;
  wire  dmOuter__EVAL_19;
  wire [3:0] dmi2tl__EVAL;
  wire  dmi2tl__EVAL_0;
  wire [1:0] dmi2tl__EVAL_1;
  wire  dmi2tl__EVAL_2;
  wire [1:0] dmi2tl__EVAL_3;
  wire [6:0] dmi2tl__EVAL_4;
  wire  dmi2tl__EVAL_5;
  wire [2:0] dmi2tl__EVAL_6;
  wire  dmi2tl__EVAL_7;
  wire [31:0] dmi2tl__EVAL_8;
  wire  dmi2tl__EVAL_9;
  wire [8:0] dmi2tl__EVAL_10;
  wire  dmi2tl__EVAL_11;
  wire  dmi2tl__EVAL_12;
  wire [31:0] dmi2tl__EVAL_13;
  wire  dmi2tl__EVAL_14;
  wire  dmi2tl__EVAL_15;
  wire  dmi2tl__EVAL_16;
  wire [31:0] dmi2tl__EVAL_17;
  wire [31:0] dmi2tl__EVAL_18;
  SiFive__EVAL_189 dmiXbar (
    ._EVAL(dmiXbar__EVAL),
    ._EVAL_0(dmiXbar__EVAL_0),
    ._EVAL_1(dmiXbar__EVAL_1),
    ._EVAL_2(dmiXbar__EVAL_2),
    ._EVAL_3(dmiXbar__EVAL_3),
    ._EVAL_4(dmiXbar__EVAL_4),
    ._EVAL_5(dmiXbar__EVAL_5),
    ._EVAL_6(dmiXbar__EVAL_6),
    ._EVAL_7(dmiXbar__EVAL_7),
    ._EVAL_8(dmiXbar__EVAL_8),
    ._EVAL_9(dmiXbar__EVAL_9),
    ._EVAL_10(dmiXbar__EVAL_10),
    ._EVAL_11(dmiXbar__EVAL_11),
    ._EVAL_12(dmiXbar__EVAL_12),
    ._EVAL_13(dmiXbar__EVAL_13),
    ._EVAL_14(dmiXbar__EVAL_14),
    ._EVAL_15(dmiXbar__EVAL_15),
    ._EVAL_16(dmiXbar__EVAL_16),
    ._EVAL_17(dmiXbar__EVAL_17),
    ._EVAL_18(dmiXbar__EVAL_18),
    ._EVAL_19(dmiXbar__EVAL_19),
    ._EVAL_20(dmiXbar__EVAL_20),
    ._EVAL_21(dmiXbar__EVAL_21),
    ._EVAL_22(dmiXbar__EVAL_22),
    ._EVAL_23(dmiXbar__EVAL_23),
    ._EVAL_24(dmiXbar__EVAL_24),
    ._EVAL_25(dmiXbar__EVAL_25),
    ._EVAL_26(dmiXbar__EVAL_26),
    ._EVAL_27(dmiXbar__EVAL_27),
    ._EVAL_28(dmiXbar__EVAL_28),
    ._EVAL_29(dmiXbar__EVAL_29),
    ._EVAL_30(dmiXbar__EVAL_30),
    ._EVAL_31(dmiXbar__EVAL_31),
    ._EVAL_32(dmiXbar__EVAL_32),
    ._EVAL_33(dmiXbar__EVAL_33),
    ._EVAL_34(dmiXbar__EVAL_34),
    ._EVAL_35(dmiXbar__EVAL_35),
    ._EVAL_36(dmiXbar__EVAL_36),
    ._EVAL_37(dmiXbar__EVAL_37)
  );
  SiFive__EVAL_206 asource (
    ._EVAL(asource__EVAL),
    ._EVAL_0(asource__EVAL_0),
    ._EVAL_1(asource__EVAL_1),
    ._EVAL_2(asource__EVAL_2),
    ._EVAL_3(asource__EVAL_3),
    ._EVAL_4(asource__EVAL_4),
    ._EVAL_5(asource__EVAL_5),
    ._EVAL_6(asource__EVAL_6),
    ._EVAL_7(asource__EVAL_7),
    ._EVAL_8(asource__EVAL_8),
    ._EVAL_9(asource__EVAL_9),
    ._EVAL_10(asource__EVAL_10),
    ._EVAL_11(asource__EVAL_11),
    ._EVAL_12(asource__EVAL_12),
    ._EVAL_13(asource__EVAL_13),
    ._EVAL_14(asource__EVAL_14),
    ._EVAL_15(asource__EVAL_15),
    ._EVAL_16(asource__EVAL_16),
    ._EVAL_17(asource__EVAL_17),
    ._EVAL_18(asource__EVAL_18),
    ._EVAL_19(asource__EVAL_19),
    ._EVAL_20(asource__EVAL_20),
    ._EVAL_21(asource__EVAL_21),
    ._EVAL_22(asource__EVAL_22),
    ._EVAL_23(asource__EVAL_23),
    ._EVAL_24(asource__EVAL_24),
    ._EVAL_25(asource__EVAL_25),
    ._EVAL_26(asource__EVAL_26),
    ._EVAL_27(asource__EVAL_27),
    ._EVAL_28(asource__EVAL_28),
    ._EVAL_29(asource__EVAL_29),
    ._EVAL_30(asource__EVAL_30),
    ._EVAL_31(asource__EVAL_31),
    ._EVAL_32(asource__EVAL_32),
    ._EVAL_33(asource__EVAL_33),
    ._EVAL_34(asource__EVAL_34)
  );
  SiFive__EVAL_207 AsyncQueueSource (
    ._EVAL(AsyncQueueSource__EVAL),
    ._EVAL_0(AsyncQueueSource__EVAL_0),
    ._EVAL_1(AsyncQueueSource__EVAL_1),
    ._EVAL_2(AsyncQueueSource__EVAL_2),
    ._EVAL_3(AsyncQueueSource__EVAL_3),
    ._EVAL_4(AsyncQueueSource__EVAL_4),
    ._EVAL_5(AsyncQueueSource__EVAL_5),
    ._EVAL_6(AsyncQueueSource__EVAL_6),
    ._EVAL_7(AsyncQueueSource__EVAL_7),
    ._EVAL_8(AsyncQueueSource__EVAL_8),
    ._EVAL_9(AsyncQueueSource__EVAL_9),
    ._EVAL_10(AsyncQueueSource__EVAL_10),
    ._EVAL_11(AsyncQueueSource__EVAL_11),
    ._EVAL_12(AsyncQueueSource__EVAL_12),
    ._EVAL_13(AsyncQueueSource__EVAL_13),
    ._EVAL_14(AsyncQueueSource__EVAL_14),
    ._EVAL_15(AsyncQueueSource__EVAL_15),
    ._EVAL_16(AsyncQueueSource__EVAL_16)
  );
  SiFive__EVAL_195 intsource (
    ._EVAL(intsource__EVAL),
    ._EVAL_0(intsource__EVAL_0)
  );
  SiFive__EVAL_194 dmOuter (
    ._EVAL(dmOuter__EVAL),
    ._EVAL_0(dmOuter__EVAL_0),
    ._EVAL_1(dmOuter__EVAL_1),
    ._EVAL_2(dmOuter__EVAL_2),
    ._EVAL_3(dmOuter__EVAL_3),
    ._EVAL_4(dmOuter__EVAL_4),
    ._EVAL_5(dmOuter__EVAL_5),
    ._EVAL_6(dmOuter__EVAL_6),
    ._EVAL_7(dmOuter__EVAL_7),
    ._EVAL_8(dmOuter__EVAL_8),
    ._EVAL_9(dmOuter__EVAL_9),
    ._EVAL_10(dmOuter__EVAL_10),
    ._EVAL_11(dmOuter__EVAL_11),
    ._EVAL_12(dmOuter__EVAL_12),
    ._EVAL_13(dmOuter__EVAL_13),
    ._EVAL_14(dmOuter__EVAL_14),
    ._EVAL_15(dmOuter__EVAL_15),
    ._EVAL_16(dmOuter__EVAL_16),
    ._EVAL_17(dmOuter__EVAL_17),
    ._EVAL_18(dmOuter__EVAL_18),
    ._EVAL_19(dmOuter__EVAL_19)
  );
  SiFive__EVAL_190 dmi2tl (
    ._EVAL(dmi2tl__EVAL),
    ._EVAL_0(dmi2tl__EVAL_0),
    ._EVAL_1(dmi2tl__EVAL_1),
    ._EVAL_2(dmi2tl__EVAL_2),
    ._EVAL_3(dmi2tl__EVAL_3),
    ._EVAL_4(dmi2tl__EVAL_4),
    ._EVAL_5(dmi2tl__EVAL_5),
    ._EVAL_6(dmi2tl__EVAL_6),
    ._EVAL_7(dmi2tl__EVAL_7),
    ._EVAL_8(dmi2tl__EVAL_8),
    ._EVAL_9(dmi2tl__EVAL_9),
    ._EVAL_10(dmi2tl__EVAL_10),
    ._EVAL_11(dmi2tl__EVAL_11),
    ._EVAL_12(dmi2tl__EVAL_12),
    ._EVAL_13(dmi2tl__EVAL_13),
    ._EVAL_14(dmi2tl__EVAL_14),
    ._EVAL_15(dmi2tl__EVAL_15),
    ._EVAL_16(dmi2tl__EVAL_16),
    ._EVAL_17(dmi2tl__EVAL_17),
    ._EVAL_18(dmi2tl__EVAL_18)
  );
  assign dmi2tl__EVAL_4 = _EVAL_41;
  assign dmi2tl__EVAL_2 = _EVAL_2;
  assign dmiXbar__EVAL_6 = dmOuter__EVAL_16;
  assign dmiXbar__EVAL_24 = dmi2tl__EVAL_10;
  assign asource__EVAL_33 = _EVAL_11;
  assign _EVAL_16 = AsyncQueueSource__EVAL_7;
  assign asource__EVAL_34 = _EVAL;
  assign _EVAL_26 = AsyncQueueSource__EVAL_6;
  assign dmOuter__EVAL_15 = dmiXbar__EVAL_8;
  assign dmiXbar__EVAL_27 = _EVAL_31;
  assign dmOuter__EVAL_2 = _EVAL_35;
  assign _EVAL_28 = dmOuter__EVAL_19;
  assign AsyncQueueSource__EVAL_12 = _EVAL_10;
  assign dmi2tl__EVAL_7 = _EVAL_1;
  assign dmiXbar__EVAL_15 = asource__EVAL_5;
  assign dmOuter__EVAL_12 = dmiXbar__EVAL_31;
  assign dmiXbar__EVAL_9 = asource__EVAL_18;
  assign AsyncQueueSource__EVAL_1 = _EVAL_20;
  assign dmiXbar__EVAL_7 = dmi2tl__EVAL_12;
  assign dmOuter__EVAL_14 = _EVAL_31;
  assign _EVAL_25 = asource__EVAL_0;
  assign _EVAL_17 = intsource__EVAL;
  assign dmiXbar__EVAL_14 = asource__EVAL_22;
  assign dmiXbar__EVAL_20 = dmi2tl__EVAL_17;
  assign _EVAL_13 = asource__EVAL_4;
  assign dmOuter__EVAL_8 = dmiXbar__EVAL_35;
  assign _EVAL_6 = asource__EVAL_25;
  assign _EVAL_38 = AsyncQueueSource__EVAL_11;
  assign _EVAL_32 = dmi2tl__EVAL_3;
  assign AsyncQueueSource__EVAL_0 = _EVAL_39;
  assign dmiXbar__EVAL_18 = dmi2tl__EVAL;
  assign asource__EVAL_27 = dmiXbar__EVAL_2;
  assign asource__EVAL_14 = dmiXbar__EVAL_4;
  assign _EVAL_18 = asource__EVAL_8;
  assign dmiXbar__EVAL_26 = dmOuter__EVAL_11;
  assign _EVAL_30 = asource__EVAL_19;
  assign dmOuter__EVAL_13 = dmiXbar__EVAL_19;
  assign dmiXbar__EVAL_1 = dmOuter__EVAL_17;
  assign _EVAL_3 = AsyncQueueSource__EVAL_3;
  assign dmiXbar__EVAL_22 = asource__EVAL_17;
  assign _EVAL_8 = asource__EVAL_28;
  assign asource__EVAL_9 = dmiXbar__EVAL_33;
  assign _EVAL_37 = asource__EVAL_2;
  assign asource__EVAL_11 = _EVAL_24;
  assign dmi2tl__EVAL_16 = dmiXbar__EVAL_12;
  assign _EVAL_34 = AsyncQueueSource__EVAL_8;
  assign _EVAL_0 = dmi2tl__EVAL_0;
  assign asource__EVAL_7 = _EVAL_27;
  assign _EVAL_5 = dmi2tl__EVAL_8;
  assign AsyncQueueSource__EVAL = dmOuter__EVAL_5;
  assign dmOuter__EVAL_9 = dmiXbar__EVAL_17;
  assign dmiXbar__EVAL_29 = dmi2tl__EVAL_6;
  assign asource__EVAL_30 = _EVAL_12;
  assign dmi2tl__EVAL_15 = dmiXbar__EVAL_23;
  assign dmiXbar__EVAL_10 = asource__EVAL_6;
  assign dmiXbar__EVAL_5 = dmOuter__EVAL_7;
  assign asource__EVAL_26 = dmiXbar__EVAL_37;
  assign _EVAL_23 = asource__EVAL_31;
  assign asource__EVAL_29 = _EVAL_15;
  assign dmiXbar__EVAL_3 = dmi2tl__EVAL_5;
  assign intsource__EVAL_0 = dmOuter__EVAL_18;
  assign dmiXbar__EVAL_0 = asource__EVAL_23;
  assign _EVAL_9 = AsyncQueueSource__EVAL_9;
  assign AsyncQueueSource__EVAL_5 = dmOuter__EVAL_3;
  assign asource__EVAL_10 = _EVAL_14;
  assign AsyncQueueSource__EVAL_14 = _EVAL_36;
  assign _EVAL_40 = dmi2tl__EVAL_9;
  assign _EVAL_21 = asource__EVAL_1;
  assign asource__EVAL_16 = dmiXbar__EVAL_30;
  assign asource__EVAL_20 = _EVAL_36;
  assign AsyncQueueSource__EVAL_13 = dmOuter__EVAL_6;
  assign dmi2tl__EVAL_18 = dmiXbar__EVAL_11;
  assign dmi2tl__EVAL_14 = dmiXbar__EVAL_34;
  assign dmOuter__EVAL_1 = dmiXbar__EVAL_28;
  assign dmOuter__EVAL_4 = _EVAL_36;
  assign dmiXbar__EVAL = asource__EVAL_32;
  assign asource__EVAL_12 = _EVAL_31;
  assign dmiXbar__EVAL_25 = asource__EVAL_15;
  assign _EVAL_22 = AsyncQueueSource__EVAL_2;
  assign dmiXbar__EVAL_13 = asource__EVAL_3;
  assign _EVAL_7 = asource__EVAL;
  assign dmi2tl__EVAL_13 = _EVAL_29;
  assign AsyncQueueSource__EVAL_4 = _EVAL_31;
  assign dmi2tl__EVAL_1 = _EVAL_4;
  assign AsyncQueueSource__EVAL_10 = dmOuter__EVAL;
  assign dmiXbar__EVAL_36 = _EVAL_36;
  assign AsyncQueueSource__EVAL_16 = dmOuter__EVAL_10;
  assign asource__EVAL_21 = dmiXbar__EVAL_16;
  assign dmi2tl__EVAL_11 = dmiXbar__EVAL_21;
  assign asource__EVAL_13 = _EVAL_19;
  assign dmiXbar__EVAL_32 = asource__EVAL_24;
  assign _EVAL_33 = dmOuter__EVAL_0;
endmodule
