//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_118(
  output        _EVAL,
  output [2:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  output [3:0]  _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  output [6:0]  _EVAL_10,
  output [29:0] _EVAL_11,
  input  [6:0]  _EVAL_12,
  output [31:0] _EVAL_13,
  input  [2:0]  _EVAL_14,
  output [2:0]  _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [29:0] _EVAL_17,
  input  [31:0] _EVAL_18,
  input         _EVAL_19,
  input  [3:0]  _EVAL_20
);
  reg  _EVAL_25 [0:1];
  reg [31:0] _RAND_0;
  wire  _EVAL_25__EVAL_26_data;
  wire  _EVAL_25__EVAL_26_addr;
  wire  _EVAL_25__EVAL_27_data;
  wire  _EVAL_25__EVAL_27_addr;
  wire  _EVAL_25__EVAL_27_mask;
  wire  _EVAL_25__EVAL_27_en;
  reg [6:0] _EVAL_29 [0:1];
  reg [31:0] _RAND_1;
  wire [6:0] _EVAL_29__EVAL_30_data;
  wire  _EVAL_29__EVAL_30_addr;
  wire [6:0] _EVAL_29__EVAL_31_data;
  wire  _EVAL_29__EVAL_31_addr;
  wire  _EVAL_29__EVAL_31_mask;
  wire  _EVAL_29__EVAL_31_en;
  reg [29:0] _EVAL_34 [0:1];
  reg [31:0] _RAND_2;
  wire [29:0] _EVAL_34__EVAL_35_data;
  wire  _EVAL_34__EVAL_35_addr;
  wire [29:0] _EVAL_34__EVAL_36_data;
  wire  _EVAL_34__EVAL_36_addr;
  wire  _EVAL_34__EVAL_36_mask;
  wire  _EVAL_34__EVAL_36_en;
  reg [2:0] _EVAL_38 [0:1];
  reg [31:0] _RAND_3;
  wire [2:0] _EVAL_38__EVAL_39_data;
  wire  _EVAL_38__EVAL_39_addr;
  wire [2:0] _EVAL_38__EVAL_40_data;
  wire  _EVAL_38__EVAL_40_addr;
  wire  _EVAL_38__EVAL_40_mask;
  wire  _EVAL_38__EVAL_40_en;
  reg [31:0] _EVAL_41 [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] _EVAL_41__EVAL_42_data;
  wire  _EVAL_41__EVAL_42_addr;
  wire [31:0] _EVAL_41__EVAL_43_data;
  wire  _EVAL_41__EVAL_43_addr;
  wire  _EVAL_41__EVAL_43_mask;
  wire  _EVAL_41__EVAL_43_en;
  reg [3:0] _EVAL_46 [0:1];
  reg [31:0] _RAND_5;
  wire [3:0] _EVAL_46__EVAL_47_data;
  wire  _EVAL_46__EVAL_47_addr;
  wire [3:0] _EVAL_46__EVAL_48_data;
  wire  _EVAL_46__EVAL_48_addr;
  wire  _EVAL_46__EVAL_48_mask;
  wire  _EVAL_46__EVAL_48_en;
  reg [2:0] _EVAL_53 [0:1];
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_53__EVAL_54_data;
  wire  _EVAL_53__EVAL_54_addr;
  wire [2:0] _EVAL_53__EVAL_55_data;
  wire  _EVAL_53__EVAL_55_addr;
  wire  _EVAL_53__EVAL_55_mask;
  wire  _EVAL_53__EVAL_55_en;
  reg [3:0] _EVAL_59 [0:1];
  reg [31:0] _RAND_7;
  wire [3:0] _EVAL_59__EVAL_60_data;
  wire  _EVAL_59__EVAL_60_addr;
  wire [3:0] _EVAL_59__EVAL_61_data;
  wire  _EVAL_59__EVAL_61_addr;
  wire  _EVAL_59__EVAL_61_mask;
  wire  _EVAL_59__EVAL_61_en;
  reg  _EVAL_33;
  reg [31:0] _RAND_8;
  reg  _EVAL_50;
  reg [31:0] _RAND_9;
  reg  _EVAL_58;
  reg [31:0] _RAND_10;
  wire  _EVAL_22;
  wire  _EVAL_57;
  wire  _EVAL_52;
  wire  _EVAL_49;
  wire  _EVAL_21;
  wire  _EVAL_44;
  wire  _EVAL_37;
  wire  _EVAL_51;
  wire  _EVAL_23;
  assign _EVAL_25__EVAL_26_addr = _EVAL_50;
  assign _EVAL_25__EVAL_26_data = _EVAL_25[_EVAL_25__EVAL_26_addr];
  assign _EVAL_25__EVAL_27_data = _EVAL_19;
  assign _EVAL_25__EVAL_27_addr = _EVAL_58;
  assign _EVAL_25__EVAL_27_mask = 1'h1;
  assign _EVAL_25__EVAL_27_en = _EVAL & _EVAL_8;
  assign _EVAL_29__EVAL_30_addr = _EVAL_50;
  assign _EVAL_29__EVAL_30_data = _EVAL_29[_EVAL_29__EVAL_30_addr];
  assign _EVAL_29__EVAL_31_data = _EVAL_12;
  assign _EVAL_29__EVAL_31_addr = _EVAL_58;
  assign _EVAL_29__EVAL_31_mask = 1'h1;
  assign _EVAL_29__EVAL_31_en = _EVAL & _EVAL_8;
  assign _EVAL_34__EVAL_35_addr = _EVAL_50;
  assign _EVAL_34__EVAL_35_data = _EVAL_34[_EVAL_34__EVAL_35_addr];
  assign _EVAL_34__EVAL_36_data = _EVAL_17;
  assign _EVAL_34__EVAL_36_addr = _EVAL_58;
  assign _EVAL_34__EVAL_36_mask = 1'h1;
  assign _EVAL_34__EVAL_36_en = _EVAL & _EVAL_8;
  assign _EVAL_38__EVAL_39_addr = _EVAL_50;
  assign _EVAL_38__EVAL_39_data = _EVAL_38[_EVAL_38__EVAL_39_addr];
  assign _EVAL_38__EVAL_40_data = _EVAL_5;
  assign _EVAL_38__EVAL_40_addr = _EVAL_58;
  assign _EVAL_38__EVAL_40_mask = 1'h1;
  assign _EVAL_38__EVAL_40_en = _EVAL & _EVAL_8;
  assign _EVAL_41__EVAL_42_addr = _EVAL_50;
  assign _EVAL_41__EVAL_42_data = _EVAL_41[_EVAL_41__EVAL_42_addr];
  assign _EVAL_41__EVAL_43_data = _EVAL_18;
  assign _EVAL_41__EVAL_43_addr = _EVAL_58;
  assign _EVAL_41__EVAL_43_mask = 1'h1;
  assign _EVAL_41__EVAL_43_en = _EVAL & _EVAL_8;
  assign _EVAL_46__EVAL_47_addr = _EVAL_50;
  assign _EVAL_46__EVAL_47_data = _EVAL_46[_EVAL_46__EVAL_47_addr];
  assign _EVAL_46__EVAL_48_data = _EVAL_1;
  assign _EVAL_46__EVAL_48_addr = _EVAL_58;
  assign _EVAL_46__EVAL_48_mask = 1'h1;
  assign _EVAL_46__EVAL_48_en = _EVAL & _EVAL_8;
  assign _EVAL_53__EVAL_54_addr = _EVAL_50;
  assign _EVAL_53__EVAL_54_data = _EVAL_53[_EVAL_53__EVAL_54_addr];
  assign _EVAL_53__EVAL_55_data = _EVAL_14;
  assign _EVAL_53__EVAL_55_addr = _EVAL_58;
  assign _EVAL_53__EVAL_55_mask = 1'h1;
  assign _EVAL_53__EVAL_55_en = _EVAL & _EVAL_8;
  assign _EVAL_59__EVAL_60_addr = _EVAL_50;
  assign _EVAL_59__EVAL_60_data = _EVAL_59[_EVAL_59__EVAL_60_addr];
  assign _EVAL_59__EVAL_61_data = _EVAL_20;
  assign _EVAL_59__EVAL_61_addr = _EVAL_58;
  assign _EVAL_59__EVAL_61_mask = 1'h1;
  assign _EVAL_59__EVAL_61_en = _EVAL & _EVAL_8;
  assign _EVAL_22 = _EVAL & _EVAL_8;
  assign _EVAL_57 = _EVAL_58 + 1'h1;
  assign _EVAL_52 = _EVAL_33 == 1'h0;
  assign _EVAL_49 = _EVAL_58 == _EVAL_50;
  assign _EVAL_21 = _EVAL_49 & _EVAL_33;
  assign _EVAL_44 = _EVAL_49 & _EVAL_52;
  assign _EVAL_37 = _EVAL_2 & _EVAL_9;
  assign _EVAL_51 = _EVAL_50 + 1'h1;
  assign _EVAL_23 = _EVAL_22 != _EVAL_37;
  assign _EVAL_15 = _EVAL_53__EVAL_54_data;
  assign _EVAL_16 = _EVAL_46__EVAL_47_data;
  assign _EVAL_4 = _EVAL_25__EVAL_26_data;
  assign _EVAL_7 = _EVAL_59__EVAL_60_data;
  assign _EVAL_9 = _EVAL_44 == 1'h0;
  assign _EVAL_0 = _EVAL_38__EVAL_39_data;
  assign _EVAL_13 = _EVAL_41__EVAL_42_data;
  assign _EVAL_11 = _EVAL_34__EVAL_35_data;
  assign _EVAL = _EVAL_21 == 1'h0;
  assign _EVAL_10 = _EVAL_29__EVAL_30_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_25[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_29[initvar] = _RAND_1[6:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_34[initvar] = _RAND_2[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_38[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_41[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_46[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_53[initvar] = _RAND_6[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_59[initvar] = _RAND_7[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_33 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_50 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_58 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if(_EVAL_25__EVAL_27_en & _EVAL_25__EVAL_27_mask) begin
      _EVAL_25[_EVAL_25__EVAL_27_addr] <= _EVAL_25__EVAL_27_data;
    end
    if(_EVAL_29__EVAL_31_en & _EVAL_29__EVAL_31_mask) begin
      _EVAL_29[_EVAL_29__EVAL_31_addr] <= _EVAL_29__EVAL_31_data;
    end
    if(_EVAL_34__EVAL_36_en & _EVAL_34__EVAL_36_mask) begin
      _EVAL_34[_EVAL_34__EVAL_36_addr] <= _EVAL_34__EVAL_36_data;
    end
    if(_EVAL_38__EVAL_40_en & _EVAL_38__EVAL_40_mask) begin
      _EVAL_38[_EVAL_38__EVAL_40_addr] <= _EVAL_38__EVAL_40_data;
    end
    if(_EVAL_41__EVAL_43_en & _EVAL_41__EVAL_43_mask) begin
      _EVAL_41[_EVAL_41__EVAL_43_addr] <= _EVAL_41__EVAL_43_data;
    end
    if(_EVAL_46__EVAL_48_en & _EVAL_46__EVAL_48_mask) begin
      _EVAL_46[_EVAL_46__EVAL_48_addr] <= _EVAL_46__EVAL_48_data;
    end
    if(_EVAL_53__EVAL_55_en & _EVAL_53__EVAL_55_mask) begin
      _EVAL_53[_EVAL_53__EVAL_55_addr] <= _EVAL_53__EVAL_55_data;
    end
    if(_EVAL_59__EVAL_61_en & _EVAL_59__EVAL_61_mask) begin
      _EVAL_59[_EVAL_59__EVAL_61_addr] <= _EVAL_59__EVAL_61_data;
    end
    if (_EVAL_6) begin
      _EVAL_33 <= 1'h0;
    end else begin
      if (_EVAL_23) begin
        _EVAL_33 <= _EVAL_22;
      end
    end
    if (_EVAL_6) begin
      _EVAL_50 <= 1'h0;
    end else begin
      if (_EVAL_37) begin
        _EVAL_50 <= _EVAL_51;
      end
    end
    if (_EVAL_6) begin
      _EVAL_58 <= 1'h0;
    end else begin
      if (_EVAL_22) begin
        _EVAL_58 <= _EVAL_57;
      end
    end
  end
endmodule
