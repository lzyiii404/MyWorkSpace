//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_57_assert(
  input  [1:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13
);
  wire [31:0] plusarg_reader_out;
  reg [7:0] _EVAL_22;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_29;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_49;
  reg [31:0] _RAND_2;
  reg  _EVAL_50;
  reg [31:0] _RAND_3;
  reg  _EVAL_64;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_95;
  reg [31:0] _RAND_5;
  reg [1:0] _EVAL_111;
  reg [31:0] _RAND_6;
  reg [7:0] _EVAL_123;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_136;
  reg [31:0] _RAND_8;
  reg [7:0] _EVAL_163;
  reg [31:0] _RAND_9;
  reg  _EVAL_171;
  reg [31:0] _RAND_10;
  reg [7:0] _EVAL_175;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_192;
  reg [31:0] _RAND_12;
  reg [3:0] _EVAL_230;
  reg [31:0] _RAND_13;
  wire [22:0] _EVAL_193;
  wire [7:0] _EVAL_74;
  wire [7:0] _EVAL_99;
  wire [31:0] _EVAL_128;
  wire  _EVAL_81;
  wire  _EVAL_232;
  wire [22:0] _EVAL_26;
  wire [7:0] _EVAL_127;
  wire  _EVAL_27;
  wire  _EVAL_139;
  wire  _EVAL_235;
  wire [1:0] _EVAL_150;
  wire  _EVAL_200;
  wire  _EVAL_248;
  wire  _EVAL_17;
  wire  _EVAL_59;
  wire  _EVAL_141;
  wire  _EVAL_207;
  wire  _EVAL_164;
  wire  _EVAL_183;
  wire  _EVAL_158;
  wire  _EVAL_78;
  wire  _EVAL_166;
  wire  _EVAL_54;
  wire  _EVAL_80;
  wire [31:0] _EVAL_209;
  wire [32:0] _EVAL_144;
  wire [32:0] _EVAL_204;
  wire [32:0] _EVAL_23;
  wire  _EVAL_110;
  wire [31:0] _EVAL_90;
  wire [32:0] _EVAL_96;
  wire [32:0] _EVAL_221;
  wire [32:0] _EVAL_58;
  wire  _EVAL_212;
  wire  _EVAL_69;
  wire [31:0] _EVAL_122;
  wire [32:0] _EVAL_214;
  wire [32:0] _EVAL_63;
  wire [32:0] _EVAL_180;
  wire  _EVAL_182;
  wire  _EVAL_129;
  wire [31:0] _EVAL_151;
  wire [32:0] _EVAL_70;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_244;
  wire  _EVAL_233;
  wire  _EVAL_229;
  wire [32:0] _EVAL_93;
  wire [32:0] _EVAL_20;
  wire [32:0] _EVAL_145;
  wire  _EVAL_16;
  wire  _EVAL_223;
  wire [31:0] _EVAL_219;
  wire [32:0] _EVAL_135;
  wire [32:0] _EVAL_112;
  wire [32:0] _EVAL_14;
  wire  _EVAL_60;
  wire  _EVAL_126;
  wire [31:0] _EVAL_224;
  wire [32:0] _EVAL_198;
  wire [32:0] _EVAL_92;
  wire [32:0] _EVAL_234;
  wire  _EVAL_117;
  wire  _EVAL_132;
  wire  _EVAL_238;
  wire  _EVAL_47;
  wire  _EVAL_240;
  wire  _EVAL_30;
  wire [7:0] _EVAL_91;
  wire [7:0] _EVAL_157;
  wire  _EVAL_170;
  wire  _EVAL_21;
  wire  _EVAL_218;
  wire  _EVAL_124;
  wire  _EVAL_86;
  wire  _EVAL_191;
  wire [31:0] _EVAL_153;
  wire [32:0] _EVAL_173;
  wire [32:0] _EVAL_84;
  wire [32:0] _EVAL_185;
  wire  _EVAL_137;
  wire  _EVAL_168;
  wire [31:0] _EVAL_53;
  wire [32:0] _EVAL_205;
  wire [32:0] _EVAL_42;
  wire [32:0] _EVAL_249;
  wire  _EVAL_113;
  wire  _EVAL_105;
  wire  _EVAL_85;
  wire  _EVAL_40;
  wire  _EVAL_149;
  wire  _EVAL_215;
  wire  _EVAL_15;
  wire [1:0] _EVAL_206;
  wire  _EVAL_125;
  wire  _EVAL_134;
  wire  _EVAL_188;
  wire  _EVAL_174;
  wire  _EVAL_41;
  wire  _EVAL_82;
  wire  _EVAL_242;
  wire  _EVAL_138;
  wire  _EVAL_56;
  wire  _EVAL_118;
  wire  _EVAL_33;
  wire  _EVAL_208;
  wire [31:0] _EVAL_246;
  wire  _EVAL_156;
  wire  _EVAL_48;
  wire  _EVAL_36;
  wire  _EVAL_176;
  wire  _EVAL_19;
  wire  _EVAL_34;
  wire  _EVAL_31;
  wire  _EVAL_222;
  wire  _EVAL_190;
  wire  _EVAL_140;
  wire [7:0] _EVAL_226;
  wire  _EVAL_44;
  wire  _EVAL_24;
  wire  _EVAL_203;
  wire  _EVAL_245;
  wire  _EVAL_195;
  wire  _EVAL_243;
  wire  _EVAL_220;
  wire  _EVAL_202;
  wire  _EVAL_179;
  wire  _EVAL_43;
  wire  _EVAL_160;
  wire  _EVAL_101;
  wire  _EVAL_186;
  wire  _EVAL_216;
  wire  _EVAL_148;
  wire  _EVAL_250;
  wire [7:0] _EVAL_142;
  wire  _EVAL_109;
  wire  _EVAL_131;
  wire  _EVAL_94;
  wire  _EVAL_154;
  wire  _EVAL_228;
  wire  _EVAL_217;
  wire  _EVAL_167;
  wire  _EVAL_102;
  wire  _EVAL_107;
  wire  _EVAL_51;
  wire  _EVAL_87;
  wire  _EVAL_227;
  wire  _EVAL_119;
  wire  _EVAL_239;
  wire  _EVAL_199;
  wire  _EVAL_52;
  wire  _EVAL_210;
  wire  _EVAL_196;
  wire [7:0] _EVAL_165;
  wire  _EVAL_147;
  wire  _EVAL_35;
  wire  _EVAL_62;
  wire  _EVAL_65;
  wire  _EVAL_55;
  wire  _EVAL_120;
  wire  _EVAL_38;
  wire  _EVAL_152;
  wire [31:0] _EVAL_37;
  wire  _EVAL_177;
  wire  _EVAL_211;
  wire  _EVAL_100;
  wire  _EVAL_72;
  wire  _EVAL_213;
  wire  _EVAL_25;
  wire  _EVAL_241;
  wire  _EVAL_98;
  wire  _EVAL_61;
  wire  _EVAL_79;
  wire  _EVAL_32;
  wire  _EVAL_187;
  wire  _EVAL_184;
  wire  _EVAL_133;
  wire  _EVAL_68;
  wire  _EVAL_108;
  wire  _EVAL_130;
  wire  _EVAL_28;
  wire  _EVAL_161;
  wire  _EVAL_106;
  wire  _EVAL_116;
  wire  _EVAL_236;
  wire  _EVAL_162;
  wire  _EVAL_197;
  wire  _EVAL_143;
  wire  _EVAL_225;
  wire  _EVAL_121;
  wire  _EVAL_83;
  wire  _EVAL_194;
  wire  _EVAL_169;
  wire  _EVAL_66;
  wire  _EVAL_18;
  wire  _EVAL_114;
  wire  _EVAL_77;
  wire  _EVAL_247;
  wire  _EVAL_189;
  wire  _EVAL_146;
  wire  _EVAL_88;
  wire  _EVAL_103;
  wire  _EVAL_46;
  wire  _EVAL_89;
  wire  _EVAL_104;
  wire  _EVAL_67;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_193 = 23'hff << _EVAL_2;
  assign _EVAL_74 = _EVAL_193[7:0];
  assign _EVAL_99 = ~ _EVAL_74;
  assign _EVAL_128 = {{24'd0}, _EVAL_99};
  assign _EVAL_81 = _EVAL <= 2'h2;
  assign _EVAL_232 = _EVAL_8 == _EVAL_136;
  assign _EVAL_26 = 23'hff << _EVAL_8;
  assign _EVAL_127 = _EVAL_26[7:0];
  assign _EVAL_27 = _EVAL_11 & _EVAL_10;
  assign _EVAL_139 = _EVAL_123 == 8'h0;
  assign _EVAL_235 = _EVAL_27 & _EVAL_139;
  assign _EVAL_150 = _EVAL_235 ? 2'h1 : 2'h0;
  assign _EVAL_200 = _EVAL_150[0];
  assign _EVAL_248 = _EVAL_200 | _EVAL_50;
  assign _EVAL_17 = _EVAL_248 | _EVAL_4;
  assign _EVAL_59 = _EVAL_50 == 1'h0;
  assign _EVAL_141 = plusarg_reader_out == 32'h0;
  assign _EVAL_207 = _EVAL_59 | _EVAL_141;
  assign _EVAL_164 = _EVAL_192 < plusarg_reader_out;
  assign _EVAL_183 = _EVAL_207 | _EVAL_164;
  assign _EVAL_158 = _EVAL_183 | _EVAL_4;
  assign _EVAL_78 = _EVAL_158 == 1'h0;
  assign _EVAL_166 = _EVAL_5[2];
  assign _EVAL_54 = _EVAL_166 == 1'h0;
  assign _EVAL_80 = _EVAL_7 <= 3'h6;
  assign _EVAL_209 = _EVAL_3 ^ 32'h40000000;
  assign _EVAL_144 = {1'b0,$signed(_EVAL_209)};
  assign _EVAL_204 = $signed(_EVAL_144) & $signed(-33'sh2000);
  assign _EVAL_23 = $signed(_EVAL_204);
  assign _EVAL_110 = $signed(_EVAL_23) == $signed(33'sh0);
  assign _EVAL_90 = _EVAL_3 ^ 32'h80000000;
  assign _EVAL_96 = {1'b0,$signed(_EVAL_90)};
  assign _EVAL_221 = $signed(_EVAL_96) & $signed(-33'sh20000);
  assign _EVAL_58 = $signed(_EVAL_221);
  assign _EVAL_212 = $signed(_EVAL_58) == $signed(33'sh0);
  assign _EVAL_69 = _EVAL_110 | _EVAL_212;
  assign _EVAL_122 = _EVAL_3 ^ 32'hc000000;
  assign _EVAL_214 = {1'b0,$signed(_EVAL_122)};
  assign _EVAL_63 = $signed(_EVAL_214) & $signed(-33'sh4000000);
  assign _EVAL_180 = $signed(_EVAL_63);
  assign _EVAL_182 = $signed(_EVAL_180) == $signed(33'sh0);
  assign _EVAL_129 = _EVAL_69 | _EVAL_182;
  assign _EVAL_151 = _EVAL_3 ^ 32'h2000000;
  assign _EVAL_70 = {1'b0,$signed(_EVAL_151)};
  assign _EVAL_172 = $signed(_EVAL_70) & $signed(-33'sh10000);
  assign _EVAL_244 = $signed(_EVAL_172);
  assign _EVAL_233 = $signed(_EVAL_244) == $signed(33'sh0);
  assign _EVAL_229 = _EVAL_129 | _EVAL_233;
  assign _EVAL_93 = {1'b0,$signed(_EVAL_3)};
  assign _EVAL_20 = $signed(_EVAL_93) & $signed(-33'sh5000);
  assign _EVAL_145 = $signed(_EVAL_20);
  assign _EVAL_16 = $signed(_EVAL_145) == $signed(33'sh0);
  assign _EVAL_223 = _EVAL_229 | _EVAL_16;
  assign _EVAL_219 = _EVAL_3 ^ 32'h1800000;
  assign _EVAL_135 = {1'b0,$signed(_EVAL_219)};
  assign _EVAL_112 = $signed(_EVAL_135) & $signed(-33'sh8000);
  assign _EVAL_14 = $signed(_EVAL_112);
  assign _EVAL_60 = $signed(_EVAL_14) == $signed(33'sh0);
  assign _EVAL_126 = _EVAL_223 | _EVAL_60;
  assign _EVAL_224 = _EVAL_3 ^ 32'h3000;
  assign _EVAL_198 = {1'b0,$signed(_EVAL_224)};
  assign _EVAL_92 = $signed(_EVAL_198) & $signed(-33'sh1000);
  assign _EVAL_234 = $signed(_EVAL_92);
  assign _EVAL_117 = $signed(_EVAL_234) == $signed(33'sh0);
  assign _EVAL_132 = _EVAL_13 == 1'h0;
  assign _EVAL_238 = _EVAL_132 | _EVAL_9;
  assign _EVAL_47 = _EVAL_0 & _EVAL_6;
  assign _EVAL_240 = _EVAL_22 == 8'h0;
  assign _EVAL_30 = _EVAL_7[0];
  assign _EVAL_91 = ~ _EVAL_127;
  assign _EVAL_157 = _EVAL_22 - 8'h1;
  assign _EVAL_170 = _EVAL != 2'h2;
  assign _EVAL_21 = _EVAL_170 | _EVAL_4;
  assign _EVAL_218 = _EVAL_132 | _EVAL_4;
  assign _EVAL_124 = _EVAL_2 == _EVAL_230;
  assign _EVAL_86 = _EVAL_7 == 3'h5;
  assign _EVAL_191 = _EVAL_2 <= 4'h6;
  assign _EVAL_153 = _EVAL_3 ^ 32'h1900000;
  assign _EVAL_173 = {1'b0,$signed(_EVAL_153)};
  assign _EVAL_84 = $signed(_EVAL_173) & $signed(-33'sh2000);
  assign _EVAL_185 = $signed(_EVAL_84);
  assign _EVAL_137 = $signed(_EVAL_185) == $signed(33'sh0);
  assign _EVAL_168 = _EVAL_126 | _EVAL_137;
  assign _EVAL_53 = _EVAL_3 ^ 32'h20000000;
  assign _EVAL_205 = {1'b0,$signed(_EVAL_53)};
  assign _EVAL_42 = $signed(_EVAL_205) & $signed(-33'sh2000);
  assign _EVAL_249 = $signed(_EVAL_42);
  assign _EVAL_113 = $signed(_EVAL_249) == $signed(33'sh0);
  assign _EVAL_105 = _EVAL_168 | _EVAL_113;
  assign _EVAL_85 = _EVAL_191 & _EVAL_105;
  assign _EVAL_40 = _EVAL_47 & _EVAL_240;
  assign _EVAL_149 = _EVAL_7 == 3'h6;
  assign _EVAL_215 = _EVAL_149 == 1'h0;
  assign _EVAL_15 = _EVAL_40 & _EVAL_215;
  assign _EVAL_206 = _EVAL_15 ? 2'h1 : 2'h0;
  assign _EVAL_125 = _EVAL_13 == _EVAL_171;
  assign _EVAL_134 = _EVAL_125 | _EVAL_4;
  assign _EVAL_188 = _EVAL_134 == 1'h0;
  assign _EVAL_174 = _EVAL_12 == _EVAL_64;
  assign _EVAL_41 = _EVAL_174 | _EVAL_4;
  assign _EVAL_82 = _EVAL_5 == 3'h6;
  assign _EVAL_242 = _EVAL_10 & _EVAL_82;
  assign _EVAL_138 = _EVAL_6 & _EVAL_86;
  assign _EVAL_56 = _EVAL_175 == 8'h0;
  assign _EVAL_118 = _EVAL_7 == _EVAL_49;
  assign _EVAL_33 = _EVAL_5 == 3'h0;
  assign _EVAL_208 = _EVAL_163 == 8'h0;
  assign _EVAL_246 = _EVAL_3 & _EVAL_128;
  assign _EVAL_156 = _EVAL_246 == 32'h0;
  assign _EVAL_48 = _EVAL_5 == 3'h4;
  assign _EVAL_36 = _EVAL_10 & _EVAL_48;
  assign _EVAL_176 = _EVAL == _EVAL_111;
  assign _EVAL_19 = _EVAL_176 | _EVAL_4;
  assign _EVAL_34 = _EVAL_19 == 1'h0;
  assign _EVAL_31 = _EVAL == 2'h0;
  assign _EVAL_222 = _EVAL_31 | _EVAL_4;
  assign _EVAL_190 = _EVAL_238 | _EVAL_4;
  assign _EVAL_140 = _EVAL_190 == 1'h0;
  assign _EVAL_226 = _EVAL_175 - 8'h1;
  assign _EVAL_44 = _EVAL_80 | _EVAL_4;
  assign _EVAL_24 = _EVAL_44 == 1'h0;
  assign _EVAL_203 = _EVAL_117 | _EVAL_182;
  assign _EVAL_245 = _EVAL_203 | _EVAL_233;
  assign _EVAL_195 = _EVAL_245 | _EVAL_16;
  assign _EVAL_243 = _EVAL_195 | _EVAL_60;
  assign _EVAL_220 = _EVAL_243 | _EVAL_137;
  assign _EVAL_202 = _EVAL_220 | _EVAL_113;
  assign _EVAL_179 = _EVAL_7 == 3'h1;
  assign _EVAL_43 = _EVAL_6 & _EVAL_179;
  assign _EVAL_160 = _EVAL_2 <= 4'h8;
  assign _EVAL_101 = _EVAL_160 & _EVAL_117;
  assign _EVAL_186 = _EVAL_101 | _EVAL_4;
  assign _EVAL_216 = _EVAL_186 == 1'h0;
  assign _EVAL_148 = _EVAL_124 | _EVAL_4;
  assign _EVAL_250 = _EVAL_148 == 1'h0;
  assign _EVAL_142 = _EVAL_163 - 8'h1;
  assign _EVAL_109 = _EVAL_191 & _EVAL_212;
  assign _EVAL_131 = _EVAL_109 | _EVAL_4;
  assign _EVAL_94 = _EVAL_2 <= 4'h2;
  assign _EVAL_154 = _EVAL_94 & _EVAL_202;
  assign _EVAL_228 = _EVAL_154 | _EVAL_4;
  assign _EVAL_217 = _EVAL_5 == _EVAL_95;
  assign _EVAL_167 = _EVAL_156 | _EVAL_4;
  assign _EVAL_102 = _EVAL_167 == 1'h0;
  assign _EVAL_107 = _EVAL_59 | _EVAL_4;
  assign _EVAL_51 = _EVAL_107 == 1'h0;
  assign _EVAL_87 = _EVAL_5 == 3'h7;
  assign _EVAL_227 = _EVAL_10 & _EVAL_87;
  assign _EVAL_119 = _EVAL_5 == 3'h3;
  assign _EVAL_239 = _EVAL_56 == 1'h0;
  assign _EVAL_199 = _EVAL_10 & _EVAL_239;
  assign _EVAL_52 = _EVAL_4 == 1'h0;
  assign _EVAL_210 = _EVAL_27 & _EVAL_56;
  assign _EVAL_196 = _EVAL_232 | _EVAL_4;
  assign _EVAL_165 = _EVAL_123 - 8'h1;
  assign _EVAL_147 = _EVAL_7 == 3'h0;
  assign _EVAL_35 = _EVAL_6 & _EVAL_147;
  assign _EVAL_62 = _EVAL_206[0];
  assign _EVAL_65 = ~ _EVAL_62;
  assign _EVAL_55 = _EVAL_5 == 3'h1;
  assign _EVAL_120 = _EVAL_85 | _EVAL_101;
  assign _EVAL_38 = _EVAL_120 | _EVAL_4;
  assign _EVAL_152 = _EVAL_38 == 1'h0;
  assign _EVAL_37 = _EVAL_192 + 32'h1;
  assign _EVAL_177 = _EVAL_81 | _EVAL_4;
  assign _EVAL_211 = _EVAL_5 == 3'h5;
  assign _EVAL_100 = _EVAL_9 == 1'h0;
  assign _EVAL_72 = _EVAL_100 | _EVAL_4;
  assign _EVAL_213 = _EVAL_72 == 1'h0;
  assign _EVAL_25 = _EVAL_10 & _EVAL_55;
  assign _EVAL_241 = _EVAL_7 == 3'h2;
  assign _EVAL_98 = _EVAL_6 & _EVAL_241;
  assign _EVAL_61 = _EVAL_3 == _EVAL_29;
  assign _EVAL_79 = _EVAL_61 | _EVAL_4;
  assign _EVAL_32 = _EVAL_79 == 1'h0;
  assign _EVAL_187 = _EVAL_200 != _EVAL_62;
  assign _EVAL_184 = _EVAL_200 == 1'h0;
  assign _EVAL_133 = _EVAL_187 | _EVAL_184;
  assign _EVAL_68 = _EVAL_133 | _EVAL_4;
  assign _EVAL_108 = _EVAL_7 == 3'h4;
  assign _EVAL_130 = _EVAL_6 & _EVAL_108;
  assign _EVAL_28 = _EVAL_10 & _EVAL_33;
  assign _EVAL_161 = _EVAL_131 == 1'h0;
  assign _EVAL_106 = _EVAL_21 == 1'h0;
  assign _EVAL_116 = _EVAL_5 == 3'h2;
  assign _EVAL_236 = _EVAL_27 | _EVAL_47;
  assign _EVAL_162 = _EVAL_218 == 1'h0;
  assign _EVAL_197 = _EVAL_17 == 1'h0;
  assign _EVAL_143 = _EVAL_208 == 1'h0;
  assign _EVAL_225 = _EVAL_6 & _EVAL_143;
  assign _EVAL_121 = _EVAL_47 & _EVAL_208;
  assign _EVAL_83 = _EVAL_10 & _EVAL_119;
  assign _EVAL_194 = _EVAL_68 == 1'h0;
  assign _EVAL_169 = _EVAL_118 | _EVAL_4;
  assign _EVAL_66 = _EVAL_10 & _EVAL_211;
  assign _EVAL_18 = _EVAL_217 | _EVAL_4;
  assign _EVAL_114 = _EVAL_41 == 1'h0;
  assign _EVAL_77 = _EVAL_169 == 1'h0;
  assign _EVAL_247 = _EVAL_228 == 1'h0;
  assign _EVAL_189 = _EVAL_10 & _EVAL_116;
  assign _EVAL_146 = _EVAL_6 & _EVAL_149;
  assign _EVAL_88 = _EVAL_196 == 1'h0;
  assign _EVAL_103 = _EVAL_222 == 1'h0;
  assign _EVAL_46 = _EVAL_50 | _EVAL_200;
  assign _EVAL_89 = _EVAL_177 == 1'h0;
  assign _EVAL_104 = _EVAL_18 == 1'h0;
  assign _EVAL_67 = _EVAL_46 & _EVAL_65;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_29 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_49 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_50 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_64 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_95 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_111 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_123 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_136 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_163 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_171 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_175 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_192 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_230 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_1) begin
    if (_EVAL_4) begin
      _EVAL_22 <= 8'h0;
    end else begin
      if (_EVAL_47) begin
        if (_EVAL_240) begin
          if (_EVAL_30) begin
            _EVAL_22 <= _EVAL_91;
          end else begin
            _EVAL_22 <= 8'h0;
          end
        end else begin
          _EVAL_22 <= _EVAL_157;
        end
      end
    end
    if (_EVAL_210) begin
      _EVAL_29 <= _EVAL_3;
    end
    if (_EVAL_121) begin
      _EVAL_49 <= _EVAL_7;
    end
    if (_EVAL_4) begin
      _EVAL_50 <= 1'h0;
    end else begin
      _EVAL_50 <= _EVAL_67;
    end
    if (_EVAL_121) begin
      _EVAL_64 <= _EVAL_12;
    end
    if (_EVAL_210) begin
      _EVAL_95 <= _EVAL_5;
    end
    if (_EVAL_121) begin
      _EVAL_111 <= _EVAL;
    end
    if (_EVAL_4) begin
      _EVAL_123 <= 8'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_139) begin
          if (_EVAL_54) begin
            _EVAL_123 <= _EVAL_99;
          end else begin
            _EVAL_123 <= 8'h0;
          end
        end else begin
          _EVAL_123 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_121) begin
      _EVAL_136 <= _EVAL_8;
    end
    if (_EVAL_4) begin
      _EVAL_163 <= 8'h0;
    end else begin
      if (_EVAL_47) begin
        if (_EVAL_208) begin
          if (_EVAL_30) begin
            _EVAL_163 <= _EVAL_91;
          end else begin
            _EVAL_163 <= 8'h0;
          end
        end else begin
          _EVAL_163 <= _EVAL_142;
        end
      end
    end
    if (_EVAL_121) begin
      _EVAL_171 <= _EVAL_13;
    end
    if (_EVAL_4) begin
      _EVAL_175 <= 8'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_56) begin
          if (_EVAL_54) begin
            _EVAL_175 <= _EVAL_99;
          end else begin
            _EVAL_175 <= 8'h0;
          end
        end else begin
          _EVAL_175 <= _EVAL_226;
        end
      end
    end
    if (_EVAL_4) begin
      _EVAL_192 <= 32'h0;
    end else begin
      if (_EVAL_236) begin
        _EVAL_192 <= 32'h0;
      end else begin
        _EVAL_192 <= _EVAL_37;
      end
    end
    if (_EVAL_210) begin
      _EVAL_230 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aba5c87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26bf0517)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3caeb5c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87910c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aab5b251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f78d4d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(289e9728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c11a534f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc74add)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddaf159d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a8c9219)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61ce576b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a29c4c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f08085d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0a4351c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45a60689)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e11b361)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd9bbc86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1713f12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7af43b14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64303b39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92464967)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(168727a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(100831f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c36b3229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d69fe8c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26a7eb75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55ba73cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8856b367)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33d05e5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59bbd623)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cf84de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(505dfc94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff4da08d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83fc6776)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa2068bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc7b686)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50e12691)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a724b6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fc5d0cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1be1846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8451c46d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(571d360a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15f279d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ac25b35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26db2826)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59184d9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
