//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_119(
  output        _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output [2:0]  _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  output [6:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input  [31:0] _EVAL_11,
  output [1:0]  _EVAL_12,
  output [3:0]  _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  input  [6:0]  _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18,
  output        _EVAL_19,
  output [31:0] _EVAL_20
);
  reg  _EVAL_23 [0:1];
  reg [31:0] _RAND_0;
  wire  _EVAL_23__EVAL_24_data;
  wire  _EVAL_23__EVAL_24_addr;
  wire  _EVAL_23__EVAL_25_data;
  wire  _EVAL_23__EVAL_25_addr;
  wire  _EVAL_23__EVAL_25_mask;
  wire  _EVAL_23__EVAL_25_en;
  reg [6:0] _EVAL_27 [0:1];
  reg [31:0] _RAND_1;
  wire [6:0] _EVAL_27__EVAL_28_data;
  wire  _EVAL_27__EVAL_28_addr;
  wire [6:0] _EVAL_27__EVAL_29_data;
  wire  _EVAL_27__EVAL_29_addr;
  wire  _EVAL_27__EVAL_29_mask;
  wire  _EVAL_27__EVAL_29_en;
  reg [31:0] _EVAL_30 [0:1];
  reg [31:0] _RAND_2;
  wire [31:0] _EVAL_30__EVAL_31_data;
  wire  _EVAL_30__EVAL_31_addr;
  wire [31:0] _EVAL_30__EVAL_32_data;
  wire  _EVAL_30__EVAL_32_addr;
  wire  _EVAL_30__EVAL_32_mask;
  wire  _EVAL_30__EVAL_32_en;
  reg [3:0] _EVAL_35 [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] _EVAL_35__EVAL_36_data;
  wire  _EVAL_35__EVAL_36_addr;
  wire [3:0] _EVAL_35__EVAL_37_data;
  wire  _EVAL_35__EVAL_37_addr;
  wire  _EVAL_35__EVAL_37_mask;
  wire  _EVAL_35__EVAL_37_en;
  reg  _EVAL_44 [0:1];
  reg [31:0] _RAND_4;
  wire  _EVAL_44__EVAL_45_data;
  wire  _EVAL_44__EVAL_45_addr;
  wire  _EVAL_44__EVAL_46_data;
  wire  _EVAL_44__EVAL_46_addr;
  wire  _EVAL_44__EVAL_46_mask;
  wire  _EVAL_44__EVAL_46_en;
  reg  _EVAL_49 [0:1];
  reg [31:0] _RAND_5;
  wire  _EVAL_49__EVAL_50_data;
  wire  _EVAL_49__EVAL_50_addr;
  wire  _EVAL_49__EVAL_51_data;
  wire  _EVAL_49__EVAL_51_addr;
  wire  _EVAL_49__EVAL_51_mask;
  wire  _EVAL_49__EVAL_51_en;
  reg [1:0] _EVAL_52 [0:1];
  reg [31:0] _RAND_6;
  wire [1:0] _EVAL_52__EVAL_53_data;
  wire  _EVAL_52__EVAL_53_addr;
  wire [1:0] _EVAL_52__EVAL_54_data;
  wire  _EVAL_52__EVAL_54_addr;
  wire  _EVAL_52__EVAL_54_mask;
  wire  _EVAL_52__EVAL_54_en;
  reg [2:0] _EVAL_57 [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire [2:0] _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  reg  _EVAL_21;
  reg [31:0] _RAND_8;
  reg  _EVAL_22;
  reg [31:0] _RAND_9;
  reg  _EVAL_33;
  reg [31:0] _RAND_10;
  wire  _EVAL_42;
  wire  _EVAL_61;
  wire  _EVAL_26;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_48;
  wire  _EVAL_34;
  wire  _EVAL_55;
  wire  _EVAL_60;
  assign _EVAL_23__EVAL_24_addr = _EVAL_21;
  assign _EVAL_23__EVAL_24_data = _EVAL_23[_EVAL_23__EVAL_24_addr];
  assign _EVAL_23__EVAL_25_data = _EVAL_5;
  assign _EVAL_23__EVAL_25_addr = _EVAL_22;
  assign _EVAL_23__EVAL_25_mask = 1'h1;
  assign _EVAL_23__EVAL_25_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_27__EVAL_28_addr = _EVAL_21;
  assign _EVAL_27__EVAL_28_data = _EVAL_27[_EVAL_27__EVAL_28_addr];
  assign _EVAL_27__EVAL_29_data = _EVAL_16;
  assign _EVAL_27__EVAL_29_addr = _EVAL_22;
  assign _EVAL_27__EVAL_29_mask = 1'h1;
  assign _EVAL_27__EVAL_29_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_30__EVAL_31_addr = _EVAL_21;
  assign _EVAL_30__EVAL_31_data = _EVAL_30[_EVAL_30__EVAL_31_addr];
  assign _EVAL_30__EVAL_32_data = _EVAL_11;
  assign _EVAL_30__EVAL_32_addr = _EVAL_22;
  assign _EVAL_30__EVAL_32_mask = 1'h1;
  assign _EVAL_30__EVAL_32_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_35__EVAL_36_addr = _EVAL_21;
  assign _EVAL_35__EVAL_36_data = _EVAL_35[_EVAL_35__EVAL_36_addr];
  assign _EVAL_35__EVAL_37_data = _EVAL_8;
  assign _EVAL_35__EVAL_37_addr = _EVAL_22;
  assign _EVAL_35__EVAL_37_mask = 1'h1;
  assign _EVAL_35__EVAL_37_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_44__EVAL_45_addr = _EVAL_21;
  assign _EVAL_44__EVAL_45_data = _EVAL_44[_EVAL_44__EVAL_45_addr];
  assign _EVAL_44__EVAL_46_data = _EVAL_15;
  assign _EVAL_44__EVAL_46_addr = _EVAL_22;
  assign _EVAL_44__EVAL_46_mask = 1'h1;
  assign _EVAL_44__EVAL_46_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_49__EVAL_50_addr = _EVAL_21;
  assign _EVAL_49__EVAL_50_data = _EVAL_49[_EVAL_49__EVAL_50_addr];
  assign _EVAL_49__EVAL_51_data = _EVAL_1;
  assign _EVAL_49__EVAL_51_addr = _EVAL_22;
  assign _EVAL_49__EVAL_51_mask = 1'h1;
  assign _EVAL_49__EVAL_51_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_52__EVAL_53_addr = _EVAL_21;
  assign _EVAL_52__EVAL_53_data = _EVAL_52[_EVAL_52__EVAL_53_addr];
  assign _EVAL_52__EVAL_54_data = _EVAL_6;
  assign _EVAL_52__EVAL_54_addr = _EVAL_22;
  assign _EVAL_52__EVAL_54_mask = 1'h1;
  assign _EVAL_52__EVAL_54_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_57__EVAL_58_addr = _EVAL_21;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_18;
  assign _EVAL_57__EVAL_59_addr = _EVAL_22;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_19 & _EVAL_10;
  assign _EVAL_42 = _EVAL_22 == _EVAL_21;
  assign _EVAL_61 = _EVAL_19 & _EVAL_10;
  assign _EVAL_26 = _EVAL_33 == 1'h0;
  assign _EVAL_40 = _EVAL_42 & _EVAL_26;
  assign _EVAL_41 = _EVAL_4 & _EVAL_9;
  assign _EVAL_48 = _EVAL_61 != _EVAL_41;
  assign _EVAL_34 = _EVAL_21 + 1'h1;
  assign _EVAL_55 = _EVAL_22 + 1'h1;
  assign _EVAL_60 = _EVAL_42 & _EVAL_33;
  assign _EVAL_19 = _EVAL_60 == 1'h0;
  assign _EVAL_7 = _EVAL_27__EVAL_28_data;
  assign _EVAL = _EVAL_44__EVAL_45_data;
  assign _EVAL_20 = _EVAL_30__EVAL_31_data;
  assign _EVAL_13 = _EVAL_35__EVAL_36_data;
  assign _EVAL_14 = _EVAL_49__EVAL_50_data;
  assign _EVAL_9 = _EVAL_40 == 1'h0;
  assign _EVAL_3 = _EVAL_23__EVAL_24_data;
  assign _EVAL_2 = _EVAL_57__EVAL_58_data;
  assign _EVAL_12 = _EVAL_52__EVAL_53_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_23[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_27[initvar] = _RAND_1[6:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_30[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_35[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_44[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_49[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_52[initvar] = _RAND_6[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_21 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_22 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_33 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_17) begin
    if(_EVAL_23__EVAL_25_en & _EVAL_23__EVAL_25_mask) begin
      _EVAL_23[_EVAL_23__EVAL_25_addr] <= _EVAL_23__EVAL_25_data;
    end
    if(_EVAL_27__EVAL_29_en & _EVAL_27__EVAL_29_mask) begin
      _EVAL_27[_EVAL_27__EVAL_29_addr] <= _EVAL_27__EVAL_29_data;
    end
    if(_EVAL_30__EVAL_32_en & _EVAL_30__EVAL_32_mask) begin
      _EVAL_30[_EVAL_30__EVAL_32_addr] <= _EVAL_30__EVAL_32_data;
    end
    if(_EVAL_35__EVAL_37_en & _EVAL_35__EVAL_37_mask) begin
      _EVAL_35[_EVAL_35__EVAL_37_addr] <= _EVAL_35__EVAL_37_data;
    end
    if(_EVAL_44__EVAL_46_en & _EVAL_44__EVAL_46_mask) begin
      _EVAL_44[_EVAL_44__EVAL_46_addr] <= _EVAL_44__EVAL_46_data;
    end
    if(_EVAL_49__EVAL_51_en & _EVAL_49__EVAL_51_mask) begin
      _EVAL_49[_EVAL_49__EVAL_51_addr] <= _EVAL_49__EVAL_51_data;
    end
    if(_EVAL_52__EVAL_54_en & _EVAL_52__EVAL_54_mask) begin
      _EVAL_52[_EVAL_52__EVAL_54_addr] <= _EVAL_52__EVAL_54_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if (_EVAL_0) begin
      _EVAL_21 <= 1'h0;
    end else begin
      if (_EVAL_41) begin
        _EVAL_21 <= _EVAL_34;
      end
    end
    if (_EVAL_0) begin
      _EVAL_22 <= 1'h0;
    end else begin
      if (_EVAL_61) begin
        _EVAL_22 <= _EVAL_55;
      end
    end
    if (_EVAL_0) begin
      _EVAL_33 <= 1'h0;
    end else begin
      if (_EVAL_48) begin
        _EVAL_33 <= _EVAL_61;
      end
    end
  end
endmodule
