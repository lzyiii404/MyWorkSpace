//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_114(
  output [31:0] _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  output [3:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  output [29:0] _EVAL_4,
  input  [31:0] _EVAL_5,
  input  [3:0]  _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output [31:0] _EVAL_9,
  input         _EVAL_10,
  input  [6:0]  _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [29:0] _EVAL_16,
  output [2:0]  _EVAL_17,
  output [6:0]  _EVAL_18,
  input  [3:0]  _EVAL_19,
  input  [3:0]  _EVAL_20,
  output [6:0]  _EVAL_21,
  input         _EVAL_22,
  input  [6:0]  _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  output [2:0]  _EVAL_27,
  output [3:0]  _EVAL_28,
  input         _EVAL_29,
  input  [2:0]  _EVAL_30,
  output [1:0]  _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  output [3:0]  _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [2:0]  _EVAL_38,
  input  [2:0]  _EVAL_39,
  input         _EVAL_40
);
  assign _EVAL_27 = _EVAL_30;
  assign _EVAL_31 = _EVAL_1;
  assign _EVAL_8 = _EVAL_40;
  assign _EVAL_4 = _EVAL_16;
  assign _EVAL_21 = _EVAL_23;
  assign _EVAL_38 = _EVAL_15;
  assign _EVAL_24 = _EVAL_0;
  assign _EVAL_9 = _EVAL_5;
  assign _EVAL_13 = _EVAL_29;
  assign _EVAL_18 = _EVAL_11;
  assign _EVAL_28 = _EVAL_19;
  assign _EVAL_33 = _EVAL_36;
  assign _EVAL_17 = _EVAL_39;
  assign _EVAL_35 = _EVAL_6;
  assign _EVAL_32 = _EVAL_37;
  assign _EVAL = _EVAL_3;
  assign _EVAL_25 = _EVAL_10;
  assign _EVAL_26 = _EVAL_12;
  assign _EVAL_2 = _EVAL_20;
  assign _EVAL_7 = _EVAL_34;
endmodule
