//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_262(
  output [31:0] _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  output [2:0]  _EVAL_2,
  output [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input  [63:0] _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  input  [7:0]  _EVAL_19,
  output [2:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output        _EVAL_22,
  input  [24:0] _EVAL_23,
  output [63:0] _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  output [3:0]  _EVAL_27,
  output [2:0]  _EVAL_28,
  output [24:0] _EVAL_29,
  output [2:0]  _EVAL_30,
  output        _EVAL_31,
  output [2:0]  _EVAL_32
);
  wire [2:0] Repeater__EVAL;
  wire [2:0] Repeater__EVAL_0;
  wire [24:0] Repeater__EVAL_1;
  wire  Repeater__EVAL_2;
  wire [24:0] Repeater__EVAL_3;
  wire [63:0] Repeater__EVAL_4;
  wire [2:0] Repeater__EVAL_5;
  wire [7:0] Repeater__EVAL_6;
  wire  Repeater__EVAL_7;
  wire [63:0] Repeater__EVAL_8;
  wire  Repeater__EVAL_9;
  wire [2:0] Repeater__EVAL_10;
  wire [2:0] Repeater__EVAL_11;
  wire  Repeater__EVAL_12;
  wire  Repeater__EVAL_13;
  wire [2:0] Repeater__EVAL_14;
  wire  Repeater__EVAL_15;
  wire [2:0] Repeater__EVAL_16;
  wire  Repeater__EVAL_17;
  wire [2:0] Repeater__EVAL_18;
  wire  Repeater__EVAL_19;
  wire  Repeater__EVAL_20;
  wire [7:0] Repeater__EVAL_21;
  reg  _EVAL_59;
  reg [31:0] _RAND_0;
  reg  _EVAL_75;
  reg [31:0] _RAND_1;
  reg [31:0] _EVAL_78;
  reg [31:0] _RAND_2;
  wire [9:0] _EVAL_53;
  wire [2:0] _EVAL_63;
  wire [2:0] _EVAL_73;
  wire  _EVAL_76;
  wire  _EVAL_60;
  wire  _EVAL_35;
  wire  _EVAL_58;
  wire  _EVAL_37;
  wire [2:0] _EVAL_42;
  wire [7:0] _EVAL_79;
  wire [2:0] _EVAL_67;
  wire [9:0] _EVAL_81;
  wire [2:0] _EVAL_51;
  wire [2:0] _EVAL_64;
  wire  _EVAL_70;
  wire  _EVAL_50;
  wire [31:0] _EVAL_66;
  wire [31:0] _EVAL_47;
  wire [63:0] _EVAL_43;
  wire  _EVAL_82;
  wire  _EVAL_69;
  wire  _EVAL_80;
  wire  _EVAL_40;
  wire  _EVAL_74;
  wire  _EVAL_34;
  wire [24:0] _EVAL_39;
  wire  _EVAL_48;
  wire  _EVAL_33;
  wire  _EVAL_52;
  wire  _EVAL_41;
  wire [31:0] _EVAL_57;
  wire [31:0] _EVAL_61;
  wire [3:0] _EVAL_36;
  wire  _EVAL_56;
  wire  _EVAL_55;
  wire  _EVAL_68;
  wire  _EVAL_38;
  wire  _EVAL_72;
  wire [31:0] _EVAL_77;
  wire  _EVAL_46;
  wire [3:0] _EVAL_49;
  SiFive__EVAL_261 Repeater (
    ._EVAL(Repeater__EVAL),
    ._EVAL_0(Repeater__EVAL_0),
    ._EVAL_1(Repeater__EVAL_1),
    ._EVAL_2(Repeater__EVAL_2),
    ._EVAL_3(Repeater__EVAL_3),
    ._EVAL_4(Repeater__EVAL_4),
    ._EVAL_5(Repeater__EVAL_5),
    ._EVAL_6(Repeater__EVAL_6),
    ._EVAL_7(Repeater__EVAL_7),
    ._EVAL_8(Repeater__EVAL_8),
    ._EVAL_9(Repeater__EVAL_9),
    ._EVAL_10(Repeater__EVAL_10),
    ._EVAL_11(Repeater__EVAL_11),
    ._EVAL_12(Repeater__EVAL_12),
    ._EVAL_13(Repeater__EVAL_13),
    ._EVAL_14(Repeater__EVAL_14),
    ._EVAL_15(Repeater__EVAL_15),
    ._EVAL_16(Repeater__EVAL_16),
    ._EVAL_17(Repeater__EVAL_17),
    ._EVAL_18(Repeater__EVAL_18),
    ._EVAL_19(Repeater__EVAL_19),
    ._EVAL_20(Repeater__EVAL_20),
    ._EVAL_21(Repeater__EVAL_21)
  );
  assign _EVAL_53 = 10'h7 << _EVAL_21;
  assign _EVAL_63 = _EVAL_53[2:0];
  assign _EVAL_73 = ~ _EVAL_63;
  assign _EVAL_76 = _EVAL_73[2:2];
  assign _EVAL_60 = _EVAL_75 == _EVAL_76;
  assign _EVAL_35 = _EVAL_13[0];
  assign _EVAL_58 = _EVAL_35 == 1'h0;
  assign _EVAL_37 = _EVAL_60 | _EVAL_58;
  assign _EVAL_42 = Repeater__EVAL_18;
  assign _EVAL_79 = Repeater__EVAL_6;
  assign _EVAL_67 = Repeater__EVAL_10;
  assign _EVAL_81 = 10'h7 << _EVAL_67;
  assign _EVAL_51 = _EVAL_81[2:0];
  assign _EVAL_64 = ~ _EVAL_51;
  assign _EVAL_70 = _EVAL_64[2:2];
  assign _EVAL_50 = _EVAL_59 == _EVAL_70;
  assign _EVAL_66 = Repeater__EVAL_4[63:32];
  assign _EVAL_47 = _EVAL_16[31:0];
  assign _EVAL_43 = {_EVAL_66,_EVAL_47};
  assign _EVAL_82 = _EVAL_37 == 1'h0;
  assign _EVAL_69 = _EVAL_8 | _EVAL_82;
  assign _EVAL_80 = _EVAL_69 & _EVAL_4;
  assign _EVAL_40 = _EVAL_75 + 1'h1;
  assign _EVAL_74 = _EVAL_42[2];
  assign _EVAL_34 = _EVAL_74 == 1'h0;
  assign _EVAL_39 = Repeater__EVAL_1;
  assign _EVAL_48 = _EVAL_39[2];
  assign _EVAL_33 = _EVAL_48 | _EVAL_59;
  assign _EVAL_52 = _EVAL_75 & _EVAL_76;
  assign _EVAL_41 = _EVAL_52 == 1'h0;
  assign _EVAL_57 = _EVAL_41 ? _EVAL_1 : _EVAL_78;
  assign _EVAL_61 = _EVAL_43[31:0];
  assign _EVAL_36 = _EVAL_79[3:0];
  assign _EVAL_56 = _EVAL_34 == 1'h0;
  assign _EVAL_55 = Repeater__EVAL_15;
  assign _EVAL_68 = _EVAL_6 & _EVAL_55;
  assign _EVAL_38 = _EVAL_50 | _EVAL_56;
  assign _EVAL_72 = _EVAL_59 + 1'h1;
  assign _EVAL_77 = _EVAL_43[63:32];
  assign _EVAL_46 = _EVAL_80 & _EVAL_82;
  assign _EVAL_49 = _EVAL_79[7:4];
  assign Repeater__EVAL_13 = _EVAL_6;
  assign Repeater__EVAL_0 = _EVAL_7;
  assign _EVAL_22 = Repeater__EVAL_7;
  assign _EVAL_27 = _EVAL_33 ? _EVAL_49 : _EVAL_36;
  assign Repeater__EVAL_8 = _EVAL_16;
  assign Repeater__EVAL_17 = _EVAL_38 == 1'h0;
  assign Repeater__EVAL_9 = _EVAL_17;
  assign _EVAL_20 = Repeater__EVAL_10;
  assign _EVAL_30 = Repeater__EVAL_18;
  assign Repeater__EVAL = _EVAL_5;
  assign _EVAL_29 = Repeater__EVAL_1;
  assign _EVAL_3 = Repeater__EVAL_5;
  assign Repeater__EVAL_21 = _EVAL_19;
  assign _EVAL_32 = _EVAL_13;
  assign Repeater__EVAL_3 = _EVAL_23;
  assign _EVAL_28 = _EVAL_14;
  assign _EVAL_24 = {_EVAL_1,_EVAL_57};
  assign Repeater__EVAL_20 = _EVAL_26;
  assign _EVAL_18 = _EVAL_21;
  assign _EVAL_10 = _EVAL_4 & _EVAL_37;
  assign Repeater__EVAL_19 = _EVAL_12;
  assign Repeater__EVAL_2 = _EVAL_15;
  assign _EVAL_31 = _EVAL_8 | _EVAL_82;
  assign Repeater__EVAL_16 = _EVAL_9;
  assign _EVAL_0 = Repeater__EVAL_12;
  assign _EVAL_11 = Repeater__EVAL_15;
  assign Repeater__EVAL_11 = _EVAL_25;
  assign _EVAL = _EVAL_33 ? _EVAL_77 : _EVAL_61;
  assign _EVAL_2 = Repeater__EVAL_14;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_59 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_75 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_78 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_26) begin
    if (_EVAL_17) begin
      _EVAL_59 <= 1'h0;
    end else begin
      if (_EVAL_68) begin
        if (_EVAL_38) begin
          _EVAL_59 <= 1'h0;
        end else begin
          _EVAL_59 <= _EVAL_72;
        end
      end
    end
    if (_EVAL_17) begin
      _EVAL_75 <= 1'h0;
    end else begin
      if (_EVAL_80) begin
        if (_EVAL_37) begin
          _EVAL_75 <= 1'h0;
        end else begin
          _EVAL_75 <= _EVAL_40;
        end
      end
    end
    if (_EVAL_46) begin
      if (_EVAL_41) begin
        _EVAL_78 <= _EVAL_1;
      end
    end
  end
endmodule
