//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
bind SiFive__EVAL_2 SiFive__EVAL_2_assert SiFive__EVAL_2_assert_0 (.*);
bind SiFive__EVAL_4 SiFive__EVAL_4_assert SiFive__EVAL_4_assert_0 (.*);
bind SiFive__EVAL_6 SiFive__EVAL_6_assert SiFive__EVAL_6_assert_0 (.*);
bind SiFive__EVAL_8 SiFive__EVAL_8_assert SiFive__EVAL_8_assert_0 (.*);
bind SiFive__EVAL_10 SiFive__EVAL_10_assert SiFive__EVAL_10_assert_0 (.*);
bind SiFive__EVAL_12 SiFive__EVAL_12_assert SiFive__EVAL_12_assert_0 (.*);
bind SiFive__EVAL_14 SiFive__EVAL_14_assert SiFive__EVAL_14_assert_0 (.*);
bind SiFive__EVAL_16 SiFive__EVAL_16_assert SiFive__EVAL_16_assert_0 (.*);
bind SiFive__EVAL_20 SiFive__EVAL_20_assert SiFive__EVAL_20_assert_0 (.*);
bind SiFive__EVAL_28 SiFive__EVAL_28_assert SiFive__EVAL_28_assert_0 (.*);
bind SiFive__EVAL_33 SiFive__EVAL_33_assert SiFive__EVAL_33_assert_0 (.*);
bind SiFive__EVAL_36 SiFive__EVAL_36_assert SiFive__EVAL_36_assert_0 (.*);
bind SiFive__EVAL_38 SiFive__EVAL_38_assert SiFive__EVAL_38_assert_0 (.*);
bind SiFive__EVAL_43 SiFive__EVAL_43_assert SiFive__EVAL_43_assert_0 (.*);
bind SiFive__EVAL_47 SiFive__EVAL_47_assert SiFive__EVAL_47_assert_0 (.*);
bind SiFive__EVAL_52 SiFive__EVAL_52_assert SiFive__EVAL_52_assert_0 (.*);
bind SiFive__EVAL_54 SiFive__EVAL_54_assert SiFive__EVAL_54_assert_0 (.*);
bind SiFive__EVAL_56 SiFive__EVAL_56_assert SiFive__EVAL_56_assert_0 (.*);
bind SiFive__EVAL_59 SiFive__EVAL_59_assert SiFive__EVAL_59_assert_0 (.*);
bind SiFive__EVAL_62 SiFive__EVAL_62_assert SiFive__EVAL_62_assert_0 (.*);
bind SiFive__EVAL_64 SiFive__EVAL_64_assert SiFive__EVAL_64_assert_0 (.*);
bind SiFive__EVAL_66 SiFive__EVAL_66_assert SiFive__EVAL_66_assert_0 (.*);
bind SiFive__EVAL_69 SiFive__EVAL_69_assert SiFive__EVAL_69_assert_0 (.*);
bind SiFive__EVAL_71 SiFive__EVAL_71_assert SiFive__EVAL_71_assert_0 (.*);
bind SiFive__EVAL_73 SiFive__EVAL_73_assert SiFive__EVAL_73_assert_0 (.*);
bind SiFive__EVAL_84 SiFive__EVAL_84_assert SiFive__EVAL_84_assert_0 (.*);
bind SiFive__EVAL_87 SiFive__EVAL_87_assert SiFive__EVAL_87_assert_0 (.*);
bind SiFive__EVAL_92 SiFive__EVAL_92_assert SiFive__EVAL_92_assert_0 (.*);
bind SiFive__EVAL_94 SiFive__EVAL_94_assert SiFive__EVAL_94_assert_0 (.*);
bind SiFive__EVAL_99 SiFive__EVAL_99_assert SiFive__EVAL_99_assert_0 (.*);
bind SiFive__EVAL_101 SiFive__EVAL_101_assert SiFive__EVAL_101_assert_0 (.*);
bind SiFive__EVAL_103 SiFive__EVAL_103_assert SiFive__EVAL_103_assert_0 (.*);
bind SiFive__EVAL_105 SiFive__EVAL_105_assert SiFive__EVAL_105_assert_0 (.*);
bind SiFive__EVAL_108 SiFive__EVAL_108_assert SiFive__EVAL_108_assert_0 (.*);
bind SiFive__EVAL_112 SiFive__EVAL_112_assert SiFive__EVAL_112_assert_0 (.*);
bind SiFive__EVAL_114 SiFive__EVAL_114_assert SiFive__EVAL_114_assert_0 (.*);
bind SiFive__EVAL_116 SiFive__EVAL_116_assert SiFive__EVAL_116_assert_0 (.*);
bind SiFive__EVAL_120 SiFive__EVAL_120_assert SiFive__EVAL_120_assert_0 (.*);
bind SiFive__EVAL_122 SiFive__EVAL_122_assert SiFive__EVAL_122_assert_0 (.*);
bind SiFive__EVAL_125 SiFive__EVAL_125_assert SiFive__EVAL_125_assert_0 (.*);
bind SiFive__EVAL_128 SiFive__EVAL_128_assert SiFive__EVAL_128_assert_0 (.*);
bind SiFive__EVAL_132 SiFive__EVAL_132_assert SiFive__EVAL_132_assert_0 (.*);
bind SiFive__EVAL_136 SiFive__EVAL_136_assert SiFive__EVAL_136_assert_0 (.*);
bind SiFive__EVAL_140 SiFive__EVAL_140_assert SiFive__EVAL_140_assert_0 (.*);
bind SiFive__EVAL_144 SiFive__EVAL_144_assert SiFive__EVAL_144_assert_0 (.*);
bind SiFive__EVAL_146 SiFive__EVAL_146_assert SiFive__EVAL_146_assert_0 (.*);
bind SiFive__EVAL_147 SiFive__EVAL_147_assert SiFive__EVAL_147_assert_0 (.*);
bind SiFive__EVAL_149 SiFive__EVAL_149_assert SiFive__EVAL_149_assert_0 (.*);
bind SiFive__EVAL_151 SiFive__EVAL_151_assert SiFive__EVAL_151_assert_0 (.*);
bind SiFive__EVAL_155 SiFive__EVAL_155_assert SiFive__EVAL_155_assert_0 (.*);
bind SiFive__EVAL_157 SiFive__EVAL_157_assert SiFive__EVAL_157_assert_0 (.*);
bind SiFive__EVAL_161 SiFive__EVAL_161_assert SiFive__EVAL_161_assert_0 (.*);
bind SiFive__EVAL_167 SiFive__EVAL_167_assert SiFive__EVAL_167_assert_0 (.*);
bind SiFive__EVAL_171 SiFive__EVAL_171_assert SiFive__EVAL_171_assert_0 (.*);
bind SiFive__EVAL_173 SiFive__EVAL_173_assert SiFive__EVAL_173_assert_0 (.*);
bind SiFive__EVAL_175 SiFive__EVAL_175_assert SiFive__EVAL_175_assert_0 (.*);
bind SiFive__EVAL_179 SiFive__EVAL_179_assert SiFive__EVAL_179_assert_0 (.*);
bind SiFive__EVAL_185 SiFive__EVAL_185_assert SiFive__EVAL_185_assert_0 (.*);
bind SiFive__EVAL_187 SiFive__EVAL_187_assert SiFive__EVAL_187_assert_0 (.*);
bind SiFive__EVAL_189 SiFive__EVAL_189_assert SiFive__EVAL_189_assert_0 (.*);
bind SiFive__EVAL_194 SiFive__EVAL_194_assert SiFive__EVAL_194_assert_0 (.*);
bind SiFive__EVAL_206 SiFive__EVAL_206_assert SiFive__EVAL_206_assert_0 (.*);
bind SiFive__EVAL_210 SiFive__EVAL_210_assert SiFive__EVAL_210_assert_0 (.*);
bind SiFive__EVAL_213 SiFive__EVAL_213_assert SiFive__EVAL_213_assert_0 (.*);
bind SiFive__EVAL_217 SiFive__EVAL_217_assert SiFive__EVAL_217_assert_0 (.*);
bind SiFive__EVAL_225 SiFive__EVAL_225_assert SiFive__EVAL_225_assert_0 (.*);
bind SiFive__EVAL_226 SiFive__EVAL_226_assert SiFive__EVAL_226_assert_0 (.*);
bind SiFive__EVAL_228 SiFive__EVAL_228_assert SiFive__EVAL_228_assert_0 (.*);
bind SiFive__EVAL_234 SiFive__EVAL_234_assert SiFive__EVAL_234_assert_0 (.*);
bind SiFive__EVAL_236 SiFive__EVAL_236_assert SiFive__EVAL_236_assert_0 (.*);
bind SiFive__EVAL_240 SiFive__EVAL_240_assert SiFive__EVAL_240_assert_0 (.*);
bind SiFive__EVAL_243 SiFive__EVAL_243_assert SiFive__EVAL_243_assert_0 (.*);
bind SiFive__EVAL_246 SiFive__EVAL_246_assert SiFive__EVAL_246_assert_0 (.*);
bind SiFive__EVAL_249 SiFive__EVAL_249_assert SiFive__EVAL_249_assert_0 (.*);
bind SiFive__EVAL_251 SiFive__EVAL_251_assert SiFive__EVAL_251_assert_0 (.*);
bind SiFive__EVAL_253 SiFive__EVAL_253_assert SiFive__EVAL_253_assert_0 (.*);
bind SiFive__EVAL_256 SiFive__EVAL_256_assert SiFive__EVAL_256_assert_0 (.*);
bind SiFive__EVAL_259 SiFive__EVAL_259_assert SiFive__EVAL_259_assert_0 (.*);
bind SiFive__EVAL_262 SiFive__EVAL_262_assert SiFive__EVAL_262_assert_0 (.*);
bind SiFive__EVAL_264 SiFive__EVAL_264_assert SiFive__EVAL_264_assert_0 (.*);
bind SiFive__EVAL_266 SiFive__EVAL_266_assert SiFive__EVAL_266_assert_0 (.*);
bind SiFive__EVAL_268 SiFive__EVAL_268_assert SiFive__EVAL_268_assert_0 (.*);
bind SiFive__EVAL_269 SiFive__EVAL_269_assert SiFive__EVAL_269_assert_0 (.*);
bind SiFive__EVAL_270 SiFive__EVAL_270_assert SiFive__EVAL_270_assert_0 (.*);
bind SiFive__EVAL_271 SiFive__EVAL_271_assert SiFive__EVAL_271_assert_0 (.*);
bind SiFive__EVAL_272 SiFive__EVAL_272_assert SiFive__EVAL_272_assert_0 (.*);
bind SiFive__EVAL_273 SiFive__EVAL_273_assert SiFive__EVAL_273_assert_0 (.*);
bind SiFive__EVAL_275 SiFive__EVAL_275_assert SiFive__EVAL_275_assert_0 (.*);
bind SiFive__EVAL_276 SiFive__EVAL_276_assert SiFive__EVAL_276_assert_0 (.*);
bind SiFive__EVAL_303 SiFive__EVAL_303_assert SiFive__EVAL_303_assert_0 (.*);
bind SiFive__EVAL_304 SiFive__EVAL_304_assert SiFive__EVAL_304_assert_0 (.*);
bind SiFive__EVAL_307 SiFive__EVAL_307_assert SiFive__EVAL_307_assert_0 (.*);
bind SiFive_TLTestIndicator SiFive_TLTestIndicator_assert SiFive_TLTestIndicator_assert_0 (.*);
bind SiFive__EVAL_318 SiFive__EVAL_318_assert SiFive__EVAL_318_assert_0 (.*);
bind SiFive__EVAL_319 SiFive__EVAL_319_assert SiFive__EVAL_319_assert_0 (.*);
bind SiFive__EVAL_320 SiFive__EVAL_320_assert SiFive__EVAL_320_assert_0 (.*);
bind SiFive__EVAL_322 SiFive__EVAL_322_assert SiFive__EVAL_322_assert_0 (.*);
bind SiFive__EVAL_324 SiFive__EVAL_324_assert SiFive__EVAL_324_assert_0 (.*);
bind SiFive__EVAL_326 SiFive__EVAL_326_assert SiFive__EVAL_326_assert_0 (.*);
bind SiFive__EVAL_327 SiFive__EVAL_327_assert SiFive__EVAL_327_assert_0 (.*);
bind SiFive__EVAL_328 SiFive__EVAL_328_assert SiFive__EVAL_328_assert_0 (.*);
bind SiFive__EVAL_329 SiFive__EVAL_329_assert SiFive__EVAL_329_assert_0 (.*);
bind SiFive__EVAL_331 SiFive__EVAL_331_assert SiFive__EVAL_331_assert_0 (.*);
bind SiFive__EVAL_332 SiFive__EVAL_332_assert SiFive__EVAL_332_assert_0 (.*);
bind SiFive__EVAL_334 SiFive__EVAL_334_assert SiFive__EVAL_334_assert_0 (.*);
bind SiFive__EVAL_335 SiFive__EVAL_335_assert SiFive__EVAL_335_assert_0 (.*);