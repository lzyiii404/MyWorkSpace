//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_320_assert(
  input         _EVAL_0,
  input         _EVAL_3,
  input  [31:0] _EVAL_8,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_17,
  input         _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [6:0]  _EVAL_21,
  input         _EVAL_22,
  input  [2:0]  _EVAL_23,
  input         _EVAL_24,
  input  [2:0]  _EVAL_30,
  input         _EVAL_33,
  input  [2:0]  _EVAL_37,
  input         _EVAL_39,
  input  [6:0]  _EVAL_46,
  input         _EVAL_47,
  input  [7:0]  _EVAL_49,
  input  [31:0] _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input  [25:0] _EVAL_69,
  input         _EVAL_101,
  input  [1:0]  _EVAL_384,
  input         _EVAL_194,
  input  [2:0]  _EVAL_231,
  input         _EVAL_78,
  input         _EVAL_65,
  input         _EVAL_59,
  input  [1:0]  _EVAL_250,
  input         _EVAL_75,
  input         _EVAL_89,
  input         _EVAL_378,
  input         _EVAL_118,
  input         _EVAL_294,
  input         _EVAL_402,
  input         _EVAL_373,
  input         _EVAL_326,
  input         _EVAL_91,
  input         _EVAL_92,
  input         _EVAL_376,
  input  [81:0] _EVAL_225
);
  wire [31:0] TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire [2:0] TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire [1:0] TLMonitor__EVAL_3;
  wire [31:0] TLMonitor__EVAL_4;
  wire [2:0] TLMonitor__EVAL_5;
  wire [2:0] TLMonitor__EVAL_6;
  wire [6:0] TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire  TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire  TLMonitor__EVAL_15;
  wire [2:0] TLMonitor__EVAL_16;
  wire  TLMonitor__EVAL_17;
  wire [2:0] TLMonitor__EVAL_18;
  wire  TLMonitor__EVAL_19;
  wire  TLMonitor__EVAL_20;
  wire  TLMonitor__EVAL_21;
  wire [2:0] TLMonitor__EVAL_22;
  wire [7:0] TLMonitor__EVAL_23;
  wire  TLMonitor__EVAL_24;
  wire [6:0] TLMonitor__EVAL_25;
  wire  TLMonitor__EVAL_26;
  wire [31:0] TLMonitor__EVAL_27;
  wire [1:0] TLMonitor__EVAL_28;
  wire  TLMonitor__EVAL_29;
  wire  TLMonitor__EVAL_30;
  wire [2:0] TLMonitor__EVAL_31;
  wire [6:0] TLMonitor__EVAL_32;
  wire  _EVAL_138;
  wire  _EVAL_221;
  wire  _EVAL_406;
  wire  _EVAL_217;
  wire  _EVAL_168;
  wire  _EVAL_109;
  wire  _EVAL_283;
  wire  _EVAL_327;
  wire  _EVAL_214;
  wire  _EVAL_241;
  wire  _EVAL_295;
  wire  _EVAL_165;
  wire  _EVAL_249;
  wire  _EVAL_390;
  wire  _EVAL_333;
  wire  _EVAL_134;
  wire  _EVAL_414;
  wire  _EVAL_71;
  wire  _EVAL_210;
  wire  _EVAL_86;
  wire  _EVAL_396;
  wire  _EVAL_317;
  wire  _EVAL_132;
  wire  _EVAL_296;
  wire  _EVAL_265;
  wire  _EVAL_170;
  wire  _EVAL_287;
  wire  _EVAL_392;
  wire  _EVAL_364;
  wire  _EVAL_252;
  wire  _EVAL_298;
  wire  _EVAL_381;
  wire  _EVAL_398;
  wire  _EVAL_185;
  wire  _EVAL_290;
  wire  _EVAL_226;
  wire  _EVAL_303;
  wire  _EVAL_338;
  SiFive__EVAL_316_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18),
    ._EVAL_19(TLMonitor__EVAL_19),
    ._EVAL_20(TLMonitor__EVAL_20),
    ._EVAL_21(TLMonitor__EVAL_21),
    ._EVAL_22(TLMonitor__EVAL_22),
    ._EVAL_23(TLMonitor__EVAL_23),
    ._EVAL_24(TLMonitor__EVAL_24),
    ._EVAL_25(TLMonitor__EVAL_25),
    ._EVAL_26(TLMonitor__EVAL_26),
    ._EVAL_27(TLMonitor__EVAL_27),
    ._EVAL_28(TLMonitor__EVAL_28),
    ._EVAL_29(TLMonitor__EVAL_29),
    ._EVAL_30(TLMonitor__EVAL_30),
    ._EVAL_31(TLMonitor__EVAL_31),
    ._EVAL_32(TLMonitor__EVAL_32)
  );
  assign _EVAL_138 = _EVAL_65 == 1'h0;
  assign _EVAL_221 = _EVAL_59 == 1'h0;
  assign _EVAL_406 = _EVAL_138 | _EVAL_221;
  assign _EVAL_217 = _EVAL_194 == 1'h0;
  assign _EVAL_168 = _EVAL_65 | _EVAL_59;
  assign _EVAL_109 = _EVAL_168 | _EVAL_194;
  assign _EVAL_283 = _EVAL_11 == 3'h0;
  assign _EVAL_327 = _EVAL_373 == 1'h0;
  assign _EVAL_214 = _EVAL_118 == 1'h0;
  assign _EVAL_241 = _EVAL_327 | _EVAL_214;
  assign _EVAL_295 = _EVAL_241 | _EVAL_19;
  assign _EVAL_165 = _EVAL_373 | _EVAL_118;
  assign _EVAL_249 = _EVAL_92 == 1'h0;
  assign _EVAL_390 = _EVAL_249 | _EVAL_165;
  assign _EVAL_333 = _EVAL_390 | _EVAL_19;
  assign _EVAL_134 = _EVAL_168 == 1'h0;
  assign _EVAL_414 = _EVAL_134 | _EVAL_217;
  assign _EVAL_71 = _EVAL_22 == 1'h0;
  assign _EVAL_210 = _EVAL_71 | _EVAL_89;
  assign _EVAL_86 = _EVAL_378 == 1'h0;
  assign _EVAL_396 = _EVAL_250 != 2'h0;
  assign _EVAL_317 = _EVAL_231 == 3'h6;
  assign _EVAL_132 = _EVAL_396 | _EVAL_317;
  assign _EVAL_296 = _EVAL_86 | _EVAL_132;
  assign _EVAL_265 = _EVAL_296 | _EVAL_19;
  assign _EVAL_170 = _EVAL_78 == 1'h0;
  assign _EVAL_287 = _EVAL_170 | _EVAL_109;
  assign _EVAL_392 = _EVAL_406 & _EVAL_414;
  assign _EVAL_364 = _EVAL_333 == 1'h0;
  assign _EVAL_252 = _EVAL_265 == 1'h0;
  assign _EVAL_298 = _EVAL_392 | _EVAL_19;
  assign _EVAL_381 = _EVAL_298 == 1'h0;
  assign _EVAL_398 = _EVAL_287 | _EVAL_19;
  assign _EVAL_185 = _EVAL_210 | _EVAL_283;
  assign _EVAL_290 = _EVAL_185 | _EVAL_19;
  assign _EVAL_226 = _EVAL_295 == 1'h0;
  assign _EVAL_303 = _EVAL_398 == 1'h0;
  assign _EVAL_338 = _EVAL_290 == 1'h0;
  assign TLMonitor__EVAL_6 = _EVAL_225[76:74];
  assign TLMonitor__EVAL_5 = _EVAL_37;
  assign TLMonitor__EVAL = {_EVAL_69, 6'h0};
  assign TLMonitor__EVAL_16 = _EVAL_30;
  assign TLMonitor__EVAL_31 = _EVAL_12;
  assign TLMonitor__EVAL_15 = _EVAL_52;
  assign TLMonitor__EVAL_29 = _EVAL_47;
  assign TLMonitor__EVAL_17 = _EVAL_53;
  assign TLMonitor__EVAL_2 = _EVAL_225[0];
  assign TLMonitor__EVAL_4 = _EVAL_8;
  assign TLMonitor__EVAL_21 = _EVAL_3;
  assign TLMonitor__EVAL_25 = _EVAL_225[73:67];
  assign TLMonitor__EVAL_26 = _EVAL_33;
  assign TLMonitor__EVAL_0 = _EVAL_101;
  assign TLMonitor__EVAL_18 = _EVAL_20;
  assign TLMonitor__EVAL_30 = _EVAL_19;
  assign TLMonitor__EVAL_28 = _EVAL_225[78:77];
  assign TLMonitor__EVAL_24 = _EVAL_294 & _EVAL_402;
  assign TLMonitor__EVAL_22 = _EVAL_17;
  assign TLMonitor__EVAL_9 = _EVAL_39;
  assign TLMonitor__EVAL_1 = _EVAL_225[81:79];
  assign TLMonitor__EVAL_19 = _EVAL_326 | _EVAL_91;
  assign TLMonitor__EVAL_10 = _EVAL_0;
  assign TLMonitor__EVAL_8 = _EVAL_24;
  assign TLMonitor__EVAL_14 = _EVAL_10;
  assign TLMonitor__EVAL_20 = _EVAL_225[66];
  assign TLMonitor__EVAL_7 = _EVAL_46;
  assign TLMonitor__EVAL_13 = _EVAL_225[65];
  assign TLMonitor__EVAL_32 = _EVAL_21;
  assign TLMonitor__EVAL_11 = _EVAL_23;
  assign TLMonitor__EVAL_27 = _EVAL_51;
  assign TLMonitor__EVAL_23 = _EVAL_49;
  assign TLMonitor__EVAL_12 = _EVAL_75 ? _EVAL_92 : _EVAL_376;
  assign TLMonitor__EVAL_3 = _EVAL_384;
  always @(posedge _EVAL_33) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_381) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(185a3b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21984a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_381) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
