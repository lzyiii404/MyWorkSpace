//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_4(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  output [3:0]  _EVAL_1,
  output [31:0] _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  input  [31:0] _EVAL_6,
  output        _EVAL_7,
  input  [63:0] _EVAL_8,
  output [31:0] _EVAL_9,
  input  [7:0]  _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output [63:0] _EVAL_13,
  output [1:0]  _EVAL_14,
  output        _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [2:0]  _EVAL_18,
  input  [1:0]  _EVAL_19,
  input  [3:0]  _EVAL_20,
  output        _EVAL_21,
  output [1:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  output [3:0]  _EVAL_32,
  input         _EVAL_33,
  input  [63:0] _EVAL_34,
  input  [31:0] _EVAL_35,
  output [3:0]  _EVAL_36,
  input         _EVAL_37,
  output [2:0]  _EVAL_38,
  input  [63:0] _EVAL_39,
  output [2:0]  _EVAL_40,
  output        _EVAL_41,
  output [3:0]  _EVAL_42,
  output [2:0]  _EVAL_43,
  input  [2:0]  _EVAL_44,
  output [2:0]  _EVAL_45,
  input  [31:0] _EVAL_46,
  input  [3:0]  _EVAL_47,
  output        _EVAL_48,
  output [31:0] _EVAL_49,
  input         _EVAL_50,
  input  [3:0]  _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input  [3:0]  _EVAL_54,
  input  [2:0]  _EVAL_55,
  output [63:0] _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  output        _EVAL_59,
  output [63:0] _EVAL_60,
  input         _EVAL_61,
  input         _EVAL_62,
  output [2:0]  _EVAL_63,
  output [3:0]  _EVAL_64,
  input  [3:0]  _EVAL_65,
  output        _EVAL_66,
  output [7:0]  _EVAL_67,
  input  [2:0]  _EVAL_68,
  input  [1:0]  _EVAL_69,
  input         _EVAL_70
);
  assign _EVAL_28 = _EVAL_24;
  assign _EVAL_16 = _EVAL_65;
  assign _EVAL_41 = _EVAL_23;
  assign _EVAL_21 = _EVAL_50;
  assign _EVAL_38 = _EVAL_44;
  assign _EVAL_64 = _EVAL_54;
  assign _EVAL_7 = _EVAL_5;
  assign _EVAL_36 = _EVAL_51;
  assign _EVAL_3 = _EVAL_58;
  assign _EVAL_14 = _EVAL_69;
  assign _EVAL_66 = _EVAL;
  assign _EVAL_32 = _EVAL_20;
  assign _EVAL_13 = _EVAL_39;
  assign _EVAL_40 = _EVAL_68;
  assign _EVAL_1 = _EVAL_0;
  assign _EVAL_42 = _EVAL_47;
  assign _EVAL_56 = _EVAL_8;
  assign _EVAL_49 = _EVAL_6;
  assign _EVAL_45 = _EVAL_55;
  assign _EVAL_30 = _EVAL_33;
  assign _EVAL_11 = _EVAL_70;
  assign _EVAL_22 = _EVAL_19;
  assign _EVAL_2 = _EVAL_46;
  assign _EVAL_15 = _EVAL_26;
  assign _EVAL_43 = _EVAL_17;
  assign _EVAL_4 = _EVAL_37;
  assign _EVAL_60 = _EVAL_34;
  assign _EVAL_67 = _EVAL_10;
  assign _EVAL_25 = _EVAL_27;
  assign _EVAL_29 = _EVAL_52;
  assign _EVAL_12 = _EVAL_31;
  assign _EVAL_48 = _EVAL_61;
  assign _EVAL_63 = _EVAL_18;
  assign _EVAL_59 = _EVAL_57;
  assign _EVAL_9 = _EVAL_35;
endmodule
