//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_305(
  output        _EVAL,
  input         _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input  [3:0]  _EVAL_4,
  input  [4:0]  _EVAL_5,
  input  [31:0] _EVAL_6,
  input         _EVAL_7,
  output [31:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  output [4:0]  _EVAL_11
);
  reg [32:0] _EVAL_21;
  reg [63:0] _RAND_0;
  reg [5:0] _EVAL_63;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_66;
  reg [31:0] _RAND_2;
  reg  _EVAL_144;
  reg [31:0] _RAND_3;
  reg  _EVAL_191;
  reg [31:0] _RAND_4;
  reg [65:0] _EVAL_196;
  reg [95:0] _RAND_5;
  reg [4:0] _EVAL_224;
  reg [31:0] _RAND_6;
  reg  _EVAL_229;
  reg [31:0] _RAND_7;
  wire [31:0] _EVAL_208;
  wire [15:0] _EVAL_236;
  wire [7:0] _EVAL_202;
  wire [3:0] _EVAL_109;
  wire  _EVAL_95;
  wire  _EVAL_58;
  wire  _EVAL_187;
  wire  _EVAL_152;
  wire [1:0] _EVAL_73;
  wire [1:0] _EVAL_178;
  wire [3:0] _EVAL_113;
  wire  _EVAL_249;
  wire  _EVAL_75;
  wire  _EVAL_61;
  wire [1:0] _EVAL_222;
  wire [1:0] _EVAL_184;
  wire [1:0] _EVAL_112;
  wire  _EVAL_120;
  wire  _EVAL_64;
  wire  _EVAL_102;
  wire  _EVAL_129;
  wire  _EVAL_39;
  wire  _EVAL_251;
  wire [15:0] _EVAL_218;
  wire [7:0] _EVAL_135;
  wire [3:0] _EVAL_53;
  wire  _EVAL_90;
  wire  _EVAL_246;
  wire [32:0] _EVAL_29;
  wire [32:0] _EVAL_124;
  wire  _EVAL_116;
  wire  _EVAL_242;
  wire  _EVAL_248;
  wire [7:0] _EVAL_240;
  wire [3:0] _EVAL_43;
  wire  _EVAL_49;
  wire  _EVAL_126;
  wire  _EVAL_131;
  wire [1:0] _EVAL_85;
  wire [1:0] _EVAL_230;
  wire  _EVAL_141;
  wire [31:0] _EVAL_183;
  wire  _EVAL_139;
  wire [31:0] _EVAL_15;
  wire [31:0] _EVAL_206;
  wire [31:0] _EVAL_179;
  wire [31:0] _EVAL_34;
  wire [15:0] _EVAL_149;
  wire [7:0] _EVAL_168;
  wire [3:0] _EVAL_19;
  wire  _EVAL_103;
  wire  _EVAL_195;
  wire [1:0] _EVAL_57;
  wire  _EVAL_197;
  wire [1:0] _EVAL_50;
  wire  _EVAL_27;
  wire  _EVAL_160;
  wire [3:0] _EVAL_154;
  wire  _EVAL_100;
  wire  _EVAL_33;
  wire  _EVAL_93;
  wire  _EVAL_198;
  wire [1:0] _EVAL_81;
  wire [1:0] _EVAL_150;
  wire  _EVAL_193;
  wire [1:0] _EVAL_13;
  wire [1:0] _EVAL_215;
  wire [1:0] _EVAL_201;
  wire [15:0] _EVAL_204;
  wire [7:0] _EVAL_238;
  wire [3:0] _EVAL_71;
  wire  _EVAL_134;
  wire [7:0] _EVAL_127;
  wire [3:0] _EVAL_114;
  wire  _EVAL_170;
  wire  _EVAL_241;
  wire  _EVAL_67;
  wire [1:0] _EVAL_16;
  wire [1:0] _EVAL_220;
  wire  _EVAL_32;
  wire [2:0] _EVAL_45;
  wire [7:0] _EVAL_188;
  wire [3:0] _EVAL_177;
  wire  _EVAL_55;
  wire  _EVAL_74;
  wire  _EVAL_153;
  wire  _EVAL_80;
  wire [1:0] _EVAL_223;
  wire [1:0] _EVAL_72;
  wire [3:0] _EVAL_65;
  wire  _EVAL_115;
  wire  _EVAL_245;
  wire  _EVAL_247;
  wire [1:0] _EVAL_12;
  wire [1:0] _EVAL_156;
  wire [1:0] _EVAL_221;
  wire [2:0] _EVAL_244;
  wire [2:0] _EVAL_186;
  wire [3:0] _EVAL_203;
  wire  _EVAL_47;
  wire [2:0] _EVAL_123;
  wire  _EVAL_138;
  wire [3:0] _EVAL_54;
  wire  _EVAL_24;
  wire  _EVAL_128;
  wire  _EVAL_14;
  wire [1:0] _EVAL_99;
  wire [1:0] _EVAL_190;
  wire [1:0] _EVAL_48;
  wire [2:0] _EVAL_158;
  wire [2:0] _EVAL_125;
  wire [3:0] _EVAL_59;
  wire [3:0] _EVAL_97;
  wire [4:0] _EVAL_36;
  wire  _EVAL_108;
  wire [7:0] _EVAL_137;
  wire  _EVAL_205;
  wire [3:0] _EVAL_173;
  wire  _EVAL_88;
  wire  _EVAL_161;
  wire  _EVAL_219;
  wire  _EVAL_239;
  wire [1:0] _EVAL_20;
  wire [1:0] _EVAL_194;
  wire [3:0] _EVAL_143;
  wire  _EVAL_98;
  wire  _EVAL_107;
  wire  _EVAL_44;
  wire [1:0] _EVAL_151;
  wire [1:0] _EVAL_76;
  wire [1:0] _EVAL_225;
  wire [2:0] _EVAL_92;
  wire [3:0] _EVAL_216;
  wire  _EVAL_213;
  wire  _EVAL_212;
  wire  _EVAL_142;
  wire  _EVAL_22;
  wire [1:0] _EVAL_145;
  wire [1:0] _EVAL_87;
  wire [1:0] _EVAL_185;
  wire [2:0] _EVAL_166;
  wire [2:0] _EVAL_42;
  wire [3:0] _EVAL_79;
  wire  _EVAL_140;
  wire  _EVAL_101;
  wire [3:0] _EVAL_30;
  wire  _EVAL_172;
  wire  _EVAL_104;
  wire  _EVAL_169;
  wire [1:0] _EVAL_17;
  wire [1:0] _EVAL_232;
  wire [1:0] _EVAL_62;
  wire [2:0] _EVAL_147;
  wire  _EVAL_86;
  wire  _EVAL_192;
  wire  _EVAL_40;
  wire [1:0] _EVAL_176;
  wire [1:0] _EVAL_110;
  wire [3:0] _EVAL_227;
  wire  _EVAL_189;
  wire  _EVAL_165;
  wire  _EVAL_182;
  wire [1:0] _EVAL_83;
  wire [1:0] _EVAL_18;
  wire [1:0] _EVAL_180;
  wire [2:0] _EVAL_35;
  wire [2:0] _EVAL_119;
  wire [3:0] _EVAL_157;
  wire [3:0] _EVAL_122;
  wire [4:0] _EVAL_70;
  wire [4:0] _EVAL_77;
  wire [4:0] _EVAL_228;
  wire  _EVAL_38;
  wire [3:0] _EVAL_60;
  wire  _EVAL_133;
  wire [3:0] _EVAL_209;
  wire  _EVAL_163;
  wire  _EVAL_181;
  wire  _EVAL_234;
  wire  _EVAL_167;
  wire  _EVAL_96;
  wire  _EVAL_231;
  wire  _EVAL_226;
  wire  _EVAL_69;
  wire [31:0] _EVAL_243;
  wire [31:0] _EVAL_23;
  wire [64:0] _EVAL_174;
  wire [15:0] _EVAL_233;
  wire [62:0] _EVAL_52;
  wire [15:0] _EVAL_250;
  wire [15:0] _EVAL_214;
  wire [32:0] _EVAL_121;
  wire  _EVAL_200;
  wire  _EVAL_118;
  wire [15:0] _EVAL_78;
  wire  _EVAL_159;
  wire [62:0] _EVAL_56;
  wire [64:0] _EVAL_91;
  wire  _EVAL_207;
  wire  _EVAL_155;
  wire  _EVAL_148;
  wire  _EVAL_162;
  wire [5:0] _EVAL_199;
  wire [15:0] _EVAL_217;
  wire [15:0] _EVAL_68;
  wire [31:0] _EVAL_175;
  assign _EVAL_208 = _EVAL_196[31:0];
  assign _EVAL_236 = _EVAL_208[31:16];
  assign _EVAL_202 = _EVAL_236[15:8];
  assign _EVAL_109 = _EVAL_202[7:4];
  assign _EVAL_95 = _EVAL_109 != 4'h0;
  assign _EVAL_58 = _EVAL_109[3];
  assign _EVAL_187 = _EVAL_109[2];
  assign _EVAL_152 = _EVAL_109[1];
  assign _EVAL_73 = _EVAL_187 ? 2'h2 : {{1'd0}, _EVAL_152};
  assign _EVAL_178 = _EVAL_58 ? 2'h3 : _EVAL_73;
  assign _EVAL_113 = _EVAL_202[3:0];
  assign _EVAL_249 = _EVAL_113[3];
  assign _EVAL_75 = _EVAL_113[2];
  assign _EVAL_61 = _EVAL_113[1];
  assign _EVAL_222 = _EVAL_75 ? 2'h2 : {{1'd0}, _EVAL_61};
  assign _EVAL_184 = _EVAL_249 ? 2'h3 : _EVAL_222;
  assign _EVAL_112 = _EVAL_95 ? _EVAL_178 : _EVAL_184;
  assign _EVAL_120 = _EVAL_0 & _EVAL_3;
  assign _EVAL_64 = _EVAL_120 | _EVAL_9;
  assign _EVAL_102 = _EVAL_66 == 3'h3;
  assign _EVAL_129 = _EVAL_63 == 6'h20;
  assign _EVAL_39 = _EVAL_66 == 3'h5;
  assign _EVAL_251 = _EVAL_66 == 3'h1;
  assign _EVAL_218 = _EVAL_208[15:0];
  assign _EVAL_135 = _EVAL_218[15:8];
  assign _EVAL_53 = _EVAL_135[3:0];
  assign _EVAL_90 = _EVAL_53[2];
  assign _EVAL_246 = _EVAL_63 == 6'h0;
  assign _EVAL_29 = _EVAL_196[64:32];
  assign _EVAL_124 = _EVAL_29 - _EVAL_21;
  assign _EVAL_116 = _EVAL_124[32];
  assign _EVAL_242 = _EVAL_116 == 1'h0;
  assign _EVAL_248 = _EVAL_246 & _EVAL_242;
  assign _EVAL_240 = _EVAL_218[7:0];
  assign _EVAL_43 = _EVAL_240[7:4];
  assign _EVAL_49 = _EVAL_43[3];
  assign _EVAL_126 = _EVAL_43[2];
  assign _EVAL_131 = _EVAL_43[1];
  assign _EVAL_85 = _EVAL_126 ? 2'h2 : {{1'd0}, _EVAL_131};
  assign _EVAL_230 = _EVAL_49 ? 2'h3 : _EVAL_85;
  assign _EVAL_141 = _EVAL_202 != 8'h0;
  assign _EVAL_183 = _EVAL_21[31:0];
  assign _EVAL_139 = _EVAL_196[31];
  assign _EVAL_15 = _EVAL_196[64:33];
  assign _EVAL_206 = _EVAL_229 ? _EVAL_15 : _EVAL_208;
  assign _EVAL_179 = 32'h0 - _EVAL_206;
  assign _EVAL_34 = _EVAL_124[31:0];
  assign _EVAL_149 = _EVAL_183[31:16];
  assign _EVAL_168 = _EVAL_149[7:0];
  assign _EVAL_19 = _EVAL_168[3:0];
  assign _EVAL_103 = _EVAL_19[2];
  assign _EVAL_195 = _EVAL_19[1];
  assign _EVAL_57 = _EVAL_103 ? 2'h2 : {{1'd0}, _EVAL_195};
  assign _EVAL_197 = _EVAL_19[3];
  assign _EVAL_50 = _EVAL_197 ? 2'h3 : _EVAL_57;
  assign _EVAL_27 = _EVAL_53[3];
  assign _EVAL_160 = _EVAL_21[31];
  assign _EVAL_154 = _EVAL_135[7:4];
  assign _EVAL_100 = _EVAL_154 != 4'h0;
  assign _EVAL_33 = _EVAL_154[3];
  assign _EVAL_93 = _EVAL_154[2];
  assign _EVAL_198 = _EVAL_154[1];
  assign _EVAL_81 = _EVAL_93 ? 2'h2 : {{1'd0}, _EVAL_198};
  assign _EVAL_150 = _EVAL_33 ? 2'h3 : _EVAL_81;
  assign _EVAL_193 = _EVAL_53[1];
  assign _EVAL_13 = _EVAL_90 ? 2'h2 : {{1'd0}, _EVAL_193};
  assign _EVAL_215 = _EVAL_27 ? 2'h3 : _EVAL_13;
  assign _EVAL_201 = _EVAL_100 ? _EVAL_150 : _EVAL_215;
  assign _EVAL_204 = _EVAL_183[15:0];
  assign _EVAL_238 = _EVAL_204[7:0];
  assign _EVAL_71 = _EVAL_238[7:4];
  assign _EVAL_134 = _EVAL_71[2];
  assign _EVAL_127 = _EVAL_204[15:8];
  assign _EVAL_114 = _EVAL_127[7:4];
  assign _EVAL_170 = _EVAL_114[3];
  assign _EVAL_241 = _EVAL_114[2];
  assign _EVAL_67 = _EVAL_114[1];
  assign _EVAL_16 = _EVAL_241 ? 2'h2 : {{1'd0}, _EVAL_67};
  assign _EVAL_220 = _EVAL_170 ? 2'h3 : _EVAL_16;
  assign _EVAL_32 = _EVAL_236 != 16'h0;
  assign _EVAL_45 = {_EVAL_95,_EVAL_112};
  assign _EVAL_188 = _EVAL_236[7:0];
  assign _EVAL_177 = _EVAL_188[7:4];
  assign _EVAL_55 = _EVAL_177 != 4'h0;
  assign _EVAL_74 = _EVAL_177[3];
  assign _EVAL_153 = _EVAL_177[2];
  assign _EVAL_80 = _EVAL_177[1];
  assign _EVAL_223 = _EVAL_153 ? 2'h2 : {{1'd0}, _EVAL_80};
  assign _EVAL_72 = _EVAL_74 ? 2'h3 : _EVAL_223;
  assign _EVAL_65 = _EVAL_188[3:0];
  assign _EVAL_115 = _EVAL_65[3];
  assign _EVAL_245 = _EVAL_65[2];
  assign _EVAL_247 = _EVAL_65[1];
  assign _EVAL_12 = _EVAL_245 ? 2'h2 : {{1'd0}, _EVAL_247};
  assign _EVAL_156 = _EVAL_115 ? 2'h3 : _EVAL_12;
  assign _EVAL_221 = _EVAL_55 ? _EVAL_72 : _EVAL_156;
  assign _EVAL_244 = {_EVAL_55,_EVAL_221};
  assign _EVAL_186 = _EVAL_141 ? _EVAL_45 : _EVAL_244;
  assign _EVAL_203 = {_EVAL_141,_EVAL_186};
  assign _EVAL_47 = _EVAL_135 != 8'h0;
  assign _EVAL_123 = {_EVAL_100,_EVAL_201};
  assign _EVAL_138 = _EVAL_43 != 4'h0;
  assign _EVAL_54 = _EVAL_240[3:0];
  assign _EVAL_24 = _EVAL_54[3];
  assign _EVAL_128 = _EVAL_54[2];
  assign _EVAL_14 = _EVAL_54[1];
  assign _EVAL_99 = _EVAL_128 ? 2'h2 : {{1'd0}, _EVAL_14};
  assign _EVAL_190 = _EVAL_24 ? 2'h3 : _EVAL_99;
  assign _EVAL_48 = _EVAL_138 ? _EVAL_230 : _EVAL_190;
  assign _EVAL_158 = {_EVAL_138,_EVAL_48};
  assign _EVAL_125 = _EVAL_47 ? _EVAL_123 : _EVAL_158;
  assign _EVAL_59 = {_EVAL_47,_EVAL_125};
  assign _EVAL_97 = _EVAL_32 ? _EVAL_203 : _EVAL_59;
  assign _EVAL_36 = {_EVAL_32,_EVAL_97};
  assign _EVAL_108 = _EVAL_149 != 16'h0;
  assign _EVAL_137 = _EVAL_149[15:8];
  assign _EVAL_205 = _EVAL_137 != 8'h0;
  assign _EVAL_173 = _EVAL_137[7:4];
  assign _EVAL_88 = _EVAL_173 != 4'h0;
  assign _EVAL_161 = _EVAL_173[3];
  assign _EVAL_219 = _EVAL_173[2];
  assign _EVAL_239 = _EVAL_173[1];
  assign _EVAL_20 = _EVAL_219 ? 2'h2 : {{1'd0}, _EVAL_239};
  assign _EVAL_194 = _EVAL_161 ? 2'h3 : _EVAL_20;
  assign _EVAL_143 = _EVAL_137[3:0];
  assign _EVAL_98 = _EVAL_143[3];
  assign _EVAL_107 = _EVAL_143[2];
  assign _EVAL_44 = _EVAL_143[1];
  assign _EVAL_151 = _EVAL_107 ? 2'h2 : {{1'd0}, _EVAL_44};
  assign _EVAL_76 = _EVAL_98 ? 2'h3 : _EVAL_151;
  assign _EVAL_225 = _EVAL_88 ? _EVAL_194 : _EVAL_76;
  assign _EVAL_92 = {_EVAL_88,_EVAL_225};
  assign _EVAL_216 = _EVAL_168[7:4];
  assign _EVAL_213 = _EVAL_216 != 4'h0;
  assign _EVAL_212 = _EVAL_216[3];
  assign _EVAL_142 = _EVAL_216[2];
  assign _EVAL_22 = _EVAL_216[1];
  assign _EVAL_145 = _EVAL_142 ? 2'h2 : {{1'd0}, _EVAL_22};
  assign _EVAL_87 = _EVAL_212 ? 2'h3 : _EVAL_145;
  assign _EVAL_185 = _EVAL_213 ? _EVAL_87 : _EVAL_50;
  assign _EVAL_166 = {_EVAL_213,_EVAL_185};
  assign _EVAL_42 = _EVAL_205 ? _EVAL_92 : _EVAL_166;
  assign _EVAL_79 = {_EVAL_205,_EVAL_42};
  assign _EVAL_140 = _EVAL_127 != 8'h0;
  assign _EVAL_101 = _EVAL_114 != 4'h0;
  assign _EVAL_30 = _EVAL_127[3:0];
  assign _EVAL_172 = _EVAL_30[3];
  assign _EVAL_104 = _EVAL_30[2];
  assign _EVAL_169 = _EVAL_30[1];
  assign _EVAL_17 = _EVAL_104 ? 2'h2 : {{1'd0}, _EVAL_169};
  assign _EVAL_232 = _EVAL_172 ? 2'h3 : _EVAL_17;
  assign _EVAL_62 = _EVAL_101 ? _EVAL_220 : _EVAL_232;
  assign _EVAL_147 = {_EVAL_101,_EVAL_62};
  assign _EVAL_86 = _EVAL_71 != 4'h0;
  assign _EVAL_192 = _EVAL_71[3];
  assign _EVAL_40 = _EVAL_71[1];
  assign _EVAL_176 = _EVAL_134 ? 2'h2 : {{1'd0}, _EVAL_40};
  assign _EVAL_110 = _EVAL_192 ? 2'h3 : _EVAL_176;
  assign _EVAL_227 = _EVAL_238[3:0];
  assign _EVAL_189 = _EVAL_227[3];
  assign _EVAL_165 = _EVAL_227[2];
  assign _EVAL_182 = _EVAL_227[1];
  assign _EVAL_83 = _EVAL_165 ? 2'h2 : {{1'd0}, _EVAL_182};
  assign _EVAL_18 = _EVAL_189 ? 2'h3 : _EVAL_83;
  assign _EVAL_180 = _EVAL_86 ? _EVAL_110 : _EVAL_18;
  assign _EVAL_35 = {_EVAL_86,_EVAL_180};
  assign _EVAL_119 = _EVAL_140 ? _EVAL_147 : _EVAL_35;
  assign _EVAL_157 = {_EVAL_140,_EVAL_119};
  assign _EVAL_122 = _EVAL_108 ? _EVAL_79 : _EVAL_157;
  assign _EVAL_70 = {_EVAL_108,_EVAL_122};
  assign _EVAL_77 = _EVAL_36 - _EVAL_70;
  assign _EVAL_228 = ~ _EVAL_77;
  assign _EVAL_38 = _EVAL_228 >= 5'h1;
  assign _EVAL_60 = _EVAL_4 & 4'h2;
  assign _EVAL_133 = _EVAL_60 == 4'h2;
  assign _EVAL_209 = _EVAL_4 & 4'h1;
  assign _EVAL_163 = _EVAL_209 == 4'h0;
  assign _EVAL_181 = _EVAL_6[31];
  assign _EVAL_234 = _EVAL_163 & _EVAL_181;
  assign _EVAL_167 = _EVAL_1[31];
  assign _EVAL_96 = _EVAL_163 & _EVAL_167;
  assign _EVAL_231 = _EVAL_234 != _EVAL_96;
  assign _EVAL_226 = _EVAL_248 == 1'h0;
  assign _EVAL_69 = _EVAL_246 & _EVAL_226;
  assign _EVAL_243 = _EVAL_196[63:32];
  assign _EVAL_23 = _EVAL_116 ? _EVAL_243 : _EVAL_34;
  assign _EVAL_174 = {_EVAL_23,_EVAL_208,_EVAL_242};
  assign _EVAL_233 = _EVAL_6[31:16];
  assign _EVAL_52 = {{31'd0}, _EVAL_208};
  assign _EVAL_250 = _EVAL_1[31:16];
  assign _EVAL_214 = _EVAL_1[15:0];
  assign _EVAL_121 = {_EVAL_96,_EVAL_250,_EVAL_214};
  assign _EVAL_200 = _EVAL_234 | _EVAL_96;
  assign _EVAL_118 = _EVAL_69 & _EVAL_38;
  assign _EVAL_78 = _EVAL_206[15:0];
  assign _EVAL_159 = _EVAL_66 == 3'h7;
  assign _EVAL_56 = _EVAL_52 << _EVAL_228;
  assign _EVAL_91 = _EVAL_118 ? {{2'd0}, _EVAL_56} : _EVAL_174;
  assign _EVAL_207 = _EVAL & _EVAL_2;
  assign _EVAL_155 = _EVAL_66 == 3'h6;
  assign _EVAL_148 = _EVAL_144 == 1'h0;
  assign _EVAL_162 = _EVAL_248 & _EVAL_148;
  assign _EVAL_199 = _EVAL_63 + 6'h1;
  assign _EVAL_217 = _EVAL_206[31:16];
  assign _EVAL_68 = _EVAL_6[15:0];
  assign _EVAL_175 = {_EVAL_233,_EVAL_68};
  assign _EVAL_3 = _EVAL_155 | _EVAL_159;
  assign _EVAL = _EVAL_66 == 3'h0;
  assign _EVAL_8 = {_EVAL_217,_EVAL_78};
  assign _EVAL_11 = _EVAL_224;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _EVAL_21 = _RAND_0[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_63 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_66 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_144 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_191 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  _EVAL_196 = _RAND_5[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_224 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_229 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_7) begin
    if (_EVAL_207) begin
      _EVAL_21 <= _EVAL_121;
    end else begin
      if (_EVAL_251) begin
        if (_EVAL_160) begin
          _EVAL_21 <= _EVAL_124;
        end
      end
    end
    if (_EVAL_207) begin
      _EVAL_63 <= 6'h0;
    end else begin
      if (_EVAL_102) begin
        if (_EVAL_118) begin
          _EVAL_63 <= {{1'd0}, _EVAL_228};
        end else begin
          _EVAL_63 <= _EVAL_199;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_66 <= 3'h0;
    end else begin
      if (_EVAL_207) begin
        if (_EVAL_200) begin
          _EVAL_66 <= 3'h1;
        end else begin
          _EVAL_66 <= 3'h3;
        end
      end else begin
        if (_EVAL_64) begin
          _EVAL_66 <= 3'h0;
        end else begin
          if (_EVAL_102) begin
            if (_EVAL_129) begin
              if (_EVAL_191) begin
                _EVAL_66 <= 3'h5;
              end else begin
                _EVAL_66 <= 3'h7;
              end
            end else begin
              if (_EVAL_39) begin
                _EVAL_66 <= 3'h7;
              end else begin
                if (_EVAL_251) begin
                  _EVAL_66 <= 3'h3;
                end
              end
            end
          end else begin
            if (_EVAL_39) begin
              _EVAL_66 <= 3'h7;
            end else begin
              if (_EVAL_251) begin
                _EVAL_66 <= 3'h3;
              end
            end
          end
        end
      end
    end
    if (_EVAL_207) begin
      _EVAL_144 <= _EVAL_133;
    end
    if (_EVAL_207) begin
      if (_EVAL_133) begin
        _EVAL_191 <= _EVAL_234;
      end else begin
        _EVAL_191 <= _EVAL_231;
      end
    end else begin
      if (_EVAL_102) begin
        if (_EVAL_162) begin
          _EVAL_191 <= 1'h0;
        end
      end
    end
    if (_EVAL_207) begin
      _EVAL_196 <= {{34'd0}, _EVAL_175};
    end else begin
      if (_EVAL_102) begin
        _EVAL_196 <= {{1'd0}, _EVAL_91};
      end else begin
        if (_EVAL_39) begin
          _EVAL_196 <= {{34'd0}, _EVAL_179};
        end else begin
          if (_EVAL_251) begin
            if (_EVAL_139) begin
              _EVAL_196 <= {{34'd0}, _EVAL_179};
            end
          end
        end
      end
    end
    if (_EVAL_207) begin
      _EVAL_224 <= _EVAL_5;
    end
    if (_EVAL_207) begin
      _EVAL_229 <= 1'h0;
    end else begin
      if (_EVAL_102) begin
        if (_EVAL_129) begin
          _EVAL_229 <= _EVAL_144;
        end else begin
          if (_EVAL_39) begin
            _EVAL_229 <= 1'h0;
          end
        end
      end else begin
        if (_EVAL_39) begin
          _EVAL_229 <= 1'h0;
        end
      end
    end
  end
endmodule
