//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_244_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [24:0] _EVAL_4,
  input         _EVAL_5,
  input  [6:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [6:0]  _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [3:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_15;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_24;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_46;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_73;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_85;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_116;
  reg [31:0] _RAND_5;
  reg [3:0] _EVAL_195;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_211;
  reg [31:0] _RAND_7;
  reg [24:0] _EVAL_216;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_223;
  reg [31:0] _RAND_9;
  reg [6:0] _EVAL_240;
  reg [31:0] _RAND_10;
  reg [72:0] _EVAL_259;
  reg [95:0] _RAND_11;
  reg [6:0] _EVAL_284;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_286;
  reg [31:0] _RAND_13;
  wire  _EVAL_63;
  wire  _EVAL_62;
  wire [12:0] _EVAL_129;
  wire [5:0] _EVAL_215;
  wire [5:0] _EVAL_56;
  wire [3:0] _EVAL_258;
  wire [3:0] _EVAL_253;
  wire [24:0] _EVAL_276;
  wire [25:0] _EVAL_283;
  wire [25:0] _EVAL_138;
  wire [25:0] _EVAL_27;
  wire  _EVAL_115;
  wire  _EVAL_152;
  wire  _EVAL_279;
  wire [127:0] _EVAL_65;
  wire [127:0] _EVAL_130;
  wire [72:0] _EVAL_232;
  wire  _EVAL_113;
  wire  _EVAL_292;
  wire [3:0] _EVAL_68;
  wire  _EVAL_213;
  wire  _EVAL_72;
  wire  _EVAL_51;
  wire  _EVAL_263;
  wire  _EVAL_228;
  wire  _EVAL_61;
  wire  _EVAL_230;
  wire  _EVAL_79;
  wire  _EVAL_256;
  wire  _EVAL_167;
  wire [1:0] _EVAL_144;
  wire [1:0] _EVAL_207;
  wire  _EVAL_169;
  wire  _EVAL_50;
  wire  _EVAL_188;
  wire  _EVAL_209;
  wire  _EVAL_25;
  wire [3:0] _EVAL_174;
  wire  _EVAL_67;
  wire  _EVAL_41;
  wire  _EVAL_187;
  wire [3:0] _EVAL_43;
  wire [3:0] _EVAL_120;
  wire  _EVAL_236;
  wire  _EVAL_89;
  wire  _EVAL_219;
  wire  _EVAL_175;
  wire  _EVAL_275;
  wire  _EVAL_19;
  wire  _EVAL_238;
  wire [2:0] _EVAL_212;
  wire  _EVAL_86;
  wire  _EVAL_206;
  wire  _EVAL_53;
  wire  _EVAL_250;
  wire  _EVAL_178;
  wire  _EVAL_98;
  wire  _EVAL_59;
  wire  _EVAL_70;
  wire  _EVAL_163;
  wire  _EVAL_166;
  wire  _EVAL_21;
  wire  _EVAL_190;
  wire  _EVAL_121;
  wire  _EVAL_108;
  wire  _EVAL_76;
  wire  _EVAL_45;
  wire  _EVAL_199;
  wire  _EVAL_31;
  wire  _EVAL_134;
  wire  _EVAL_109;
  wire  _EVAL_52;
  wire  _EVAL_269;
  wire  _EVAL_139;
  wire  _EVAL_106;
  wire  _EVAL_288;
  wire [2:0] _EVAL_28;
  wire  _EVAL_34;
  wire  _EVAL_100;
  wire  _EVAL_243;
  wire  _EVAL_176;
  wire  _EVAL_137;
  wire  _EVAL_48;
  wire  _EVAL_162;
  wire  _EVAL_42;
  wire  _EVAL_290;
  wire  _EVAL_66;
  wire  _EVAL_164;
  wire  _EVAL_40;
  wire  _EVAL_241;
  wire  _EVAL_202;
  wire [3:0] _EVAL_171;
  wire [3:0] _EVAL_118;
  wire [3:0] _EVAL_97;
  wire  _EVAL_191;
  wire  _EVAL_149;
  wire [72:0] _EVAL_177;
  wire  _EVAL_57;
  wire  _EVAL_270;
  wire  _EVAL_148;
  wire  _EVAL_155;
  wire  _EVAL_17;
  wire  _EVAL_102;
  wire [127:0] _EVAL_126;
  wire [127:0] _EVAL_194;
  wire [72:0] _EVAL_272;
  wire [72:0] _EVAL_165;
  wire [72:0] _EVAL_135;
  wire  _EVAL_231;
  wire [72:0] _EVAL_145;
  wire  _EVAL_39;
  wire  _EVAL_239;
  wire  _EVAL_142;
  wire  _EVAL_92;
  wire  _EVAL_88;
  wire  _EVAL_16;
  wire  _EVAL_257;
  wire  _EVAL_225;
  wire  _EVAL_103;
  wire  _EVAL_29;
  wire  _EVAL_136;
  wire  _EVAL_26;
  wire  _EVAL_110;
  wire  _EVAL_172;
  wire  _EVAL_104;
  wire  _EVAL_227;
  wire  _EVAL_244;
  wire [3:0] _EVAL_271;
  wire  _EVAL_93;
  wire  _EVAL_180;
  wire  _EVAL_222;
  wire  _EVAL_168;
  wire  _EVAL_37;
  wire  _EVAL_281;
  wire  _EVAL_185;
  wire  _EVAL_261;
  wire  _EVAL_60;
  wire  _EVAL_122;
  wire  _EVAL_132;
  wire  _EVAL_226;
  wire  _EVAL_252;
  wire  _EVAL_87;
  wire  _EVAL_33;
  wire  _EVAL_183;
  wire  _EVAL_274;
  wire  _EVAL_214;
  wire  _EVAL_147;
  wire  _EVAL_255;
  wire  _EVAL_99;
  wire  _EVAL_90;
  wire  _EVAL_143;
  wire  _EVAL_234;
  wire [31:0] _EVAL_248;
  wire  _EVAL_184;
  wire  _EVAL_36;
  wire  _EVAL_217;
  wire  _EVAL_30;
  wire [12:0] _EVAL_267;
  wire [5:0] _EVAL_208;
  wire [5:0] _EVAL_260;
  wire [24:0] _EVAL_265;
  wire [24:0] _EVAL_112;
  wire  _EVAL_111;
  wire  _EVAL_245;
  wire [72:0] _EVAL_233;
  wire [3:0] _EVAL_204;
  wire [3:0] _EVAL_128;
  wire  _EVAL_22;
  wire  _EVAL_181;
  wire  _EVAL_71;
  wire  _EVAL_44;
  wire  _EVAL_198;
  wire  _EVAL_119;
  wire  _EVAL_123;
  wire  _EVAL_249;
  wire  _EVAL_80;
  wire  _EVAL_84;
  wire  _EVAL_224;
  wire  _EVAL_156;
  wire  _EVAL_203;
  wire  _EVAL_158;
  wire  _EVAL_146;
  wire  _EVAL_196;
  wire  _EVAL_131;
  wire  _EVAL_264;
  wire  _EVAL_23;
  wire  _EVAL_179;
  wire  _EVAL_200;
  wire  _EVAL_273;
  wire [72:0] _EVAL_133;
  wire  _EVAL_83;
  wire  _EVAL_220;
  wire  _EVAL_154;
  wire  _EVAL_197;
  wire  _EVAL_170;
  wire  _EVAL_277;
  wire  _EVAL_193;
  wire  _EVAL_278;
  wire  _EVAL_54;
  wire  _EVAL_221;
  wire  _EVAL_55;
  wire  _EVAL_38;
  wire  _EVAL_282;
  wire  _EVAL_74;
  wire  _EVAL_82;
  wire  _EVAL_47;
  wire  _EVAL_289;
  wire  _EVAL_242;
  wire  _EVAL_161;
  wire  _EVAL_280;
  wire  _EVAL_125;
  wire  _EVAL_95;
  wire  _EVAL_205;
  wire  _EVAL_254;
  wire  _EVAL_107;
  wire  _EVAL_20;
  wire  _EVAL_32;
  wire  _EVAL_262;
  wire  _EVAL_140;
  wire  _EVAL_69;
  wire  _EVAL_189;
  wire  _EVAL_287;
  wire  _EVAL_91;
  wire  _EVAL_247;
  wire  _EVAL_49;
  wire  _EVAL_246;
  wire  _EVAL_285;
  wire  _EVAL_124;
  wire  _EVAL_77;
  wire  _EVAL_157;
  wire  _EVAL_141;
  wire  _EVAL_173;
  wire  _EVAL_186;
  wire  _EVAL_201;
  wire  _EVAL_151;
  wire  _EVAL_150;
  wire  _EVAL_58;
  wire  _EVAL_153;
  wire  _EVAL_266;
  wire  _EVAL_218;
  wire  _EVAL_160;
  wire  _EVAL_101;
  wire  _EVAL_229;
  wire  _EVAL_210;
  wire  _EVAL_127;
  wire  _EVAL_81;
  wire  _EVAL_114;
  wire  _EVAL_268;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_63 = _EVAL_211 == 4'h0;
  assign _EVAL_62 = _EVAL_1[0];
  assign _EVAL_129 = 13'h3f << _EVAL_13;
  assign _EVAL_215 = _EVAL_129[5:0];
  assign _EVAL_56 = ~ _EVAL_215;
  assign _EVAL_258 = _EVAL_56[5:2];
  assign _EVAL_253 = _EVAL_211 - 4'h1;
  assign _EVAL_276 = _EVAL_4 ^ 25'h1900000;
  assign _EVAL_283 = {1'b0,$signed(_EVAL_276)};
  assign _EVAL_138 = $signed(_EVAL_283) & $signed(-26'sh2000);
  assign _EVAL_27 = $signed(_EVAL_138);
  assign _EVAL_115 = _EVAL_8 & _EVAL;
  assign _EVAL_152 = _EVAL_46 == 4'h0;
  assign _EVAL_279 = _EVAL_115 & _EVAL_152;
  assign _EVAL_65 = 128'h1 << _EVAL_6;
  assign _EVAL_130 = _EVAL_279 ? _EVAL_65 : 128'h0;
  assign _EVAL_232 = _EVAL_130[72:0];
  assign _EVAL_113 = _EVAL_232 != 73'h0;
  assign _EVAL_292 = _EVAL_113 == 1'h0;
  assign _EVAL_68 = _EVAL_195 - 4'h1;
  assign _EVAL_213 = _EVAL_259 != 73'h0;
  assign _EVAL_72 = _EVAL_213 == 1'h0;
  assign _EVAL_51 = plusarg_reader_out == 32'h0;
  assign _EVAL_263 = _EVAL_72 | _EVAL_51;
  assign _EVAL_228 = _EVAL_24 < plusarg_reader_out;
  assign _EVAL_61 = _EVAL_263 | _EVAL_228;
  assign _EVAL_230 = _EVAL_61 | _EVAL_5;
  assign _EVAL_79 = _EVAL_230 == 1'h0;
  assign _EVAL_256 = _EVAL_3 >= 3'h2;
  assign _EVAL_167 = _EVAL_3[0];
  assign _EVAL_144 = 2'h1 << _EVAL_167;
  assign _EVAL_207 = _EVAL_144 | 2'h1;
  assign _EVAL_169 = _EVAL_207[1];
  assign _EVAL_50 = _EVAL_4[1];
  assign _EVAL_188 = _EVAL_50 == 1'h0;
  assign _EVAL_209 = _EVAL_169 & _EVAL_188;
  assign _EVAL_25 = _EVAL_256 | _EVAL_209;
  assign _EVAL_174 = _EVAL_116 - 4'h1;
  assign _EVAL_67 = _EVAL_1 <= 3'h6;
  assign _EVAL_41 = _EVAL_67 | _EVAL_5;
  assign _EVAL_187 = _EVAL_41 == 1'h0;
  assign _EVAL_43 = ~ _EVAL_14;
  assign _EVAL_120 = _EVAL_6[6:3];
  assign _EVAL_236 = _EVAL_120 == 4'h0;
  assign _EVAL_89 = _EVAL_195 == 4'h0;
  assign _EVAL_219 = _EVAL_89 == 1'h0;
  assign _EVAL_175 = _EVAL_6 == 7'h48;
  assign _EVAL_275 = _EVAL_6 == 7'h40;
  assign _EVAL_19 = _EVAL_175 | _EVAL_275;
  assign _EVAL_238 = _EVAL_120 == 4'h8;
  assign _EVAL_212 = _EVAL_6[2:0];
  assign _EVAL_86 = 3'h1 <= _EVAL_212;
  assign _EVAL_206 = _EVAL_238 & _EVAL_86;
  assign _EVAL_53 = _EVAL_19 | _EVAL_206;
  assign _EVAL_250 = _EVAL_6 == 7'h20;
  assign _EVAL_178 = _EVAL_53 | _EVAL_250;
  assign _EVAL_98 = _EVAL_178 | _EVAL_236;
  assign _EVAL_59 = _EVAL_120 == 4'h1;
  assign _EVAL_70 = _EVAL_98 | _EVAL_59;
  assign _EVAL_163 = _EVAL_120 == 4'h2;
  assign _EVAL_166 = _EVAL_70 | _EVAL_163;
  assign _EVAL_21 = _EVAL_9 == _EVAL_15;
  assign _EVAL_190 = _EVAL_169 & _EVAL_50;
  assign _EVAL_121 = _EVAL_256 | _EVAL_190;
  assign _EVAL_108 = _EVAL_207[0];
  assign _EVAL_76 = _EVAL_4[0];
  assign _EVAL_45 = _EVAL_50 & _EVAL_76;
  assign _EVAL_199 = _EVAL_108 & _EVAL_45;
  assign _EVAL_31 = _EVAL_121 | _EVAL_199;
  assign _EVAL_134 = _EVAL_115 & _EVAL_89;
  assign _EVAL_109 = _EVAL_11 == _EVAL_240;
  assign _EVAL_52 = _EVAL_0 == _EVAL_73;
  assign _EVAL_269 = _EVAL_9[2];
  assign _EVAL_139 = _EVAL_269 == 1'h0;
  assign _EVAL_106 = _EVAL_1 == 3'h1;
  assign _EVAL_288 = _EVAL_9 == 3'h2;
  assign _EVAL_28 = _EVAL_11[2:0];
  assign _EVAL_34 = _EVAL_3 <= 3'h2;
  assign _EVAL_100 = _EVAL_13 == _EVAL_85;
  assign _EVAL_243 = _EVAL_100 | _EVAL_5;
  assign _EVAL_176 = _EVAL_12 == 1'h0;
  assign _EVAL_137 = _EVAL_76 == 1'h0;
  assign _EVAL_48 = _EVAL_50 & _EVAL_137;
  assign _EVAL_162 = _EVAL_108 & _EVAL_48;
  assign _EVAL_42 = _EVAL_121 | _EVAL_162;
  assign _EVAL_290 = _EVAL_188 & _EVAL_76;
  assign _EVAL_66 = _EVAL_108 & _EVAL_290;
  assign _EVAL_164 = _EVAL_25 | _EVAL_66;
  assign _EVAL_40 = _EVAL_188 & _EVAL_137;
  assign _EVAL_241 = _EVAL_108 & _EVAL_40;
  assign _EVAL_202 = _EVAL_25 | _EVAL_241;
  assign _EVAL_171 = {_EVAL_31,_EVAL_42,_EVAL_164,_EVAL_202};
  assign _EVAL_118 = ~ _EVAL_171;
  assign _EVAL_97 = _EVAL_14 & _EVAL_118;
  assign _EVAL_191 = _EVAL_97 == 4'h0;
  assign _EVAL_149 = _EVAL_9 == 3'h3;
  assign _EVAL_177 = _EVAL_259 | _EVAL_232;
  assign _EVAL_57 = _EVAL_7 & _EVAL_2;
  assign _EVAL_270 = _EVAL_116 == 4'h0;
  assign _EVAL_148 = _EVAL_57 & _EVAL_270;
  assign _EVAL_155 = _EVAL_1 == 3'h6;
  assign _EVAL_17 = _EVAL_155 == 1'h0;
  assign _EVAL_102 = _EVAL_148 & _EVAL_17;
  assign _EVAL_126 = 128'h1 << _EVAL_11;
  assign _EVAL_194 = _EVAL_102 ? _EVAL_126 : 128'h0;
  assign _EVAL_272 = _EVAL_194[72:0];
  assign _EVAL_165 = ~ _EVAL_272;
  assign _EVAL_135 = _EVAL_177 & _EVAL_165;
  assign _EVAL_231 = _EVAL_2 & _EVAL_106;
  assign _EVAL_145 = _EVAL_232 | _EVAL_259;
  assign _EVAL_39 = _EVAL_9 == 3'h7;
  assign _EVAL_239 = _EVAL_0 <= 3'h3;
  assign _EVAL_142 = _EVAL_243 == 1'h0;
  assign _EVAL_92 = _EVAL_3 <= 3'h6;
  assign _EVAL_88 = $signed(_EVAL_27) == $signed(26'sh0);
  assign _EVAL_16 = _EVAL_92 & _EVAL_88;
  assign _EVAL_257 = _EVAL_16 | _EVAL_5;
  assign _EVAL_225 = _EVAL_257 == 1'h0;
  assign _EVAL_103 = _EVAL_9 == 3'h6;
  assign _EVAL_29 = _EVAL & _EVAL_103;
  assign _EVAL_136 = _EVAL_34 & _EVAL_88;
  assign _EVAL_26 = _EVAL_136 | _EVAL_5;
  assign _EVAL_110 = _EVAL_0 <= 3'h4;
  assign _EVAL_172 = _EVAL_110 | _EVAL_5;
  assign _EVAL_104 = _EVAL_11 == 7'h48;
  assign _EVAL_227 = _EVAL_11 == 7'h40;
  assign _EVAL_244 = _EVAL_104 | _EVAL_227;
  assign _EVAL_271 = _EVAL_11[6:3];
  assign _EVAL_93 = _EVAL_271 == 4'h8;
  assign _EVAL_180 = 3'h1 <= _EVAL_28;
  assign _EVAL_222 = _EVAL_93 & _EVAL_180;
  assign _EVAL_168 = _EVAL_244 | _EVAL_222;
  assign _EVAL_37 = _EVAL_11 == 7'h20;
  assign _EVAL_281 = _EVAL_168 | _EVAL_37;
  assign _EVAL_185 = _EVAL_271 == 4'h0;
  assign _EVAL_261 = _EVAL_281 | _EVAL_185;
  assign _EVAL_60 = _EVAL_271 == 4'h1;
  assign _EVAL_122 = _EVAL_261 | _EVAL_60;
  assign _EVAL_132 = _EVAL_271 == 4'h2;
  assign _EVAL_226 = _EVAL_122 | _EVAL_132;
  assign _EVAL_252 = _EVAL_271 == 4'h3;
  assign _EVAL_87 = _EVAL_226 | _EVAL_252;
  assign _EVAL_33 = _EVAL_191 | _EVAL_5;
  assign _EVAL_183 = _EVAL_13 >= 3'h2;
  assign _EVAL_274 = 3'h6 == _EVAL_3;
  assign _EVAL_214 = _EVAL_275 ? _EVAL_274 : 1'h0;
  assign _EVAL_147 = _EVAL_0 == 3'h0;
  assign _EVAL_255 = _EVAL_147 | _EVAL_5;
  assign _EVAL_99 = _EVAL_43 == 4'h0;
  assign _EVAL_90 = _EVAL_99 | _EVAL_5;
  assign _EVAL_143 = _EVAL_33 == 1'h0;
  assign _EVAL_234 = _EVAL_115 | _EVAL_57;
  assign _EVAL_248 = _EVAL_24 + 32'h1;
  assign _EVAL_184 = _EVAL_0 <= 3'h2;
  assign _EVAL_36 = _EVAL_184 | _EVAL_5;
  assign _EVAL_217 = _EVAL_36 == 1'h0;
  assign _EVAL_30 = _EVAL_21 | _EVAL_5;
  assign _EVAL_267 = 13'h3f << _EVAL_3;
  assign _EVAL_208 = _EVAL_267[5:0];
  assign _EVAL_260 = ~ _EVAL_208;
  assign _EVAL_265 = {{19'd0}, _EVAL_260};
  assign _EVAL_112 = _EVAL_4 & _EVAL_265;
  assign _EVAL_111 = _EVAL_120 == 4'h3;
  assign _EVAL_245 = _EVAL_1 == _EVAL_223;
  assign _EVAL_233 = _EVAL_259 >> _EVAL_6;
  assign _EVAL_204 = _EVAL_260[5:2];
  assign _EVAL_128 = _EVAL_46 - 4'h1;
  assign _EVAL_22 = _EVAL & _EVAL_219;
  assign _EVAL_181 = _EVAL_1 == 3'h4;
  assign _EVAL_71 = _EVAL_14 == _EVAL_171;
  assign _EVAL_44 = _EVAL_109 | _EVAL_5;
  assign _EVAL_198 = _EVAL_256 | _EVAL_5;
  assign _EVAL_119 = _EVAL_9 == 3'h1;
  assign _EVAL_123 = _EVAL & _EVAL_119;
  assign _EVAL_249 = _EVAL_52 | _EVAL_5;
  assign _EVAL_80 = _EVAL_249 == 1'h0;
  assign _EVAL_84 = _EVAL_232 != _EVAL_272;
  assign _EVAL_224 = _EVAL_84 | _EVAL_292;
  assign _EVAL_156 = _EVAL_9 == 3'h4;
  assign _EVAL_203 = _EVAL & _EVAL_156;
  assign _EVAL_158 = _EVAL_87 | _EVAL_5;
  assign _EVAL_146 = _EVAL_158 == 1'h0;
  assign _EVAL_196 = _EVAL_233[0];
  assign _EVAL_131 = _EVAL_44 == 1'h0;
  assign _EVAL_264 = _EVAL_9 == 3'h5;
  assign _EVAL_23 = _EVAL_214 | _EVAL_5;
  assign _EVAL_179 = _EVAL_255 == 1'h0;
  assign _EVAL_200 = _EVAL_71 | _EVAL_5;
  assign _EVAL_273 = _EVAL_63 == 1'h0;
  assign _EVAL_133 = _EVAL_145 >> _EVAL_11;
  assign _EVAL_83 = _EVAL_133[0];
  assign _EVAL_220 = _EVAL_9 == 3'h0;
  assign _EVAL_154 = _EVAL & _EVAL_220;
  assign _EVAL_197 = _EVAL_196 == 1'h0;
  assign _EVAL_170 = _EVAL_197 | _EVAL_5;
  assign _EVAL_277 = _EVAL_1 == 3'h5;
  assign _EVAL_193 = _EVAL_2 & _EVAL_277;
  assign _EVAL_278 = _EVAL_176 | _EVAL_5;
  assign _EVAL_54 = _EVAL_278 == 1'h0;
  assign _EVAL_221 = _EVAL_1 == 3'h2;
  assign _EVAL_55 = _EVAL_245 | _EVAL_5;
  assign _EVAL_38 = _EVAL_55 == 1'h0;
  assign _EVAL_282 = _EVAL_198 == 1'h0;
  assign _EVAL_74 = _EVAL_30 == 1'h0;
  assign _EVAL_82 = _EVAL_0 != 3'h0;
  assign _EVAL_47 = _EVAL_82 | _EVAL_5;
  assign _EVAL_289 = _EVAL_47 == 1'h0;
  assign _EVAL_242 = _EVAL_90 == 1'h0;
  assign _EVAL_161 = _EVAL_166 | _EVAL_111;
  assign _EVAL_280 = _EVAL_161 | _EVAL_5;
  assign _EVAL_125 = _EVAL_112 == 25'h0;
  assign _EVAL_95 = _EVAL_183 | _EVAL_5;
  assign _EVAL_205 = _EVAL_95 == 1'h0;
  assign _EVAL_254 = _EVAL_2 & _EVAL_155;
  assign _EVAL_107 = _EVAL_23 == 1'h0;
  assign _EVAL_20 = _EVAL_83 | _EVAL_5;
  assign _EVAL_32 = _EVAL_125 | _EVAL_5;
  assign _EVAL_262 = _EVAL_280 == 1'h0;
  assign _EVAL_140 = _EVAL_1 == 3'h0;
  assign _EVAL_69 = _EVAL_2 & _EVAL_140;
  assign _EVAL_189 = _EVAL_4 == _EVAL_216;
  assign _EVAL_287 = _EVAL_2 & _EVAL_221;
  assign _EVAL_91 = _EVAL & _EVAL_39;
  assign _EVAL_247 = _EVAL_239 | _EVAL_5;
  assign _EVAL_49 = _EVAL_189 | _EVAL_5;
  assign _EVAL_246 = _EVAL_6 == _EVAL_284;
  assign _EVAL_285 = _EVAL_246 | _EVAL_5;
  assign _EVAL_124 = _EVAL_3 == _EVAL_286;
  assign _EVAL_77 = _EVAL_124 | _EVAL_5;
  assign _EVAL_157 = _EVAL_77 == 1'h0;
  assign _EVAL_141 = _EVAL & _EVAL_288;
  assign _EVAL_173 = _EVAL_2 & _EVAL_273;
  assign _EVAL_186 = _EVAL_224 | _EVAL_5;
  assign _EVAL_201 = _EVAL_170 == 1'h0;
  assign _EVAL_151 = _EVAL_285 == 1'h0;
  assign _EVAL_150 = _EVAL_26 == 1'h0;
  assign _EVAL_58 = _EVAL_49 == 1'h0;
  assign _EVAL_153 = _EVAL_2 & _EVAL_181;
  assign _EVAL_266 = _EVAL_5 == 1'h0;
  assign _EVAL_218 = _EVAL_172 == 1'h0;
  assign _EVAL_160 = _EVAL_32 == 1'h0;
  assign _EVAL_101 = _EVAL_200 == 1'h0;
  assign _EVAL_229 = _EVAL_247 == 1'h0;
  assign _EVAL_210 = _EVAL_57 & _EVAL_63;
  assign _EVAL_127 = _EVAL & _EVAL_149;
  assign _EVAL_81 = _EVAL & _EVAL_264;
  assign _EVAL_114 = _EVAL_20 == 1'h0;
  assign _EVAL_268 = _EVAL_186 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_15 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_24 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_46 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_73 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_85 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_116 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_195 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_211 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_216 = _RAND_8[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_223 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_240 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {3{`RANDOM}};
  _EVAL_259 = _RAND_11[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_284 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_286 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_10) begin
    if (_EVAL_134) begin
      _EVAL_15 <= _EVAL_9;
    end
    if (_EVAL_5) begin
      _EVAL_24 <= 32'h0;
    end else begin
      if (_EVAL_234) begin
        _EVAL_24 <= 32'h0;
      end else begin
        _EVAL_24 <= _EVAL_248;
      end
    end
    if (_EVAL_5) begin
      _EVAL_46 <= 4'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_152) begin
          if (_EVAL_139) begin
            _EVAL_46 <= _EVAL_204;
          end else begin
            _EVAL_46 <= 4'h0;
          end
        end else begin
          _EVAL_46 <= _EVAL_128;
        end
      end
    end
    if (_EVAL_134) begin
      _EVAL_73 <= _EVAL_0;
    end
    if (_EVAL_210) begin
      _EVAL_85 <= _EVAL_13;
    end
    if (_EVAL_5) begin
      _EVAL_116 <= 4'h0;
    end else begin
      if (_EVAL_57) begin
        if (_EVAL_270) begin
          if (_EVAL_62) begin
            _EVAL_116 <= _EVAL_258;
          end else begin
            _EVAL_116 <= 4'h0;
          end
        end else begin
          _EVAL_116 <= _EVAL_174;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_195 <= 4'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_89) begin
          if (_EVAL_139) begin
            _EVAL_195 <= _EVAL_204;
          end else begin
            _EVAL_195 <= 4'h0;
          end
        end else begin
          _EVAL_195 <= _EVAL_68;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_211 <= 4'h0;
    end else begin
      if (_EVAL_57) begin
        if (_EVAL_63) begin
          if (_EVAL_62) begin
            _EVAL_211 <= _EVAL_258;
          end else begin
            _EVAL_211 <= 4'h0;
          end
        end else begin
          _EVAL_211 <= _EVAL_253;
        end
      end
    end
    if (_EVAL_134) begin
      _EVAL_216 <= _EVAL_4;
    end
    if (_EVAL_210) begin
      _EVAL_223 <= _EVAL_1;
    end
    if (_EVAL_210) begin
      _EVAL_240 <= _EVAL_11;
    end
    if (_EVAL_5) begin
      _EVAL_259 <= 73'h0;
    end else begin
      _EVAL_259 <= _EVAL_135;
    end
    if (_EVAL_134) begin
      _EVAL_284 <= _EVAL_6;
    end
    if (_EVAL_134) begin
      _EVAL_286 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d3367d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2adc913d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e233ca4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bba2eaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55e34dde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39fc802)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40c8866a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6b0b275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31e4a0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4da9c14b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce59452e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f97c4ba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2321fde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af013701)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b57b2d5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15e0e3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(115233eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7157c27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4579deb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(974e15b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a00a2a32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddfbff61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62b4f3d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bd27b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca9795fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31fab4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f149eb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa3343b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30f000b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5d6ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c206e30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86c1bb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cf1e6cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0a4966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4dedbd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3be5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36e9c690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f5ff776)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f99a1378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2887ee8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb61257a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e95e33e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c88a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed51617)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d4a918f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bbc0109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d589178c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e170d38e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fdab1ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27c7eb09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48a2ec51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8f6c484)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da732404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac3ac19e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c37f875a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0fe2111)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b70c55a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b26ee2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af19f0d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2718e257)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43971b33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaad7346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348fdae4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a1ab953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61396fc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71b6e8d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f78c6c7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f744d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63460ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfea3da9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44fb6fe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c92a34eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
