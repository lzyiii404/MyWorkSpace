//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_239_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [3:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_68;
  reg [31:0] _RAND_0;
  reg  _EVAL_85;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_98;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_108;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_113;
  reg [31:0] _RAND_4;
  reg [31:0] _EVAL_136;
  reg [31:0] _RAND_5;
  reg [4:0] _EVAL_140;
  reg [31:0] _RAND_6;
  reg  _EVAL_146;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_165;
  reg [31:0] _RAND_8;
  reg  _EVAL_176;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_186;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_192;
  reg [31:0] _RAND_11;
  wire  _EVAL_20;
  wire  _EVAL_97;
  wire  _EVAL_92;
  wire  _EVAL_152;
  wire  _EVAL_168;
  wire  _EVAL_49;
  wire  _EVAL_181;
  wire  _EVAL_169;
  wire  _EVAL_141;
  wire  _EVAL_38;
  wire [1:0] _EVAL_115;
  wire  _EVAL_103;
  wire  _EVAL_143;
  wire  _EVAL_64;
  wire  _EVAL_117;
  wire [31:0] _EVAL_191;
  wire [32:0] _EVAL_21;
  wire [31:0] _EVAL_51;
  wire [32:0] _EVAL_53;
  wire  _EVAL_82;
  wire  _EVAL_153;
  wire [22:0] _EVAL_123;
  wire [7:0] _EVAL_173;
  wire [7:0] _EVAL_175;
  wire  _EVAL_28;
  wire  _EVAL_182;
  wire  _EVAL_84;
  wire  _EVAL_112;
  wire  _EVAL_145;
  wire [31:0] _EVAL_17;
  wire [32:0] _EVAL_61;
  wire [32:0] _EVAL_35;
  wire [32:0] _EVAL_44;
  wire  _EVAL_27;
  wire [31:0] _EVAL_157;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_129;
  wire [32:0] _EVAL_14;
  wire  _EVAL_124;
  wire  _EVAL_130;
  wire [31:0] _EVAL_88;
  wire [32:0] _EVAL_111;
  wire [32:0] _EVAL_73;
  wire [32:0] _EVAL_170;
  wire  _EVAL_90;
  wire  _EVAL_131;
  wire [31:0] _EVAL_121;
  wire [32:0] _EVAL_48;
  wire [32:0] _EVAL_114;
  wire [32:0] _EVAL_36;
  wire  _EVAL_172;
  wire  _EVAL_72;
  wire [32:0] _EVAL_80;
  wire [32:0] _EVAL_57;
  wire [32:0] _EVAL_106;
  wire  _EVAL_26;
  wire  _EVAL_107;
  wire  _EVAL_63;
  wire [32:0] _EVAL_11;
  wire [32:0] _EVAL_139;
  wire  _EVAL_58;
  wire  _EVAL_91;
  wire [32:0] _EVAL_138;
  wire [32:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_77;
  wire [31:0] _EVAL_29;
  wire [32:0] _EVAL_156;
  wire [32:0] _EVAL_158;
  wire [32:0] _EVAL_69;
  wire  _EVAL_13;
  wire  _EVAL_101;
  wire [31:0] _EVAL_16;
  wire [32:0] _EVAL_137;
  wire [32:0] _EVAL_122;
  wire [32:0] _EVAL_41;
  wire  _EVAL_56;
  wire  _EVAL_184;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [4:0] _EVAL_190;
  wire  _EVAL_151;
  wire [4:0] _EVAL_100;
  wire [4:0] _EVAL_42;
  wire  _EVAL_178;
  wire  _EVAL_66;
  wire  _EVAL_118;
  wire [1:0] _EVAL_81;
  wire  _EVAL_110;
  wire  _EVAL_22;
  wire  _EVAL_104;
  wire  _EVAL_128;
  wire [31:0] _EVAL_164;
  wire  _EVAL_183;
  wire  _EVAL_171;
  wire  _EVAL_43;
  wire  _EVAL_179;
  wire  _EVAL_167;
  wire  _EVAL_196;
  wire  _EVAL_125;
  wire  _EVAL_166;
  wire  _EVAL_198;
  wire  _EVAL_142;
  wire  _EVAL_154;
  wire  _EVAL_149;
  wire  _EVAL_134;
  wire  _EVAL_105;
  wire  _EVAL_189;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_65;
  wire  _EVAL_197;
  wire  _EVAL_95;
  wire  _EVAL_18;
  wire  _EVAL_132;
  wire  _EVAL_34;
  wire  _EVAL_94;
  wire  _EVAL_67;
  wire [4:0] _EVAL_12;
  wire  _EVAL_193;
  wire  _EVAL_19;
  wire  _EVAL_86;
  wire  _EVAL_31;
  wire  _EVAL_96;
  wire  _EVAL_93;
  wire  _EVAL_71;
  wire  _EVAL_23;
  wire  _EVAL_40;
  wire  _EVAL_194;
  wire  _EVAL_187;
  wire  _EVAL_119;
  wire [4:0] _EVAL_174;
  wire  _EVAL_75;
  wire  _EVAL_133;
  wire  _EVAL_188;
  wire  _EVAL_127;
  wire  _EVAL_78;
  wire  _EVAL_102;
  wire  _EVAL_55;
  wire  _EVAL_70;
  wire  _EVAL_33;
  wire  _EVAL_87;
  wire  _EVAL_15;
  wire  _EVAL_62;
  wire  _EVAL_54;
  wire  _EVAL_24;
  wire  _EVAL_109;
  wire  _EVAL_159;
  wire  _EVAL_155;
  wire [31:0] _EVAL_83;
  wire  _EVAL_47;
  wire  _EVAL_126;
  wire  _EVAL_76;
  wire  _EVAL_25;
  wire  _EVAL_37;
  wire  _EVAL_39;
  wire  _EVAL_99;
  wire  _EVAL_160;
  wire  _EVAL_185;
  wire  _EVAL_52;
  wire  _EVAL_74;
  wire  _EVAL_177;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_20 = _EVAL_4 == 3'h1;
  assign _EVAL_97 = _EVAL_186 == 5'h0;
  assign _EVAL_92 = _EVAL_97 == 1'h0;
  assign _EVAL_152 = _EVAL_7 != 2'h2;
  assign _EVAL_168 = _EVAL_152 | _EVAL_0;
  assign _EVAL_49 = _EVAL_113 == 5'h0;
  assign _EVAL_181 = _EVAL_9 & _EVAL_49;
  assign _EVAL_169 = _EVAL_4 == 3'h6;
  assign _EVAL_141 = _EVAL_169 == 1'h0;
  assign _EVAL_38 = _EVAL_181 & _EVAL_141;
  assign _EVAL_115 = _EVAL_38 ? 2'h1 : 2'h0;
  assign _EVAL_103 = _EVAL_115[0];
  assign _EVAL_143 = _EVAL_176 == 1'h0;
  assign _EVAL_64 = _EVAL_143 | _EVAL_0;
  assign _EVAL_117 = _EVAL_64 == 1'h0;
  assign _EVAL_191 = _EVAL_10 ^ 32'h1800000;
  assign _EVAL_21 = {1'b0,$signed(_EVAL_191)};
  assign _EVAL_51 = _EVAL_10 ^ 32'h1900000;
  assign _EVAL_53 = {1'b0,$signed(_EVAL_51)};
  assign _EVAL_82 = _EVAL_4 <= 3'h6;
  assign _EVAL_153 = _EVAL_82 | _EVAL_0;
  assign _EVAL_123 = 23'hff << _EVAL_1;
  assign _EVAL_173 = _EVAL_123[7:0];
  assign _EVAL_175 = ~ _EVAL_173;
  assign _EVAL_28 = _EVAL_153 == 1'h0;
  assign _EVAL_182 = _EVAL_7 == _EVAL_165;
  assign _EVAL_84 = _EVAL_98 == 5'h0;
  assign _EVAL_112 = _EVAL_84 == 1'h0;
  assign _EVAL_145 = _EVAL_3 & _EVAL_112;
  assign _EVAL_17 = _EVAL_10 ^ 32'h40000000;
  assign _EVAL_61 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_35 = $signed(_EVAL_61) & $signed(-33'sh2000);
  assign _EVAL_44 = $signed(_EVAL_35);
  assign _EVAL_27 = $signed(_EVAL_44) == $signed(33'sh0);
  assign _EVAL_157 = _EVAL_10 ^ 32'h80000000;
  assign _EVAL_150 = {1'b0,$signed(_EVAL_157)};
  assign _EVAL_129 = $signed(_EVAL_150) & $signed(-33'sh20000);
  assign _EVAL_14 = $signed(_EVAL_129);
  assign _EVAL_124 = $signed(_EVAL_14) == $signed(33'sh0);
  assign _EVAL_130 = _EVAL_27 | _EVAL_124;
  assign _EVAL_88 = _EVAL_10 ^ 32'hc000000;
  assign _EVAL_111 = {1'b0,$signed(_EVAL_88)};
  assign _EVAL_73 = $signed(_EVAL_111) & $signed(-33'sh4000000);
  assign _EVAL_170 = $signed(_EVAL_73);
  assign _EVAL_90 = $signed(_EVAL_170) == $signed(33'sh0);
  assign _EVAL_131 = _EVAL_130 | _EVAL_90;
  assign _EVAL_121 = _EVAL_10 ^ 32'h2000000;
  assign _EVAL_48 = {1'b0,$signed(_EVAL_121)};
  assign _EVAL_114 = $signed(_EVAL_48) & $signed(-33'sh10000);
  assign _EVAL_36 = $signed(_EVAL_114);
  assign _EVAL_172 = $signed(_EVAL_36) == $signed(33'sh0);
  assign _EVAL_72 = _EVAL_131 | _EVAL_172;
  assign _EVAL_80 = {1'b0,$signed(_EVAL_10)};
  assign _EVAL_57 = $signed(_EVAL_80) & $signed(-33'sh5000);
  assign _EVAL_106 = $signed(_EVAL_57);
  assign _EVAL_26 = $signed(_EVAL_106) == $signed(33'sh0);
  assign _EVAL_107 = _EVAL_72 | _EVAL_26;
  assign _EVAL_63 = _EVAL_168 == 1'h0;
  assign _EVAL_11 = $signed(_EVAL_21) & $signed(-33'sh8000);
  assign _EVAL_139 = $signed(_EVAL_11);
  assign _EVAL_58 = $signed(_EVAL_139) == $signed(33'sh0);
  assign _EVAL_91 = _EVAL_107 | _EVAL_58;
  assign _EVAL_138 = $signed(_EVAL_53) & $signed(-33'sh2000);
  assign _EVAL_147 = $signed(_EVAL_138);
  assign _EVAL_148 = $signed(_EVAL_147) == $signed(33'sh0);
  assign _EVAL_77 = _EVAL_91 | _EVAL_148;
  assign _EVAL_29 = _EVAL_10 ^ 32'h20000000;
  assign _EVAL_156 = {1'b0,$signed(_EVAL_29)};
  assign _EVAL_158 = $signed(_EVAL_156) & $signed(-33'sh2000);
  assign _EVAL_69 = $signed(_EVAL_158);
  assign _EVAL_13 = $signed(_EVAL_69) == $signed(33'sh0);
  assign _EVAL_101 = _EVAL_77 | _EVAL_13;
  assign _EVAL_16 = _EVAL_10 ^ 32'h3000;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_122 = $signed(_EVAL_137) & $signed(-33'sh1000);
  assign _EVAL_41 = $signed(_EVAL_122);
  assign _EVAL_56 = $signed(_EVAL_41) == $signed(33'sh0);
  assign _EVAL_184 = _EVAL_101 | _EVAL_56;
  assign _EVAL_45 = _EVAL_184 | _EVAL_0;
  assign _EVAL_46 = _EVAL_45 == 1'h0;
  assign _EVAL_190 = _EVAL_140 - 5'h1;
  assign _EVAL_151 = _EVAL_4[0];
  assign _EVAL_100 = _EVAL_175[7:3];
  assign _EVAL_42 = _EVAL_113 - 5'h1;
  assign _EVAL_178 = _EVAL & _EVAL_3;
  assign _EVAL_66 = _EVAL_140 == 5'h0;
  assign _EVAL_118 = _EVAL_178 & _EVAL_66;
  assign _EVAL_81 = _EVAL_118 ? 2'h1 : 2'h0;
  assign _EVAL_110 = _EVAL_81[0];
  assign _EVAL_22 = _EVAL_110 | _EVAL_176;
  assign _EVAL_104 = _EVAL_22 | _EVAL_0;
  assign _EVAL_128 = _EVAL_104 == 1'h0;
  assign _EVAL_164 = _EVAL_10 & 32'h3f;
  assign _EVAL_183 = _EVAL_164 == 32'h0;
  assign _EVAL_171 = _EVAL_110 != _EVAL_103;
  assign _EVAL_43 = _EVAL_110 == 1'h0;
  assign _EVAL_179 = _EVAL_171 | _EVAL_43;
  assign _EVAL_167 = _EVAL_179 | _EVAL_0;
  assign _EVAL_196 = _EVAL_6 == 1'h0;
  assign _EVAL_125 = _EVAL_196 | _EVAL_0;
  assign _EVAL_166 = _EVAL_7 <= 2'h2;
  assign _EVAL_198 = plusarg_reader_out == 32'h0;
  assign _EVAL_142 = ~ _EVAL_103;
  assign _EVAL_154 = _EVAL_8 == 1'h0;
  assign _EVAL_149 = _EVAL_154 | _EVAL_0;
  assign _EVAL_134 = _EVAL_149 == 1'h0;
  assign _EVAL_105 = _EVAL_7 == 2'h0;
  assign _EVAL_189 = _EVAL_196 | _EVAL_8;
  assign _EVAL_59 = _EVAL_6 == _EVAL_85;
  assign _EVAL_60 = _EVAL_59 | _EVAL_0;
  assign _EVAL_65 = _EVAL_60 == 1'h0;
  assign _EVAL_197 = _EVAL_4 == 3'h5;
  assign _EVAL_95 = _EVAL_183 | _EVAL_0;
  assign _EVAL_18 = _EVAL_95 == 1'h0;
  assign _EVAL_132 = _EVAL_105 | _EVAL_0;
  assign _EVAL_34 = _EVAL_132 == 1'h0;
  assign _EVAL_94 = _EVAL_189 | _EVAL_0;
  assign _EVAL_67 = _EVAL_94 == 1'h0;
  assign _EVAL_12 = _EVAL_98 - 5'h1;
  assign _EVAL_193 = _EVAL_176 | _EVAL_110;
  assign _EVAL_19 = _EVAL_182 | _EVAL_0;
  assign _EVAL_86 = _EVAL_4 == 3'h0;
  assign _EVAL_31 = _EVAL_9 & _EVAL_86;
  assign _EVAL_96 = _EVAL_1 >= 4'h3;
  assign _EVAL_93 = _EVAL_96 | _EVAL_0;
  assign _EVAL_71 = _EVAL_10 == _EVAL_192;
  assign _EVAL_23 = _EVAL_71 | _EVAL_0;
  assign _EVAL_40 = _EVAL_23 == 1'h0;
  assign _EVAL_194 = _EVAL_5 == _EVAL_146;
  assign _EVAL_187 = _EVAL_194 | _EVAL_0;
  assign _EVAL_119 = _EVAL_93 == 1'h0;
  assign _EVAL_174 = _EVAL_186 - 5'h1;
  assign _EVAL_75 = _EVAL_1 == _EVAL_68;
  assign _EVAL_133 = _EVAL_75 | _EVAL_0;
  assign _EVAL_188 = _EVAL_133 == 1'h0;
  assign _EVAL_127 = _EVAL_143 | _EVAL_198;
  assign _EVAL_78 = _EVAL_136 < plusarg_reader_out;
  assign _EVAL_102 = _EVAL_127 | _EVAL_78;
  assign _EVAL_55 = _EVAL_102 | _EVAL_0;
  assign _EVAL_70 = _EVAL_55 == 1'h0;
  assign _EVAL_33 = _EVAL_125 == 1'h0;
  assign _EVAL_87 = _EVAL_166 | _EVAL_0;
  assign _EVAL_15 = _EVAL_19 == 1'h0;
  assign _EVAL_62 = _EVAL_9 & _EVAL_197;
  assign _EVAL_54 = _EVAL_178 | _EVAL_9;
  assign _EVAL_24 = _EVAL_4 == 3'h4;
  assign _EVAL_109 = _EVAL_9 & _EVAL_24;
  assign _EVAL_159 = _EVAL_9 & _EVAL_92;
  assign _EVAL_155 = _EVAL_9 & _EVAL_97;
  assign _EVAL_83 = _EVAL_136 + 32'h1;
  assign _EVAL_47 = _EVAL_187 == 1'h0;
  assign _EVAL_126 = _EVAL_9 & _EVAL_20;
  assign _EVAL_76 = _EVAL_4 == 3'h2;
  assign _EVAL_25 = _EVAL_9 & _EVAL_76;
  assign _EVAL_37 = _EVAL_87 == 1'h0;
  assign _EVAL_39 = _EVAL_4 == _EVAL_108;
  assign _EVAL_99 = _EVAL_39 | _EVAL_0;
  assign _EVAL_160 = _EVAL_99 == 1'h0;
  assign _EVAL_185 = _EVAL_9 & _EVAL_169;
  assign _EVAL_52 = _EVAL_193 & _EVAL_142;
  assign _EVAL_74 = _EVAL_178 & _EVAL_84;
  assign _EVAL_177 = _EVAL_167 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_68 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_85 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_98 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_108 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_113 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_136 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_140 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_146 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_165 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_176 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_186 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_192 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_155) begin
      _EVAL_68 <= _EVAL_1;
    end
    if (_EVAL_155) begin
      _EVAL_85 <= _EVAL_6;
    end
    if (_EVAL_0) begin
      _EVAL_98 <= 5'h0;
    end else begin
      if (_EVAL_178) begin
        if (_EVAL_84) begin
          _EVAL_98 <= 5'h0;
        end else begin
          _EVAL_98 <= _EVAL_12;
        end
      end
    end
    if (_EVAL_155) begin
      _EVAL_108 <= _EVAL_4;
    end
    if (_EVAL_0) begin
      _EVAL_113 <= 5'h0;
    end else begin
      if (_EVAL_9) begin
        if (_EVAL_49) begin
          if (_EVAL_151) begin
            _EVAL_113 <= _EVAL_100;
          end else begin
            _EVAL_113 <= 5'h0;
          end
        end else begin
          _EVAL_113 <= _EVAL_42;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_136 <= 32'h0;
    end else begin
      if (_EVAL_54) begin
        _EVAL_136 <= 32'h0;
      end else begin
        _EVAL_136 <= _EVAL_83;
      end
    end
    if (_EVAL_0) begin
      _EVAL_140 <= 5'h0;
    end else begin
      if (_EVAL_178) begin
        if (_EVAL_66) begin
          _EVAL_140 <= 5'h0;
        end else begin
          _EVAL_140 <= _EVAL_190;
        end
      end
    end
    if (_EVAL_155) begin
      _EVAL_146 <= _EVAL_5;
    end
    if (_EVAL_155) begin
      _EVAL_165 <= _EVAL_7;
    end
    if (_EVAL_0) begin
      _EVAL_176 <= 1'h0;
    end else begin
      _EVAL_176 <= _EVAL_52;
    end
    if (_EVAL_0) begin
      _EVAL_186 <= 5'h0;
    end else begin
      if (_EVAL_9) begin
        if (_EVAL_97) begin
          if (_EVAL_151) begin
            _EVAL_186 <= _EVAL_100;
          end else begin
            _EVAL_186 <= 5'h0;
          end
        end else begin
          _EVAL_186 <= _EVAL_174;
        end
      end
    end
    if (_EVAL_74) begin
      _EVAL_192 <= _EVAL_10;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e39f6578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8c66ba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f9a4af1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce594e1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf9f9f05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65f68e46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5f1bab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71f1faf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70687f32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ff19ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccd4d8fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7ffea41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15e56f7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17c9becd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc993a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a97b0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67c3c708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e552d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10604e32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5910deb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcf2e9bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(965a4b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27005f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8432b23a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d489700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e2d2dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(470d89f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9940759)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b7acce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60377c9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2611c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
