//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_2(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  input         _EVAL_1,
  output [6:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  output [6:0]  _EVAL_4,
  output [7:0]  _EVAL_5,
  output [3:0]  _EVAL_6,
  output [2:0]  _EVAL_7,
  output [2:0]  _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  input  [2:0]  _EVAL_11,
  output [31:0] _EVAL_12,
  input  [31:0] _EVAL_13,
  output [2:0]  _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output [2:0]  _EVAL_17,
  output [2:0]  _EVAL_18,
  output [63:0] _EVAL_19,
  input  [6:0]  _EVAL_20,
  input  [63:0] _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output [6:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  output [3:0]  _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  input  [1:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input  [6:0]  _EVAL_34,
  output [2:0]  _EVAL_35,
  input         _EVAL_36,
  output [2:0]  _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input  [3:0]  _EVAL_40,
  output [2:0]  _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  input  [2:0]  _EVAL_45,
  output        _EVAL_46,
  input  [63:0] _EVAL_47,
  input  [2:0]  _EVAL_48,
  input         _EVAL_49,
  output        _EVAL_50,
  input         _EVAL_51,
  output [63:0] _EVAL_52,
  output [31:0] _EVAL_53,
  input         _EVAL_54,
  output [29:0] _EVAL_55,
  input  [3:0]  _EVAL_56,
  output        _EVAL_57,
  output [2:0]  _EVAL_58,
  input  [1:0]  _EVAL_59,
  input         _EVAL_60,
  input  [2:0]  _EVAL_61,
  input  [2:0]  _EVAL_62,
  output        _EVAL_63,
  output        _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  input  [7:0]  _EVAL_67,
  input  [1:0]  _EVAL_68,
  input  [31:0] _EVAL_69,
  output [63:0] _EVAL_70,
  input  [3:0]  _EVAL_71,
  output        _EVAL_72,
  output        _EVAL_73,
  input         _EVAL_74,
  output [2:0]  _EVAL_75,
  input  [63:0] _EVAL_76,
  input  [3:0]  _EVAL_77,
  output        _EVAL_78,
  input  [63:0] _EVAL_79,
  output [1:0]  _EVAL_80,
  output        _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  input  [6:0]  _EVAL_85,
  output        _EVAL_86,
  output [63:0] _EVAL_87,
  output [7:0]  _EVAL_88,
  output [5:0]  _EVAL_89,
  input  [2:0]  _EVAL_90,
  input         _EVAL_91,
  output        _EVAL_92,
  output [7:0]  _EVAL_93,
  output [63:0] _EVAL_94,
  input  [3:0]  _EVAL_95,
  output        _EVAL_96,
  output        _EVAL_97,
  input  [2:0]  _EVAL_98,
  input         _EVAL_99,
  input         _EVAL_100,
  input         _EVAL_101,
  output [3:0]  _EVAL_102,
  input         _EVAL_103,
  output [3:0]  _EVAL_104,
  output        _EVAL_105,
  output        _EVAL_106,
  output        _EVAL_107,
  output [2:0]  _EVAL_108,
  output [1:0]  _EVAL_109,
  output [1:0]  _EVAL_110,
  output [63:0] _EVAL_111,
  input  [63:0] _EVAL_112,
  input         _EVAL_113,
  input  [31:0] _EVAL_114,
  output        _EVAL_115,
  output [30:0] _EVAL_116,
  input  [3:0]  _EVAL_117,
  input  [2:0]  _EVAL_118,
  input  [63:0] _EVAL_119,
  output        _EVAL_120,
  input  [7:0]  _EVAL_121,
  input         _EVAL_122,
  input         _EVAL_123,
  input         _EVAL_124,
  output [6:0]  _EVAL_125,
  input         _EVAL_126,
  input  [5:0]  _EVAL_127,
  output [2:0]  _EVAL_128
);
  reg [2:0] _EVAL_131;
  reg [31:0] _RAND_0;
  reg  _EVAL_193;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_202;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_211;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_223;
  reg [31:0] _RAND_4;
  reg  _EVAL_242;
  reg [31:0] _RAND_5;
  reg [1:0] _EVAL_253;
  reg [31:0] _RAND_6;
  reg  _EVAL_273;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_278;
  reg [31:0] _RAND_8;
  reg  _EVAL_318;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_321;
  reg [31:0] _RAND_10;
  reg  _EVAL_324;
  reg [31:0] _RAND_11;
  reg  _EVAL_409;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_432;
  reg [31:0] _RAND_13;
  reg  _EVAL_433;
  reg [31:0] _RAND_14;
  reg  _EVAL_458;
  reg [31:0] _RAND_15;
  reg [1:0] _EVAL_486;
  reg [31:0] _RAND_16;
  reg [4:0] _EVAL_508;
  reg [31:0] _RAND_17;
  reg  _EVAL_567;
  reg [31:0] _RAND_18;
  reg  _EVAL_574;
  reg [31:0] _RAND_19;
  reg  _EVAL_613;
  reg [31:0] _RAND_20;
  reg  _EVAL_619;
  reg [31:0] _RAND_21;
  wire  _EVAL_501;
  wire [32:0] _EVAL_513;
  wire [32:0] _EVAL_312;
  wire [32:0] _EVAL_585;
  wire  _EVAL_461;
  wire  _EVAL_500;
  wire [32:0] _EVAL_533;
  wire [32:0] _EVAL_276;
  wire [32:0] _EVAL_234;
  wire  _EVAL_505;
  wire  _EVAL_538;
  wire  _EVAL_366;
  wire  _EVAL_628;
  wire  _EVAL_244;
  wire  _EVAL_445;
  wire  _EVAL_381;
  wire [31:0] _EVAL_323;
  wire [32:0] _EVAL_622;
  wire [32:0] _EVAL_602;
  wire [32:0] _EVAL_308;
  wire  _EVAL_153;
  wire  _EVAL_210;
  wire [22:0] _EVAL_272;
  wire [7:0] _EVAL_469;
  wire [7:0] _EVAL_420;
  wire [2:0] _EVAL_402;
  wire  _EVAL_201;
  wire  _EVAL_416;
  wire [2:0] _EVAL_541;
  wire  _EVAL_224;
  wire  _EVAL_277;
  wire [2:0] _EVAL_512;
  wire  _EVAL_293;
  wire  _EVAL_164;
  wire [2:0] _EVAL_261;
  wire [2:0] _EVAL_334;
  wire [2:0] _EVAL_499;
  wire [5:0] _EVAL_236;
  wire [4:0] _EVAL_150;
  wire [5:0] _EVAL_418;
  wire  _EVAL_610;
  wire [1:0] _EVAL_441;
  wire  _EVAL_491;
  wire  _EVAL_403;
  wire [1:0] _EVAL_426;
  wire [1:0] _EVAL_296;
  wire [3:0] _EVAL_478;
  wire [2:0] _EVAL_399;
  wire [3:0] _EVAL_181;
  wire [3:0] _EVAL_596;
  wire [2:0] _EVAL_382;
  wire [3:0] _EVAL_477;
  wire [3:0] _EVAL_415;
  wire [3:0] _EVAL_481;
  wire [1:0] _EVAL_145;
  wire [1:0] _EVAL_454;
  wire [1:0] _EVAL_337;
  wire [1:0] _EVAL_397;
  wire [1:0] _EVAL_136;
  wire [2:0] _EVAL_480;
  wire [1:0] _EVAL_171;
  wire [1:0] _EVAL_190;
  wire [31:0] _EVAL_262;
  wire [32:0] _EVAL_226;
  wire [32:0] _EVAL_355;
  wire [32:0] _EVAL_392;
  wire  _EVAL_249;
  wire  _EVAL_525;
  wire [31:0] _EVAL_496;
  wire [32:0] _EVAL_372;
  wire [32:0] _EVAL_564;
  wire [32:0] _EVAL_571;
  wire  _EVAL_615;
  wire  _EVAL_137;
  wire  _EVAL_178;
  wire [31:0] _EVAL_186;
  wire [32:0] _EVAL_365;
  wire [32:0] _EVAL_265;
  wire [32:0] _EVAL_266;
  wire  _EVAL_600;
  wire  _EVAL_142;
  wire [1:0] _EVAL_229;
  wire  _EVAL_373;
  wire [5:0] _EVAL_175;
  wire [3:0] _EVAL_487;
  wire [5:0] _EVAL_459;
  wire [5:0] _EVAL_280;
  wire [4:0] _EVAL_268;
  wire [5:0] _EVAL_221;
  wire [5:0] _EVAL_309;
  wire [5:0] _EVAL_146;
  wire [2:0] _EVAL_603;
  wire [2:0] _EVAL_322;
  wire [2:0] _EVAL_450;
  wire [2:0] _EVAL_274;
  wire  _EVAL_594;
  wire  _EVAL_435;
  wire  _EVAL_161;
  wire  _EVAL_520;
  wire  _EVAL_562;
  wire  _EVAL_460;
  wire [22:0] _EVAL_182;
  wire [7:0] _EVAL_453;
  wire [7:0] _EVAL_383;
  wire  _EVAL_184;
  wire  _EVAL_297;
  wire [1:0] _EVAL_140;
  wire [1:0] _EVAL_447;
  wire [1:0] _EVAL_475;
  wire [3:0] _EVAL_588;
  wire [2:0] _EVAL_356;
  wire  _EVAL_160;
  wire  _EVAL_436;
  wire [22:0] _EVAL_401;
  wire [7:0] _EVAL_431;
  wire [7:0] _EVAL_605;
  wire [4:0] _EVAL_172;
  wire [4:0] _EVAL_389;
  wire [4:0] _EVAL_540;
  wire  _EVAL_446;
  wire  _EVAL_479;
  wire  _EVAL_568;
  wire  _EVAL_414;
  wire [4:0] _EVAL_346;
  wire [4:0] _EVAL_183;
  wire [4:0] _EVAL_177;
  wire [4:0] _EVAL_377;
  wire  _EVAL_517;
  wire [1:0] _EVAL_452;
  wire [1:0] _EVAL_255;
  wire [3:0] _EVAL_618;
  wire [2:0] _EVAL_302;
  wire [3:0] _EVAL_314;
  wire [3:0] _EVAL_144;
  wire [2:0] _EVAL_404;
  wire [3:0] _EVAL_492;
  wire [3:0] _EVAL_300;
  wire [3:0] _EVAL_287;
  wire [1:0] _EVAL_609;
  wire [1:0] _EVAL_154;
  wire [1:0] _EVAL_173;
  wire [1:0] _EVAL_188;
  wire  _EVAL_582;
  wire  _EVAL_341;
  wire  _EVAL_621;
  wire [6:0] _EVAL_497;
  wire [6:0] _EVAL_561;
  wire [121:0] _EVAL_529;
  wire [121:0] _EVAL_316;
  wire  _EVAL_400;
  wire  _EVAL_166;
  wire  _EVAL_176;
  wire [6:0] _EVAL_271;
  wire [121:0] _EVAL_521;
  wire [121:0] _EVAL_546;
  wire [121:0] _EVAL_345;
  wire  _EVAL_370;
  wire  _EVAL_206;
  wire  _EVAL_214;
  wire  _EVAL_509;
  wire  _EVAL_200;
  wire  _EVAL_319;
  wire  _EVAL_537;
  wire  _EVAL_472;
  wire  _EVAL_374;
  wire  _EVAL_130;
  wire  _EVAL_148;
  wire  _EVAL_379;
  wire  _EVAL_483;
  wire  _EVAL_215;
  wire  _EVAL_290;
  wire  _EVAL_625;
  wire  _EVAL_591;
  wire  _EVAL_359;
  wire  _EVAL_554;
  wire  _EVAL_573;
  wire  _EVAL_428;
  wire  _EVAL_199;
  wire  _EVAL_209;
  wire  _EVAL_256;
  wire [4:0] _EVAL_163;
  wire [4:0] _EVAL_451;
  wire [1:0] _EVAL_132;
  wire [4:0] _EVAL_299;
  wire  _EVAL_326;
  wire [3:0] _EVAL_336;
  wire [3:0] _EVAL_343;
  wire [3:0] _EVAL_231;
  wire [2:0] _EVAL_134;
  wire [3:0] _EVAL_471;
  wire [3:0] _EVAL_557;
  wire [3:0] _EVAL_463;
  wire [1:0] _EVAL_257;
  wire [1:0] _EVAL_289;
  wire [1:0] _EVAL_553;
  wire [1:0] _EVAL_230;
  wire [1:0] _EVAL_456;
  wire  _EVAL_158;
  wire  _EVAL_547;
  wire  _EVAL_180;
  wire  _EVAL_283;
  wire  _EVAL_443;
  wire  _EVAL_248;
  wire [4:0] _EVAL_129;
  wire [4:0] _EVAL_398;
  wire  _EVAL_327;
  wire  _EVAL_282;
  wire  _EVAL_539;
  wire  _EVAL_135;
  wire  _EVAL_419;
  wire [4:0] _EVAL_468;
  wire [2:0] _EVAL_620;
  wire [2:0] _EVAL_507;
  wire [2:0] _EVAL_335;
  wire [5:0] _EVAL_522;
  wire [4:0] _EVAL_353;
  wire [5:0] _EVAL_310;
  wire [5:0] _EVAL_412;
  wire [3:0] _EVAL_207;
  wire [5:0] _EVAL_387;
  wire [5:0] _EVAL_320;
  wire [4:0] _EVAL_608;
  wire [5:0] _EVAL_331;
  wire [5:0] _EVAL_213;
  wire [5:0] _EVAL_330;
  wire [2:0] _EVAL_587;
  wire [2:0] _EVAL_169;
  wire [3:0] _EVAL_294;
  wire [2:0] _EVAL_368;
  wire [2:0] _EVAL_284;
  wire [4:0] _EVAL_208;
  wire [2:0] _EVAL_246;
  wire [2:0] _EVAL_504;
  wire [2:0] _EVAL_344;
  wire  _EVAL_565;
  wire  _EVAL_563;
  wire  _EVAL_203;
  wire [3:0] _EVAL_576;
  wire [20:0] _EVAL_250;
  wire [5:0] _EVAL_216;
  wire [5:0] _EVAL_580;
  wire [2:0] _EVAL_578;
  wire [2:0] _EVAL_592;
  wire [2:0] _EVAL_581;
  wire  _EVAL_386;
  wire  _EVAL_490;
  wire [3:0] _EVAL_225;
  wire [20:0] _EVAL_473;
  wire [5:0] _EVAL_270;
  wire [5:0] _EVAL_254;
  wire  _EVAL_498;
  wire [4:0] _EVAL_228;
  wire [82:0] _EVAL_306;
  wire  _EVAL_222;
  wire  _EVAL_251;
  wire  _EVAL_198;
  wire  _EVAL_275;
  wire  _EVAL_376;
  wire  _EVAL_523;
  wire [4:0] _EVAL_219;
  wire  _EVAL_194;
  wire  _EVAL_422;
  wire [4:0] _EVAL_577;
  wire [4:0] _EVAL_307;
  wire  _EVAL_442;
  wire  _EVAL_364;
  wire  _EVAL_349;
  wire  _EVAL_348;
  wire  _EVAL_133;
  wire [4:0] _EVAL_362;
  wire [4:0] _EVAL_332;
  wire  _EVAL_267;
  wire  _EVAL_503;
  wire  _EVAL_360;
  wire  _EVAL_185;
  wire [121:0] _EVAL_558;
  wire  _EVAL_339;
  wire [82:0] _EVAL_626;
  wire  _EVAL_288;
  wire [82:0] _EVAL_485;
  wire [82:0] _EVAL_515;
  wire [82:0] _EVAL_559;
  wire  _EVAL_524;
  wire [82:0] _EVAL_434;
  wire [82:0] _EVAL_555;
  wire [82:0] _EVAL_396;
  wire  _EVAL_239;
  wire  _EVAL_196;
  wire  _EVAL_217;
  wire  _EVAL_488;
  wire  _EVAL_425;
  wire  _EVAL_187;
  wire  _EVAL_506;
  wire [4:0] _EVAL_241;
  wire [4:0] _EVAL_298;
  wire [4:0] _EVAL_474;
  wire [2:0] _EVAL_351;
  wire [1:0] _EVAL_511;
  wire [1:0] _EVAL_484;
  wire [4:0] _EVAL_162;
  wire  _EVAL_410;
  wire [4:0] _EVAL_590;
  wire [2:0] _EVAL_179;
  wire [4:0] _EVAL_357;
  wire  _EVAL_220;
  wire  _EVAL_227;
  wire  _EVAL_139;
  wire  _EVAL_566;
  wire [2:0] _EVAL_338;
  wire [2:0] _EVAL_449;
  wire [2:0] _EVAL_531;
  wire [2:0] _EVAL_495;
  wire  _EVAL_519;
  wire  _EVAL_593;
  wire [2:0] _EVAL_354;
  wire [1:0] _EVAL_192;
  wire [1:0] _EVAL_240;
  wire  _EVAL_384;
  wire [121:0] _EVAL_313;
  wire [121:0] _EVAL_394;
  wire [31:0] _EVAL_439;
  wire  _EVAL_437;
  wire [82:0] _EVAL_624;
  wire [2:0] _EVAL_548;
  wire [3:0] _EVAL_380;
  wire [2:0] _EVAL_575;
  wire [2:0] _EVAL_502;
  wire [4:0] _EVAL_589;
  wire  _EVAL_358;
  wire  _EVAL_157;
  wire  _EVAL_149;
  wire  _EVAL_612;
  wire  _EVAL_466;
  wire  _EVAL_604;
  wire  _EVAL_536;
  wire  _EVAL_350;
  wire [2:0] _EVAL_204;
  wire [2:0] _EVAL_584;
  wire  _EVAL_407;
  wire  _EVAL_421;
  wire  _EVAL_385;
  wire  _EVAL_311;
  wire [4:0] _EVAL_627;
  wire [4:0] _EVAL_467;
  wire [121:0] _EVAL_601;
  wire  _EVAL_550;
  wire [121:0] _EVAL_281;
  wire [121:0] _EVAL_245;
  wire [6:0] _EVAL_235;
  wire  _EVAL_347;
  wire  _EVAL_464;
  wire  _EVAL_406;
  wire  _EVAL_340;
  wire  _EVAL_598;
  wire  _EVAL_417;
  wire  _EVAL_333;
  wire  _EVAL_325;
  wire  _EVAL_408;
  wire [2:0] _EVAL_371;
  wire [2:0] _EVAL_607;
  wire [2:0] _EVAL_514;
  wire [4:0] _EVAL_361;
  wire [4:0] _EVAL_532;
  wire  _EVAL_595;
  wire [4:0] _EVAL_388;
  wire [4:0] _EVAL_526;
  wire  _EVAL_159;
  wire  _EVAL_597;
  wire [2:0] _EVAL_151;
  wire  _EVAL_342;
  wire  _EVAL_569;
  wire [82:0] _EVAL_405;
  wire  _EVAL_430;
  wire [82:0] _EVAL_189;
  wire [82:0] _EVAL_455;
  wire [82:0] _EVAL_614;
  wire  _EVAL_518;
  wire  _EVAL_378;
  wire  _EVAL_243;
  wire  _EVAL_476;
  wire  _EVAL_263;
  wire [6:0] _EVAL_170;
  wire [31:0] _EVAL_191;
  wire [6:0] _EVAL_247;
  wire  _EVAL_429;
  wire  _EVAL_623;
  wire  _EVAL_424;
  wire [3:0] _EVAL_391;
  assign _EVAL_501 = _EVAL_223 == 5'h0;
  assign _EVAL_513 = {1'b0,$signed(_EVAL_33)};
  assign _EVAL_312 = $signed(_EVAL_513) & $signed(33'shc0000000);
  assign _EVAL_585 = $signed(_EVAL_312);
  assign _EVAL_461 = $signed(_EVAL_585) == $signed(33'sh0);
  assign _EVAL_500 = _EVAL_54 & _EVAL_461;
  assign _EVAL_533 = {1'b0,$signed(_EVAL_13)};
  assign _EVAL_276 = $signed(_EVAL_533) & $signed(33'shc0000000);
  assign _EVAL_234 = $signed(_EVAL_276);
  assign _EVAL_505 = $signed(_EVAL_234) == $signed(33'sh0);
  assign _EVAL_538 = _EVAL_84 & _EVAL_505;
  assign _EVAL_366 = _EVAL_500 | _EVAL_538;
  assign _EVAL_628 = _EVAL_433 ? _EVAL_500 : 1'h0;
  assign _EVAL_244 = _EVAL_619 ? _EVAL_538 : 1'h0;
  assign _EVAL_445 = _EVAL_628 | _EVAL_244;
  assign _EVAL_381 = _EVAL_501 ? _EVAL_366 : _EVAL_445;
  assign _EVAL_323 = _EVAL_13 ^ 32'h80000000;
  assign _EVAL_622 = {1'b0,$signed(_EVAL_323)};
  assign _EVAL_602 = $signed(_EVAL_622) & $signed(33'shc0000000);
  assign _EVAL_308 = $signed(_EVAL_602);
  assign _EVAL_153 = $signed(_EVAL_308) == $signed(33'sh0);
  assign _EVAL_210 = _EVAL_84 & _EVAL_153;
  assign _EVAL_272 = 23'hff << _EVAL_95;
  assign _EVAL_469 = _EVAL_272[7:0];
  assign _EVAL_420 = ~ _EVAL_469;
  assign _EVAL_402 = _EVAL_20[6:4];
  assign _EVAL_201 = _EVAL_402 == 3'h4;
  assign _EVAL_416 = _EVAL_126 & _EVAL_201;
  assign _EVAL_541 = _EVAL_85[6:4];
  assign _EVAL_224 = _EVAL_541 == 3'h4;
  assign _EVAL_277 = _EVAL_39 & _EVAL_224;
  assign _EVAL_512 = _EVAL_34[6:4];
  assign _EVAL_293 = _EVAL_512 == 3'h4;
  assign _EVAL_164 = _EVAL_123 & _EVAL_293;
  assign _EVAL_261 = {_EVAL_416,_EVAL_277,_EVAL_164};
  assign _EVAL_334 = ~ _EVAL_131;
  assign _EVAL_499 = _EVAL_261 & _EVAL_334;
  assign _EVAL_236 = {_EVAL_499,_EVAL_416,_EVAL_277,_EVAL_164};
  assign _EVAL_150 = _EVAL_236[5:1];
  assign _EVAL_418 = {{1'd0}, _EVAL_150};
  assign _EVAL_610 = _EVAL_501 & _EVAL_49;
  assign _EVAL_441 = {_EVAL_538,_EVAL_500};
  assign _EVAL_491 = _EVAL_441 != 2'h0;
  assign _EVAL_403 = _EVAL_610 & _EVAL_491;
  assign _EVAL_426 = ~ _EVAL_278;
  assign _EVAL_296 = _EVAL_441 & _EVAL_426;
  assign _EVAL_478 = {_EVAL_296,_EVAL_538,_EVAL_500};
  assign _EVAL_399 = _EVAL_478[3:1];
  assign _EVAL_181 = {{1'd0}, _EVAL_399};
  assign _EVAL_596 = _EVAL_478 | _EVAL_181;
  assign _EVAL_382 = _EVAL_596[3:1];
  assign _EVAL_477 = {{1'd0}, _EVAL_382};
  assign _EVAL_415 = {_EVAL_278, 2'h0};
  assign _EVAL_481 = _EVAL_477 | _EVAL_415;
  assign _EVAL_145 = _EVAL_481[3:2];
  assign _EVAL_454 = _EVAL_481[1:0];
  assign _EVAL_337 = _EVAL_145 & _EVAL_454;
  assign _EVAL_397 = ~ _EVAL_337;
  assign _EVAL_136 = _EVAL_397 & _EVAL_441;
  assign _EVAL_480 = {_EVAL_136, 1'h0};
  assign _EVAL_171 = _EVAL_480[1:0];
  assign _EVAL_190 = _EVAL_136 | _EVAL_171;
  assign _EVAL_262 = _EVAL_33 ^ 32'h40000000;
  assign _EVAL_226 = {1'b0,$signed(_EVAL_262)};
  assign _EVAL_355 = $signed(_EVAL_226) & $signed(33'shc0000000);
  assign _EVAL_392 = $signed(_EVAL_355);
  assign _EVAL_249 = $signed(_EVAL_392) == $signed(33'sh0);
  assign _EVAL_525 = _EVAL_54 & _EVAL_249;
  assign _EVAL_496 = _EVAL_13 ^ 32'h40000000;
  assign _EVAL_372 = {1'b0,$signed(_EVAL_496)};
  assign _EVAL_564 = $signed(_EVAL_372) & $signed(33'shc0000000);
  assign _EVAL_571 = $signed(_EVAL_564);
  assign _EVAL_615 = $signed(_EVAL_571) == $signed(33'sh0);
  assign _EVAL_137 = _EVAL_84 & _EVAL_615;
  assign _EVAL_178 = _EVAL_525 | _EVAL_137;
  assign _EVAL_186 = _EVAL_33 ^ 32'h80000000;
  assign _EVAL_365 = {1'b0,$signed(_EVAL_186)};
  assign _EVAL_265 = $signed(_EVAL_365) & $signed(33'shc0000000);
  assign _EVAL_266 = $signed(_EVAL_265);
  assign _EVAL_600 = $signed(_EVAL_266) == $signed(33'sh0);
  assign _EVAL_142 = _EVAL_54 & _EVAL_600;
  assign _EVAL_229 = {_EVAL_210,_EVAL_142};
  assign _EVAL_373 = _EVAL_229 != 2'h0;
  assign _EVAL_175 = _EVAL_236 | _EVAL_418;
  assign _EVAL_487 = _EVAL_175[5:2];
  assign _EVAL_459 = {{2'd0}, _EVAL_487};
  assign _EVAL_280 = _EVAL_175 | _EVAL_459;
  assign _EVAL_268 = _EVAL_280[5:1];
  assign _EVAL_221 = {{1'd0}, _EVAL_268};
  assign _EVAL_309 = {_EVAL_131, 3'h0};
  assign _EVAL_146 = _EVAL_221 | _EVAL_309;
  assign _EVAL_603 = _EVAL_146[5:3];
  assign _EVAL_322 = _EVAL_146[2:0];
  assign _EVAL_450 = _EVAL_603 & _EVAL_322;
  assign _EVAL_274 = ~ _EVAL_450;
  assign _EVAL_594 = _EVAL_274[0];
  assign _EVAL_435 = _EVAL_594 & _EVAL_164;
  assign _EVAL_161 = _EVAL_274[1];
  assign _EVAL_520 = _EVAL_161 & _EVAL_277;
  assign _EVAL_562 = _EVAL_274[2];
  assign _EVAL_460 = _EVAL_562 & _EVAL_416;
  assign _EVAL_182 = 23'hff << _EVAL_117;
  assign _EVAL_453 = _EVAL_182[7:0];
  assign _EVAL_383 = ~ _EVAL_453;
  assign _EVAL_184 = _EVAL_397[0];
  assign _EVAL_297 = _EVAL_184 & _EVAL_500;
  assign _EVAL_140 = {_EVAL_137,_EVAL_525};
  assign _EVAL_447 = ~ _EVAL_486;
  assign _EVAL_475 = _EVAL_140 & _EVAL_447;
  assign _EVAL_588 = {_EVAL_475,_EVAL_137,_EVAL_525};
  assign _EVAL_356 = _EVAL_588[3:1];
  assign _EVAL_160 = _EVAL_61[2];
  assign _EVAL_436 = _EVAL_160 == 1'h0;
  assign _EVAL_401 = 23'hff << _EVAL_40;
  assign _EVAL_431 = _EVAL_401[7:0];
  assign _EVAL_605 = ~ _EVAL_431;
  assign _EVAL_172 = _EVAL_605[7:3];
  assign _EVAL_389 = _EVAL_436 ? _EVAL_172 : 5'h0;
  assign _EVAL_540 = _EVAL_297 ? _EVAL_389 : 5'h0;
  assign _EVAL_446 = _EVAL_397[1];
  assign _EVAL_479 = _EVAL_446 & _EVAL_538;
  assign _EVAL_568 = _EVAL_45[2];
  assign _EVAL_414 = _EVAL_568 == 1'h0;
  assign _EVAL_346 = _EVAL_383[7:3];
  assign _EVAL_183 = _EVAL_414 ? _EVAL_346 : 5'h0;
  assign _EVAL_177 = _EVAL_479 ? _EVAL_183 : 5'h0;
  assign _EVAL_377 = _EVAL_540 | _EVAL_177;
  assign _EVAL_517 = _EVAL_432 == 5'h0;
  assign _EVAL_452 = ~ _EVAL_253;
  assign _EVAL_255 = _EVAL_229 & _EVAL_452;
  assign _EVAL_618 = {_EVAL_255,_EVAL_210,_EVAL_142};
  assign _EVAL_302 = _EVAL_618[3:1];
  assign _EVAL_314 = {{1'd0}, _EVAL_302};
  assign _EVAL_144 = _EVAL_618 | _EVAL_314;
  assign _EVAL_404 = _EVAL_144[3:1];
  assign _EVAL_492 = {{1'd0}, _EVAL_404};
  assign _EVAL_300 = {_EVAL_253, 2'h0};
  assign _EVAL_287 = _EVAL_492 | _EVAL_300;
  assign _EVAL_609 = _EVAL_287[3:2];
  assign _EVAL_154 = _EVAL_287[1:0];
  assign _EVAL_173 = _EVAL_609 & _EVAL_154;
  assign _EVAL_188 = ~ _EVAL_173;
  assign _EVAL_582 = _EVAL_188[0];
  assign _EVAL_341 = _EVAL_582 & _EVAL_142;
  assign _EVAL_621 = _EVAL_517 ? _EVAL_341 : _EVAL_613;
  assign _EVAL_497 = {{3'd0}, _EVAL_71};
  assign _EVAL_561 = _EVAL_497 | 7'h40;
  assign _EVAL_529 = {_EVAL_61,_EVAL_90,_EVAL_40,_EVAL_561,_EVAL_33,_EVAL_67,_EVAL_76,_EVAL_42};
  assign _EVAL_316 = _EVAL_621 ? _EVAL_529 : 122'h0;
  assign _EVAL_400 = _EVAL_188[1];
  assign _EVAL_166 = _EVAL_400 & _EVAL_210;
  assign _EVAL_176 = _EVAL_517 ? _EVAL_166 : _EVAL_574;
  assign _EVAL_271 = {{1'd0}, _EVAL_127};
  assign _EVAL_521 = {_EVAL_45,_EVAL_3,_EVAL_117,_EVAL_271,_EVAL_13,_EVAL_121,_EVAL_79,_EVAL_15};
  assign _EVAL_546 = _EVAL_176 ? _EVAL_521 : 122'h0;
  assign _EVAL_345 = _EVAL_316 | _EVAL_546;
  assign _EVAL_370 = _EVAL_34[6:6];
  assign _EVAL_206 = _EVAL_370 == 1'h0;
  assign _EVAL_214 = _EVAL_123 & _EVAL_206;
  assign _EVAL_509 = _EVAL_324 ? _EVAL_214 : 1'h0;
  assign _EVAL_200 = _EVAL_85[6:6];
  assign _EVAL_319 = _EVAL_200 == 1'h0;
  assign _EVAL_537 = _EVAL_39 & _EVAL_319;
  assign _EVAL_472 = _EVAL_193 ? _EVAL_537 : 1'h0;
  assign _EVAL_374 = _EVAL_509 | _EVAL_472;
  assign _EVAL_130 = _EVAL_20[6:6];
  assign _EVAL_148 = _EVAL_130 == 1'h0;
  assign _EVAL_379 = _EVAL_126 & _EVAL_148;
  assign _EVAL_483 = _EVAL_242 ? _EVAL_379 : 1'h0;
  assign _EVAL_215 = _EVAL_374 | _EVAL_483;
  assign _EVAL_290 = _EVAL_321 == 5'h0;
  assign _EVAL_625 = _EVAL_164 | _EVAL_277;
  assign _EVAL_591 = _EVAL_625 | _EVAL_416;
  assign _EVAL_359 = _EVAL_273 ? _EVAL_164 : 1'h0;
  assign _EVAL_554 = _EVAL_409 ? _EVAL_277 : 1'h0;
  assign _EVAL_573 = _EVAL_359 | _EVAL_554;
  assign _EVAL_428 = _EVAL_567 ? _EVAL_416 : 1'h0;
  assign _EVAL_199 = _EVAL_573 | _EVAL_428;
  assign _EVAL_209 = _EVAL_290 ? _EVAL_591 : _EVAL_199;
  assign _EVAL_256 = _EVAL_38 & _EVAL_209;
  assign _EVAL_163 = {{4'd0}, _EVAL_256};
  assign _EVAL_451 = _EVAL_321 - _EVAL_163;
  assign _EVAL_132 = _EVAL_188 & _EVAL_229;
  assign _EVAL_299 = _EVAL_166 ? _EVAL_183 : 5'h0;
  assign _EVAL_326 = _EVAL_290 ? _EVAL_562 : _EVAL_567;
  assign _EVAL_336 = _EVAL_345[115:112];
  assign _EVAL_343 = {{1'd0}, _EVAL_356};
  assign _EVAL_231 = _EVAL_588 | _EVAL_343;
  assign _EVAL_134 = _EVAL_231[3:1];
  assign _EVAL_471 = {{1'd0}, _EVAL_134};
  assign _EVAL_557 = {_EVAL_486, 2'h0};
  assign _EVAL_463 = _EVAL_471 | _EVAL_557;
  assign _EVAL_257 = _EVAL_463[3:2];
  assign _EVAL_289 = _EVAL_463[1:0];
  assign _EVAL_553 = _EVAL_257 & _EVAL_289;
  assign _EVAL_230 = ~ _EVAL_553;
  assign _EVAL_456 = _EVAL_230 & _EVAL_140;
  assign _EVAL_158 = _EVAL_142 | _EVAL_210;
  assign _EVAL_547 = _EVAL_613 ? _EVAL_142 : 1'h0;
  assign _EVAL_180 = _EVAL_574 ? _EVAL_210 : 1'h0;
  assign _EVAL_283 = _EVAL_547 | _EVAL_180;
  assign _EVAL_443 = _EVAL_517 ? _EVAL_158 : _EVAL_283;
  assign _EVAL_248 = _EVAL_83 & _EVAL_443;
  assign _EVAL_129 = {{4'd0}, _EVAL_248};
  assign _EVAL_398 = _EVAL_432 - _EVAL_129;
  assign _EVAL_327 = _EVAL_508 == 5'h0;
  assign _EVAL_282 = _EVAL_214 | _EVAL_537;
  assign _EVAL_539 = _EVAL_282 | _EVAL_379;
  assign _EVAL_135 = _EVAL_327 ? _EVAL_539 : _EVAL_215;
  assign _EVAL_419 = _EVAL_60 & _EVAL_135;
  assign _EVAL_468 = {{4'd0}, _EVAL_419};
  assign _EVAL_620 = {_EVAL_379,_EVAL_537,_EVAL_214};
  assign _EVAL_507 = ~ _EVAL_211;
  assign _EVAL_335 = _EVAL_620 & _EVAL_507;
  assign _EVAL_522 = {_EVAL_335,_EVAL_379,_EVAL_537,_EVAL_214};
  assign _EVAL_353 = _EVAL_522[5:1];
  assign _EVAL_310 = {{1'd0}, _EVAL_353};
  assign _EVAL_412 = _EVAL_522 | _EVAL_310;
  assign _EVAL_207 = _EVAL_412[5:2];
  assign _EVAL_387 = {{2'd0}, _EVAL_207};
  assign _EVAL_320 = _EVAL_412 | _EVAL_387;
  assign _EVAL_608 = _EVAL_320[5:1];
  assign _EVAL_331 = {{1'd0}, _EVAL_608};
  assign _EVAL_213 = {_EVAL_211, 3'h0};
  assign _EVAL_330 = _EVAL_331 | _EVAL_213;
  assign _EVAL_587 = _EVAL_330[2:0];
  assign _EVAL_169 = _EVAL_274 & _EVAL_261;
  assign _EVAL_294 = {_EVAL_169, 1'h0};
  assign _EVAL_368 = _EVAL_294[2:0];
  assign _EVAL_284 = _EVAL_169 | _EVAL_368;
  assign _EVAL_208 = {_EVAL_284, 2'h0};
  assign _EVAL_246 = _EVAL_330[5:3];
  assign _EVAL_504 = _EVAL_246 & _EVAL_587;
  assign _EVAL_344 = ~ _EVAL_504;
  assign _EVAL_565 = _EVAL_344[0];
  assign _EVAL_563 = _EVAL_565 & _EVAL_214;
  assign _EVAL_203 = _EVAL_118[0];
  assign _EVAL_576 = {{1'd0}, _EVAL_48};
  assign _EVAL_250 = 21'h3f << _EVAL_576;
  assign _EVAL_216 = _EVAL_250[5:0];
  assign _EVAL_580 = ~ _EVAL_216;
  assign _EVAL_578 = _EVAL_580[5:3];
  assign _EVAL_592 = _EVAL_203 ? _EVAL_578 : 3'h0;
  assign _EVAL_581 = _EVAL_563 ? _EVAL_592 : 3'h0;
  assign _EVAL_386 = _EVAL_501 ? _EVAL_446 : _EVAL_619;
  assign _EVAL_490 = _EVAL_49 & _EVAL_386;
  assign _EVAL_225 = {{1'd0}, _EVAL_22};
  assign _EVAL_473 = 21'h3f << _EVAL_225;
  assign _EVAL_270 = _EVAL_473[5:0];
  assign _EVAL_254 = ~ _EVAL_270;
  assign _EVAL_498 = _EVAL_344[2];
  assign _EVAL_228 = _EVAL_508 - _EVAL_468;
  assign _EVAL_306 = {_EVAL_118,2'h0,_EVAL_576,_EVAL_34,1'h0,_EVAL_99,_EVAL_21,_EVAL};
  assign _EVAL_222 = _EVAL_327 ? _EVAL_565 : _EVAL_324;
  assign _EVAL_251 = _EVAL_60 & _EVAL_222;
  assign _EVAL_198 = _EVAL_202 == 5'h0;
  assign _EVAL_275 = _EVAL_198 & _EVAL_100;
  assign _EVAL_376 = _EVAL_230[0];
  assign _EVAL_523 = _EVAL_376 & _EVAL_525;
  assign _EVAL_219 = _EVAL_523 ? _EVAL_389 : 5'h0;
  assign _EVAL_194 = _EVAL_230[1];
  assign _EVAL_422 = _EVAL_194 & _EVAL_137;
  assign _EVAL_577 = _EVAL_422 ? _EVAL_183 : 5'h0;
  assign _EVAL_307 = _EVAL_219 | _EVAL_577;
  assign _EVAL_442 = _EVAL_458 ? _EVAL_525 : 1'h0;
  assign _EVAL_364 = _EVAL_318 ? _EVAL_137 : 1'h0;
  assign _EVAL_349 = _EVAL_442 | _EVAL_364;
  assign _EVAL_348 = _EVAL_198 ? _EVAL_178 : _EVAL_349;
  assign _EVAL_133 = _EVAL_100 & _EVAL_348;
  assign _EVAL_362 = {{4'd0}, _EVAL_133};
  assign _EVAL_332 = _EVAL_202 - _EVAL_362;
  assign _EVAL_267 = _EVAL_517 ? _EVAL_400 : _EVAL_574;
  assign _EVAL_503 = _EVAL_83 & _EVAL_267;
  assign _EVAL_360 = _EVAL_153 ? _EVAL_503 : 1'h0;
  assign _EVAL_185 = _EVAL_501 ? _EVAL_479 : _EVAL_619;
  assign _EVAL_558 = _EVAL_185 ? _EVAL_521 : 122'h0;
  assign _EVAL_339 = _EVAL_290 ? _EVAL_435 : _EVAL_273;
  assign _EVAL_626 = _EVAL_339 ? _EVAL_306 : 83'h0;
  assign _EVAL_288 = _EVAL_290 ? _EVAL_520 : _EVAL_409;
  assign _EVAL_485 = {_EVAL_11,_EVAL_59,_EVAL_225,_EVAL_85,_EVAL_74,_EVAL_24,_EVAL_47,_EVAL_124};
  assign _EVAL_515 = _EVAL_288 ? _EVAL_485 : 83'h0;
  assign _EVAL_559 = _EVAL_626 | _EVAL_515;
  assign _EVAL_524 = _EVAL_290 ? _EVAL_460 : _EVAL_567;
  assign _EVAL_434 = {_EVAL_98,_EVAL_68,_EVAL_95,_EVAL_20,_EVAL_91,_EVAL_43,_EVAL_112,_EVAL_23};
  assign _EVAL_555 = _EVAL_524 ? _EVAL_434 : 83'h0;
  assign _EVAL_396 = _EVAL_559 | _EVAL_555;
  assign _EVAL_239 = _EVAL_517 ? _EVAL_582 : _EVAL_613;
  assign _EVAL_196 = _EVAL_83 & _EVAL_239;
  assign _EVAL_217 = _EVAL_327 ? _EVAL_498 : _EVAL_242;
  assign _EVAL_488 = _EVAL_60 & _EVAL_217;
  assign _EVAL_425 = _EVAL_148 ? _EVAL_488 : 1'h0;
  assign _EVAL_187 = _EVAL_498 & _EVAL_379;
  assign _EVAL_506 = _EVAL_98[0];
  assign _EVAL_241 = _EVAL_420[7:3];
  assign _EVAL_298 = _EVAL_506 ? _EVAL_241 : 5'h0;
  assign _EVAL_474 = _EVAL_187 ? _EVAL_298 : 5'h0;
  assign _EVAL_351 = {_EVAL_132, 1'h0};
  assign _EVAL_511 = _EVAL_351[1:0];
  assign _EVAL_484 = _EVAL_132 | _EVAL_511;
  assign _EVAL_162 = _EVAL_460 ? _EVAL_298 : 5'h0;
  assign _EVAL_410 = _EVAL_49 & _EVAL_381;
  assign _EVAL_590 = {{4'd0}, _EVAL_410};
  assign _EVAL_179 = _EVAL_208[2:0];
  assign _EVAL_357 = _EVAL_223 - _EVAL_590;
  assign _EVAL_220 = _EVAL_327 & _EVAL_60;
  assign _EVAL_227 = _EVAL_344[1];
  assign _EVAL_139 = _EVAL_227 & _EVAL_537;
  assign _EVAL_566 = _EVAL_11[0];
  assign _EVAL_338 = _EVAL_254[5:3];
  assign _EVAL_449 = _EVAL_566 ? _EVAL_338 : 3'h0;
  assign _EVAL_531 = _EVAL_139 ? _EVAL_449 : 3'h0;
  assign _EVAL_495 = _EVAL_581 | _EVAL_531;
  assign _EVAL_519 = _EVAL_198 ? _EVAL_523 : _EVAL_458;
  assign _EVAL_593 = _EVAL_140 != 2'h0;
  assign _EVAL_354 = {_EVAL_456, 1'h0};
  assign _EVAL_192 = _EVAL_354[1:0];
  assign _EVAL_240 = _EVAL_456 | _EVAL_192;
  assign _EVAL_384 = _EVAL_501 ? _EVAL_297 : _EVAL_433;
  assign _EVAL_313 = _EVAL_384 ? _EVAL_529 : 122'h0;
  assign _EVAL_394 = _EVAL_313 | _EVAL_558;
  assign _EVAL_439 = _EVAL_394[104:73];
  assign _EVAL_437 = _EVAL_327 ? _EVAL_187 : _EVAL_242;
  assign _EVAL_624 = _EVAL_437 ? _EVAL_434 : 83'h0;
  assign _EVAL_548 = _EVAL_344 & _EVAL_620;
  assign _EVAL_380 = {_EVAL_548, 1'h0};
  assign _EVAL_575 = _EVAL_380[2:0];
  assign _EVAL_502 = _EVAL_548 | _EVAL_575;
  assign _EVAL_589 = {_EVAL_502, 2'h0};
  assign _EVAL_358 = _EVAL_290 ? _EVAL_594 : _EVAL_273;
  assign _EVAL_157 = _EVAL_327 ? _EVAL_227 : _EVAL_193;
  assign _EVAL_149 = _EVAL_60 & _EVAL_157;
  assign _EVAL_612 = _EVAL_319 ? _EVAL_149 : 1'h0;
  assign _EVAL_466 = _EVAL_501 ? _EVAL_184 : _EVAL_433;
  assign _EVAL_604 = _EVAL_49 & _EVAL_466;
  assign _EVAL_536 = _EVAL_620 != 3'h0;
  assign _EVAL_350 = _EVAL_220 & _EVAL_536;
  assign _EVAL_204 = _EVAL_589[2:0];
  assign _EVAL_584 = _EVAL_502 | _EVAL_204;
  assign _EVAL_407 = _EVAL_198 ? _EVAL_194 : _EVAL_318;
  assign _EVAL_421 = _EVAL_100 & _EVAL_407;
  assign _EVAL_385 = _EVAL_615 ? _EVAL_421 : 1'h0;
  assign _EVAL_311 = _EVAL_385 | _EVAL_360;
  assign _EVAL_627 = _EVAL_341 ? _EVAL_389 : 5'h0;
  assign _EVAL_467 = _EVAL_627 | _EVAL_299;
  assign _EVAL_601 = _EVAL_519 ? _EVAL_529 : 122'h0;
  assign _EVAL_550 = _EVAL_198 ? _EVAL_422 : _EVAL_318;
  assign _EVAL_281 = _EVAL_550 ? _EVAL_521 : 122'h0;
  assign _EVAL_245 = _EVAL_601 | _EVAL_281;
  assign _EVAL_235 = _EVAL_396[73:67];
  assign _EVAL_347 = _EVAL_327 ? _EVAL_563 : _EVAL_324;
  assign _EVAL_464 = _EVAL_517 & _EVAL_83;
  assign _EVAL_406 = _EVAL_464 & _EVAL_373;
  assign _EVAL_340 = _EVAL_290 ? _EVAL_161 : _EVAL_409;
  assign _EVAL_598 = _EVAL_38 & _EVAL_340;
  assign _EVAL_417 = _EVAL_224 ? _EVAL_598 : 1'h0;
  assign _EVAL_333 = _EVAL_198 ? _EVAL_376 : _EVAL_458;
  assign _EVAL_325 = _EVAL_100 & _EVAL_333;
  assign _EVAL_408 = _EVAL_249 ? _EVAL_325 : 1'h0;
  assign _EVAL_371 = _EVAL_435 ? _EVAL_592 : 3'h0;
  assign _EVAL_607 = _EVAL_520 ? _EVAL_449 : 3'h0;
  assign _EVAL_514 = _EVAL_371 | _EVAL_607;
  assign _EVAL_361 = {{2'd0}, _EVAL_514};
  assign _EVAL_532 = _EVAL_361 | _EVAL_162;
  assign _EVAL_595 = _EVAL_261 != 3'h0;
  assign _EVAL_388 = {{2'd0}, _EVAL_495};
  assign _EVAL_526 = _EVAL_388 | _EVAL_474;
  assign _EVAL_159 = _EVAL_290 & _EVAL_38;
  assign _EVAL_597 = _EVAL_159 & _EVAL_595;
  assign _EVAL_151 = _EVAL_284 | _EVAL_179;
  assign _EVAL_342 = _EVAL_600 ? _EVAL_196 : 1'h0;
  assign _EVAL_569 = _EVAL_408 | _EVAL_342;
  assign _EVAL_405 = _EVAL_347 ? _EVAL_306 : 83'h0;
  assign _EVAL_430 = _EVAL_327 ? _EVAL_139 : _EVAL_193;
  assign _EVAL_189 = _EVAL_430 ? _EVAL_485 : 83'h0;
  assign _EVAL_455 = _EVAL_405 | _EVAL_189;
  assign _EVAL_614 = _EVAL_455 | _EVAL_624;
  assign _EVAL_518 = _EVAL_275 & _EVAL_593;
  assign _EVAL_378 = _EVAL_461 ? _EVAL_604 : 1'h0;
  assign _EVAL_243 = _EVAL_505 ? _EVAL_490 : 1'h0;
  assign _EVAL_476 = _EVAL_38 & _EVAL_326;
  assign _EVAL_263 = _EVAL_201 ? _EVAL_476 : 1'h0;
  assign _EVAL_170 = _EVAL_614[73:67];
  assign _EVAL_191 = _EVAL_245[104:73];
  assign _EVAL_247 = {{3'd0}, _EVAL_56};
  assign _EVAL_429 = _EVAL_38 & _EVAL_358;
  assign _EVAL_623 = _EVAL_293 ? _EVAL_429 : 1'h0;
  assign _EVAL_424 = _EVAL_206 ? _EVAL_251 : 1'h0;
  assign _EVAL_391 = _EVAL_245[115:112];
  assign _EVAL_64 = _EVAL_569 | _EVAL_378;
  assign _EVAL_70 = _EVAL_394[64:1];
  assign _EVAL_87 = _EVAL_245[64:1];
  assign _EVAL_110 = _EVAL_396[79:78];
  assign _EVAL_29 = _EVAL_417 | _EVAL_612;
  assign _EVAL_80 = _EVAL_31;
  assign _EVAL_41 = _EVAL_394[121:119];
  assign _EVAL_63 = _EVAL_113;
  assign _EVAL_4 = _EVAL_394[111:105];
  assign _EVAL_96 = _EVAL_290 ? _EVAL_591 : _EVAL_199;
  assign _EVAL_108 = _EVAL_32;
  assign _EVAL_7 = _EVAL_614[82:80];
  assign _EVAL_65 = _EVAL_311 | _EVAL_243;
  assign _EVAL_2 = _EVAL_245[111:105];
  assign _EVAL_27 = _EVAL_114;
  assign _EVAL_19 = _EVAL_119;
  assign _EVAL_5 = _EVAL_394[72:65];
  assign _EVAL_58 = _EVAL_336[2:0];
  assign _EVAL_89 = _EVAL_170[5:0];
  assign _EVAL_72 = _EVAL_396[65];
  assign _EVAL_73 = _EVAL_517 ? _EVAL_158 : _EVAL_283;
  assign _EVAL_25 = _EVAL_82;
  assign _EVAL_120 = _EVAL_103;
  assign _EVAL_35 = _EVAL_245[118:116];
  assign _EVAL_115 = _EVAL_345[0];
  assign _EVAL_57 = _EVAL_614[0];
  assign _EVAL_66 = _EVAL_614[65];
  assign _EVAL_78 = _EVAL_245[0];
  assign _EVAL_93 = _EVAL_245[72:65];
  assign _EVAL_88 = _EVAL_345[72:65];
  assign _EVAL_8 = _EVAL_345[121:119];
  assign _EVAL_105 = _EVAL_198 ? _EVAL_178 : _EVAL_349;
  assign _EVAL_128 = _EVAL_396[82:80];
  assign _EVAL_28 = _EVAL_235[3:0];
  assign _EVAL_106 = _EVAL_9;
  assign _EVAL_6 = _EVAL_614[77:74];
  assign _EVAL_55 = _EVAL_439[29:0];
  assign _EVAL_26 = _EVAL_345[111:105];
  assign _EVAL_16 = _EVAL_396[0];
  assign _EVAL_10 = _EVAL_122;
  assign _EVAL_104 = _EVAL_396[77:74];
  assign _EVAL_107 = _EVAL_36;
  assign _EVAL_37 = _EVAL_77[2:0];
  assign _EVAL_53 = _EVAL_345[104:73];
  assign _EVAL_94 = _EVAL_345[64:1];
  assign _EVAL_30 = _EVAL_501 ? _EVAL_366 : _EVAL_445;
  assign _EVAL_14 = _EVAL_245[121:119];
  assign _EVAL_81 = _EVAL_396[66];
  assign _EVAL_109 = _EVAL_614[79:78];
  assign _EVAL_12 = _EVAL_69;
  assign _EVAL_125 = _EVAL_247 | 7'h40;
  assign _EVAL_18 = _EVAL_345[118:116];
  assign _EVAL_17 = _EVAL_62;
  assign _EVAL_46 = _EVAL_623 | _EVAL_424;
  assign _EVAL_44 = _EVAL_327 ? _EVAL_539 : _EVAL_215;
  assign _EVAL_102 = _EVAL_394[115:112];
  assign _EVAL_116 = _EVAL_191[30:0];
  assign _EVAL_86 = _EVAL_263 | _EVAL_425;
  assign _EVAL_111 = _EVAL_396[64:1];
  assign _EVAL_97 = _EVAL_614[66];
  assign _EVAL_50 = _EVAL_1;
  assign _EVAL_75 = _EVAL_394[118:116];
  assign _EVAL_52 = _EVAL_614[64:1];
  assign _EVAL_92 = _EVAL_394[0];
  assign _EVAL_0 = _EVAL_391[2:0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_131 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_193 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_202 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_211 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_223 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_242 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_253 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_273 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_278 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_318 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_321 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_324 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_409 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_432 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_433 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_458 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_486 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_508 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_567 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_574 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_613 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_619 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_101) begin
    if (_EVAL_51) begin
      _EVAL_131 <= 3'h7;
    end else begin
      if (_EVAL_597) begin
        _EVAL_131 <= _EVAL_151;
      end
    end
    if (_EVAL_51) begin
      _EVAL_193 <= 1'h0;
    end else begin
      if (_EVAL_327) begin
        _EVAL_193 <= _EVAL_139;
      end
    end
    if (_EVAL_51) begin
      _EVAL_202 <= 5'h0;
    end else begin
      if (_EVAL_275) begin
        _EVAL_202 <= _EVAL_307;
      end else begin
        _EVAL_202 <= _EVAL_332;
      end
    end
    if (_EVAL_51) begin
      _EVAL_211 <= 3'h7;
    end else begin
      if (_EVAL_350) begin
        _EVAL_211 <= _EVAL_584;
      end
    end
    if (_EVAL_51) begin
      _EVAL_223 <= 5'h0;
    end else begin
      if (_EVAL_610) begin
        _EVAL_223 <= _EVAL_377;
      end else begin
        _EVAL_223 <= _EVAL_357;
      end
    end
    if (_EVAL_51) begin
      _EVAL_242 <= 1'h0;
    end else begin
      if (_EVAL_327) begin
        _EVAL_242 <= _EVAL_187;
      end
    end
    if (_EVAL_51) begin
      _EVAL_253 <= 2'h3;
    end else begin
      if (_EVAL_406) begin
        _EVAL_253 <= _EVAL_484;
      end
    end
    if (_EVAL_51) begin
      _EVAL_273 <= 1'h0;
    end else begin
      if (_EVAL_290) begin
        _EVAL_273 <= _EVAL_435;
      end
    end
    if (_EVAL_51) begin
      _EVAL_278 <= 2'h3;
    end else begin
      if (_EVAL_403) begin
        _EVAL_278 <= _EVAL_190;
      end
    end
    if (_EVAL_51) begin
      _EVAL_318 <= 1'h0;
    end else begin
      if (_EVAL_198) begin
        _EVAL_318 <= _EVAL_422;
      end
    end
    if (_EVAL_51) begin
      _EVAL_321 <= 5'h0;
    end else begin
      if (_EVAL_159) begin
        _EVAL_321 <= _EVAL_532;
      end else begin
        _EVAL_321 <= _EVAL_451;
      end
    end
    if (_EVAL_51) begin
      _EVAL_324 <= 1'h0;
    end else begin
      if (_EVAL_327) begin
        _EVAL_324 <= _EVAL_563;
      end
    end
    if (_EVAL_51) begin
      _EVAL_409 <= 1'h0;
    end else begin
      if (_EVAL_290) begin
        _EVAL_409 <= _EVAL_520;
      end
    end
    if (_EVAL_51) begin
      _EVAL_432 <= 5'h0;
    end else begin
      if (_EVAL_464) begin
        _EVAL_432 <= _EVAL_467;
      end else begin
        _EVAL_432 <= _EVAL_398;
      end
    end
    if (_EVAL_51) begin
      _EVAL_433 <= 1'h0;
    end else begin
      if (_EVAL_501) begin
        _EVAL_433 <= _EVAL_297;
      end
    end
    if (_EVAL_51) begin
      _EVAL_458 <= 1'h0;
    end else begin
      if (_EVAL_198) begin
        _EVAL_458 <= _EVAL_523;
      end
    end
    if (_EVAL_51) begin
      _EVAL_486 <= 2'h3;
    end else begin
      if (_EVAL_518) begin
        _EVAL_486 <= _EVAL_240;
      end
    end
    if (_EVAL_51) begin
      _EVAL_508 <= 5'h0;
    end else begin
      if (_EVAL_220) begin
        _EVAL_508 <= _EVAL_526;
      end else begin
        _EVAL_508 <= _EVAL_228;
      end
    end
    if (_EVAL_51) begin
      _EVAL_567 <= 1'h0;
    end else begin
      if (_EVAL_290) begin
        _EVAL_567 <= _EVAL_460;
      end
    end
    if (_EVAL_51) begin
      _EVAL_574 <= 1'h0;
    end else begin
      if (_EVAL_517) begin
        _EVAL_574 <= _EVAL_166;
      end
    end
    if (_EVAL_51) begin
      _EVAL_613 <= 1'h0;
    end else begin
      if (_EVAL_517) begin
        _EVAL_613 <= _EVAL_341;
      end
    end
    if (_EVAL_51) begin
      _EVAL_619 <= 1'h0;
    end else begin
      if (_EVAL_501) begin
        _EVAL_619 <= _EVAL_479;
      end
    end
  end
endmodule
