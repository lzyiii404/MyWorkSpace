//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_39(
  input         _EVAL,
  input         _EVAL_0,
  output [30:0] _EVAL_1,
  output        _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  input  [3:0]  _EVAL_8,
  output [2:0]  _EVAL_9,
  output [3:0]  _EVAL_10,
  input  [31:0] _EVAL_11,
  output [2:0]  _EVAL_12,
  output [1:0]  _EVAL_13,
  output [30:0] _EVAL_14,
  input  [1:0]  _EVAL_15,
  input         _EVAL_16,
  output [3:0]  _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  output [3:0]  _EVAL_20,
  output        _EVAL_21,
  output        _EVAL_22,
  output [2:0]  _EVAL_23,
  output [6:0]  _EVAL_24,
  input         _EVAL_25,
  output [3:0]  _EVAL_26,
  output        _EVAL_27,
  input         _EVAL_28,
  output [3:0]  _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  output [3:0]  _EVAL_32,
  output        _EVAL_33,
  output [7:0]  _EVAL_34,
  input         _EVAL_35,
  output        _EVAL_36,
  input         _EVAL_37,
  output [1:0]  _EVAL_38,
  input  [6:0]  _EVAL_39,
  output [2:0]  _EVAL_40,
  output [2:0]  _EVAL_41,
  input         _EVAL_42,
  input  [1:0]  _EVAL_43,
  output [31:0] _EVAL_44,
  input  [30:0] _EVAL_45,
  output [3:0]  _EVAL_46,
  input  [3:0]  _EVAL_47,
  input  [7:0]  _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input  [2:0]  _EVAL_51,
  output [63:0] _EVAL_52,
  input  [63:0] _EVAL_53,
  output [7:0]  _EVAL_54,
  output [2:0]  _EVAL_55
);
  wire  axi4index__EVAL;
  wire  axi4index__EVAL_0;
  wire [31:0] axi4index__EVAL_1;
  wire [10:0] axi4index__EVAL_2;
  wire [3:0] axi4index__EVAL_3;
  wire [10:0] axi4index__EVAL_4;
  wire  axi4index__EVAL_5;
  wire  axi4index__EVAL_6;
  wire [3:0] axi4index__EVAL_7;
  wire [3:0] axi4index__EVAL_8;
  wire [3:0] axi4index__EVAL_9;
  wire  axi4index__EVAL_10;
  wire  axi4index__EVAL_11;
  wire [7:0] axi4index__EVAL_12;
  wire  axi4index__EVAL_13;
  wire [10:0] axi4index__EVAL_14;
  wire [3:0] axi4index__EVAL_15;
  wire [10:0] axi4index__EVAL_16;
  wire [10:0] axi4index__EVAL_17;
  wire [1:0] axi4index__EVAL_18;
  wire  axi4index__EVAL_19;
  wire [3:0] axi4index__EVAL_20;
  wire [3:0] axi4index__EVAL_21;
  wire  axi4index__EVAL_22;
  wire [2:0] axi4index__EVAL_23;
  wire  axi4index__EVAL_24;
  wire  axi4index__EVAL_25;
  wire [31:0] axi4index__EVAL_26;
  wire [7:0] axi4index__EVAL_27;
  wire  axi4index__EVAL_28;
  wire [2:0] axi4index__EVAL_29;
  wire  axi4index__EVAL_30;
  wire  axi4index__EVAL_31;
  wire [1:0] axi4index__EVAL_32;
  wire [3:0] axi4index__EVAL_33;
  wire [2:0] axi4index__EVAL_34;
  wire  axi4index__EVAL_35;
  wire [3:0] axi4index__EVAL_36;
  wire [31:0] axi4index__EVAL_37;
  wire [30:0] axi4index__EVAL_38;
  wire  axi4index__EVAL_39;
  wire [30:0] axi4index__EVAL_40;
  wire  axi4index__EVAL_41;
  wire  axi4index__EVAL_42;
  wire [3:0] axi4index__EVAL_43;
  wire [10:0] axi4index__EVAL_44;
  wire [2:0] axi4index__EVAL_45;
  wire [3:0] axi4index__EVAL_46;
  wire [3:0] axi4index__EVAL_47;
  wire  axi4index__EVAL_48;
  wire [1:0] axi4index__EVAL_49;
  wire [1:0] axi4index__EVAL_50;
  wire [2:0] axi4index__EVAL_51;
  wire [7:0] axi4index__EVAL_52;
  wire [2:0] axi4index__EVAL_53;
  wire [1:0] axi4index__EVAL_54;
  wire [30:0] axi4index__EVAL_55;
  wire [1:0] axi4index__EVAL_56;
  wire [2:0] axi4index__EVAL_57;
  wire [1:0] axi4index__EVAL_58;
  wire [3:0] axi4index__EVAL_59;
  wire  axi4index__EVAL_60;
  wire [10:0] axi4index__EVAL_61;
  wire [2:0] axi4index__EVAL_62;
  wire [3:0] axi4index__EVAL_63;
  wire [30:0] axi4index__EVAL_64;
  wire  axi4index__EVAL_65;
  wire  axi4index__EVAL_66;
  wire [2:0] axi4index__EVAL_67;
  wire  axi4index__EVAL_68;
  wire [2:0] axi4index__EVAL_69;
  wire  axi4index__EVAL_70;
  wire [1:0] axi4index__EVAL_71;
  wire  axi4index__EVAL_72;
  wire [7:0] axi4index__EVAL_73;
  wire [2:0] axi4index__EVAL_74;
  wire  axi4index__EVAL_75;
  wire [10:0] axi4index__EVAL_76;
  wire  axi4index__EVAL_77;
  wire  axi4index__EVAL_78;
  wire [2:0] axi4index__EVAL_79;
  wire [31:0] axi4index__EVAL_80;
  wire [3:0] axi4deint__EVAL;
  wire [10:0] axi4deint__EVAL_0;
  wire [31:0] axi4deint__EVAL_1;
  wire  axi4deint__EVAL_2;
  wire  axi4deint__EVAL_3;
  wire [7:0] axi4deint__EVAL_4;
  wire [1:0] axi4deint__EVAL_5;
  wire  axi4deint__EVAL_6;
  wire [2:0] axi4deint__EVAL_7;
  wire  axi4deint__EVAL_8;
  wire [2:0] axi4deint__EVAL_9;
  wire [7:0] axi4deint__EVAL_10;
  wire [3:0] axi4deint__EVAL_11;
  wire  axi4deint__EVAL_12;
  wire [3:0] axi4deint__EVAL_13;
  wire [3:0] axi4deint__EVAL_14;
  wire  axi4deint__EVAL_15;
  wire  axi4deint__EVAL_16;
  wire [3:0] axi4deint__EVAL_17;
  wire [3:0] axi4deint__EVAL_18;
  wire  axi4deint__EVAL_19;
  wire  axi4deint__EVAL_20;
  wire  axi4deint__EVAL_21;
  wire [30:0] axi4deint__EVAL_22;
  wire  axi4deint__EVAL_23;
  wire [10:0] axi4deint__EVAL_24;
  wire  axi4deint__EVAL_25;
  wire  axi4deint__EVAL_26;
  wire  axi4deint__EVAL_27;
  wire [10:0] axi4deint__EVAL_28;
  wire  axi4deint__EVAL_29;
  wire [31:0] axi4deint__EVAL_30;
  wire [31:0] axi4deint__EVAL_31;
  wire [10:0] axi4deint__EVAL_32;
  wire  axi4deint__EVAL_33;
  wire  axi4deint__EVAL_34;
  wire [30:0] axi4deint__EVAL_35;
  wire [3:0] axi4deint__EVAL_36;
  wire  axi4deint__EVAL_37;
  wire  axi4deint__EVAL_38;
  wire [1:0] axi4deint__EVAL_39;
  wire  axi4deint__EVAL_40;
  wire [3:0] axi4deint__EVAL_41;
  wire [3:0] axi4deint__EVAL_42;
  wire [10:0] axi4deint__EVAL_43;
  wire  axi4deint__EVAL_44;
  wire  axi4deint__EVAL_45;
  wire [3:0] axi4deint__EVAL_46;
  wire [1:0] axi4deint__EVAL_47;
  wire  axi4deint__EVAL_48;
  wire [1:0] axi4deint__EVAL_49;
  wire [1:0] axi4deint__EVAL_50;
  wire [3:0] axi4deint__EVAL_51;
  wire [30:0] axi4deint__EVAL_52;
  wire  axi4deint__EVAL_53;
  wire [3:0] axi4deint__EVAL_54;
  wire [31:0] axi4deint__EVAL_55;
  wire [7:0] axi4deint__EVAL_56;
  wire [10:0] axi4deint__EVAL_57;
  wire [3:0] axi4deint__EVAL_58;
  wire [3:0] axi4deint__EVAL_59;
  wire [2:0] axi4deint__EVAL_60;
  wire [7:0] axi4deint__EVAL_61;
  wire [2:0] axi4deint__EVAL_62;
  wire [3:0] axi4deint__EVAL_63;
  wire [2:0] axi4deint__EVAL_64;
  wire  axi4deint__EVAL_65;
  wire  axi4deint__EVAL_66;
  wire [3:0] axi4deint__EVAL_67;
  wire [2:0] axi4deint__EVAL_68;
  wire [1:0] axi4deint__EVAL_69;
  wire [3:0] axi4deint__EVAL_70;
  wire [2:0] axi4deint__EVAL_71;
  wire [1:0] axi4deint__EVAL_72;
  wire [10:0] axi4deint__EVAL_73;
  wire [30:0] axi4deint__EVAL_74;
  wire  axi4deint__EVAL_75;
  wire  axi4deint__EVAL_76;
  wire  axi4deint__EVAL_77;
  wire [2:0] axi4deint__EVAL_78;
  wire [3:0] axi4deint__EVAL_79;
  wire [1:0] axi4deint__EVAL_80;
  wire  axi4deint__EVAL_81;
  wire [10:0] axi4deint__EVAL_82;
  wire  axi4yank__EVAL;
  wire [3:0] axi4yank__EVAL_0;
  wire [7:0] axi4yank__EVAL_1;
  wire  axi4yank__EVAL_2;
  wire [2:0] axi4yank__EVAL_3;
  wire  axi4yank__EVAL_4;
  wire [3:0] axi4yank__EVAL_5;
  wire  axi4yank__EVAL_6;
  wire  axi4yank__EVAL_7;
  wire [1:0] axi4yank__EVAL_8;
  wire  axi4yank__EVAL_9;
  wire [2:0] axi4yank__EVAL_10;
  wire [1:0] axi4yank__EVAL_11;
  wire  axi4yank__EVAL_12;
  wire [1:0] axi4yank__EVAL_13;
  wire [3:0] axi4yank__EVAL_14;
  wire [7:0] axi4yank__EVAL_15;
  wire [3:0] axi4yank__EVAL_16;
  wire  axi4yank__EVAL_17;
  wire [3:0] axi4yank__EVAL_18;
  wire  axi4yank__EVAL_19;
  wire  axi4yank__EVAL_20;
  wire [3:0] axi4yank__EVAL_21;
  wire [31:0] axi4yank__EVAL_22;
  wire [1:0] axi4yank__EVAL_23;
  wire  axi4yank__EVAL_24;
  wire  axi4yank__EVAL_25;
  wire  axi4yank__EVAL_26;
  wire [2:0] axi4yank__EVAL_27;
  wire  axi4yank__EVAL_28;
  wire [3:0] axi4yank__EVAL_29;
  wire  axi4yank__EVAL_30;
  wire [2:0] axi4yank__EVAL_31;
  wire  axi4yank__EVAL_32;
  wire [30:0] axi4yank__EVAL_33;
  wire  axi4yank__EVAL_34;
  wire [3:0] axi4yank__EVAL_35;
  wire  axi4yank__EVAL_36;
  wire [3:0] axi4yank__EVAL_37;
  wire [3:0] axi4yank__EVAL_38;
  wire [30:0] axi4yank__EVAL_39;
  wire [2:0] axi4yank__EVAL_40;
  wire [2:0] axi4yank__EVAL_41;
  wire [30:0] axi4yank__EVAL_42;
  wire  axi4yank__EVAL_43;
  wire [1:0] axi4yank__EVAL_44;
  wire [1:0] axi4yank__EVAL_45;
  wire  axi4yank__EVAL_46;
  wire [7:0] axi4yank__EVAL_47;
  wire  axi4yank__EVAL_48;
  wire [1:0] axi4yank__EVAL_49;
  wire [3:0] axi4yank__EVAL_50;
  wire [10:0] axi4yank__EVAL_51;
  wire [3:0] axi4yank__EVAL_52;
  wire [31:0] axi4yank__EVAL_53;
  wire  axi4yank__EVAL_54;
  wire [10:0] axi4yank__EVAL_55;
  wire  axi4yank__EVAL_56;
  wire [7:0] axi4yank__EVAL_57;
  wire  axi4yank__EVAL_58;
  wire  axi4yank__EVAL_59;
  wire [10:0] axi4yank__EVAL_60;
  wire [30:0] axi4yank__EVAL_61;
  wire  axi4yank__EVAL_62;
  wire  axi4yank__EVAL_63;
  wire [31:0] axi4yank__EVAL_64;
  wire  axi4yank__EVAL_65;
  wire [31:0] axi4yank__EVAL_66;
  wire  axi4yank__EVAL_67;
  wire [2:0] axi4yank__EVAL_68;
  wire [3:0] axi4yank__EVAL_69;
  wire [3:0] axi4yank__EVAL_70;
  wire [3:0] axi4yank__EVAL_71;
  wire [3:0] axi4yank__EVAL_72;
  wire [2:0] axi4yank__EVAL_73;
  wire [3:0] axi4yank__EVAL_74;
  wire [3:0] axi4yank__EVAL_75;
  wire  axi4yank__EVAL_76;
  wire [10:0] axi4yank__EVAL_77;
  wire [1:0] axi4yank__EVAL_78;
  wire  widget__EVAL;
  wire  widget__EVAL_0;
  wire [2:0] widget__EVAL_1;
  wire  widget__EVAL_2;
  wire  widget__EVAL_3;
  wire [3:0] widget__EVAL_4;
  wire [63:0] widget__EVAL_5;
  wire [2:0] widget__EVAL_6;
  wire  widget__EVAL_7;
  wire [6:0] widget__EVAL_8;
  wire [7:0] widget__EVAL_9;
  wire [6:0] widget__EVAL_10;
  wire [31:0] widget__EVAL_11;
  wire [6:0] widget__EVAL_12;
  wire [30:0] widget__EVAL_13;
  wire  widget__EVAL_14;
  wire [2:0] widget__EVAL_15;
  wire  widget__EVAL_16;
  wire  widget__EVAL_17;
  wire  widget__EVAL_18;
  wire  widget__EVAL_19;
  wire  widget__EVAL_20;
  wire  widget__EVAL_21;
  wire [2:0] widget__EVAL_22;
  wire [30:0] widget__EVAL_23;
  wire [6:0] widget__EVAL_24;
  wire  widget__EVAL_25;
  wire  widget__EVAL_26;
  wire  widget__EVAL_27;
  wire [2:0] widget__EVAL_28;
  wire [2:0] widget__EVAL_29;
  wire [63:0] widget__EVAL_30;
  wire [2:0] widget__EVAL_31;
  wire [2:0] widget__EVAL_32;
  wire [31:0] widget__EVAL_33;
  wire [2:0] widget__EVAL_34;
  wire  widget__EVAL_35;
  wire [2:0] widget__EVAL_36;
  wire  tl2axi4__EVAL;
  wire [2:0] tl2axi4__EVAL_0;
  wire  tl2axi4__EVAL_1;
  wire  tl2axi4__EVAL_2;
  wire [7:0] tl2axi4__EVAL_3;
  wire [1:0] tl2axi4__EVAL_4;
  wire [1:0] tl2axi4__EVAL_5;
  wire [3:0] tl2axi4__EVAL_6;
  wire [2:0] tl2axi4__EVAL_7;
  wire  tl2axi4__EVAL_8;
  wire  tl2axi4__EVAL_9;
  wire [2:0] tl2axi4__EVAL_10;
  wire [3:0] tl2axi4__EVAL_11;
  wire [6:0] tl2axi4__EVAL_12;
  wire  tl2axi4__EVAL_13;
  wire [2:0] tl2axi4__EVAL_14;
  wire  tl2axi4__EVAL_15;
  wire [1:0] tl2axi4__EVAL_16;
  wire [3:0] tl2axi4__EVAL_17;
  wire  tl2axi4__EVAL_18;
  wire  tl2axi4__EVAL_19;
  wire [3:0] tl2axi4__EVAL_20;
  wire [30:0] tl2axi4__EVAL_21;
  wire [10:0] tl2axi4__EVAL_22;
  wire [2:0] tl2axi4__EVAL_23;
  wire  tl2axi4__EVAL_24;
  wire  tl2axi4__EVAL_25;
  wire [31:0] tl2axi4__EVAL_26;
  wire  tl2axi4__EVAL_27;
  wire  tl2axi4__EVAL_28;
  wire [10:0] tl2axi4__EVAL_29;
  wire [7:0] tl2axi4__EVAL_30;
  wire  tl2axi4__EVAL_31;
  wire [31:0] tl2axi4__EVAL_32;
  wire [2:0] tl2axi4__EVAL_33;
  wire  tl2axi4__EVAL_34;
  wire [31:0] tl2axi4__EVAL_35;
  wire [2:0] tl2axi4__EVAL_36;
  wire [2:0] tl2axi4__EVAL_37;
  wire [31:0] tl2axi4__EVAL_38;
  wire [2:0] tl2axi4__EVAL_39;
  wire  tl2axi4__EVAL_40;
  wire [6:0] tl2axi4__EVAL_41;
  wire [3:0] tl2axi4__EVAL_42;
  wire [30:0] tl2axi4__EVAL_43;
  wire [3:0] tl2axi4__EVAL_44;
  wire [2:0] tl2axi4__EVAL_45;
  wire [2:0] tl2axi4__EVAL_46;
  wire  tl2axi4__EVAL_47;
  wire  tl2axi4__EVAL_48;
  wire  tl2axi4__EVAL_49;
  wire  tl2axi4__EVAL_50;
  wire [10:0] tl2axi4__EVAL_51;
  wire [1:0] tl2axi4__EVAL_52;
  wire  tl2axi4__EVAL_53;
  wire  tl2axi4__EVAL_54;
  wire [30:0] tl2axi4__EVAL_55;
  wire [10:0] tl2axi4__EVAL_56;
  wire [2:0] tl2axi4__EVAL_57;
  wire [2:0] tl2axi4__EVAL_58;
  wire  tl2axi4__EVAL_59;
  wire  buffer__EVAL;
  wire  buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire [2:0] buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [2:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [63:0] buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire [63:0] buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire [2:0] buffer__EVAL_13;
  wire [2:0] buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire [30:0] buffer__EVAL_17;
  wire [6:0] buffer__EVAL_18;
  wire [63:0] buffer__EVAL_19;
  wire [2:0] buffer__EVAL_20;
  wire [2:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire [6:0] buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire [2:0] buffer__EVAL_26;
  wire [2:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire [7:0] buffer__EVAL_29;
  wire [6:0] buffer__EVAL_30;
  wire [6:0] buffer__EVAL_31;
  wire [63:0] buffer__EVAL_32;
  wire [2:0] buffer__EVAL_33;
  wire [30:0] buffer__EVAL_34;
  wire [2:0] buffer__EVAL_35;
  wire [7:0] buffer__EVAL_36;
  wire [31:0] axi4buf__EVAL;
  wire [3:0] axi4buf__EVAL_0;
  wire [3:0] axi4buf__EVAL_1;
  wire [1:0] axi4buf__EVAL_2;
  wire [1:0] axi4buf__EVAL_3;
  wire  axi4buf__EVAL_4;
  wire [3:0] axi4buf__EVAL_5;
  wire [30:0] axi4buf__EVAL_6;
  wire [1:0] axi4buf__EVAL_7;
  wire  axi4buf__EVAL_8;
  wire [3:0] axi4buf__EVAL_9;
  wire [3:0] axi4buf__EVAL_10;
  wire  axi4buf__EVAL_11;
  wire  axi4buf__EVAL_12;
  wire  axi4buf__EVAL_13;
  wire  axi4buf__EVAL_14;
  wire [30:0] axi4buf__EVAL_15;
  wire [3:0] axi4buf__EVAL_16;
  wire  axi4buf__EVAL_17;
  wire  axi4buf__EVAL_18;
  wire [7:0] axi4buf__EVAL_19;
  wire [3:0] axi4buf__EVAL_20;
  wire [3:0] axi4buf__EVAL_21;
  wire  axi4buf__EVAL_22;
  wire [31:0] axi4buf__EVAL_23;
  wire [3:0] axi4buf__EVAL_24;
  wire [3:0] axi4buf__EVAL_25;
  wire [1:0] axi4buf__EVAL_26;
  wire [2:0] axi4buf__EVAL_27;
  wire [31:0] axi4buf__EVAL_28;
  wire  axi4buf__EVAL_29;
  wire  axi4buf__EVAL_30;
  wire  axi4buf__EVAL_31;
  wire [7:0] axi4buf__EVAL_32;
  wire [3:0] axi4buf__EVAL_33;
  wire [3:0] axi4buf__EVAL_34;
  wire [3:0] axi4buf__EVAL_35;
  wire [2:0] axi4buf__EVAL_36;
  wire [7:0] axi4buf__EVAL_37;
  wire  axi4buf__EVAL_38;
  wire  axi4buf__EVAL_39;
  wire [2:0] axi4buf__EVAL_40;
  wire  axi4buf__EVAL_41;
  wire [3:0] axi4buf__EVAL_42;
  wire  axi4buf__EVAL_43;
  wire [2:0] axi4buf__EVAL_44;
  wire  axi4buf__EVAL_45;
  wire  axi4buf__EVAL_46;
  wire [3:0] axi4buf__EVAL_47;
  wire  axi4buf__EVAL_48;
  wire [3:0] axi4buf__EVAL_49;
  wire [2:0] axi4buf__EVAL_50;
  wire [1:0] axi4buf__EVAL_51;
  wire [7:0] axi4buf__EVAL_52;
  wire [30:0] axi4buf__EVAL_53;
  wire [2:0] axi4buf__EVAL_54;
  wire  axi4buf__EVAL_55;
  wire  axi4buf__EVAL_56;
  wire  axi4buf__EVAL_57;
  wire  axi4buf__EVAL_58;
  wire  axi4buf__EVAL_59;
  wire [1:0] axi4buf__EVAL_60;
  wire  axi4buf__EVAL_61;
  wire [31:0] axi4buf__EVAL_62;
  wire  axi4buf__EVAL_63;
  wire  axi4buf__EVAL_64;
  wire [3:0] axi4buf__EVAL_65;
  wire  axi4buf__EVAL_66;
  wire [1:0] axi4buf__EVAL_67;
  wire  axi4buf__EVAL_68;
  wire [30:0] axi4buf__EVAL_69;
  wire [2:0] axi4buf__EVAL_70;
  wire  axi4buf__EVAL_71;
  wire [1:0] axi4buf__EVAL_72;
  wire [3:0] axi4buf__EVAL_73;
  wire [2:0] axi4buf__EVAL_74;
  SiFive__EVAL_29 axi4index (
    ._EVAL(axi4index__EVAL),
    ._EVAL_0(axi4index__EVAL_0),
    ._EVAL_1(axi4index__EVAL_1),
    ._EVAL_2(axi4index__EVAL_2),
    ._EVAL_3(axi4index__EVAL_3),
    ._EVAL_4(axi4index__EVAL_4),
    ._EVAL_5(axi4index__EVAL_5),
    ._EVAL_6(axi4index__EVAL_6),
    ._EVAL_7(axi4index__EVAL_7),
    ._EVAL_8(axi4index__EVAL_8),
    ._EVAL_9(axi4index__EVAL_9),
    ._EVAL_10(axi4index__EVAL_10),
    ._EVAL_11(axi4index__EVAL_11),
    ._EVAL_12(axi4index__EVAL_12),
    ._EVAL_13(axi4index__EVAL_13),
    ._EVAL_14(axi4index__EVAL_14),
    ._EVAL_15(axi4index__EVAL_15),
    ._EVAL_16(axi4index__EVAL_16),
    ._EVAL_17(axi4index__EVAL_17),
    ._EVAL_18(axi4index__EVAL_18),
    ._EVAL_19(axi4index__EVAL_19),
    ._EVAL_20(axi4index__EVAL_20),
    ._EVAL_21(axi4index__EVAL_21),
    ._EVAL_22(axi4index__EVAL_22),
    ._EVAL_23(axi4index__EVAL_23),
    ._EVAL_24(axi4index__EVAL_24),
    ._EVAL_25(axi4index__EVAL_25),
    ._EVAL_26(axi4index__EVAL_26),
    ._EVAL_27(axi4index__EVAL_27),
    ._EVAL_28(axi4index__EVAL_28),
    ._EVAL_29(axi4index__EVAL_29),
    ._EVAL_30(axi4index__EVAL_30),
    ._EVAL_31(axi4index__EVAL_31),
    ._EVAL_32(axi4index__EVAL_32),
    ._EVAL_33(axi4index__EVAL_33),
    ._EVAL_34(axi4index__EVAL_34),
    ._EVAL_35(axi4index__EVAL_35),
    ._EVAL_36(axi4index__EVAL_36),
    ._EVAL_37(axi4index__EVAL_37),
    ._EVAL_38(axi4index__EVAL_38),
    ._EVAL_39(axi4index__EVAL_39),
    ._EVAL_40(axi4index__EVAL_40),
    ._EVAL_41(axi4index__EVAL_41),
    ._EVAL_42(axi4index__EVAL_42),
    ._EVAL_43(axi4index__EVAL_43),
    ._EVAL_44(axi4index__EVAL_44),
    ._EVAL_45(axi4index__EVAL_45),
    ._EVAL_46(axi4index__EVAL_46),
    ._EVAL_47(axi4index__EVAL_47),
    ._EVAL_48(axi4index__EVAL_48),
    ._EVAL_49(axi4index__EVAL_49),
    ._EVAL_50(axi4index__EVAL_50),
    ._EVAL_51(axi4index__EVAL_51),
    ._EVAL_52(axi4index__EVAL_52),
    ._EVAL_53(axi4index__EVAL_53),
    ._EVAL_54(axi4index__EVAL_54),
    ._EVAL_55(axi4index__EVAL_55),
    ._EVAL_56(axi4index__EVAL_56),
    ._EVAL_57(axi4index__EVAL_57),
    ._EVAL_58(axi4index__EVAL_58),
    ._EVAL_59(axi4index__EVAL_59),
    ._EVAL_60(axi4index__EVAL_60),
    ._EVAL_61(axi4index__EVAL_61),
    ._EVAL_62(axi4index__EVAL_62),
    ._EVAL_63(axi4index__EVAL_63),
    ._EVAL_64(axi4index__EVAL_64),
    ._EVAL_65(axi4index__EVAL_65),
    ._EVAL_66(axi4index__EVAL_66),
    ._EVAL_67(axi4index__EVAL_67),
    ._EVAL_68(axi4index__EVAL_68),
    ._EVAL_69(axi4index__EVAL_69),
    ._EVAL_70(axi4index__EVAL_70),
    ._EVAL_71(axi4index__EVAL_71),
    ._EVAL_72(axi4index__EVAL_72),
    ._EVAL_73(axi4index__EVAL_73),
    ._EVAL_74(axi4index__EVAL_74),
    ._EVAL_75(axi4index__EVAL_75),
    ._EVAL_76(axi4index__EVAL_76),
    ._EVAL_77(axi4index__EVAL_77),
    ._EVAL_78(axi4index__EVAL_78),
    ._EVAL_79(axi4index__EVAL_79),
    ._EVAL_80(axi4index__EVAL_80)
  );
  SiFive__EVAL_20 axi4deint (
    ._EVAL(axi4deint__EVAL),
    ._EVAL_0(axi4deint__EVAL_0),
    ._EVAL_1(axi4deint__EVAL_1),
    ._EVAL_2(axi4deint__EVAL_2),
    ._EVAL_3(axi4deint__EVAL_3),
    ._EVAL_4(axi4deint__EVAL_4),
    ._EVAL_5(axi4deint__EVAL_5),
    ._EVAL_6(axi4deint__EVAL_6),
    ._EVAL_7(axi4deint__EVAL_7),
    ._EVAL_8(axi4deint__EVAL_8),
    ._EVAL_9(axi4deint__EVAL_9),
    ._EVAL_10(axi4deint__EVAL_10),
    ._EVAL_11(axi4deint__EVAL_11),
    ._EVAL_12(axi4deint__EVAL_12),
    ._EVAL_13(axi4deint__EVAL_13),
    ._EVAL_14(axi4deint__EVAL_14),
    ._EVAL_15(axi4deint__EVAL_15),
    ._EVAL_16(axi4deint__EVAL_16),
    ._EVAL_17(axi4deint__EVAL_17),
    ._EVAL_18(axi4deint__EVAL_18),
    ._EVAL_19(axi4deint__EVAL_19),
    ._EVAL_20(axi4deint__EVAL_20),
    ._EVAL_21(axi4deint__EVAL_21),
    ._EVAL_22(axi4deint__EVAL_22),
    ._EVAL_23(axi4deint__EVAL_23),
    ._EVAL_24(axi4deint__EVAL_24),
    ._EVAL_25(axi4deint__EVAL_25),
    ._EVAL_26(axi4deint__EVAL_26),
    ._EVAL_27(axi4deint__EVAL_27),
    ._EVAL_28(axi4deint__EVAL_28),
    ._EVAL_29(axi4deint__EVAL_29),
    ._EVAL_30(axi4deint__EVAL_30),
    ._EVAL_31(axi4deint__EVAL_31),
    ._EVAL_32(axi4deint__EVAL_32),
    ._EVAL_33(axi4deint__EVAL_33),
    ._EVAL_34(axi4deint__EVAL_34),
    ._EVAL_35(axi4deint__EVAL_35),
    ._EVAL_36(axi4deint__EVAL_36),
    ._EVAL_37(axi4deint__EVAL_37),
    ._EVAL_38(axi4deint__EVAL_38),
    ._EVAL_39(axi4deint__EVAL_39),
    ._EVAL_40(axi4deint__EVAL_40),
    ._EVAL_41(axi4deint__EVAL_41),
    ._EVAL_42(axi4deint__EVAL_42),
    ._EVAL_43(axi4deint__EVAL_43),
    ._EVAL_44(axi4deint__EVAL_44),
    ._EVAL_45(axi4deint__EVAL_45),
    ._EVAL_46(axi4deint__EVAL_46),
    ._EVAL_47(axi4deint__EVAL_47),
    ._EVAL_48(axi4deint__EVAL_48),
    ._EVAL_49(axi4deint__EVAL_49),
    ._EVAL_50(axi4deint__EVAL_50),
    ._EVAL_51(axi4deint__EVAL_51),
    ._EVAL_52(axi4deint__EVAL_52),
    ._EVAL_53(axi4deint__EVAL_53),
    ._EVAL_54(axi4deint__EVAL_54),
    ._EVAL_55(axi4deint__EVAL_55),
    ._EVAL_56(axi4deint__EVAL_56),
    ._EVAL_57(axi4deint__EVAL_57),
    ._EVAL_58(axi4deint__EVAL_58),
    ._EVAL_59(axi4deint__EVAL_59),
    ._EVAL_60(axi4deint__EVAL_60),
    ._EVAL_61(axi4deint__EVAL_61),
    ._EVAL_62(axi4deint__EVAL_62),
    ._EVAL_63(axi4deint__EVAL_63),
    ._EVAL_64(axi4deint__EVAL_64),
    ._EVAL_65(axi4deint__EVAL_65),
    ._EVAL_66(axi4deint__EVAL_66),
    ._EVAL_67(axi4deint__EVAL_67),
    ._EVAL_68(axi4deint__EVAL_68),
    ._EVAL_69(axi4deint__EVAL_69),
    ._EVAL_70(axi4deint__EVAL_70),
    ._EVAL_71(axi4deint__EVAL_71),
    ._EVAL_72(axi4deint__EVAL_72),
    ._EVAL_73(axi4deint__EVAL_73),
    ._EVAL_74(axi4deint__EVAL_74),
    ._EVAL_75(axi4deint__EVAL_75),
    ._EVAL_76(axi4deint__EVAL_76),
    ._EVAL_77(axi4deint__EVAL_77),
    ._EVAL_78(axi4deint__EVAL_78),
    ._EVAL_79(axi4deint__EVAL_79),
    ._EVAL_80(axi4deint__EVAL_80),
    ._EVAL_81(axi4deint__EVAL_81),
    ._EVAL_82(axi4deint__EVAL_82)
  );
  SiFive__EVAL_28 axi4yank (
    ._EVAL(axi4yank__EVAL),
    ._EVAL_0(axi4yank__EVAL_0),
    ._EVAL_1(axi4yank__EVAL_1),
    ._EVAL_2(axi4yank__EVAL_2),
    ._EVAL_3(axi4yank__EVAL_3),
    ._EVAL_4(axi4yank__EVAL_4),
    ._EVAL_5(axi4yank__EVAL_5),
    ._EVAL_6(axi4yank__EVAL_6),
    ._EVAL_7(axi4yank__EVAL_7),
    ._EVAL_8(axi4yank__EVAL_8),
    ._EVAL_9(axi4yank__EVAL_9),
    ._EVAL_10(axi4yank__EVAL_10),
    ._EVAL_11(axi4yank__EVAL_11),
    ._EVAL_12(axi4yank__EVAL_12),
    ._EVAL_13(axi4yank__EVAL_13),
    ._EVAL_14(axi4yank__EVAL_14),
    ._EVAL_15(axi4yank__EVAL_15),
    ._EVAL_16(axi4yank__EVAL_16),
    ._EVAL_17(axi4yank__EVAL_17),
    ._EVAL_18(axi4yank__EVAL_18),
    ._EVAL_19(axi4yank__EVAL_19),
    ._EVAL_20(axi4yank__EVAL_20),
    ._EVAL_21(axi4yank__EVAL_21),
    ._EVAL_22(axi4yank__EVAL_22),
    ._EVAL_23(axi4yank__EVAL_23),
    ._EVAL_24(axi4yank__EVAL_24),
    ._EVAL_25(axi4yank__EVAL_25),
    ._EVAL_26(axi4yank__EVAL_26),
    ._EVAL_27(axi4yank__EVAL_27),
    ._EVAL_28(axi4yank__EVAL_28),
    ._EVAL_29(axi4yank__EVAL_29),
    ._EVAL_30(axi4yank__EVAL_30),
    ._EVAL_31(axi4yank__EVAL_31),
    ._EVAL_32(axi4yank__EVAL_32),
    ._EVAL_33(axi4yank__EVAL_33),
    ._EVAL_34(axi4yank__EVAL_34),
    ._EVAL_35(axi4yank__EVAL_35),
    ._EVAL_36(axi4yank__EVAL_36),
    ._EVAL_37(axi4yank__EVAL_37),
    ._EVAL_38(axi4yank__EVAL_38),
    ._EVAL_39(axi4yank__EVAL_39),
    ._EVAL_40(axi4yank__EVAL_40),
    ._EVAL_41(axi4yank__EVAL_41),
    ._EVAL_42(axi4yank__EVAL_42),
    ._EVAL_43(axi4yank__EVAL_43),
    ._EVAL_44(axi4yank__EVAL_44),
    ._EVAL_45(axi4yank__EVAL_45),
    ._EVAL_46(axi4yank__EVAL_46),
    ._EVAL_47(axi4yank__EVAL_47),
    ._EVAL_48(axi4yank__EVAL_48),
    ._EVAL_49(axi4yank__EVAL_49),
    ._EVAL_50(axi4yank__EVAL_50),
    ._EVAL_51(axi4yank__EVAL_51),
    ._EVAL_52(axi4yank__EVAL_52),
    ._EVAL_53(axi4yank__EVAL_53),
    ._EVAL_54(axi4yank__EVAL_54),
    ._EVAL_55(axi4yank__EVAL_55),
    ._EVAL_56(axi4yank__EVAL_56),
    ._EVAL_57(axi4yank__EVAL_57),
    ._EVAL_58(axi4yank__EVAL_58),
    ._EVAL_59(axi4yank__EVAL_59),
    ._EVAL_60(axi4yank__EVAL_60),
    ._EVAL_61(axi4yank__EVAL_61),
    ._EVAL_62(axi4yank__EVAL_62),
    ._EVAL_63(axi4yank__EVAL_63),
    ._EVAL_64(axi4yank__EVAL_64),
    ._EVAL_65(axi4yank__EVAL_65),
    ._EVAL_66(axi4yank__EVAL_66),
    ._EVAL_67(axi4yank__EVAL_67),
    ._EVAL_68(axi4yank__EVAL_68),
    ._EVAL_69(axi4yank__EVAL_69),
    ._EVAL_70(axi4yank__EVAL_70),
    ._EVAL_71(axi4yank__EVAL_71),
    ._EVAL_72(axi4yank__EVAL_72),
    ._EVAL_73(axi4yank__EVAL_73),
    ._EVAL_74(axi4yank__EVAL_74),
    ._EVAL_75(axi4yank__EVAL_75),
    ._EVAL_76(axi4yank__EVAL_76),
    ._EVAL_77(axi4yank__EVAL_77),
    ._EVAL_78(axi4yank__EVAL_78)
  );
  SiFive__EVAL_36 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36)
  );
  SiFive__EVAL_33 tl2axi4 (
    ._EVAL(tl2axi4__EVAL),
    ._EVAL_0(tl2axi4__EVAL_0),
    ._EVAL_1(tl2axi4__EVAL_1),
    ._EVAL_2(tl2axi4__EVAL_2),
    ._EVAL_3(tl2axi4__EVAL_3),
    ._EVAL_4(tl2axi4__EVAL_4),
    ._EVAL_5(tl2axi4__EVAL_5),
    ._EVAL_6(tl2axi4__EVAL_6),
    ._EVAL_7(tl2axi4__EVAL_7),
    ._EVAL_8(tl2axi4__EVAL_8),
    ._EVAL_9(tl2axi4__EVAL_9),
    ._EVAL_10(tl2axi4__EVAL_10),
    ._EVAL_11(tl2axi4__EVAL_11),
    ._EVAL_12(tl2axi4__EVAL_12),
    ._EVAL_13(tl2axi4__EVAL_13),
    ._EVAL_14(tl2axi4__EVAL_14),
    ._EVAL_15(tl2axi4__EVAL_15),
    ._EVAL_16(tl2axi4__EVAL_16),
    ._EVAL_17(tl2axi4__EVAL_17),
    ._EVAL_18(tl2axi4__EVAL_18),
    ._EVAL_19(tl2axi4__EVAL_19),
    ._EVAL_20(tl2axi4__EVAL_20),
    ._EVAL_21(tl2axi4__EVAL_21),
    ._EVAL_22(tl2axi4__EVAL_22),
    ._EVAL_23(tl2axi4__EVAL_23),
    ._EVAL_24(tl2axi4__EVAL_24),
    ._EVAL_25(tl2axi4__EVAL_25),
    ._EVAL_26(tl2axi4__EVAL_26),
    ._EVAL_27(tl2axi4__EVAL_27),
    ._EVAL_28(tl2axi4__EVAL_28),
    ._EVAL_29(tl2axi4__EVAL_29),
    ._EVAL_30(tl2axi4__EVAL_30),
    ._EVAL_31(tl2axi4__EVAL_31),
    ._EVAL_32(tl2axi4__EVAL_32),
    ._EVAL_33(tl2axi4__EVAL_33),
    ._EVAL_34(tl2axi4__EVAL_34),
    ._EVAL_35(tl2axi4__EVAL_35),
    ._EVAL_36(tl2axi4__EVAL_36),
    ._EVAL_37(tl2axi4__EVAL_37),
    ._EVAL_38(tl2axi4__EVAL_38),
    ._EVAL_39(tl2axi4__EVAL_39),
    ._EVAL_40(tl2axi4__EVAL_40),
    ._EVAL_41(tl2axi4__EVAL_41),
    ._EVAL_42(tl2axi4__EVAL_42),
    ._EVAL_43(tl2axi4__EVAL_43),
    ._EVAL_44(tl2axi4__EVAL_44),
    ._EVAL_45(tl2axi4__EVAL_45),
    ._EVAL_46(tl2axi4__EVAL_46),
    ._EVAL_47(tl2axi4__EVAL_47),
    ._EVAL_48(tl2axi4__EVAL_48),
    ._EVAL_49(tl2axi4__EVAL_49),
    ._EVAL_50(tl2axi4__EVAL_50),
    ._EVAL_51(tl2axi4__EVAL_51),
    ._EVAL_52(tl2axi4__EVAL_52),
    ._EVAL_53(tl2axi4__EVAL_53),
    ._EVAL_54(tl2axi4__EVAL_54),
    ._EVAL_55(tl2axi4__EVAL_55),
    ._EVAL_56(tl2axi4__EVAL_56),
    ._EVAL_57(tl2axi4__EVAL_57),
    ._EVAL_58(tl2axi4__EVAL_58),
    ._EVAL_59(tl2axi4__EVAL_59)
  );
  SiFive__EVAL_38 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36)
  );
  SiFive__EVAL_24 axi4buf (
    ._EVAL(axi4buf__EVAL),
    ._EVAL_0(axi4buf__EVAL_0),
    ._EVAL_1(axi4buf__EVAL_1),
    ._EVAL_2(axi4buf__EVAL_2),
    ._EVAL_3(axi4buf__EVAL_3),
    ._EVAL_4(axi4buf__EVAL_4),
    ._EVAL_5(axi4buf__EVAL_5),
    ._EVAL_6(axi4buf__EVAL_6),
    ._EVAL_7(axi4buf__EVAL_7),
    ._EVAL_8(axi4buf__EVAL_8),
    ._EVAL_9(axi4buf__EVAL_9),
    ._EVAL_10(axi4buf__EVAL_10),
    ._EVAL_11(axi4buf__EVAL_11),
    ._EVAL_12(axi4buf__EVAL_12),
    ._EVAL_13(axi4buf__EVAL_13),
    ._EVAL_14(axi4buf__EVAL_14),
    ._EVAL_15(axi4buf__EVAL_15),
    ._EVAL_16(axi4buf__EVAL_16),
    ._EVAL_17(axi4buf__EVAL_17),
    ._EVAL_18(axi4buf__EVAL_18),
    ._EVAL_19(axi4buf__EVAL_19),
    ._EVAL_20(axi4buf__EVAL_20),
    ._EVAL_21(axi4buf__EVAL_21),
    ._EVAL_22(axi4buf__EVAL_22),
    ._EVAL_23(axi4buf__EVAL_23),
    ._EVAL_24(axi4buf__EVAL_24),
    ._EVAL_25(axi4buf__EVAL_25),
    ._EVAL_26(axi4buf__EVAL_26),
    ._EVAL_27(axi4buf__EVAL_27),
    ._EVAL_28(axi4buf__EVAL_28),
    ._EVAL_29(axi4buf__EVAL_29),
    ._EVAL_30(axi4buf__EVAL_30),
    ._EVAL_31(axi4buf__EVAL_31),
    ._EVAL_32(axi4buf__EVAL_32),
    ._EVAL_33(axi4buf__EVAL_33),
    ._EVAL_34(axi4buf__EVAL_34),
    ._EVAL_35(axi4buf__EVAL_35),
    ._EVAL_36(axi4buf__EVAL_36),
    ._EVAL_37(axi4buf__EVAL_37),
    ._EVAL_38(axi4buf__EVAL_38),
    ._EVAL_39(axi4buf__EVAL_39),
    ._EVAL_40(axi4buf__EVAL_40),
    ._EVAL_41(axi4buf__EVAL_41),
    ._EVAL_42(axi4buf__EVAL_42),
    ._EVAL_43(axi4buf__EVAL_43),
    ._EVAL_44(axi4buf__EVAL_44),
    ._EVAL_45(axi4buf__EVAL_45),
    ._EVAL_46(axi4buf__EVAL_46),
    ._EVAL_47(axi4buf__EVAL_47),
    ._EVAL_48(axi4buf__EVAL_48),
    ._EVAL_49(axi4buf__EVAL_49),
    ._EVAL_50(axi4buf__EVAL_50),
    ._EVAL_51(axi4buf__EVAL_51),
    ._EVAL_52(axi4buf__EVAL_52),
    ._EVAL_53(axi4buf__EVAL_53),
    ._EVAL_54(axi4buf__EVAL_54),
    ._EVAL_55(axi4buf__EVAL_55),
    ._EVAL_56(axi4buf__EVAL_56),
    ._EVAL_57(axi4buf__EVAL_57),
    ._EVAL_58(axi4buf__EVAL_58),
    ._EVAL_59(axi4buf__EVAL_59),
    ._EVAL_60(axi4buf__EVAL_60),
    ._EVAL_61(axi4buf__EVAL_61),
    ._EVAL_62(axi4buf__EVAL_62),
    ._EVAL_63(axi4buf__EVAL_63),
    ._EVAL_64(axi4buf__EVAL_64),
    ._EVAL_65(axi4buf__EVAL_65),
    ._EVAL_66(axi4buf__EVAL_66),
    ._EVAL_67(axi4buf__EVAL_67),
    ._EVAL_68(axi4buf__EVAL_68),
    ._EVAL_69(axi4buf__EVAL_69),
    ._EVAL_70(axi4buf__EVAL_70),
    ._EVAL_71(axi4buf__EVAL_71),
    ._EVAL_72(axi4buf__EVAL_72),
    ._EVAL_73(axi4buf__EVAL_73),
    ._EVAL_74(axi4buf__EVAL_74)
  );
  assign buffer__EVAL_7 = _EVAL_49;
  assign axi4index__EVAL_58 = tl2axi4__EVAL_5;
  assign tl2axi4__EVAL_9 = axi4index__EVAL_72;
  assign _EVAL_6 = axi4buf__EVAL_64;
  assign axi4buf__EVAL_54 = axi4yank__EVAL_68;
  assign axi4yank__EVAL_43 = axi4buf__EVAL_41;
  assign axi4index__EVAL_6 = axi4deint__EVAL_40;
  assign axi4buf__EVAL_57 = _EVAL_42;
  assign tl2axi4__EVAL_23 = axi4index__EVAL_57;
  assign buffer__EVAL_12 = _EVAL_37;
  assign axi4buf__EVAL_48 = _EVAL_4;
  assign buffer__EVAL_2 = widget__EVAL;
  assign _EVAL_9 = axi4buf__EVAL_36;
  assign widget__EVAL_10 = tl2axi4__EVAL_12;
  assign _EVAL_29 = axi4buf__EVAL_20;
  assign tl2axi4__EVAL_47 = axi4index__EVAL_65;
  assign axi4deint__EVAL_57 = axi4index__EVAL_2;
  assign axi4deint__EVAL_21 = axi4index__EVAL_11;
  assign axi4index__EVAL_34 = tl2axi4__EVAL_37;
  assign axi4index__EVAL_37 = tl2axi4__EVAL_26;
  assign axi4yank__EVAL_27 = axi4deint__EVAL_7;
  assign _EVAL_46 = axi4buf__EVAL_0;
  assign axi4deint__EVAL = axi4index__EVAL_7;
  assign buffer__EVAL_27 = widget__EVAL_36;
  assign axi4buf__EVAL_32 = axi4yank__EVAL_1;
  assign axi4buf__EVAL_65 = axi4yank__EVAL_52;
  assign axi4deint__EVAL_58 = axi4yank__EVAL_50;
  assign tl2axi4__EVAL_19 = widget__EVAL_20;
  assign axi4deint__EVAL_43 = axi4index__EVAL_16;
  assign axi4deint__EVAL_61 = axi4index__EVAL_73;
  assign axi4index__EVAL_44 = tl2axi4__EVAL_29;
  assign axi4deint__EVAL_42 = axi4index__EVAL_33;
  assign axi4yank__EVAL_31 = axi4deint__EVAL_78;
  assign axi4index__EVAL_60 = tl2axi4__EVAL_1;
  assign axi4index__EVAL_74 = tl2axi4__EVAL_57;
  assign axi4yank__EVAL_47 = axi4deint__EVAL_56;
  assign widget__EVAL_2 = tl2axi4__EVAL_25;
  assign axi4index__EVAL_42 = tl2axi4__EVAL_50;
  assign axi4index__EVAL_36 = tl2axi4__EVAL_17;
  assign tl2axi4__EVAL_7 = widget__EVAL_22;
  assign axi4index__EVAL_63 = tl2axi4__EVAL_42;
  assign _EVAL_22 = axi4buf__EVAL_56;
  assign _EVAL_38 = axi4buf__EVAL_72;
  assign axi4deint__EVAL_79 = axi4index__EVAL_20;
  assign tl2axi4__EVAL_15 = _EVAL_37;
  assign axi4index__EVAL_47 = tl2axi4__EVAL_6;
  assign tl2axi4__EVAL_59 = axi4index__EVAL_41;
  assign axi4index__EVAL_75 = tl2axi4__EVAL_40;
  assign axi4yank__EVAL_53 = axi4buf__EVAL_23;
  assign axi4index__EVAL_10 = tl2axi4__EVAL_49;
  assign axi4index__EVAL_22 = axi4deint__EVAL_8;
  assign axi4index__EVAL_51 = tl2axi4__EVAL_46;
  assign axi4buf__EVAL_9 = axi4yank__EVAL_72;
  assign axi4deint__EVAL_69 = axi4index__EVAL_18;
  assign axi4index__EVAL_35 = tl2axi4__EVAL_31;
  assign tl2axi4__EVAL_39 = widget__EVAL_6;
  assign axi4index__EVAL_15 = axi4deint__EVAL_41;
  assign _EVAL_34 = axi4buf__EVAL_37;
  assign widget__EVAL_26 = buffer__EVAL_15;
  assign _EVAL_54 = axi4buf__EVAL_52;
  assign axi4index__EVAL_5 = axi4deint__EVAL_66;
  assign tl2axi4__EVAL_58 = widget__EVAL_15;
  assign tl2axi4__EVAL_16 = axi4index__EVAL_49;
  assign tl2axi4__EVAL_48 = axi4index__EVAL_77;
  assign _EVAL_36 = buffer__EVAL_25;
  assign axi4yank__EVAL_37 = axi4deint__EVAL_59;
  assign axi4index__EVAL_25 = tl2axi4__EVAL_2;
  assign axi4yank__EVAL_35 = axi4buf__EVAL_34;
  assign axi4index__EVAL_4 = axi4deint__EVAL_0;
  assign widget__EVAL_13 = buffer__EVAL_34;
  assign axi4yank__EVAL_69 = axi4deint__EVAL_18;
  assign _EVAL_14 = axi4buf__EVAL_6;
  assign axi4yank__EVAL_8 = axi4deint__EVAL_50;
  assign axi4yank__EVAL_58 = axi4deint__EVAL_37;
  assign widget__EVAL_29 = buffer__EVAL_33;
  assign axi4yank__EVAL_63 = axi4deint__EVAL_2;
  assign axi4deint__EVAL_76 = _EVAL_37;
  assign buffer__EVAL_1 = _EVAL_25;
  assign axi4deint__EVAL_47 = axi4yank__EVAL_49;
  assign axi4buf__EVAL_59 = _EVAL_0;
  assign axi4yank__EVAL_61 = axi4deint__EVAL_35;
  assign axi4index__EVAL_1 = axi4deint__EVAL_55;
  assign axi4deint__EVAL_23 = axi4yank__EVAL_32;
  assign widget__EVAL_9 = buffer__EVAL_36;
  assign axi4buf__EVAL_14 = _EVAL_37;
  assign axi4yank__EVAL_65 = axi4deint__EVAL_20;
  assign buffer__EVAL_6 = _EVAL_5;
  assign tl2axi4__EVAL_32 = widget__EVAL_33;
  assign axi4deint__EVAL_81 = axi4yank__EVAL_67;
  assign buffer__EVAL_14 = _EVAL_3;
  assign axi4yank__EVAL_13 = axi4deint__EVAL_49;
  assign axi4index__EVAL_23 = tl2axi4__EVAL_33;
  assign axi4yank__EVAL_9 = axi4deint__EVAL_38;
  assign axi4buf__EVAL_33 = axi4yank__EVAL_75;
  assign axi4buf__EVAL_39 = axi4yank__EVAL_36;
  assign axi4yank__EVAL_29 = axi4buf__EVAL_49;
  assign widget__EVAL_21 = tl2axi4__EVAL_24;
  assign axi4deint__EVAL_51 = axi4index__EVAL_3;
  assign axi4deint__EVAL_31 = axi4yank__EVAL_66;
  assign widget__EVAL_0 = tl2axi4__EVAL_18;
  assign axi4index__EVAL_24 = axi4deint__EVAL_6;
  assign axi4buf__EVAL_51 = _EVAL_15;
  assign buffer__EVAL_16 = widget__EVAL_19;
  assign widget__EVAL_25 = tl2axi4__EVAL_8;
  assign axi4yank__EVAL_2 = axi4deint__EVAL_27;
  assign buffer__EVAL_10 = _EVAL_16;
  assign axi4buf__EVAL_28 = axi4yank__EVAL_22;
  assign axi4yank__EVAL_19 = axi4deint__EVAL_53;
  assign widget__EVAL_28 = tl2axi4__EVAL_0;
  assign axi4deint__EVAL_67 = axi4yank__EVAL_74;
  assign axi4yank__EVAL_41 = axi4deint__EVAL_60;
  assign axi4yank__EVAL_64 = axi4deint__EVAL_1;
  assign axi4yank__EVAL_51 = axi4deint__EVAL_28;
  assign axi4buf__EVAL_2 = axi4yank__EVAL_78;
  assign axi4yank__EVAL_46 = _EVAL_37;
  assign axi4deint__EVAL_74 = axi4index__EVAL_38;
  assign axi4buf__EVAL_1 = _EVAL_47;
  assign axi4index__EVAL_69 = tl2axi4__EVAL_45;
  assign axi4index__EVAL_14 = tl2axi4__EVAL_56;
  assign tl2axi4__EVAL_38 = axi4index__EVAL_80;
  assign _EVAL_30 = axi4buf__EVAL_31;
  assign axi4deint__EVAL_15 = axi4index__EVAL_0;
  assign _EVAL_7 = buffer__EVAL_23;
  assign axi4buf__EVAL_62 = _EVAL_11;
  assign buffer__EVAL_29 = _EVAL_48;
  assign widget__EVAL_16 = _EVAL_37;
  assign axi4buf__EVAL_43 = axi4yank__EVAL_4;
  assign axi4buf__EVAL_47 = axi4yank__EVAL_38;
  assign axi4deint__EVAL_62 = axi4index__EVAL_53;
  assign axi4yank__EVAL_40 = axi4deint__EVAL_64;
  assign buffer__EVAL_24 = widget__EVAL_12;
  assign widget__EVAL_18 = _EVAL_25;
  assign tl2axi4__EVAL_22 = axi4index__EVAL_76;
  assign axi4index__EVAL_21 = tl2axi4__EVAL_20;
  assign tl2axi4__EVAL_13 = widget__EVAL_3;
  assign buffer__EVAL_0 = widget__EVAL_17;
  assign tl2axi4__EVAL_34 = widget__EVAL_35;
  assign axi4yank__EVAL_14 = axi4deint__EVAL_46;
  assign axi4index__EVAL_40 = tl2axi4__EVAL_55;
  assign buffer__EVAL_5 = widget__EVAL_14;
  assign axi4deint__EVAL_17 = axi4index__EVAL_43;
  assign axi4index__EVAL_56 = tl2axi4__EVAL_52;
  assign axi4deint__EVAL_26 = axi4index__EVAL_39;
  assign axi4deint__EVAL_45 = axi4yank__EVAL_56;
  assign _EVAL_1 = axi4buf__EVAL_69;
  assign _EVAL_23 = axi4buf__EVAL_40;
  assign axi4buf__EVAL_17 = axi4yank__EVAL_20;
  assign axi4index__EVAL_17 = axi4deint__EVAL_32;
  assign buffer__EVAL_4 = _EVAL;
  assign axi4buf__EVAL_13 = axi4yank__EVAL_7;
  assign axi4buf__EVAL_16 = _EVAL_8;
  assign tl2axi4__EVAL_4 = axi4index__EVAL_54;
  assign axi4deint__EVAL_9 = axi4index__EVAL_67;
  assign axi4deint__EVAL_71 = axi4index__EVAL_79;
  assign axi4yank__EVAL_33 = axi4deint__EVAL_52;
  assign axi4index__EVAL_27 = tl2axi4__EVAL_3;
  assign buffer__EVAL_21 = _EVAL_51;
  assign axi4buf__EVAL_12 = _EVAL_25;
  assign axi4deint__EVAL_73 = axi4yank__EVAL_55;
  assign axi4deint__EVAL_77 = axi4yank__EVAL_54;
  assign buffer__EVAL_17 = _EVAL_45;
  assign tl2axi4__EVAL_27 = axi4index__EVAL_30;
  assign axi4yank__EVAL_24 = axi4buf__EVAL_68;
  assign axi4yank__EVAL_18 = axi4deint__EVAL_36;
  assign axi4index__EVAL_19 = tl2axi4__EVAL_28;
  assign axi4deint__EVAL_10 = axi4index__EVAL_52;
  assign widget__EVAL_34 = buffer__EVAL_13;
  assign axi4yank__EVAL_44 = axi4buf__EVAL_7;
  assign _EVAL_41 = axi4buf__EVAL_50;
  assign _EVAL_32 = axi4buf__EVAL_42;
  assign axi4deint__EVAL_25 = axi4index__EVAL_78;
  assign _EVAL_55 = axi4buf__EVAL_27;
  assign axi4yank__EVAL_34 = _EVAL_25;
  assign tl2axi4__EVAL = axi4index__EVAL_48;
  assign buffer__EVAL_26 = widget__EVAL_31;
  assign axi4buf__EVAL_19 = axi4yank__EVAL_57;
  assign axi4deint__EVAL_12 = axi4index__EVAL_31;
  assign axi4deint__EVAL_68 = axi4index__EVAL_29;
  assign _EVAL_27 = axi4buf__EVAL_66;
  assign axi4index__EVAL_71 = axi4deint__EVAL_72;
  assign _EVAL_44 = axi4buf__EVAL;
  assign widget__EVAL_1 = buffer__EVAL_3;
  assign _EVAL_18 = axi4buf__EVAL_71;
  assign axi4yank__EVAL_62 = axi4deint__EVAL_44;
  assign axi4yank__EVAL_30 = axi4buf__EVAL_29;
  assign _EVAL_20 = axi4buf__EVAL_24;
  assign _EVAL_52 = buffer__EVAL_8;
  assign axi4deint__EVAL_24 = axi4yank__EVAL_77;
  assign axi4yank__EVAL_15 = axi4deint__EVAL_4;
  assign buffer__EVAL_19 = widget__EVAL_30;
  assign axi4yank__EVAL_16 = axi4deint__EVAL_70;
  assign axi4buf__EVAL_22 = axi4yank__EVAL_59;
  assign _EVAL_33 = axi4buf__EVAL_45;
  assign _EVAL_24 = buffer__EVAL_30;
  assign axi4buf__EVAL_15 = axi4yank__EVAL_42;
  assign axi4yank__EVAL_25 = axi4buf__EVAL_30;
  assign axi4index__EVAL_12 = tl2axi4__EVAL_30;
  assign axi4index__EVAL_28 = tl2axi4__EVAL_53;
  assign axi4buf__EVAL_74 = axi4yank__EVAL_3;
  assign axi4buf__EVAL_8 = axi4yank__EVAL_26;
  assign _EVAL_19 = buffer__EVAL_28;
  assign axi4buf__EVAL_10 = axi4yank__EVAL_70;
  assign tl2axi4__EVAL_41 = widget__EVAL_24;
  assign axi4buf__EVAL_61 = axi4yank__EVAL_76;
  assign _EVAL_13 = axi4buf__EVAL_26;
  assign axi4buf__EVAL_70 = axi4yank__EVAL_73;
  assign axi4buf__EVAL_53 = axi4yank__EVAL_39;
  assign axi4index__EVAL_64 = tl2axi4__EVAL_21;
  assign tl2axi4__EVAL_54 = _EVAL_25;
  assign tl2axi4__EVAL_11 = widget__EVAL_4;
  assign axi4deint__EVAL_13 = axi4index__EVAL_9;
  assign axi4buf__EVAL_5 = axi4yank__EVAL_21;
  assign widget__EVAL_27 = buffer__EVAL_9;
  assign axi4yank__EVAL_17 = axi4buf__EVAL_58;
  assign axi4buf__EVAL_44 = axi4yank__EVAL_10;
  assign axi4index__EVAL_62 = tl2axi4__EVAL_14;
  assign axi4index__EVAL_8 = tl2axi4__EVAL_44;
  assign _EVAL_26 = axi4buf__EVAL_35;
  assign axi4buf__EVAL_55 = axi4yank__EVAL_48;
  assign _EVAL_17 = axi4buf__EVAL_25;
  assign axi4deint__EVAL_16 = axi4yank__EVAL_28;
  assign widget__EVAL_11 = tl2axi4__EVAL_35;
  assign axi4index__EVAL_68 = axi4deint__EVAL_75;
  assign axi4deint__EVAL_22 = axi4index__EVAL_55;
  assign axi4deint__EVAL_65 = axi4index__EVAL_66;
  assign _EVAL_21 = axi4buf__EVAL_46;
  assign axi4index__EVAL_50 = axi4deint__EVAL_5;
  assign axi4yank__EVAL_60 = axi4deint__EVAL_82;
  assign axi4yank__EVAL_12 = axi4buf__EVAL_11;
  assign _EVAL_2 = buffer__EVAL_22;
  assign axi4deint__EVAL_11 = axi4index__EVAL_59;
  assign axi4index__EVAL_70 = axi4deint__EVAL_34;
  assign _EVAL_10 = axi4buf__EVAL_21;
  assign axi4deint__EVAL_29 = axi4yank__EVAL;
  assign axi4yank__EVAL_6 = axi4deint__EVAL_48;
  assign tl2axi4__EVAL_51 = axi4index__EVAL_61;
  assign tl2axi4__EVAL_10 = axi4index__EVAL_45;
  assign _EVAL_12 = buffer__EVAL_20;
  assign axi4buf__EVAL_73 = axi4yank__EVAL_71;
  assign axi4deint__EVAL_33 = axi4index__EVAL_13;
  assign widget__EVAL_8 = buffer__EVAL_31;
  assign axi4deint__EVAL_80 = axi4index__EVAL_32;
  assign axi4deint__EVAL_30 = axi4index__EVAL_26;
  assign axi4buf__EVAL_38 = _EVAL_35;
  assign axi4yank__EVAL_5 = axi4deint__EVAL_14;
  assign axi4index__EVAL_46 = axi4deint__EVAL_54;
  assign buffer__EVAL_32 = _EVAL_53;
  assign _EVAL_40 = buffer__EVAL_35;
  assign axi4buf__EVAL_63 = _EVAL_50;
  assign buffer__EVAL_18 = _EVAL_39;
  assign widget__EVAL_5 = buffer__EVAL_11;
  assign axi4buf__EVAL_67 = _EVAL_43;
  assign widget__EVAL_32 = tl2axi4__EVAL_36;
  assign widget__EVAL_7 = buffer__EVAL;
  assign axi4buf__EVAL_60 = axi4yank__EVAL_45;
  assign axi4yank__EVAL_11 = axi4buf__EVAL_3;
  assign axi4deint__EVAL_3 = _EVAL_25;
  assign tl2axi4__EVAL_43 = widget__EVAL_23;
  assign axi4deint__EVAL_19 = axi4index__EVAL;
  assign _EVAL_31 = axi4buf__EVAL_4;
  assign axi4deint__EVAL_39 = axi4yank__EVAL_23;
  assign axi4yank__EVAL_0 = axi4deint__EVAL_63;
  assign axi4buf__EVAL_18 = _EVAL_28;
endmodule
