//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_117_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input  [6:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [29:0] _EVAL_12,
  input  [6:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [2:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [5:0] _EVAL_19;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_31;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_66;
  reg [31:0] _RAND_2;
  reg [5:0] _EVAL_79;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_83;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_85;
  reg [31:0] _RAND_5;
  reg [6:0] _EVAL_109;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_110;
  reg [31:0] _RAND_7;
  reg [29:0] _EVAL_155;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_157;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_161;
  reg [31:0] _RAND_10;
  reg  _EVAL_162;
  reg [31:0] _RAND_11;
  reg [1:0] _EVAL_169;
  reg [31:0] _RAND_12;
  reg [72:0] _EVAL_223;
  reg [95:0] _RAND_13;
  reg [2:0] _EVAL_225;
  reg [31:0] _RAND_14;
  reg [5:0] _EVAL_246;
  reg [31:0] _RAND_15;
  reg  _EVAL_316;
  reg [31:0] _RAND_16;
  wire  _EVAL_42;
  wire  _EVAL_177;
  wire  _EVAL_135;
  wire [3:0] _EVAL_170;
  wire  _EVAL_206;
  wire [2:0] _EVAL_88;
  wire  _EVAL_116;
  wire  _EVAL_61;
  wire  _EVAL_332;
  wire  _EVAL_311;
  wire  _EVAL_25;
  wire  _EVAL_186;
  wire  _EVAL_55;
  wire  _EVAL_207;
  wire  _EVAL_192;
  wire  _EVAL_364;
  wire  _EVAL_59;
  wire [1:0] _EVAL_72;
  wire [1:0] _EVAL_90;
  wire  _EVAL_262;
  wire  _EVAL_307;
  wire  _EVAL_65;
  wire  _EVAL_335;
  wire  _EVAL_54;
  wire [30:0] _EVAL_43;
  wire [30:0] _EVAL_194;
  wire [30:0] _EVAL_199;
  wire  _EVAL_341;
  wire  _EVAL_232;
  wire  _EVAL_240;
  wire  _EVAL_298;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_165;
  wire [29:0] _EVAL_39;
  wire [30:0] _EVAL_112;
  wire [3:0] _EVAL_114;
  wire [29:0] _EVAL_64;
  wire [30:0] _EVAL_357;
  wire [30:0] _EVAL_82;
  wire [30:0] _EVAL_208;
  wire  _EVAL_358;
  wire [30:0] _EVAL_99;
  wire [30:0] _EVAL_49;
  wire  _EVAL_330;
  wire  _EVAL_138;
  wire  _EVAL_159;
  wire  _EVAL_297;
  wire [29:0] _EVAL_271;
  wire [30:0] _EVAL_185;
  wire [30:0] _EVAL_160;
  wire [30:0] _EVAL_68;
  wire  _EVAL_344;
  wire  _EVAL_156;
  wire [29:0] _EVAL_36;
  wire [30:0] _EVAL_180;
  wire [30:0] _EVAL_264;
  wire [30:0] _EVAL_53;
  wire  _EVAL_267;
  wire  _EVAL_184;
  wire [29:0] _EVAL_69;
  wire [30:0] _EVAL_293;
  wire [30:0] _EVAL_242;
  wire [30:0] _EVAL_292;
  wire  _EVAL_77;
  wire  _EVAL_189;
  wire  _EVAL_203;
  wire  _EVAL_171;
  wire  _EVAL_323;
  wire  _EVAL_356;
  wire  _EVAL_62;
  wire  _EVAL_277;
  wire  _EVAL_57;
  wire  _EVAL_179;
  wire [29:0] _EVAL_351;
  wire [30:0] _EVAL_283;
  wire [30:0] _EVAL_152;
  wire [30:0] _EVAL_322;
  wire  _EVAL_128;
  wire  _EVAL_256;
  wire  _EVAL_211;
  wire  _EVAL_362;
  wire  _EVAL_336;
  wire  _EVAL_280;
  wire  _EVAL_93;
  wire  _EVAL_98;
  wire [31:0] _EVAL_241;
  wire  _EVAL_150;
  wire  _EVAL_346;
  wire  _EVAL_96;
  wire  _EVAL_129;
  wire  _EVAL_236;
  wire  _EVAL_350;
  wire  _EVAL_244;
  wire  _EVAL_302;
  wire  _EVAL_305;
  wire  _EVAL_318;
  wire  _EVAL_361;
  wire  _EVAL_123;
  wire  _EVAL_95;
  wire [127:0] _EVAL_331;
  wire [127:0] _EVAL_228;
  wire [72:0] _EVAL_266;
  wire [72:0] _EVAL_313;
  wire [72:0] _EVAL_202;
  wire  _EVAL_288;
  wire  _EVAL_91;
  wire  _EVAL_120;
  wire  _EVAL_259;
  wire  _EVAL_248;
  wire  _EVAL_349;
  wire  _EVAL_260;
  wire  _EVAL_213;
  wire  _EVAL_196;
  wire  _EVAL_193;
  wire  _EVAL_343;
  wire  _EVAL_294;
  wire  _EVAL_75;
  wire  _EVAL_295;
  wire  _EVAL_47;
  wire  _EVAL_272;
  wire  _EVAL_253;
  wire  _EVAL_268;
  wire [72:0] _EVAL_153;
  wire  _EVAL_278;
  wire  _EVAL_360;
  wire  _EVAL_26;
  wire  _EVAL_130;
  wire  _EVAL_34;
  wire  _EVAL_317;
  wire  _EVAL_87;
  wire  _EVAL_78;
  wire  _EVAL_197;
  wire  _EVAL_243;
  wire  _EVAL_63;
  wire  _EVAL_127;
  wire  _EVAL_29;
  wire  _EVAL_235;
  wire  _EVAL_219;
  wire  _EVAL_354;
  wire  _EVAL_124;
  wire  _EVAL_217;
  wire  _EVAL_325;
  wire  _EVAL_178;
  wire [3:0] _EVAL_191;
  wire  _EVAL_113;
  wire [22:0] _EVAL_279;
  wire [7:0] _EVAL_276;
  wire [7:0] _EVAL_21;
  wire [5:0] _EVAL_188;
  wire  _EVAL_89;
  wire  _EVAL_198;
  wire  _EVAL_44;
  wire  _EVAL_97;
  wire  _EVAL_103;
  wire  _EVAL_201;
  wire  _EVAL_76;
  wire  _EVAL_173;
  wire [2:0] _EVAL_275;
  wire  _EVAL_359;
  wire  _EVAL_348;
  wire  _EVAL_338;
  wire  _EVAL_125;
  wire  _EVAL_140;
  wire  _EVAL_282;
  wire  _EVAL_32;
  wire [72:0] _EVAL_94;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_151;
  wire  _EVAL_106;
  wire  _EVAL_117;
  wire  _EVAL_142;
  wire  _EVAL_24;
  wire  _EVAL_299;
  wire  _EVAL_222;
  wire  _EVAL_174;
  wire  _EVAL_190;
  wire  _EVAL_333;
  wire  _EVAL_345;
  wire  _EVAL_50;
  wire  _EVAL_132;
  wire  _EVAL_334;
  wire  _EVAL_229;
  wire  _EVAL_284;
  wire  _EVAL_133;
  wire  _EVAL_340;
  wire  _EVAL_352;
  wire  _EVAL_269;
  wire  _EVAL_70;
  wire  _EVAL_33;
  wire  _EVAL_46;
  wire  _EVAL_215;
  wire  _EVAL_230;
  wire  _EVAL_239;
  wire [3:0] _EVAL_209;
  wire [3:0] _EVAL_30;
  wire  _EVAL_101;
  wire  _EVAL_270;
  wire [22:0] _EVAL_104;
  wire [7:0] _EVAL_231;
  wire [7:0] _EVAL_252;
  wire [29:0] _EVAL_111;
  wire [29:0] _EVAL_126;
  wire  _EVAL_163;
  wire  _EVAL_320;
  wire  _EVAL_210;
  wire [5:0] _EVAL_48;
  wire [5:0] _EVAL_107;
  wire  _EVAL_261;
  wire  _EVAL_314;
  wire  _EVAL_300;
  wire  _EVAL_265;
  wire  _EVAL_176;
  wire  _EVAL_290;
  wire  _EVAL_251;
  wire  _EVAL_175;
  wire  _EVAL_45;
  wire  _EVAL_23;
  wire  _EVAL_181;
  wire  _EVAL_281;
  wire  _EVAL_84;
  wire  _EVAL_339;
  wire  _EVAL_118;
  wire  _EVAL_80;
  wire [5:0] _EVAL_139;
  wire [5:0] _EVAL_28;
  wire  _EVAL_212;
  wire  _EVAL_347;
  wire  _EVAL_245;
  wire  _EVAL_81;
  wire  _EVAL_224;
  wire  _EVAL_51;
  wire  _EVAL_289;
  wire  _EVAL_187;
  wire [127:0] _EVAL_182;
  wire [127:0] _EVAL_321;
  wire [72:0] _EVAL_27;
  wire  _EVAL_20;
  wire  _EVAL_115;
  wire  _EVAL_234;
  wire  _EVAL_355;
  wire  _EVAL_154;
  wire  _EVAL_233;
  wire  _EVAL_35;
  wire  _EVAL_273;
  wire  _EVAL_324;
  wire  _EVAL_285;
  wire [5:0] _EVAL_255;
  wire  _EVAL_329;
  wire  _EVAL_131;
  wire  _EVAL_86;
  wire  _EVAL_287;
  wire  _EVAL_274;
  wire  _EVAL_52;
  wire  _EVAL_204;
  wire  _EVAL_301;
  wire  _EVAL_147;
  wire  _EVAL_250;
  wire  _EVAL_303;
  wire [3:0] _EVAL_195;
  wire  _EVAL_56;
  wire  _EVAL_37;
  wire  _EVAL_102;
  wire  _EVAL_137;
  wire  _EVAL_249;
  wire  _EVAL_41;
  wire  _EVAL_304;
  wire  _EVAL_353;
  wire  _EVAL_92;
  wire  _EVAL_257;
  wire  _EVAL_71;
  wire  _EVAL_286;
  wire  _EVAL_145;
  wire  _EVAL_148;
  wire  _EVAL_158;
  wire  _EVAL_58;
  wire  _EVAL_146;
  wire  _EVAL_74;
  wire  _EVAL_247;
  wire  _EVAL_67;
  wire  _EVAL_263;
  wire  _EVAL_296;
  wire  _EVAL_221;
  wire  _EVAL_40;
  wire  _EVAL_326;
  wire  _EVAL_214;
  wire  _EVAL_308;
  wire  _EVAL_319;
  wire  _EVAL_122;
  wire  _EVAL_342;
  wire  _EVAL_200;
  wire  _EVAL_291;
  wire  _EVAL_258;
  wire [72:0] _EVAL_121;
  wire  _EVAL_136;
  wire  _EVAL_227;
  wire  _EVAL_100;
  wire  _EVAL_108;
  wire  _EVAL_238;
  wire  _EVAL_141;
  wire [72:0] _EVAL_310;
  wire  _EVAL_218;
  wire  _EVAL_220;
  wire  _EVAL_119;
  wire  _EVAL_363;
  wire  _EVAL_366;
  wire  _EVAL_164;
  wire  _EVAL_38;
  wire  _EVAL_337;
  wire  _EVAL_144;
  wire  _EVAL_22;
  wire  _EVAL_315;
  wire  _EVAL_205;
  wire  _EVAL_143;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_42 = _EVAL_5 == 7'h48;
  assign _EVAL_177 = _EVAL_5 == 7'h40;
  assign _EVAL_135 = _EVAL_42 | _EVAL_177;
  assign _EVAL_170 = _EVAL_5[6:3];
  assign _EVAL_206 = _EVAL_170 == 4'h8;
  assign _EVAL_88 = _EVAL_5[2:0];
  assign _EVAL_116 = 3'h1 <= _EVAL_88;
  assign _EVAL_61 = _EVAL_206 & _EVAL_116;
  assign _EVAL_332 = _EVAL_135 | _EVAL_61;
  assign _EVAL_311 = _EVAL_5 == 7'h20;
  assign _EVAL_25 = _EVAL_332 | _EVAL_311;
  assign _EVAL_186 = _EVAL_170 == 4'h0;
  assign _EVAL_55 = _EVAL_25 | _EVAL_186;
  assign _EVAL_207 = _EVAL_170 == 4'h1;
  assign _EVAL_192 = _EVAL_55 | _EVAL_207;
  assign _EVAL_364 = _EVAL_3 >= 4'h2;
  assign _EVAL_59 = _EVAL_3[0];
  assign _EVAL_72 = 2'h1 << _EVAL_59;
  assign _EVAL_90 = _EVAL_72 | 2'h1;
  assign _EVAL_262 = _EVAL_90[1];
  assign _EVAL_307 = _EVAL_12[1];
  assign _EVAL_65 = _EVAL_307 == 1'h0;
  assign _EVAL_335 = _EVAL_262 & _EVAL_65;
  assign _EVAL_54 = _EVAL_364 | _EVAL_335;
  assign _EVAL_43 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_194 = $signed(_EVAL_43) & $signed(-31'sh5000);
  assign _EVAL_199 = $signed(_EVAL_194);
  assign _EVAL_341 = _EVAL_2 <= 2'h2;
  assign _EVAL_232 = _EVAL_10[2];
  assign _EVAL_240 = _EVAL_232 == 1'h0;
  assign _EVAL_298 = _EVAL_10 == 3'h6;
  assign _EVAL_166 = _EVAL_5 == _EVAL_31;
  assign _EVAL_167 = _EVAL_166 | _EVAL_11;
  assign _EVAL_165 = _EVAL_167 == 1'h0;
  assign _EVAL_39 = _EVAL_12 ^ 30'h2000000;
  assign _EVAL_112 = {1'b0,$signed(_EVAL_39)};
  assign _EVAL_114 = _EVAL_13[6:3];
  assign _EVAL_64 = _EVAL_12 ^ 30'hc000000;
  assign _EVAL_357 = {1'b0,$signed(_EVAL_64)};
  assign _EVAL_82 = $signed(_EVAL_357) & $signed(-31'sh4000000);
  assign _EVAL_208 = $signed(_EVAL_82);
  assign _EVAL_358 = $signed(_EVAL_208) == $signed(31'sh0);
  assign _EVAL_99 = $signed(_EVAL_112) & $signed(-31'sh10000);
  assign _EVAL_49 = $signed(_EVAL_99);
  assign _EVAL_330 = $signed(_EVAL_49) == $signed(31'sh0);
  assign _EVAL_138 = _EVAL_358 | _EVAL_330;
  assign _EVAL_159 = $signed(_EVAL_199) == $signed(31'sh0);
  assign _EVAL_297 = _EVAL_138 | _EVAL_159;
  assign _EVAL_271 = _EVAL_12 ^ 30'h1800000;
  assign _EVAL_185 = {1'b0,$signed(_EVAL_271)};
  assign _EVAL_160 = $signed(_EVAL_185) & $signed(-31'sh8000);
  assign _EVAL_68 = $signed(_EVAL_160);
  assign _EVAL_344 = $signed(_EVAL_68) == $signed(31'sh0);
  assign _EVAL_156 = _EVAL_297 | _EVAL_344;
  assign _EVAL_36 = _EVAL_12 ^ 30'h1900000;
  assign _EVAL_180 = {1'b0,$signed(_EVAL_36)};
  assign _EVAL_264 = $signed(_EVAL_180) & $signed(-31'sh2000);
  assign _EVAL_53 = $signed(_EVAL_264);
  assign _EVAL_267 = $signed(_EVAL_53) == $signed(31'sh0);
  assign _EVAL_184 = _EVAL_156 | _EVAL_267;
  assign _EVAL_69 = _EVAL_12 ^ 30'h20000000;
  assign _EVAL_293 = {1'b0,$signed(_EVAL_69)};
  assign _EVAL_242 = $signed(_EVAL_293) & $signed(-31'sh2000);
  assign _EVAL_292 = $signed(_EVAL_242);
  assign _EVAL_77 = $signed(_EVAL_292) == $signed(31'sh0);
  assign _EVAL_189 = _EVAL_184 | _EVAL_77;
  assign _EVAL_203 = _EVAL_13 == 7'h20;
  assign _EVAL_171 = _EVAL_2 == 2'h0;
  assign _EVAL_323 = _EVAL_171 | _EVAL_11;
  assign _EVAL_356 = _EVAL_13 == 7'h40;
  assign _EVAL_62 = 4'h6 == _EVAL_3;
  assign _EVAL_277 = _EVAL_356 ? _EVAL_62 : 1'h0;
  assign _EVAL_57 = _EVAL_364 | _EVAL_11;
  assign _EVAL_179 = _EVAL_3 <= 4'h2;
  assign _EVAL_351 = _EVAL_12 ^ 30'h3000;
  assign _EVAL_283 = {1'b0,$signed(_EVAL_351)};
  assign _EVAL_152 = $signed(_EVAL_283) & $signed(-31'sh1000);
  assign _EVAL_322 = $signed(_EVAL_152);
  assign _EVAL_128 = $signed(_EVAL_322) == $signed(31'sh0);
  assign _EVAL_256 = _EVAL_128 | _EVAL_267;
  assign _EVAL_211 = _EVAL_179 & _EVAL_256;
  assign _EVAL_362 = _EVAL_211 | _EVAL_11;
  assign _EVAL_336 = _EVAL_362 == 1'h0;
  assign _EVAL_280 = _EVAL_8 & _EVAL_6;
  assign _EVAL_93 = _EVAL_16 & _EVAL_1;
  assign _EVAL_98 = _EVAL_280 | _EVAL_93;
  assign _EVAL_241 = _EVAL_83 + 32'h1;
  assign _EVAL_150 = _EVAL_18 == 3'h4;
  assign _EVAL_346 = _EVAL_7 == 1'h0;
  assign _EVAL_96 = _EVAL_346 | _EVAL_11;
  assign _EVAL_129 = _EVAL_13 == _EVAL_109;
  assign _EVAL_236 = _EVAL_129 | _EVAL_11;
  assign _EVAL_350 = _EVAL_18 <= 3'h6;
  assign _EVAL_244 = _EVAL_350 | _EVAL_11;
  assign _EVAL_302 = _EVAL_90[0];
  assign _EVAL_305 = _EVAL_12[0];
  assign _EVAL_318 = _EVAL_65 & _EVAL_305;
  assign _EVAL_361 = _EVAL_302 & _EVAL_318;
  assign _EVAL_123 = _EVAL_157 == 6'h0;
  assign _EVAL_95 = _EVAL_280 & _EVAL_123;
  assign _EVAL_331 = 128'h1 << _EVAL_13;
  assign _EVAL_228 = _EVAL_95 ? _EVAL_331 : 128'h0;
  assign _EVAL_266 = _EVAL_228[72:0];
  assign _EVAL_313 = _EVAL_266 | _EVAL_223;
  assign _EVAL_202 = _EVAL_313 >> _EVAL_5;
  assign _EVAL_288 = _EVAL_202[0];
  assign _EVAL_91 = _EVAL_288 | _EVAL_11;
  assign _EVAL_120 = _EVAL_3 <= 4'h8;
  assign _EVAL_259 = _EVAL_120 & _EVAL_128;
  assign _EVAL_248 = _EVAL_259 | _EVAL_11;
  assign _EVAL_349 = _EVAL_248 == 1'h0;
  assign _EVAL_260 = _EVAL_10 == _EVAL_66;
  assign _EVAL_213 = _EVAL_260 | _EVAL_11;
  assign _EVAL_196 = _EVAL_213 == 1'h0;
  assign _EVAL_193 = _EVAL_18 == 3'h2;
  assign _EVAL_343 = _EVAL_17 != 3'h0;
  assign _EVAL_294 = _EVAL_10 == 3'h1;
  assign _EVAL_75 = _EVAL_170 == 4'h2;
  assign _EVAL_295 = _EVAL_192 | _EVAL_75;
  assign _EVAL_47 = _EVAL_170 == 4'h3;
  assign _EVAL_272 = _EVAL_295 | _EVAL_47;
  assign _EVAL_253 = _EVAL_18 == 3'h6;
  assign _EVAL_268 = _EVAL_253 == 1'h0;
  assign _EVAL_153 = _EVAL_223 >> _EVAL_13;
  assign _EVAL_278 = _EVAL_153[0];
  assign _EVAL_360 = _EVAL_278 == 1'h0;
  assign _EVAL_26 = _EVAL_360 | _EVAL_11;
  assign _EVAL_130 = _EVAL_9 == 1'h0;
  assign _EVAL_34 = _EVAL_130 | _EVAL_11;
  assign _EVAL_317 = _EVAL_34 == 1'h0;
  assign _EVAL_87 = _EVAL_14 >= 4'h2;
  assign _EVAL_78 = _EVAL_87 | _EVAL_11;
  assign _EVAL_197 = _EVAL_114 == 4'h3;
  assign _EVAL_243 = _EVAL_19 == 6'h0;
  assign _EVAL_63 = _EVAL_243 == 1'h0;
  assign _EVAL_127 = _EVAL_346 | _EVAL;
  assign _EVAL_29 = _EVAL_127 | _EVAL_11;
  assign _EVAL_235 = _EVAL_29 == 1'h0;
  assign _EVAL_219 = _EVAL_12 == _EVAL_155;
  assign _EVAL_354 = _EVAL_305 == 1'h0;
  assign _EVAL_124 = _EVAL_65 & _EVAL_354;
  assign _EVAL_217 = _EVAL_302 & _EVAL_124;
  assign _EVAL_325 = _EVAL_54 | _EVAL_217;
  assign _EVAL_178 = _EVAL_83 < plusarg_reader_out;
  assign _EVAL_191 = ~ _EVAL_15;
  assign _EVAL_113 = _EVAL_191 == 4'h0;
  assign _EVAL_279 = 23'hff << _EVAL_14;
  assign _EVAL_276 = _EVAL_279[7:0];
  assign _EVAL_21 = ~ _EVAL_276;
  assign _EVAL_188 = _EVAL_21[7:2];
  assign _EVAL_89 = _EVAL_3 <= 4'h6;
  assign _EVAL_198 = _EVAL_89 & _EVAL_189;
  assign _EVAL_44 = _EVAL_259 | _EVAL_198;
  assign _EVAL_97 = _EVAL_44 | _EVAL_11;
  assign _EVAL_103 = _EVAL_97 == 1'h0;
  assign _EVAL_201 = _EVAL_13 == 7'h48;
  assign _EVAL_76 = _EVAL_201 | _EVAL_356;
  assign _EVAL_173 = _EVAL_114 == 4'h8;
  assign _EVAL_275 = _EVAL_13[2:0];
  assign _EVAL_359 = 3'h1 <= _EVAL_275;
  assign _EVAL_348 = _EVAL_173 & _EVAL_359;
  assign _EVAL_338 = _EVAL_76 | _EVAL_348;
  assign _EVAL_125 = _EVAL_2 == _EVAL_169;
  assign _EVAL_140 = _EVAL_1 & _EVAL_63;
  assign _EVAL_282 = _EVAL_93 & _EVAL_243;
  assign _EVAL_32 = _EVAL_17 <= 3'h2;
  assign _EVAL_94 = _EVAL_223 | _EVAL_266;
  assign _EVAL_327 = _EVAL_262 & _EVAL_307;
  assign _EVAL_328 = _EVAL_364 | _EVAL_327;
  assign _EVAL_151 = _EVAL_307 & _EVAL_305;
  assign _EVAL_106 = _EVAL_302 & _EVAL_151;
  assign _EVAL_117 = _EVAL_328 | _EVAL_106;
  assign _EVAL_142 = _EVAL_10 == 3'h7;
  assign _EVAL_24 = _EVAL_6 & _EVAL_142;
  assign _EVAL_299 = _EVAL_18 == 3'h0;
  assign _EVAL_222 = _EVAL_1 & _EVAL_193;
  assign _EVAL_174 = _EVAL_3 == _EVAL_110;
  assign _EVAL_190 = _EVAL_174 | _EVAL_11;
  assign _EVAL_333 = _EVAL_4 == _EVAL_316;
  assign _EVAL_345 = _EVAL_333 | _EVAL_11;
  assign _EVAL_50 = _EVAL_18 == _EVAL_85;
  assign _EVAL_132 = _EVAL_50 | _EVAL_11;
  assign _EVAL_334 = _EVAL_132 == 1'h0;
  assign _EVAL_229 = _EVAL_10 == 3'h3;
  assign _EVAL_284 = _EVAL_6 & _EVAL_229;
  assign _EVAL_133 = _EVAL_79 == 6'h0;
  assign _EVAL_340 = _EVAL_133 == 1'h0;
  assign _EVAL_352 = _EVAL_10 == 3'h2;
  assign _EVAL_269 = _EVAL_6 & _EVAL_352;
  assign _EVAL_70 = _EVAL_341 | _EVAL_11;
  assign _EVAL_33 = _EVAL_18[0];
  assign _EVAL_46 = _EVAL_307 & _EVAL_354;
  assign _EVAL_215 = _EVAL_302 & _EVAL_46;
  assign _EVAL_230 = _EVAL_328 | _EVAL_215;
  assign _EVAL_239 = _EVAL_54 | _EVAL_361;
  assign _EVAL_209 = {_EVAL_117,_EVAL_230,_EVAL_239,_EVAL_325};
  assign _EVAL_30 = ~ _EVAL_209;
  assign _EVAL_101 = _EVAL_343 | _EVAL_11;
  assign _EVAL_270 = _EVAL_113 | _EVAL_11;
  assign _EVAL_104 = 23'hff << _EVAL_3;
  assign _EVAL_231 = _EVAL_104[7:0];
  assign _EVAL_252 = ~ _EVAL_231;
  assign _EVAL_111 = {{22'd0}, _EVAL_252};
  assign _EVAL_126 = _EVAL_12 & _EVAL_111;
  assign _EVAL_163 = _EVAL_126 == 30'h0;
  assign _EVAL_320 = _EVAL_163 | _EVAL_11;
  assign _EVAL_210 = _EVAL_320 == 1'h0;
  assign _EVAL_48 = _EVAL_252[7:2];
  assign _EVAL_107 = _EVAL_157 - 6'h1;
  assign _EVAL_261 = _EVAL_17 == 3'h0;
  assign _EVAL_314 = _EVAL_261 | _EVAL_11;
  assign _EVAL_300 = _EVAL_314 == 1'h0;
  assign _EVAL_265 = _EVAL_270 == 1'h0;
  assign _EVAL_176 = _EVAL_223 != 73'h0;
  assign _EVAL_290 = _EVAL_176 == 1'h0;
  assign _EVAL_251 = plusarg_reader_out == 32'h0;
  assign _EVAL_175 = _EVAL_290 | _EVAL_251;
  assign _EVAL_45 = _EVAL_236 == 1'h0;
  assign _EVAL_23 = _EVAL_338 | _EVAL_203;
  assign _EVAL_181 = _EVAL_114 == 4'h0;
  assign _EVAL_281 = _EVAL_23 | _EVAL_181;
  assign _EVAL_84 = _EVAL_114 == 4'h1;
  assign _EVAL_339 = _EVAL_281 | _EVAL_84;
  assign _EVAL_118 = _EVAL_114 == 4'h2;
  assign _EVAL_80 = _EVAL_339 | _EVAL_118;
  assign _EVAL_139 = _EVAL_19 - 6'h1;
  assign _EVAL_28 = _EVAL_79 - 6'h1;
  assign _EVAL_212 = _EVAL_32 | _EVAL_11;
  assign _EVAL_347 = _EVAL_17 <= 3'h3;
  assign _EVAL_245 = _EVAL_347 | _EVAL_11;
  assign _EVAL_81 = _EVAL_245 == 1'h0;
  assign _EVAL_224 = _EVAL_10 == 3'h0;
  assign _EVAL_51 = _EVAL_246 == 6'h0;
  assign _EVAL_289 = _EVAL_93 & _EVAL_51;
  assign _EVAL_187 = _EVAL_289 & _EVAL_268;
  assign _EVAL_182 = 128'h1 << _EVAL_5;
  assign _EVAL_321 = _EVAL_187 ? _EVAL_182 : 128'h0;
  assign _EVAL_27 = _EVAL_321[72:0];
  assign _EVAL_20 = _EVAL_266 != _EVAL_27;
  assign _EVAL_115 = _EVAL_175 | _EVAL_178;
  assign _EVAL_234 = _EVAL_115 | _EVAL_11;
  assign _EVAL_355 = _EVAL_266 != 73'h0;
  assign _EVAL_154 = _EVAL_355 == 1'h0;
  assign _EVAL_233 = _EVAL_15 == _EVAL_209;
  assign _EVAL_35 = _EVAL_17 <= 3'h4;
  assign _EVAL_273 = _EVAL_35 | _EVAL_11;
  assign _EVAL_324 = _EVAL_10 == 3'h4;
  assign _EVAL_285 = _EVAL_1 & _EVAL_253;
  assign _EVAL_255 = _EVAL_246 - 6'h1;
  assign _EVAL_329 = _EVAL_10 == 3'h5;
  assign _EVAL_131 = _EVAL_6 & _EVAL_329;
  assign _EVAL_86 = _EVAL_91 == 1'h0;
  assign _EVAL_287 = _EVAL_2 != 2'h2;
  assign _EVAL_274 = _EVAL_287 | _EVAL_11;
  assign _EVAL_52 = _EVAL_18 == 3'h5;
  assign _EVAL_204 = _EVAL_6 & _EVAL_298;
  assign _EVAL_301 = _EVAL_277 | _EVAL_11;
  assign _EVAL_147 = _EVAL_301 == 1'h0;
  assign _EVAL_250 = _EVAL_96 == 1'h0;
  assign _EVAL_303 = _EVAL_219 | _EVAL_11;
  assign _EVAL_195 = _EVAL_15 & _EVAL_30;
  assign _EVAL_56 = _EVAL_7 == _EVAL_162;
  assign _EVAL_37 = _EVAL_56 | _EVAL_11;
  assign _EVAL_102 = _EVAL_14 == _EVAL_161;
  assign _EVAL_137 = _EVAL_102 | _EVAL_11;
  assign _EVAL_249 = _EVAL_137 == 1'h0;
  assign _EVAL_41 = _EVAL == 1'h0;
  assign _EVAL_304 = _EVAL_41 | _EVAL_11;
  assign _EVAL_353 = _EVAL_304 == 1'h0;
  assign _EVAL_92 = _EVAL_190 == 1'h0;
  assign _EVAL_257 = _EVAL_17 == _EVAL_225;
  assign _EVAL_71 = _EVAL_257 | _EVAL_11;
  assign _EVAL_286 = _EVAL_6 & _EVAL_324;
  assign _EVAL_145 = _EVAL_212 == 1'h0;
  assign _EVAL_148 = _EVAL_272 | _EVAL_11;
  assign _EVAL_158 = _EVAL_148 == 1'h0;
  assign _EVAL_58 = _EVAL_57 == 1'h0;
  assign _EVAL_146 = _EVAL_80 | _EVAL_197;
  assign _EVAL_74 = _EVAL_146 | _EVAL_11;
  assign _EVAL_247 = _EVAL_273 == 1'h0;
  assign _EVAL_67 = _EVAL_234 == 1'h0;
  assign _EVAL_263 = _EVAL_6 & _EVAL_224;
  assign _EVAL_296 = _EVAL_233 | _EVAL_11;
  assign _EVAL_221 = _EVAL_296 == 1'h0;
  assign _EVAL_40 = _EVAL_18 == 3'h1;
  assign _EVAL_326 = _EVAL_1 & _EVAL_40;
  assign _EVAL_214 = _EVAL_280 & _EVAL_133;
  assign _EVAL_308 = _EVAL_20 | _EVAL_154;
  assign _EVAL_319 = _EVAL_244 == 1'h0;
  assign _EVAL_122 = _EVAL_71 == 1'h0;
  assign _EVAL_342 = _EVAL_74 == 1'h0;
  assign _EVAL_200 = _EVAL_308 | _EVAL_11;
  assign _EVAL_291 = _EVAL_200 == 1'h0;
  assign _EVAL_258 = _EVAL_78 == 1'h0;
  assign _EVAL_121 = ~ _EVAL_27;
  assign _EVAL_136 = _EVAL_125 | _EVAL_11;
  assign _EVAL_227 = _EVAL_136 == 1'h0;
  assign _EVAL_100 = _EVAL_345 == 1'h0;
  assign _EVAL_108 = _EVAL_303 == 1'h0;
  assign _EVAL_238 = _EVAL_101 == 1'h0;
  assign _EVAL_141 = _EVAL_11 == 1'h0;
  assign _EVAL_310 = _EVAL_94 & _EVAL_121;
  assign _EVAL_218 = _EVAL_274 == 1'h0;
  assign _EVAL_220 = _EVAL_195 == 4'h0;
  assign _EVAL_119 = _EVAL_220 | _EVAL_11;
  assign _EVAL_363 = _EVAL_119 == 1'h0;
  assign _EVAL_366 = _EVAL_26 == 1'h0;
  assign _EVAL_164 = _EVAL_323 == 1'h0;
  assign _EVAL_38 = _EVAL_6 & _EVAL_294;
  assign _EVAL_337 = _EVAL_1 & _EVAL_299;
  assign _EVAL_144 = _EVAL_1 & _EVAL_150;
  assign _EVAL_22 = _EVAL_1 & _EVAL_52;
  assign _EVAL_315 = _EVAL_6 & _EVAL_340;
  assign _EVAL_205 = _EVAL_70 == 1'h0;
  assign _EVAL_143 = _EVAL_37 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_19 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_31 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_66 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_79 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_83 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_85 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_109 = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_110 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_155 = _RAND_8[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_157 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_161 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_162 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_169 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {3{`RANDOM}};
  _EVAL_223 = _RAND_13[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_225 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_246 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_316 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_11) begin
      _EVAL_19 <= 6'h0;
    end else begin
      if (_EVAL_93) begin
        if (_EVAL_243) begin
          if (_EVAL_33) begin
            _EVAL_19 <= _EVAL_188;
          end else begin
            _EVAL_19 <= 6'h0;
          end
        end else begin
          _EVAL_19 <= _EVAL_139;
        end
      end
    end
    if (_EVAL_282) begin
      _EVAL_31 <= _EVAL_5;
    end
    if (_EVAL_214) begin
      _EVAL_66 <= _EVAL_10;
    end
    if (_EVAL_11) begin
      _EVAL_79 <= 6'h0;
    end else begin
      if (_EVAL_280) begin
        if (_EVAL_133) begin
          if (_EVAL_240) begin
            _EVAL_79 <= _EVAL_48;
          end else begin
            _EVAL_79 <= 6'h0;
          end
        end else begin
          _EVAL_79 <= _EVAL_28;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_83 <= 32'h0;
    end else begin
      if (_EVAL_98) begin
        _EVAL_83 <= 32'h0;
      end else begin
        _EVAL_83 <= _EVAL_241;
      end
    end
    if (_EVAL_282) begin
      _EVAL_85 <= _EVAL_18;
    end
    if (_EVAL_214) begin
      _EVAL_109 <= _EVAL_13;
    end
    if (_EVAL_214) begin
      _EVAL_110 <= _EVAL_3;
    end
    if (_EVAL_214) begin
      _EVAL_155 <= _EVAL_12;
    end
    if (_EVAL_11) begin
      _EVAL_157 <= 6'h0;
    end else begin
      if (_EVAL_280) begin
        if (_EVAL_123) begin
          if (_EVAL_240) begin
            _EVAL_157 <= _EVAL_48;
          end else begin
            _EVAL_157 <= 6'h0;
          end
        end else begin
          _EVAL_157 <= _EVAL_107;
        end
      end
    end
    if (_EVAL_282) begin
      _EVAL_161 <= _EVAL_14;
    end
    if (_EVAL_282) begin
      _EVAL_162 <= _EVAL_7;
    end
    if (_EVAL_282) begin
      _EVAL_169 <= _EVAL_2;
    end
    if (_EVAL_11) begin
      _EVAL_223 <= 73'h0;
    end else begin
      _EVAL_223 <= _EVAL_310;
    end
    if (_EVAL_214) begin
      _EVAL_225 <= _EVAL_17;
    end
    if (_EVAL_11) begin
      _EVAL_246 <= 6'h0;
    end else begin
      if (_EVAL_93) begin
        if (_EVAL_51) begin
          if (_EVAL_33) begin
            _EVAL_246 <= _EVAL_188;
          end else begin
            _EVAL_246 <= 6'h0;
          end
        end else begin
          _EVAL_246 <= _EVAL_255;
        end
      end
    end
    if (_EVAL_282) begin
      _EVAL_316 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(553ff9b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2df5bfa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a68cea46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7c773d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_336) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9993b59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14391ed5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8deca50c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e0362a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a8128b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a473f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ede844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4f3577f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(431be397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_349) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f7887d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a97e2a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5768a7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22f8c31b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd3c689a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63004937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ea55a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fcfc05a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42165537)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41ab8f4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6521103)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46b644c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb2efec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23682a43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50045a8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce57c6f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5352b887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f44194f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd145e34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dcc33c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eab393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef978bcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f42f46ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(573b8e2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86eb325d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63776452)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d8a986e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d1900e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2280750f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_336) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ffef9b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e4cf363)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44c271d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_336) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c507ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e08b0197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51f9a284)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d0bfc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28512dbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(178f26db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d59d1b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4b1c0b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4faa449d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e58c25af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8d16446)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83cf6506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfc1f03f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_349) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed121c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8213080f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f99c0fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1b9134)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f690da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95816ffb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34f7ce5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_336) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7be39bd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8215ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed1d8b82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f01ae7c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a039c27a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a880b14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5b56c2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4f66bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c95618d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1631da3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4266a674)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ff1b596)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b088fd49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4135ec3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7194b43f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86832af8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a68b74e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77244d82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b02289d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e3cd3d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfa59a4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_334) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c561d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62c61119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(535ce5e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(273d886e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
