//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_326(
  output [63:0] _EVAL,
  input         _EVAL_0,
  output [3:0]  _EVAL_1,
  input  [6:0]  _EVAL_2,
  input         _EVAL_3,
  input  [29:0] _EVAL_4,
  input  [6:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  output [2:0]  _EVAL_8,
  input  [63:0] _EVAL_9,
  output [3:0]  _EVAL_10,
  output [1:0]  _EVAL_11,
  output [29:0] _EVAL_12,
  output [2:0]  _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  input  [1:0]  _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  output [6:0]  _EVAL_19,
  input         _EVAL_20,
  output [6:0]  _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  input  [63:0] _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  input  [2:0]  _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [7:0]  _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  output [7:0]  _EVAL_36,
  output [63:0] _EVAL_37,
  input         _EVAL_38,
  output [2:0]  _EVAL_39,
  input         _EVAL_40
);
  assign _EVAL_12 = _EVAL_4;
  assign _EVAL_36 = _EVAL_33;
  assign _EVAL_17 = _EVAL_38;
  assign _EVAL_28 = _EVAL_26;
  assign _EVAL_37 = _EVAL_24;
  assign _EVAL_21 = _EVAL_2;
  assign _EVAL = _EVAL_9;
  assign _EVAL_11 = _EVAL_16;
  assign _EVAL_14 = _EVAL_40;
  assign _EVAL_13 = _EVAL_27;
  assign _EVAL_19 = _EVAL_5;
  assign _EVAL_39 = _EVAL_25;
  assign _EVAL_22 = _EVAL_35;
  assign _EVAL_15 = _EVAL_29;
  assign _EVAL_1 = _EVAL_6;
  assign _EVAL_23 = _EVAL_20;
  assign _EVAL_30 = _EVAL_3;
  assign _EVAL_8 = _EVAL_32;
  assign _EVAL_10 = _EVAL_7;
  assign _EVAL_34 = _EVAL_31;
endmodule
