//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_245_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [24:0] _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [2:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_57;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_86;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_90;
  reg [31:0] _RAND_2;
  reg [24:0] _EVAL_102;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_103;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_108;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_132;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_142;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_149;
  reg [31:0] _RAND_8;
  reg [31:0] _EVAL_169;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_183;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_185;
  reg [31:0] _RAND_11;
  reg [7:0] _EVAL_204;
  reg [31:0] _RAND_12;
  reg [3:0] _EVAL_235;
  reg [31:0] _RAND_13;
  wire  _EVAL_31;
  wire  _EVAL_220;
  wire [1:0] _EVAL_253;
  wire [1:0] _EVAL_34;
  wire  _EVAL_52;
  wire  _EVAL_186;
  wire  _EVAL_81;
  wire  _EVAL_21;
  wire  _EVAL_75;
  wire  _EVAL_26;
  wire  _EVAL_252;
  wire  _EVAL_197;
  wire  _EVAL_65;
  wire  _EVAL_157;
  wire  _EVAL_122;
  wire  _EVAL_119;
  wire  _EVAL_206;
  wire  _EVAL_242;
  wire  _EVAL_213;
  wire  _EVAL_247;
  wire  _EVAL_112;
  wire  _EVAL_66;
  wire  _EVAL_255;
  wire  _EVAL_36;
  wire  _EVAL_257;
  wire  _EVAL_37;
  wire  _EVAL_33;
  wire [12:0] _EVAL_22;
  wire [5:0] _EVAL_251;
  wire [5:0] _EVAL_41;
  wire [24:0] _EVAL_146;
  wire [24:0] _EVAL_73;
  wire  _EVAL_85;
  wire  _EVAL_82;
  wire  _EVAL_196;
  wire  _EVAL_193;
  wire  _EVAL_228;
  wire  _EVAL_100;
  wire  _EVAL_258;
  wire  _EVAL_71;
  wire  _EVAL_125;
  wire  _EVAL_246;
  wire  _EVAL_231;
  wire  _EVAL_115;
  wire  _EVAL_171;
  wire [3:0] _EVAL_249;
  wire  _EVAL_162;
  wire  _EVAL_89;
  wire  _EVAL_28;
  wire [7:0] _EVAL_194;
  wire [7:0] _EVAL_224;
  wire  _EVAL_46;
  wire  _EVAL_244;
  wire  _EVAL_61;
  wire  _EVAL_189;
  wire  _EVAL_178;
  wire [7:0] _EVAL_42;
  wire [7:0] _EVAL_83;
  wire  _EVAL_234;
  wire  _EVAL_222;
  wire  _EVAL_216;
  wire  _EVAL_24;
  wire  _EVAL_210;
  wire  _EVAL_54;
  wire [7:0] _EVAL_98;
  wire [7:0] _EVAL_129;
  wire  _EVAL_236;
  wire  _EVAL_165;
  wire [3:0] _EVAL_135;
  wire  _EVAL_151;
  wire  _EVAL_248;
  wire  _EVAL_69;
  wire [7:0] _EVAL_97;
  wire  _EVAL_177;
  wire  _EVAL_120;
  wire  _EVAL_80;
  wire  _EVAL_250;
  wire  _EVAL_200;
  wire  _EVAL_137;
  wire  _EVAL_30;
  wire  _EVAL_188;
  wire  _EVAL_43;
  wire  _EVAL_111;
  wire  _EVAL_172;
  wire  _EVAL_76;
  wire  _EVAL_239;
  wire  _EVAL_136;
  wire  _EVAL_92;
  wire  _EVAL_145;
  wire  _EVAL_192;
  wire  _EVAL_211;
  wire  _EVAL_240;
  wire  _EVAL_121;
  wire  _EVAL_214;
  wire  _EVAL_68;
  wire  _EVAL_88;
  wire  _EVAL_87;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_138;
  wire  _EVAL_110;
  wire [3:0] _EVAL_215;
  wire  _EVAL_72;
  wire  _EVAL_203;
  wire [24:0] _EVAL_101;
  wire [25:0] _EVAL_152;
  wire [25:0] _EVAL_238;
  wire [25:0] _EVAL_230;
  wire  _EVAL_49;
  wire  _EVAL_77;
  wire  _EVAL_114;
  wire  _EVAL_140;
  wire  _EVAL_182;
  wire [3:0] _EVAL_19;
  wire  _EVAL_219;
  wire  _EVAL_59;
  wire  _EVAL_217;
  wire  _EVAL_93;
  wire  _EVAL_212;
  wire  _EVAL_15;
  wire  _EVAL_170;
  wire [3:0] _EVAL_148;
  wire [3:0] _EVAL_60;
  wire  _EVAL_187;
  wire  _EVAL_180;
  wire [12:0] _EVAL_53;
  wire [5:0] _EVAL_199;
  wire [5:0] _EVAL_127;
  wire [3:0] _EVAL_96;
  wire  _EVAL_233;
  wire  _EVAL_51;
  wire  _EVAL_113;
  wire  _EVAL_64;
  wire  _EVAL_91;
  wire  _EVAL_184;
  wire  _EVAL_202;
  wire  _EVAL_159;
  wire  _EVAL_176;
  wire  _EVAL_198;
  wire  _EVAL_105;
  wire  _EVAL_168;
  wire  _EVAL_167;
  wire  _EVAL_118;
  wire  _EVAL_227;
  wire  _EVAL_84;
  wire  _EVAL_237;
  wire  _EVAL_106;
  wire  _EVAL_131;
  wire  _EVAL_143;
  wire [7:0] _EVAL_32;
  wire  _EVAL_70;
  wire  _EVAL_99;
  wire [31:0] _EVAL_218;
  wire  _EVAL_48;
  wire  _EVAL_174;
  wire  _EVAL_63;
  wire  _EVAL_209;
  wire  _EVAL_156;
  wire  _EVAL_223;
  wire [3:0] _EVAL_67;
  wire [3:0] _EVAL_221;
  wire  _EVAL_256;
  wire  _EVAL_39;
  wire  _EVAL_158;
  wire  _EVAL_161;
  wire  _EVAL_163;
  wire [3:0] _EVAL_74;
  wire  _EVAL_35;
  wire  _EVAL_241;
  wire  _EVAL_173;
  wire  _EVAL_153;
  wire  _EVAL_56;
  wire  _EVAL_208;
  wire  _EVAL_27;
  wire  _EVAL_226;
  wire  _EVAL_95;
  wire  _EVAL_179;
  wire  _EVAL_104;
  wire [7:0] _EVAL_107;
  wire  _EVAL_25;
  wire  _EVAL_40;
  wire  _EVAL_109;
  wire  _EVAL_29;
  wire  _EVAL_160;
  wire  _EVAL_245;
  wire  _EVAL_225;
  wire  _EVAL_144;
  wire  _EVAL_229;
  wire  _EVAL_175;
  wire  _EVAL_191;
  wire  _EVAL_45;
  wire  _EVAL_232;
  wire  _EVAL_117;
  wire  _EVAL_50;
  wire  _EVAL_164;
  wire  _EVAL_205;
  wire [7:0] _EVAL_141;
  wire  _EVAL_201;
  wire  _EVAL_150;
  wire  _EVAL_55;
  wire  _EVAL_181;
  wire  _EVAL_23;
  wire  _EVAL_139;
  wire  _EVAL_17;
  wire  _EVAL_130;
  wire  _EVAL_20;
  wire  _EVAL_128;
  wire  _EVAL_58;
  wire  _EVAL_124;
  wire  _EVAL_166;
  wire  _EVAL_44;
  wire  _EVAL_116;
  wire  _EVAL_195;
  wire  _EVAL_16;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_31 = _EVAL_10 >= 3'h2;
  assign _EVAL_220 = _EVAL_10[0];
  assign _EVAL_253 = 2'h1 << _EVAL_220;
  assign _EVAL_34 = _EVAL_253 | 2'h1;
  assign _EVAL_52 = _EVAL_34[1];
  assign _EVAL_186 = _EVAL_2[1];
  assign _EVAL_81 = _EVAL_186 == 1'h0;
  assign _EVAL_21 = _EVAL_52 & _EVAL_81;
  assign _EVAL_75 = _EVAL_31 | _EVAL_21;
  assign _EVAL_26 = _EVAL_34[0];
  assign _EVAL_252 = _EVAL_2[0];
  assign _EVAL_197 = _EVAL_252 == 1'h0;
  assign _EVAL_65 = _EVAL_81 & _EVAL_197;
  assign _EVAL_157 = _EVAL_26 & _EVAL_65;
  assign _EVAL_122 = _EVAL_75 | _EVAL_157;
  assign _EVAL_119 = _EVAL_7 == 3'h0;
  assign _EVAL_206 = 3'h1 <= _EVAL_7;
  assign _EVAL_242 = _EVAL_119 | _EVAL_206;
  assign _EVAL_213 = _EVAL_4 == _EVAL_132;
  assign _EVAL_247 = _EVAL_213 | _EVAL_8;
  assign _EVAL_112 = _EVAL_247 == 1'h0;
  assign _EVAL_66 = _EVAL == 3'h3;
  assign _EVAL_255 = _EVAL_5 & _EVAL_66;
  assign _EVAL_36 = _EVAL_108 == 4'h0;
  assign _EVAL_257 = _EVAL_14 <= 3'h2;
  assign _EVAL_37 = _EVAL_257 | _EVAL_8;
  assign _EVAL_33 = _EVAL_8 == 1'h0;
  assign _EVAL_22 = 13'h3f << _EVAL_10;
  assign _EVAL_251 = _EVAL_22[5:0];
  assign _EVAL_41 = ~ _EVAL_251;
  assign _EVAL_146 = {{19'd0}, _EVAL_41};
  assign _EVAL_73 = _EVAL_2 & _EVAL_146;
  assign _EVAL_85 = _EVAL_73 == 25'h0;
  assign _EVAL_82 = _EVAL_85 | _EVAL_8;
  assign _EVAL_196 = 3'h6 == _EVAL_10;
  assign _EVAL_193 = _EVAL_119 ? _EVAL_196 : 1'h0;
  assign _EVAL_228 = _EVAL_193 | _EVAL_8;
  assign _EVAL_100 = _EVAL_3 == _EVAL_183;
  assign _EVAL_258 = _EVAL_100 | _EVAL_8;
  assign _EVAL_71 = _EVAL_4 == 3'h0;
  assign _EVAL_125 = 3'h1 <= _EVAL_4;
  assign _EVAL_246 = _EVAL_71 | _EVAL_125;
  assign _EVAL_231 = _EVAL_246 | _EVAL_8;
  assign _EVAL_115 = _EVAL_11 <= 3'h6;
  assign _EVAL_171 = _EVAL_115 | _EVAL_8;
  assign _EVAL_249 = _EVAL_57 - 4'h1;
  assign _EVAL_162 = _EVAL_9 & _EVAL_5;
  assign _EVAL_89 = _EVAL_235 == 4'h0;
  assign _EVAL_28 = _EVAL_162 & _EVAL_89;
  assign _EVAL_194 = 8'h1 << _EVAL_7;
  assign _EVAL_224 = _EVAL_28 ? _EVAL_194 : 8'h0;
  assign _EVAL_46 = _EVAL_6 & _EVAL_1;
  assign _EVAL_244 = _EVAL_46 & _EVAL_36;
  assign _EVAL_61 = _EVAL_11 == 3'h6;
  assign _EVAL_189 = _EVAL_61 == 1'h0;
  assign _EVAL_178 = _EVAL_244 & _EVAL_189;
  assign _EVAL_42 = 8'h1 << _EVAL_4;
  assign _EVAL_83 = _EVAL_178 ? _EVAL_42 : 8'h0;
  assign _EVAL_234 = _EVAL_224 != _EVAL_83;
  assign _EVAL_222 = _EVAL_224 != 8'h0;
  assign _EVAL_216 = _EVAL_222 == 1'h0;
  assign _EVAL_24 = _EVAL_234 | _EVAL_216;
  assign _EVAL_210 = _EVAL_24 | _EVAL_8;
  assign _EVAL_54 = _EVAL_186 & _EVAL_252;
  assign _EVAL_98 = _EVAL_224 | _EVAL_204;
  assign _EVAL_129 = _EVAL_98 >> _EVAL_4;
  assign _EVAL_236 = _EVAL_129[0];
  assign _EVAL_165 = _EVAL_236 | _EVAL_8;
  assign _EVAL_135 = ~ _EVAL_13;
  assign _EVAL_151 = _EVAL_135 == 4'h0;
  assign _EVAL_248 = _EVAL_151 | _EVAL_8;
  assign _EVAL_69 = _EVAL_258 == 1'h0;
  assign _EVAL_97 = _EVAL_204 >> _EVAL_7;
  assign _EVAL_177 = _EVAL_97[0];
  assign _EVAL_120 = _EVAL == 3'h1;
  assign _EVAL_80 = _EVAL_5 & _EVAL_120;
  assign _EVAL_250 = _EVAL_2 == _EVAL_102;
  assign _EVAL_200 = _EVAL_250 | _EVAL_8;
  assign _EVAL_137 = _EVAL_14 != 3'h0;
  assign _EVAL_30 = _EVAL_137 | _EVAL_8;
  assign _EVAL_188 = _EVAL_30 == 1'h0;
  assign _EVAL_43 = _EVAL_204 != 8'h0;
  assign _EVAL_111 = _EVAL_43 == 1'h0;
  assign _EVAL_172 = plusarg_reader_out == 32'h0;
  assign _EVAL_76 = _EVAL_111 | _EVAL_172;
  assign _EVAL_239 = _EVAL_11 == 3'h2;
  assign _EVAL_136 = _EVAL_82 == 1'h0;
  assign _EVAL_92 = _EVAL_11 == 3'h5;
  assign _EVAL_145 = _EVAL_1 & _EVAL_92;
  assign _EVAL_192 = _EVAL_185 == 4'h0;
  assign _EVAL_211 = _EVAL_162 & _EVAL_192;
  assign _EVAL_240 = _EVAL_52 & _EVAL_186;
  assign _EVAL_121 = _EVAL_31 | _EVAL_240;
  assign _EVAL_214 = _EVAL_26 & _EVAL_54;
  assign _EVAL_68 = _EVAL_121 | _EVAL_214;
  assign _EVAL_88 = _EVAL_186 & _EVAL_197;
  assign _EVAL_87 = _EVAL_26 & _EVAL_88;
  assign _EVAL_133 = _EVAL_121 | _EVAL_87;
  assign _EVAL_134 = _EVAL_81 & _EVAL_252;
  assign _EVAL_138 = _EVAL_26 & _EVAL_134;
  assign _EVAL_110 = _EVAL_75 | _EVAL_138;
  assign _EVAL_215 = {_EVAL_68,_EVAL_133,_EVAL_110,_EVAL_122};
  assign _EVAL_72 = _EVAL_13 == _EVAL_215;
  assign _EVAL_203 = _EVAL_10 <= 3'h6;
  assign _EVAL_101 = _EVAL_2 ^ 25'h1900000;
  assign _EVAL_152 = {1'b0,$signed(_EVAL_101)};
  assign _EVAL_238 = $signed(_EVAL_152) & $signed(-26'sh2000);
  assign _EVAL_230 = $signed(_EVAL_238);
  assign _EVAL_49 = $signed(_EVAL_230) == $signed(26'sh0);
  assign _EVAL_77 = _EVAL_203 & _EVAL_49;
  assign _EVAL_114 = _EVAL_77 | _EVAL_8;
  assign _EVAL_140 = _EVAL_114 == 1'h0;
  assign _EVAL_182 = _EVAL_57 == 4'h0;
  assign _EVAL_19 = _EVAL_108 - 4'h1;
  assign _EVAL_219 = _EVAL_192 == 1'h0;
  assign _EVAL_59 = _EVAL_5 & _EVAL_219;
  assign _EVAL_217 = _EVAL_11 == _EVAL_103;
  assign _EVAL_93 = _EVAL_217 | _EVAL_8;
  assign _EVAL_212 = _EVAL_93 == 1'h0;
  assign _EVAL_15 = _EVAL[2];
  assign _EVAL_170 = _EVAL_15 == 1'h0;
  assign _EVAL_148 = _EVAL_41[5:2];
  assign _EVAL_60 = _EVAL_185 - 4'h1;
  assign _EVAL_187 = _EVAL_182 == 1'h0;
  assign _EVAL_180 = _EVAL_11[0];
  assign _EVAL_53 = 13'h3f << _EVAL_3;
  assign _EVAL_199 = _EVAL_53[5:0];
  assign _EVAL_127 = ~ _EVAL_199;
  assign _EVAL_96 = _EVAL_127[5:2];
  assign _EVAL_233 = _EVAL_14 <= 3'h4;
  assign _EVAL_51 = _EVAL_233 | _EVAL_8;
  assign _EVAL_113 = _EVAL_51 == 1'h0;
  assign _EVAL_64 = _EVAL_200 == 1'h0;
  assign _EVAL_91 = _EVAL_11 == 3'h1;
  assign _EVAL_184 = _EVAL_171 == 1'h0;
  assign _EVAL_202 = _EVAL == 3'h0;
  assign _EVAL_159 = _EVAL_177 == 1'h0;
  assign _EVAL_176 = _EVAL_159 | _EVAL_8;
  assign _EVAL_198 = _EVAL_176 == 1'h0;
  assign _EVAL_105 = _EVAL_7 == _EVAL_90;
  assign _EVAL_168 = _EVAL_105 | _EVAL_8;
  assign _EVAL_167 = _EVAL == 3'h2;
  assign _EVAL_118 = _EVAL_1 & _EVAL_187;
  assign _EVAL_227 = _EVAL_169 < plusarg_reader_out;
  assign _EVAL_84 = _EVAL_76 | _EVAL_227;
  assign _EVAL_237 = _EVAL_14 == _EVAL_86;
  assign _EVAL_106 = _EVAL_237 | _EVAL_8;
  assign _EVAL_131 = _EVAL_106 == 1'h0;
  assign _EVAL_143 = _EVAL_5 & _EVAL_202;
  assign _EVAL_32 = _EVAL_204 | _EVAL_224;
  assign _EVAL_70 = _EVAL_10 == _EVAL_142;
  assign _EVAL_99 = _EVAL_70 | _EVAL_8;
  assign _EVAL_218 = _EVAL_169 + 32'h1;
  assign _EVAL_48 = _EVAL_14 <= 3'h3;
  assign _EVAL_174 = _EVAL_48 | _EVAL_8;
  assign _EVAL_63 = _EVAL_174 == 1'h0;
  assign _EVAL_209 = _EVAL_84 | _EVAL_8;
  assign _EVAL_156 = _EVAL_209 == 1'h0;
  assign _EVAL_223 = _EVAL_1 & _EVAL_91;
  assign _EVAL_67 = ~ _EVAL_215;
  assign _EVAL_221 = _EVAL_13 & _EVAL_67;
  assign _EVAL_256 = _EVAL_0 == 1'h0;
  assign _EVAL_39 = _EVAL_3 >= 3'h2;
  assign _EVAL_158 = _EVAL_39 | _EVAL_8;
  assign _EVAL_161 = _EVAL_158 == 1'h0;
  assign _EVAL_163 = _EVAL_1 & _EVAL_61;
  assign _EVAL_74 = _EVAL_235 - 4'h1;
  assign _EVAL_35 = _EVAL_11 == 3'h0;
  assign _EVAL_241 = _EVAL_1 & _EVAL_35;
  assign _EVAL_173 = _EVAL_5 & _EVAL_167;
  assign _EVAL_153 = _EVAL_248 == 1'h0;
  assign _EVAL_56 = _EVAL == 3'h5;
  assign _EVAL_208 = _EVAL_37 == 1'h0;
  assign _EVAL_27 = _EVAL_228 == 1'h0;
  assign _EVAL_226 = _EVAL == _EVAL_149;
  assign _EVAL_95 = _EVAL_226 | _EVAL_8;
  assign _EVAL_179 = _EVAL_14 == 3'h0;
  assign _EVAL_104 = _EVAL_168 == 1'h0;
  assign _EVAL_107 = ~ _EVAL_83;
  assign _EVAL_25 = _EVAL_179 | _EVAL_8;
  assign _EVAL_40 = _EVAL == 3'h4;
  assign _EVAL_109 = _EVAL_5 & _EVAL_40;
  assign _EVAL_29 = _EVAL_10 <= 3'h2;
  assign _EVAL_160 = _EVAL_31 | _EVAL_8;
  assign _EVAL_245 = _EVAL_160 == 1'h0;
  assign _EVAL_225 = _EVAL_221 == 4'h0;
  assign _EVAL_144 = _EVAL_225 | _EVAL_8;
  assign _EVAL_229 = _EVAL_231 == 1'h0;
  assign _EVAL_175 = _EVAL_165 == 1'h0;
  assign _EVAL_191 = _EVAL_256 | _EVAL_8;
  assign _EVAL_45 = _EVAL_191 == 1'h0;
  assign _EVAL_232 = _EVAL_29 & _EVAL_49;
  assign _EVAL_117 = _EVAL == 3'h6;
  assign _EVAL_50 = _EVAL_5 & _EVAL_117;
  assign _EVAL_164 = _EVAL_242 | _EVAL_8;
  assign _EVAL_205 = _EVAL_25 == 1'h0;
  assign _EVAL_141 = _EVAL_32 & _EVAL_107;
  assign _EVAL_201 = _EVAL_72 | _EVAL_8;
  assign _EVAL_150 = _EVAL_201 == 1'h0;
  assign _EVAL_55 = _EVAL_95 == 1'h0;
  assign _EVAL_181 = _EVAL_232 | _EVAL_8;
  assign _EVAL_23 = _EVAL_181 == 1'h0;
  assign _EVAL_139 = _EVAL_11 == 3'h4;
  assign _EVAL_17 = _EVAL_164 == 1'h0;
  assign _EVAL_130 = _EVAL_144 == 1'h0;
  assign _EVAL_20 = _EVAL_46 & _EVAL_182;
  assign _EVAL_128 = _EVAL == 3'h7;
  assign _EVAL_58 = _EVAL_5 & _EVAL_128;
  assign _EVAL_124 = _EVAL_1 & _EVAL_139;
  assign _EVAL_166 = _EVAL_1 & _EVAL_239;
  assign _EVAL_44 = _EVAL_99 == 1'h0;
  assign _EVAL_116 = _EVAL_5 & _EVAL_56;
  assign _EVAL_195 = _EVAL_162 | _EVAL_46;
  assign _EVAL_16 = _EVAL_210 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_57 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_86 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_90 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_102 = _RAND_3[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_103 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_108 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_132 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_142 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_149 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_169 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_183 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_185 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_204 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_235 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_12) begin
    if (_EVAL_8) begin
      _EVAL_57 <= 4'h0;
    end else begin
      if (_EVAL_46) begin
        if (_EVAL_182) begin
          if (_EVAL_180) begin
            _EVAL_57 <= _EVAL_96;
          end else begin
            _EVAL_57 <= 4'h0;
          end
        end else begin
          _EVAL_57 <= _EVAL_249;
        end
      end
    end
    if (_EVAL_211) begin
      _EVAL_86 <= _EVAL_14;
    end
    if (_EVAL_211) begin
      _EVAL_90 <= _EVAL_7;
    end
    if (_EVAL_211) begin
      _EVAL_102 <= _EVAL_2;
    end
    if (_EVAL_20) begin
      _EVAL_103 <= _EVAL_11;
    end
    if (_EVAL_8) begin
      _EVAL_108 <= 4'h0;
    end else begin
      if (_EVAL_46) begin
        if (_EVAL_36) begin
          if (_EVAL_180) begin
            _EVAL_108 <= _EVAL_96;
          end else begin
            _EVAL_108 <= 4'h0;
          end
        end else begin
          _EVAL_108 <= _EVAL_19;
        end
      end
    end
    if (_EVAL_20) begin
      _EVAL_132 <= _EVAL_4;
    end
    if (_EVAL_211) begin
      _EVAL_142 <= _EVAL_10;
    end
    if (_EVAL_211) begin
      _EVAL_149 <= _EVAL;
    end
    if (_EVAL_8) begin
      _EVAL_169 <= 32'h0;
    end else begin
      if (_EVAL_195) begin
        _EVAL_169 <= 32'h0;
      end else begin
        _EVAL_169 <= _EVAL_218;
      end
    end
    if (_EVAL_20) begin
      _EVAL_183 <= _EVAL_3;
    end
    if (_EVAL_8) begin
      _EVAL_185 <= 4'h0;
    end else begin
      if (_EVAL_162) begin
        if (_EVAL_192) begin
          if (_EVAL_170) begin
            _EVAL_185 <= _EVAL_148;
          end else begin
            _EVAL_185 <= 4'h0;
          end
        end else begin
          _EVAL_185 <= _EVAL_60;
        end
      end
    end
    if (_EVAL_8) begin
      _EVAL_204 <= 8'h0;
    end else begin
      _EVAL_204 <= _EVAL_141;
    end
    if (_EVAL_8) begin
      _EVAL_235 <= 4'h0;
    end else begin
      if (_EVAL_162) begin
        if (_EVAL_89) begin
          if (_EVAL_170) begin
            _EVAL_235 <= _EVAL_148;
          end else begin
            _EVAL_235 <= 4'h0;
          end
        end else begin
          _EVAL_235 <= _EVAL_74;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8c5587c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59591d0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de9605c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80af9bb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5726930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ba66d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd800080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d71a284)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9b41b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8133a533)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b6c3250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a93168db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2066c729)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e80df3dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e30d0cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(857807db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cab3fbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(306c54fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41689fd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3f416fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4debc375)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6789e23d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fad7fcba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de4349b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4901c1cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddfce8f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23217040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0274f4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd5c5f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(219a1a8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c50c549)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f756129)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68294b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f47ac7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee6e8a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bc95d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7aa8fd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(414d7e91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9285b694)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4378e481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da6ea213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a24f530e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85d82508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2efb0383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42bf81ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62a0fbac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c67f00ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a30abcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5883d277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25e14a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84fadb87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8231b112)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e510268)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6389aeea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9ad0e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12d4ffe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c362178b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dd4cae7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c1b6f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d1c4a01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b50eac24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a86097e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81e7633a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cee9c7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1da8619)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(118f2e3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37d2d528)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb16395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(457d7a48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6582b998)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec264649)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(306f50d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
