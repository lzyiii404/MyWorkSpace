//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_226(
  input  [31:0] _EVAL,
  input  [31:0] _EVAL_0,
  output        _EVAL_1,
  input  [24:0] _EVAL_2,
  input  [2:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  output [1:0]  _EVAL_6,
  output [2:0]  _EVAL_7,
  output        _EVAL_8,
  output [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  output [31:0] _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  output [2:0]  _EVAL_17,
  input         _EVAL_18,
  output [2:0]  _EVAL_19,
  input  [6:0]  _EVAL_20,
  output [24:0] _EVAL_21,
  output [6:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  output        _EVAL_29,
  output [6:0]  _EVAL_30,
  input  [6:0]  _EVAL_31,
  input  [6:0]  _EVAL_32,
  output [2:0]  _EVAL_33,
  output        _EVAL_34,
  output [6:0]  _EVAL_35,
  output [3:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  output        _EVAL_38,
  output [3:0]  _EVAL_39,
  output [31:0] _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  output [24:0] _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output        _EVAL_46,
  output [31:0] _EVAL_47,
  input         _EVAL_48,
  input  [2:0]  _EVAL_49,
  input  [31:0] _EVAL_50
);
  reg  _EVAL_74;
  reg [31:0] _RAND_0;
  reg  _EVAL_78;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_99;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_140;
  reg [31:0] _RAND_3;
  wire  _EVAL_84;
  wire [1:0] _EVAL_64;
  wire [1:0] _EVAL_116;
  wire [1:0] _EVAL_93;
  wire [3:0] _EVAL_96;
  wire [2:0] _EVAL_97;
  wire [3:0] _EVAL_130;
  wire [3:0] _EVAL_60;
  wire [2:0] _EVAL_87;
  wire [3:0] _EVAL_100;
  wire [3:0] _EVAL_76;
  wire [3:0] _EVAL_56;
  wire [1:0] _EVAL_88;
  wire [1:0] _EVAL_72;
  wire [1:0] _EVAL_80;
  wire [1:0] _EVAL_115;
  wire  _EVAL_82;
  wire  _EVAL_68;
  wire [12:0] _EVAL_54;
  wire [5:0] _EVAL_92;
  wire [5:0] _EVAL_71;
  wire  _EVAL_112;
  wire  _EVAL_53;
  wire  _EVAL_131;
  wire  _EVAL_83;
  wire [49:0] _EVAL_58;
  wire [49:0] _EVAL_73;
  wire  _EVAL_123;
  wire  _EVAL_51;
  wire  _EVAL_108;
  wire  _EVAL_127;
  wire  _EVAL_134;
  wire  _EVAL_75;
  wire [3:0] _EVAL_62;
  wire [24:0] _EVAL_125;
  wire [25:0] _EVAL_111;
  wire [25:0] _EVAL_139;
  wire [25:0] _EVAL_128;
  wire  _EVAL_119;
  wire  _EVAL_136;
  wire  _EVAL_86;
  wire [12:0] _EVAL_89;
  wire [5:0] _EVAL_103;
  wire [5:0] _EVAL_65;
  wire [3:0] _EVAL_70;
  wire [3:0] _EVAL_137;
  wire [3:0] _EVAL_114;
  wire [49:0] _EVAL_81;
  wire  _EVAL_107;
  wire [1:0] _EVAL_129;
  wire [2:0] _EVAL_55;
  wire  _EVAL_106;
  wire [25:0] _EVAL_98;
  wire [25:0] _EVAL_94;
  wire [25:0] _EVAL_102;
  wire  _EVAL_122;
  wire  _EVAL_121;
  wire [3:0] _EVAL_91;
  wire [3:0] _EVAL_79;
  wire [3:0] _EVAL_138;
  wire [3:0] _EVAL_126;
  wire [3:0] _EVAL_105;
  wire  _EVAL_66;
  wire [49:0] _EVAL_67;
  wire [49:0] _EVAL_118;
  wire  _EVAL_101;
  wire  _EVAL_110;
  wire [1:0] _EVAL_69;
  wire [1:0] _EVAL_113;
  wire  _EVAL_63;
  assign _EVAL_84 = _EVAL_99 == 4'h0;
  assign _EVAL_64 = {_EVAL_44,_EVAL_42};
  assign _EVAL_116 = ~ _EVAL_140;
  assign _EVAL_93 = _EVAL_64 & _EVAL_116;
  assign _EVAL_96 = {_EVAL_93,_EVAL_44,_EVAL_42};
  assign _EVAL_97 = _EVAL_96[3:1];
  assign _EVAL_130 = {{1'd0}, _EVAL_97};
  assign _EVAL_60 = _EVAL_96 | _EVAL_130;
  assign _EVAL_87 = _EVAL_60[3:1];
  assign _EVAL_100 = {{1'd0}, _EVAL_87};
  assign _EVAL_76 = {_EVAL_140, 2'h0};
  assign _EVAL_56 = _EVAL_100 | _EVAL_76;
  assign _EVAL_88 = _EVAL_56[3:2];
  assign _EVAL_72 = _EVAL_56[1:0];
  assign _EVAL_80 = _EVAL_88 & _EVAL_72;
  assign _EVAL_115 = ~ _EVAL_80;
  assign _EVAL_82 = _EVAL_115[0];
  assign _EVAL_68 = _EVAL_84 ? _EVAL_82 : _EVAL_78;
  assign _EVAL_54 = 13'h3f << _EVAL_3;
  assign _EVAL_92 = _EVAL_54[5:0];
  assign _EVAL_71 = ~ _EVAL_92;
  assign _EVAL_112 = _EVAL_82 & _EVAL_42;
  assign _EVAL_53 = _EVAL_115[1];
  assign _EVAL_131 = _EVAL_53 & _EVAL_44;
  assign _EVAL_83 = _EVAL_84 ? _EVAL_112 : _EVAL_78;
  assign _EVAL_58 = {_EVAL_23,2'h0,_EVAL_3,_EVAL_20,2'h0,_EVAL_50,1'h0};
  assign _EVAL_73 = _EVAL_83 ? _EVAL_58 : 50'h0;
  assign _EVAL_123 = _EVAL_42 | _EVAL_44;
  assign _EVAL_51 = _EVAL_78 ? _EVAL_42 : 1'h0;
  assign _EVAL_108 = _EVAL_74 ? _EVAL_44 : 1'h0;
  assign _EVAL_127 = _EVAL_51 | _EVAL_108;
  assign _EVAL_134 = _EVAL_84 ? _EVAL_123 : _EVAL_127;
  assign _EVAL_75 = _EVAL_10 & _EVAL_134;
  assign _EVAL_62 = {{3'd0}, _EVAL_75};
  assign _EVAL_125 = _EVAL_2 ^ 25'h100000;
  assign _EVAL_111 = {1'b0,$signed(_EVAL_125)};
  assign _EVAL_139 = $signed(_EVAL_111) & $signed(26'sh100000);
  assign _EVAL_128 = $signed(_EVAL_139);
  assign _EVAL_119 = $signed(_EVAL_128) == $signed(26'sh0);
  assign _EVAL_136 = _EVAL_119 ? _EVAL_18 : 1'h0;
  assign _EVAL_86 = _EVAL_49[0];
  assign _EVAL_89 = 13'h3f << _EVAL_5;
  assign _EVAL_103 = _EVAL_89[5:0];
  assign _EVAL_65 = ~ _EVAL_103;
  assign _EVAL_70 = _EVAL_65[5:2];
  assign _EVAL_137 = _EVAL_86 ? _EVAL_70 : 4'h0;
  assign _EVAL_114 = _EVAL_131 ? _EVAL_137 : 4'h0;
  assign _EVAL_81 = {_EVAL_49,2'h0,_EVAL_5,_EVAL_32,2'h0,_EVAL,1'h0};
  assign _EVAL_107 = _EVAL_84 ? _EVAL_53 : _EVAL_74;
  assign _EVAL_129 = _EVAL_115 & _EVAL_64;
  assign _EVAL_55 = {_EVAL_129, 1'h0};
  assign _EVAL_106 = _EVAL_84 & _EVAL_10;
  assign _EVAL_98 = {1'b0,$signed(_EVAL_2)};
  assign _EVAL_94 = $signed(_EVAL_98) & $signed(26'sh100000);
  assign _EVAL_102 = $signed(_EVAL_94);
  assign _EVAL_122 = $signed(_EVAL_102) == $signed(26'sh0);
  assign _EVAL_121 = _EVAL_23[0];
  assign _EVAL_91 = _EVAL_71[5:2];
  assign _EVAL_79 = _EVAL_121 ? _EVAL_91 : 4'h0;
  assign _EVAL_138 = _EVAL_112 ? _EVAL_79 : 4'h0;
  assign _EVAL_126 = _EVAL_138 | _EVAL_114;
  assign _EVAL_105 = _EVAL_99 - _EVAL_62;
  assign _EVAL_66 = _EVAL_84 ? _EVAL_131 : _EVAL_74;
  assign _EVAL_67 = _EVAL_66 ? _EVAL_81 : 50'h0;
  assign _EVAL_118 = _EVAL_73 | _EVAL_67;
  assign _EVAL_101 = _EVAL_64 != 2'h0;
  assign _EVAL_110 = _EVAL_106 & _EVAL_101;
  assign _EVAL_69 = _EVAL_55[1:0];
  assign _EVAL_113 = _EVAL_129 | _EVAL_69;
  assign _EVAL_63 = _EVAL_122 ? _EVAL_48 : 1'h0;
  assign _EVAL_17 = _EVAL_11;
  assign _EVAL_39 = _EVAL_16;
  assign _EVAL_24 = _EVAL_118[34];
  assign _EVAL_19 = _EVAL_11;
  assign _EVAL_36 = _EVAL_16;
  assign _EVAL_13 = _EVAL_118[0];
  assign _EVAL_30 = _EVAL_31;
  assign _EVAL_40 = _EVAL_0;
  assign _EVAL_37 = _EVAL_28;
  assign _EVAL_12 = _EVAL_10 & _EVAL_68;
  assign _EVAL_21 = _EVAL_2;
  assign _EVAL_38 = _EVAL_27 & _EVAL_119;
  assign _EVAL_35 = _EVAL_31;
  assign _EVAL_6 = _EVAL_118[46:45];
  assign _EVAL_41 = _EVAL_63 | _EVAL_136;
  assign _EVAL_47 = _EVAL_0;
  assign _EVAL_29 = _EVAL_45;
  assign _EVAL_8 = _EVAL_118[33];
  assign _EVAL_14 = _EVAL_118[32:1];
  assign _EVAL_46 = _EVAL_27 & _EVAL_122;
  assign _EVAL_1 = _EVAL_84 ? _EVAL_123 : _EVAL_127;
  assign _EVAL_43 = _EVAL_2;
  assign _EVAL_4 = _EVAL_25;
  assign _EVAL_7 = _EVAL_28;
  assign _EVAL_33 = _EVAL_118[44:42];
  assign _EVAL_34 = _EVAL_10 & _EVAL_107;
  assign _EVAL_9 = _EVAL_118[49:47];
  assign _EVAL_22 = _EVAL_118[41:35];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_74 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_78 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_99 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_140 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_26) begin
    if (_EVAL_15) begin
      _EVAL_74 <= 1'h0;
    end else begin
      if (_EVAL_84) begin
        _EVAL_74 <= _EVAL_131;
      end
    end
    if (_EVAL_15) begin
      _EVAL_78 <= 1'h0;
    end else begin
      if (_EVAL_84) begin
        _EVAL_78 <= _EVAL_112;
      end
    end
    if (_EVAL_15) begin
      _EVAL_99 <= 4'h0;
    end else begin
      if (_EVAL_106) begin
        _EVAL_99 <= _EVAL_126;
      end else begin
        _EVAL_99 <= _EVAL_105;
      end
    end
    if (_EVAL_15) begin
      _EVAL_140 <= 2'h3;
    end else begin
      if (_EVAL_110) begin
        _EVAL_140 <= _EVAL_113;
      end
    end
  end
endmodule
