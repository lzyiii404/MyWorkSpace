//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_256_assert(
  input        _EVAL,
  input        _EVAL_2,
  input        _EVAL_4,
  input        _EVAL_5,
  input        _EVAL_7,
  input        _EVAL_8,
  input  [1:0] _EVAL_9,
  input        _EVAL_10,
  input        _EVAL_11,
  input        _EVAL_14,
  input        _EVAL_17,
  input        _EVAL_18,
  input  [1:0] _EVAL_21,
  input        _EVAL_23,
  input  [1:0] _EVAL_24,
  input        _EVAL_25,
  input        _EVAL_26,
  input        _EVAL_28,
  input        _EVAL_29,
  input        _EVAL_30,
  input        _EVAL_31,
  input        _EVAL_32,
  input  [1:0] _EVAL_34,
  input        _EVAL_35,
  input        _EVAL_36,
  input        _EVAL_38,
  input  [1:0] _EVAL_39,
  input        _EVAL_40,
  input  [1:0] _EVAL_41,
  input  [1:0] _EVAL_44,
  input        _EVAL_45,
  input        _EVAL_46,
  input        _EVAL_47,
  input        _EVAL_50,
  input        _EVAL_51,
  input        _EVAL_52,
  input        _EVAL_53,
  input  [1:0] _EVAL_54,
  input        _EVAL_55,
  input        _EVAL_58,
  input        _EVAL_59,
  input        _EVAL_60,
  input        _EVAL_85,
  input        _EVAL_333,
  input        _EVAL_358,
  input        _EVAL_266,
  input        _EVAL_161,
  input        _EVAL_283,
  input        _EVAL_376,
  input        _EVAL_160,
  input        _EVAL_293,
  input        _EVAL_253,
  input        _EVAL_203,
  input        _EVAL_303,
  input        _EVAL_310,
  input        _EVAL_338,
  input        _EVAL_352,
  input        _EVAL_285
);
  wire  _EVAL_189;
  wire  _EVAL_195;
  wire [2:0] _EVAL_75;
  wire  _EVAL_304;
  wire  _EVAL_234;
  wire  _EVAL_181;
  wire  _EVAL_325;
  wire [2:0] _EVAL_101;
  wire  _EVAL_120;
  wire [2:0] _EVAL_246;
  wire  _EVAL_104;
  wire [2:0] _EVAL_371;
  wire  _EVAL_364;
  wire [2:0] _EVAL_164;
  wire  _EVAL_277;
  wire  _EVAL_135;
  wire  _EVAL_172;
  wire  _EVAL_309;
  wire  _EVAL_198;
  wire  _EVAL_136;
  wire  _EVAL_206;
  wire  _EVAL_330;
  wire  _EVAL_257;
  wire  _EVAL_240;
  wire  _EVAL_93;
  wire  _EVAL_275;
  wire  _EVAL_186;
  wire  _EVAL_67;
  wire  _EVAL_347;
  wire  _EVAL_61;
  wire  _EVAL_157;
  wire  _EVAL_344;
  wire  _EVAL_134;
  wire  _EVAL_268;
  wire  _EVAL_342;
  wire  _EVAL_115;
  wire  _EVAL_138;
  wire  _EVAL_386;
  wire  _EVAL_383;
  wire  _EVAL_175;
  wire  _EVAL_81;
  wire [2:0] _EVAL_305;
  wire  _EVAL_350;
  wire  _EVAL_291;
  wire  _EVAL_256;
  wire  _EVAL_121;
  wire  _EVAL_355;
  wire  _EVAL_216;
  wire  _EVAL_308;
  wire  _EVAL_90;
  wire  _EVAL_95;
  wire  _EVAL_340;
  wire  _EVAL_262;
  wire  _EVAL_77;
  wire  _EVAL_194;
  wire  _EVAL_224;
  wire  _EVAL_375;
  wire  _EVAL_367;
  wire  _EVAL_307;
  wire  _EVAL_79;
  wire  _EVAL_382;
  wire [2:0] _EVAL_370;
  wire  _EVAL_132;
  wire  _EVAL_173;
  wire  _EVAL_239;
  wire  _EVAL_324;
  wire  _EVAL_165;
  wire  _EVAL_379;
  wire  _EVAL_141;
  wire  _EVAL_221;
  wire  _EVAL_166;
  wire  _EVAL_232;
  wire  _EVAL_247;
  wire  _EVAL_236;
  wire [2:0] _EVAL_129;
  wire  _EVAL_295;
  wire  _EVAL_200;
  wire  _EVAL_150;
  wire  _EVAL_255;
  wire  _EVAL_182;
  wire  _EVAL_226;
  wire  _EVAL_177;
  wire  _EVAL_299;
  wire  _EVAL_149;
  wire  _EVAL_201;
  wire  _EVAL_243;
  wire  _EVAL_292;
  wire  _EVAL_328;
  wire  _EVAL_204;
  wire  _EVAL_271;
  wire  _EVAL_248;
  wire  _EVAL_152;
  wire  _EVAL_123;
  wire  _EVAL_139;
  wire  _EVAL_167;
  wire  _EVAL_335;
  wire  _EVAL_214;
  wire  _EVAL_158;
  wire  _EVAL_74;
  wire  _EVAL_89;
  wire  _EVAL_332;
  wire  _EVAL_159;
  wire  _EVAL_279;
  wire  _EVAL_127;
  wire  _EVAL_106;
  wire  _EVAL_196;
  wire  _EVAL_220;
  wire  _EVAL_361;
  wire  _EVAL_112;
  wire  _EVAL_137;
  wire  _EVAL_289;
  wire  _EVAL_100;
  wire  _EVAL_341;
  wire  _EVAL_385;
  wire  _EVAL_171;
  wire  _EVAL_103;
  wire  _EVAL_296;
  wire  _EVAL_318;
  wire  _EVAL_133;
  wire  _EVAL_345;
  wire  _EVAL_306;
  wire  _EVAL_66;
  wire  _EVAL_209;
  wire  _EVAL_119;
  wire  _EVAL_265;
  wire  _EVAL_128;
  wire  _EVAL_92;
  wire  _EVAL_249;
  wire  _EVAL_144;
  wire  _EVAL_331;
  wire  _EVAL_117;
  wire  _EVAL_238;
  wire  _EVAL_346;
  wire  _EVAL_282;
  wire  _EVAL_187;
  wire  _EVAL_110;
  wire  _EVAL_228;
  wire  _EVAL_301;
  wire  _EVAL_380;
  wire  _EVAL_87;
  wire  _EVAL_348;
  wire  _EVAL_197;
  wire  _EVAL_174;
  wire  _EVAL_96;
  wire  _EVAL_300;
  wire  _EVAL_319;
  wire  _EVAL_192;
  wire  _EVAL_365;
  wire  _EVAL_337;
  wire  _EVAL_235;
  wire  _EVAL_327;
  wire  _EVAL_208;
  wire  _EVAL_199;
  wire  _EVAL_264;
  wire  _EVAL_176;
  wire  _EVAL_278;
  wire  _EVAL_180;
  wire  _EVAL_102;
  wire  _EVAL_178;
  wire  _EVAL_351;
  wire  _EVAL_65;
  assign _EVAL_189 = _EVAL_39 == 2'h0;
  assign _EVAL_195 = _EVAL_34 == 2'h2;
  assign _EVAL_75 = {_EVAL_2,_EVAL_58,_EVAL_51};
  assign _EVAL_304 = _EVAL_75 == 3'h3;
  assign _EVAL_234 = _EVAL_9 == 2'h3;
  assign _EVAL_181 = _EVAL_24 == 2'h0;
  assign _EVAL_325 = _EVAL_39 == 2'h2;
  assign _EVAL_101 = {_EVAL_7,_EVAL_10,_EVAL_14};
  assign _EVAL_120 = _EVAL_101 == 3'h1;
  assign _EVAL_246 = {_EVAL_38,_EVAL_23,_EVAL};
  assign _EVAL_104 = _EVAL_246 == 3'h0;
  assign _EVAL_371 = {_EVAL_17,_EVAL_50,_EVAL_5};
  assign _EVAL_364 = _EVAL_371 == 3'h5;
  assign _EVAL_164 = {_EVAL_29,_EVAL_40,_EVAL_8};
  assign _EVAL_277 = _EVAL_164 == 3'h4;
  assign _EVAL_135 = _EVAL_24 == 2'h1;
  assign _EVAL_172 = _EVAL_39 == 2'h1;
  assign _EVAL_309 = _EVAL_41 == 2'h3;
  assign _EVAL_198 = _EVAL_60 & _EVAL_333;
  assign _EVAL_136 = _EVAL_34 == 2'h3;
  assign _EVAL_206 = _EVAL_198 & _EVAL_136;
  assign _EVAL_330 = _EVAL_54 == 2'h3;
  assign _EVAL_257 = _EVAL_55 & _EVAL_160;
  assign _EVAL_240 = _EVAL_253 == 1'h0;
  assign _EVAL_93 = _EVAL_240 & _EVAL_333;
  assign _EVAL_275 = _EVAL_161 == 1'h0;
  assign _EVAL_186 = _EVAL_275 & _EVAL_266;
  assign _EVAL_67 = _EVAL_44 == 2'h3;
  assign _EVAL_347 = _EVAL_186 & _EVAL_67;
  assign _EVAL_61 = _EVAL_303 == 1'h0;
  assign _EVAL_157 = _EVAL_61 & _EVAL_203;
  assign _EVAL_344 = _EVAL_164 == 3'h0;
  assign _EVAL_134 = _EVAL_4 & _EVAL_266;
  assign _EVAL_268 = _EVAL_134 & _EVAL_67;
  assign _EVAL_342 = _EVAL_44 == 2'h0;
  assign _EVAL_115 = _EVAL_85 == 1'h0;
  assign _EVAL_138 = _EVAL_115 & _EVAL_285;
  assign _EVAL_386 = _EVAL_138 & _EVAL_330;
  assign _EVAL_383 = _EVAL_44 == 2'h1;
  assign _EVAL_175 = _EVAL_186 & _EVAL_383;
  assign _EVAL_81 = _EVAL_41 == 2'h1;
  assign _EVAL_305 = {_EVAL_28,_EVAL_52,_EVAL_30};
  assign _EVAL_350 = _EVAL_338 == 1'h0;
  assign _EVAL_291 = _EVAL_350 & _EVAL_310;
  assign _EVAL_256 = _EVAL_21 == 2'h1;
  assign _EVAL_121 = _EVAL_291 & _EVAL_256;
  assign _EVAL_355 = _EVAL_358 == 1'h0;
  assign _EVAL_216 = _EVAL_355 & _EVAL_352;
  assign _EVAL_308 = _EVAL_9 == 2'h1;
  assign _EVAL_90 = _EVAL_216 & _EVAL_308;
  assign _EVAL_95 = _EVAL_75 == 3'h1;
  assign _EVAL_340 = _EVAL_21 == 2'h3;
  assign _EVAL_262 = _EVAL_41 == 2'h0;
  assign _EVAL_77 = _EVAL_75 == 3'h7;
  assign _EVAL_194 = _EVAL_305 == 3'h3;
  assign _EVAL_224 = _EVAL_53 & _EVAL_203;
  assign _EVAL_375 = _EVAL_224 & _EVAL_309;
  assign _EVAL_367 = _EVAL_21 == 2'h0;
  assign _EVAL_307 = _EVAL_36 & _EVAL_285;
  assign _EVAL_79 = _EVAL_34 == 2'h1;
  assign _EVAL_382 = _EVAL_198 & _EVAL_79;
  assign _EVAL_370 = {_EVAL_32,_EVAL_47,_EVAL_25};
  assign _EVAL_132 = _EVAL_370 == 3'h1;
  assign _EVAL_173 = _EVAL_75 == 3'h5;
  assign _EVAL_239 = _EVAL_164 == 3'h1;
  assign _EVAL_324 = _EVAL_246 == 3'h3;
  assign _EVAL_165 = _EVAL_18 == 1'h0;
  assign _EVAL_379 = _EVAL_371 == 3'h7;
  assign _EVAL_141 = _EVAL_21 == 2'h2;
  assign _EVAL_221 = _EVAL_376 == 1'h0;
  assign _EVAL_166 = _EVAL_221 & _EVAL_283;
  assign _EVAL_232 = _EVAL_24 == 2'h3;
  assign _EVAL_247 = _EVAL_166 & _EVAL_232;
  assign _EVAL_236 = _EVAL_93 & _EVAL_79;
  assign _EVAL_129 = {_EVAL_11,_EVAL_46,_EVAL_26};
  assign _EVAL_295 = _EVAL_129 == 3'h7;
  assign _EVAL_200 = _EVAL_291 & _EVAL_340;
  assign _EVAL_150 = _EVAL_370 == 3'h3;
  assign _EVAL_255 = _EVAL_45 & _EVAL_352;
  assign _EVAL_182 = _EVAL_255 & _EVAL_308;
  assign _EVAL_226 = _EVAL_293 == 1'h0;
  assign _EVAL_177 = _EVAL_226 & _EVAL_160;
  assign _EVAL_299 = _EVAL_129 == 3'h3;
  assign _EVAL_149 = _EVAL_93 & _EVAL_136;
  assign _EVAL_201 = _EVAL_41 == 2'h2;
  assign _EVAL_243 = _EVAL_305 == 3'h7;
  assign _EVAL_292 = _EVAL_224 & _EVAL_201;
  assign _EVAL_328 = _EVAL_157 & _EVAL_201;
  assign _EVAL_204 = _EVAL_44 == 2'h2;
  assign _EVAL_271 = _EVAL_186 & _EVAL_204;
  assign _EVAL_248 = _EVAL_134 & _EVAL_383;
  assign _EVAL_152 = _EVAL_291 & _EVAL_141;
  assign _EVAL_123 = _EVAL_59 & _EVAL_283;
  assign _EVAL_139 = _EVAL_123 & _EVAL_232;
  assign _EVAL_167 = _EVAL_129 == 3'h4;
  assign _EVAL_335 = _EVAL_224 & _EVAL_81;
  assign _EVAL_214 = _EVAL_35 & _EVAL_310;
  assign _EVAL_158 = _EVAL_370 == 3'h4;
  assign _EVAL_74 = _EVAL_214 & _EVAL_340;
  assign _EVAL_89 = _EVAL_101 == 3'h7;
  assign _EVAL_332 = _EVAL_371 == 3'h4;
  assign _EVAL_159 = _EVAL_101 == 3'h5;
  assign _EVAL_279 = _EVAL_54 == 2'h2;
  assign _EVAL_127 = _EVAL_54 == 2'h1;
  assign _EVAL_106 = _EVAL_138 & _EVAL_127;
  assign _EVAL_196 = _EVAL_129 == 3'h0;
  assign _EVAL_220 = _EVAL_307 & _EVAL_279;
  assign _EVAL_361 = _EVAL_75 == 3'h0;
  assign _EVAL_112 = _EVAL_54 == 2'h0;
  assign _EVAL_137 = _EVAL_134 & _EVAL_204;
  assign _EVAL_289 = _EVAL_138 & _EVAL_279;
  assign _EVAL_100 = _EVAL_164 == 3'h5;
  assign _EVAL_341 = _EVAL_39 == 2'h3;
  assign _EVAL_385 = _EVAL_257 & _EVAL_341;
  assign _EVAL_171 = _EVAL_164 == 3'h7;
  assign _EVAL_103 = _EVAL_371 == 3'h1;
  assign _EVAL_296 = _EVAL_370 == 3'h0;
  assign _EVAL_318 = _EVAL_75 == 3'h4;
  assign _EVAL_133 = _EVAL_257 & _EVAL_172;
  assign _EVAL_345 = _EVAL_255 & _EVAL_234;
  assign _EVAL_306 = _EVAL_129 == 3'h1;
  assign _EVAL_66 = _EVAL_370 == 3'h7;
  assign _EVAL_209 = _EVAL_216 & _EVAL_234;
  assign _EVAL_119 = _EVAL_9 == 2'h0;
  assign _EVAL_265 = _EVAL_24 == 2'h2;
  assign _EVAL_128 = _EVAL_166 & _EVAL_265;
  assign _EVAL_92 = _EVAL_9 == 2'h2;
  assign _EVAL_249 = _EVAL_305 == 3'h1;
  assign _EVAL_144 = _EVAL_198 & _EVAL_195;
  assign _EVAL_331 = _EVAL_305 == 3'h4;
  assign _EVAL_117 = _EVAL_246 == 3'h4;
  assign _EVAL_238 = _EVAL_214 & _EVAL_256;
  assign _EVAL_346 = _EVAL_371 == 3'h0;
  assign _EVAL_282 = _EVAL_157 & _EVAL_81;
  assign _EVAL_187 = _EVAL_255 & _EVAL_92;
  assign _EVAL_110 = _EVAL_370 == 3'h5;
  assign _EVAL_228 = _EVAL_166 & _EVAL_135;
  assign _EVAL_301 = _EVAL_129 == 3'h5;
  assign _EVAL_380 = _EVAL_101 == 3'h4;
  assign _EVAL_87 = _EVAL_371 == 3'h3;
  assign _EVAL_348 = _EVAL_305 == 3'h0;
  assign _EVAL_197 = _EVAL_214 & _EVAL_141;
  assign _EVAL_174 = _EVAL_257 & _EVAL_325;
  assign _EVAL_96 = _EVAL_177 & _EVAL_325;
  assign _EVAL_300 = _EVAL_305 == 3'h5;
  assign _EVAL_319 = _EVAL_307 & _EVAL_330;
  assign _EVAL_192 = _EVAL_216 & _EVAL_92;
  assign _EVAL_365 = _EVAL_164 == 3'h3;
  assign _EVAL_337 = _EVAL_123 & _EVAL_265;
  assign _EVAL_235 = _EVAL_101 == 3'h0;
  assign _EVAL_327 = _EVAL_246 == 3'h7;
  assign _EVAL_208 = _EVAL_177 & _EVAL_172;
  assign _EVAL_199 = _EVAL_101 == 3'h3;
  assign _EVAL_264 = _EVAL_307 & _EVAL_127;
  assign _EVAL_176 = _EVAL_246 == 3'h1;
  assign _EVAL_278 = _EVAL_93 & _EVAL_195;
  assign _EVAL_180 = _EVAL_157 & _EVAL_309;
  assign _EVAL_102 = _EVAL_246 == 3'h5;
  assign _EVAL_178 = _EVAL_123 & _EVAL_135;
  assign _EVAL_351 = _EVAL_177 & _EVAL_341;
  assign _EVAL_65 = _EVAL_34 == 2'h0;
  always @(posedge _EVAL_31) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_379 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_332 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_327 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_351 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_348 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
