//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_126_assert(
  input  [2:0]  _EVAL,
  input  [1:0]  _EVAL_0,
  input  [6:0]  _EVAL_1,
  input  [6:0]  _EVAL_2,
  input         _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [13:0] _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_33;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_77;
  reg [31:0] _RAND_1;
  reg [72:0] _EVAL_89;
  reg [95:0] _RAND_2;
  reg [5:0] _EVAL_105;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_110;
  reg [31:0] _RAND_4;
  reg [13:0] _EVAL_115;
  reg [31:0] _RAND_5;
  reg [5:0] _EVAL_124;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_147;
  reg [31:0] _RAND_7;
  reg [5:0] _EVAL_152;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_163;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_169;
  reg [31:0] _RAND_10;
  reg [6:0] _EVAL_196;
  reg [31:0] _RAND_11;
  reg [3:0] _EVAL_197;
  reg [31:0] _RAND_12;
  reg  _EVAL_245;
  reg [31:0] _RAND_13;
  reg [31:0] _EVAL_259;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_298;
  reg [31:0] _RAND_15;
  reg [1:0] _EVAL_312;
  reg [31:0] _RAND_16;
  wire [72:0] _EVAL_230;
  wire  _EVAL_87;
  wire  _EVAL_194;
  wire  _EVAL_182;
  wire  _EVAL_116;
  wire [127:0] _EVAL_60;
  wire [127:0] _EVAL_246;
  wire [72:0] _EVAL_248;
  wire [72:0] _EVAL_125;
  wire [22:0] _EVAL_261;
  wire [3:0] _EVAL_291;
  wire  _EVAL_69;
  wire  _EVAL_64;
  wire  _EVAL_256;
  wire  _EVAL_43;
  wire  _EVAL_242;
  wire  _EVAL_146;
  wire  _EVAL_192;
  wire  _EVAL_305;
  wire  _EVAL_222;
  wire  _EVAL_20;
  wire  _EVAL_243;
  wire [22:0] _EVAL_94;
  wire [7:0] _EVAL_320;
  wire [7:0] _EVAL_302;
  wire [5:0] _EVAL_181;
  wire [5:0] _EVAL_287;
  wire  _EVAL_244;
  wire  _EVAL_53;
  wire  _EVAL_283;
  wire  _EVAL_106;
  wire  _EVAL_97;
  wire  _EVAL_167;
  wire  _EVAL_206;
  wire  _EVAL_257;
  wire  _EVAL_203;
  wire  _EVAL_91;
  wire  _EVAL_314;
  wire [1:0] _EVAL_299;
  wire [1:0] _EVAL_85;
  wire  _EVAL_156;
  wire  _EVAL_131;
  wire  _EVAL_216;
  wire  _EVAL_95;
  wire  _EVAL_195;
  wire  _EVAL_276;
  wire  _EVAL_325;
  wire [72:0] _EVAL_272;
  wire [72:0] _EVAL_63;
  wire  _EVAL_129;
  wire  _EVAL_311;
  wire  _EVAL_268;
  wire  _EVAL_46;
  wire [5:0] _EVAL_293;
  wire  _EVAL_285;
  wire  _EVAL_112;
  wire  _EVAL_211;
  wire  _EVAL_126;
  wire  _EVAL_19;
  wire  _EVAL_187;
  wire  _EVAL_120;
  wire  _EVAL_258;
  wire  _EVAL_149;
  wire  _EVAL_29;
  wire  _EVAL_317;
  wire [127:0] _EVAL_153;
  wire [127:0] _EVAL_238;
  wire  _EVAL_253;
  wire  _EVAL_81;
  wire  _EVAL_193;
  wire  _EVAL_40;
  wire  _EVAL_186;
  wire  _EVAL_260;
  wire  _EVAL_321;
  wire  _EVAL_67;
  wire  _EVAL_212;
  wire  _EVAL_247;
  wire  _EVAL_183;
  wire  _EVAL_290;
  wire  _EVAL_301;
  wire  _EVAL_21;
  wire  _EVAL_76;
  wire [3:0] _EVAL_159;
  wire  _EVAL_318;
  wire  _EVAL_315;
  wire [5:0] _EVAL_136;
  wire  _EVAL_171;
  wire  _EVAL_62;
  wire  _EVAL_72;
  wire  _EVAL_22;
  wire  _EVAL_143;
  wire  _EVAL_31;
  wire  _EVAL_172;
  wire  _EVAL_34;
  wire  _EVAL_270;
  wire  _EVAL_179;
  wire  _EVAL_191;
  wire  _EVAL_284;
  wire  _EVAL_188;
  wire  _EVAL_265;
  wire  _EVAL_239;
  wire  _EVAL_226;
  wire  _EVAL_264;
  wire [72:0] _EVAL_304;
  wire  _EVAL_83;
  wire  _EVAL_310;
  wire  _EVAL_263;
  wire  _EVAL_164;
  wire  _EVAL_84;
  wire [13:0] _EVAL_48;
  wire [14:0] _EVAL_58;
  wire [14:0] _EVAL_173;
  wire [14:0] _EVAL_41;
  wire  _EVAL_27;
  wire  _EVAL_223;
  wire  _EVAL_300;
  wire  _EVAL_213;
  wire  _EVAL_128;
  wire  _EVAL_56;
  wire  _EVAL_93;
  wire  _EVAL_30;
  wire  _EVAL_117;
  wire  _EVAL_205;
  wire  _EVAL_113;
  wire  _EVAL_49;
  wire  _EVAL_208;
  wire  _EVAL_119;
  wire  _EVAL_249;
  wire [3:0] _EVAL_55;
  wire  _EVAL_78;
  wire  _EVAL_54;
  wire [3:0] _EVAL_36;
  wire  _EVAL_151;
  wire [2:0] _EVAL_286;
  wire  _EVAL_38;
  wire  _EVAL_237;
  wire  _EVAL_80;
  wire  _EVAL_199;
  wire  _EVAL_303;
  wire  _EVAL_24;
  wire  _EVAL_234;
  wire  _EVAL_109;
  wire  _EVAL_219;
  wire [7:0] _EVAL_319;
  wire [7:0] _EVAL_32;
  wire [5:0] _EVAL_88;
  wire  _EVAL_292;
  wire  _EVAL_133;
  wire  _EVAL_296;
  wire  _EVAL_65;
  wire [2:0] _EVAL_184;
  wire  _EVAL_100;
  wire  _EVAL_154;
  wire  _EVAL_254;
  wire  _EVAL_150;
  wire  _EVAL_228;
  wire  _EVAL_86;
  wire [72:0] _EVAL_289;
  wire [72:0] _EVAL_103;
  wire [3:0] _EVAL_224;
  wire [3:0] _EVAL_274;
  wire  _EVAL_90;
  wire  _EVAL_231;
  wire  _EVAL_59;
  wire  _EVAL_70;
  wire  _EVAL_50;
  wire [13:0] _EVAL_209;
  wire  _EVAL_178;
  wire  _EVAL_130;
  wire  _EVAL_104;
  wire  _EVAL_297;
  wire  _EVAL_225;
  wire  _EVAL_207;
  wire  _EVAL_176;
  wire  _EVAL_139;
  wire  _EVAL_267;
  wire  _EVAL_39;
  wire  _EVAL_107;
  wire  _EVAL_294;
  wire [31:0] _EVAL_134;
  wire  _EVAL_210;
  wire  _EVAL_162;
  wire  _EVAL_57;
  wire  _EVAL_215;
  wire  _EVAL_316;
  wire  _EVAL_266;
  wire  _EVAL_190;
  wire  _EVAL_144;
  wire  _EVAL_148;
  wire  _EVAL_278;
  wire  _EVAL_170;
  wire  _EVAL_280;
  wire  _EVAL_240;
  wire  _EVAL_79;
  wire  _EVAL_111;
  wire  _EVAL_204;
  wire  _EVAL_96;
  wire  _EVAL_141;
  wire  _EVAL_44;
  wire  _EVAL_160;
  wire  _EVAL_108;
  wire  _EVAL_137;
  wire  _EVAL_326;
  wire  _EVAL_166;
  wire  _EVAL_140;
  wire  _EVAL_168;
  wire  _EVAL_123;
  wire  _EVAL_189;
  wire  _EVAL_101;
  wire  _EVAL_98;
  wire  _EVAL_324;
  wire  _EVAL_229;
  wire  _EVAL_175;
  wire  _EVAL_165;
  wire  _EVAL_271;
  wire  _EVAL_118;
  wire [13:0] _EVAL_295;
  wire  _EVAL_127;
  wire  _EVAL_217;
  wire  _EVAL_73;
  wire  _EVAL_180;
  wire  _EVAL_102;
  wire  _EVAL_232;
  wire  _EVAL_51;
  wire  _EVAL_233;
  wire  _EVAL_61;
  wire  _EVAL_308;
  wire  _EVAL_52;
  wire [5:0] _EVAL_275;
  wire  _EVAL_281;
  wire  _EVAL_251;
  wire  _EVAL_198;
  wire  _EVAL_221;
  wire  _EVAL_177;
  wire  _EVAL_45;
  wire  _EVAL_200;
  wire  _EVAL_25;
  wire  _EVAL_82;
  wire  _EVAL_47;
  wire  _EVAL_218;
  wire  _EVAL_250;
  wire  _EVAL_161;
  wire  _EVAL_174;
  wire  _EVAL_202;
  wire  _EVAL_121;
  wire  _EVAL_307;
  wire  _EVAL_66;
  wire  _EVAL_235;
  wire  _EVAL_313;
  wire  _EVAL_306;
  wire  _EVAL_323;
  wire  _EVAL_99;
  wire  _EVAL_42;
  wire  _EVAL_74;
  wire  _EVAL_155;
  wire  _EVAL_322;
  wire  _EVAL_28;
  wire  _EVAL_309;
  wire  _EVAL_269;
  wire  _EVAL_273;
  wire  _EVAL_220;
  wire  _EVAL_138;
  wire  _EVAL_185;
  wire  _EVAL_122;
  wire  _EVAL_114;
  wire  _EVAL_23;
  wire  _EVAL_201;
  wire  _EVAL_92;
  wire  _EVAL_132;
  wire  _EVAL_68;
  wire  _EVAL_241;
  wire  _EVAL_288;
  wire  _EVAL_277;
  wire  _EVAL_135;
  wire  _EVAL_71;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_230 = _EVAL_89 >> _EVAL_2;
  assign _EVAL_87 = _EVAL_230[0];
  assign _EVAL_194 = _EVAL_6 & _EVAL_14;
  assign _EVAL_182 = _EVAL_105 == 6'h0;
  assign _EVAL_116 = _EVAL_194 & _EVAL_182;
  assign _EVAL_60 = 128'h1 << _EVAL_2;
  assign _EVAL_246 = _EVAL_116 ? _EVAL_60 : 128'h0;
  assign _EVAL_248 = _EVAL_246[72:0];
  assign _EVAL_125 = _EVAL_89 | _EVAL_248;
  assign _EVAL_261 = 23'hff << _EVAL_18;
  assign _EVAL_291 = ~ _EVAL_4;
  assign _EVAL_69 = _EVAL_291 == 4'h0;
  assign _EVAL_64 = _EVAL_69 | _EVAL_5;
  assign _EVAL_256 = _EVAL_64 == 1'h0;
  assign _EVAL_43 = _EVAL_1 == 7'h48;
  assign _EVAL_242 = _EVAL_1 == 7'h40;
  assign _EVAL_146 = _EVAL_43 | _EVAL_242;
  assign _EVAL_192 = _EVAL_13 == 3'h3;
  assign _EVAL_305 = _EVAL_124 == 6'h0;
  assign _EVAL_222 = _EVAL_194 & _EVAL_305;
  assign _EVAL_20 = _EVAL_163 == 6'h0;
  assign _EVAL_243 = _EVAL[0];
  assign _EVAL_94 = 23'hff << _EVAL_7;
  assign _EVAL_320 = _EVAL_94[7:0];
  assign _EVAL_302 = ~ _EVAL_320;
  assign _EVAL_181 = _EVAL_302[7:2];
  assign _EVAL_287 = _EVAL_163 - 6'h1;
  assign _EVAL_244 = _EVAL_0 == 2'h0;
  assign _EVAL_53 = _EVAL_244 | _EVAL_5;
  assign _EVAL_283 = _EVAL_9 != 3'h0;
  assign _EVAL_106 = _EVAL_283 | _EVAL_5;
  assign _EVAL_97 = _EVAL_248 != 73'h0;
  assign _EVAL_167 = _EVAL_9 <= 3'h4;
  assign _EVAL_206 = _EVAL_12 == _EVAL_115;
  assign _EVAL_257 = _EVAL_206 | _EVAL_5;
  assign _EVAL_203 = _EVAL_0 <= 2'h2;
  assign _EVAL_91 = _EVAL_203 | _EVAL_5;
  assign _EVAL_314 = _EVAL_18[0];
  assign _EVAL_299 = 2'h1 << _EVAL_314;
  assign _EVAL_85 = _EVAL_299 | 2'h1;
  assign _EVAL_156 = _EVAL_85[0];
  assign _EVAL_131 = _EVAL_12[1];
  assign _EVAL_216 = _EVAL_131 == 1'h0;
  assign _EVAL_95 = _EVAL_12[0];
  assign _EVAL_195 = _EVAL_95 == 1'h0;
  assign _EVAL_276 = _EVAL_216 & _EVAL_195;
  assign _EVAL_325 = _EVAL_156 & _EVAL_276;
  assign _EVAL_272 = _EVAL_248 | _EVAL_89;
  assign _EVAL_63 = _EVAL_272 >> _EVAL_1;
  assign _EVAL_129 = _EVAL_63[0];
  assign _EVAL_311 = _EVAL_129 | _EVAL_5;
  assign _EVAL_268 = _EVAL_311 == 1'h0;
  assign _EVAL_46 = _EVAL == 3'h5;
  assign _EVAL_293 = _EVAL_105 - 6'h1;
  assign _EVAL_285 = _EVAL_18 >= 4'h2;
  assign _EVAL_112 = _EVAL_85[1];
  assign _EVAL_211 = _EVAL_112 & _EVAL_216;
  assign _EVAL_126 = _EVAL_285 | _EVAL_211;
  assign _EVAL_19 = _EVAL_305 == 1'h0;
  assign _EVAL_187 = _EVAL_14 & _EVAL_19;
  assign _EVAL_120 = _EVAL_8 & _EVAL_11;
  assign _EVAL_258 = _EVAL_120 & _EVAL_20;
  assign _EVAL_149 = _EVAL == 3'h6;
  assign _EVAL_29 = _EVAL_149 == 1'h0;
  assign _EVAL_317 = _EVAL_258 & _EVAL_29;
  assign _EVAL_153 = 128'h1 << _EVAL_1;
  assign _EVAL_238 = _EVAL_317 ? _EVAL_153 : 128'h0;
  assign _EVAL_253 = _EVAL == _EVAL_298;
  assign _EVAL_81 = _EVAL_253 | _EVAL_5;
  assign _EVAL_193 = _EVAL_81 == 1'h0;
  assign _EVAL_40 = _EVAL_131 & _EVAL_195;
  assign _EVAL_186 = _EVAL_156 & _EVAL_40;
  assign _EVAL_260 = _EVAL_112 & _EVAL_131;
  assign _EVAL_321 = _EVAL_285 | _EVAL_260;
  assign _EVAL_67 = _EVAL_321 | _EVAL_186;
  assign _EVAL_212 = _EVAL_131 & _EVAL_95;
  assign _EVAL_247 = _EVAL_156 & _EVAL_212;
  assign _EVAL_183 = _EVAL_321 | _EVAL_247;
  assign _EVAL_290 = _EVAL_216 & _EVAL_95;
  assign _EVAL_301 = _EVAL_156 & _EVAL_290;
  assign _EVAL_21 = _EVAL_126 | _EVAL_301;
  assign _EVAL_76 = _EVAL_126 | _EVAL_325;
  assign _EVAL_159 = {_EVAL_183,_EVAL_67,_EVAL_21,_EVAL_76};
  assign _EVAL_318 = _EVAL_2 == 7'h40;
  assign _EVAL_315 = _EVAL_18 <= 4'h2;
  assign _EVAL_136 = _EVAL_124 - 6'h1;
  assign _EVAL_171 = _EVAL_4 == _EVAL_159;
  assign _EVAL_62 = _EVAL_171 | _EVAL_5;
  assign _EVAL_72 = _EVAL_62 == 1'h0;
  assign _EVAL_22 = _EVAL_13 == 3'h0;
  assign _EVAL_143 = _EVAL_14 & _EVAL_22;
  assign _EVAL_31 = _EVAL_106 == 1'h0;
  assign _EVAL_172 = _EVAL_89 != 73'h0;
  assign _EVAL_34 = _EVAL_172 == 1'h0;
  assign _EVAL_270 = plusarg_reader_out == 32'h0;
  assign _EVAL_179 = _EVAL_34 | _EVAL_270;
  assign _EVAL_191 = _EVAL_259 < plusarg_reader_out;
  assign _EVAL_284 = _EVAL_179 | _EVAL_191;
  assign _EVAL_188 = _EVAL_13 == 3'h2;
  assign _EVAL_265 = _EVAL_14 & _EVAL_188;
  assign _EVAL_239 = _EVAL_15 == 1'h0;
  assign _EVAL_226 = _EVAL_239 | _EVAL_5;
  assign _EVAL_264 = _EVAL_226 == 1'h0;
  assign _EVAL_304 = _EVAL_238[72:0];
  assign _EVAL_83 = _EVAL_248 != _EVAL_304;
  assign _EVAL_310 = _EVAL_97 == 1'h0;
  assign _EVAL_263 = _EVAL_83 | _EVAL_310;
  assign _EVAL_164 = _EVAL_13 == 3'h4;
  assign _EVAL_84 = _EVAL_14 & _EVAL_164;
  assign _EVAL_48 = _EVAL_12 ^ 14'h3000;
  assign _EVAL_58 = {1'b0,$signed(_EVAL_48)};
  assign _EVAL_173 = $signed(_EVAL_58) & $signed(-15'sh1000);
  assign _EVAL_41 = $signed(_EVAL_173);
  assign _EVAL_27 = _EVAL_9 <= 3'h3;
  assign _EVAL_223 = _EVAL_7 == _EVAL_197;
  assign _EVAL_300 = _EVAL_223 | _EVAL_5;
  assign _EVAL_213 = _EVAL_300 == 1'h0;
  assign _EVAL_128 = _EVAL_17 == _EVAL_33;
  assign _EVAL_56 = _EVAL_128 | _EVAL_5;
  assign _EVAL_93 = _EVAL_56 == 1'h0;
  assign _EVAL_30 = _EVAL_15 == _EVAL_245;
  assign _EVAL_117 = $signed(_EVAL_41) == $signed(15'sh0);
  assign _EVAL_205 = _EVAL_315 & _EVAL_117;
  assign _EVAL_113 = _EVAL_205 | _EVAL_5;
  assign _EVAL_49 = _EVAL_9 == _EVAL_147;
  assign _EVAL_208 = _EVAL_49 | _EVAL_5;
  assign _EVAL_119 = _EVAL_13 == 3'h5;
  assign _EVAL_249 = _EVAL_14 & _EVAL_119;
  assign _EVAL_55 = _EVAL_2[6:3];
  assign _EVAL_78 = _EVAL_55 == 4'h1;
  assign _EVAL_54 = _EVAL_13[2];
  assign _EVAL_36 = _EVAL_1[6:3];
  assign _EVAL_151 = _EVAL_36 == 4'h8;
  assign _EVAL_286 = _EVAL_1[2:0];
  assign _EVAL_38 = 3'h1 <= _EVAL_286;
  assign _EVAL_237 = _EVAL_151 & _EVAL_38;
  assign _EVAL_80 = _EVAL_146 | _EVAL_237;
  assign _EVAL_199 = _EVAL_1 == 7'h20;
  assign _EVAL_303 = _EVAL_80 | _EVAL_199;
  assign _EVAL_24 = _EVAL_36 == 4'h0;
  assign _EVAL_234 = _EVAL_303 | _EVAL_24;
  assign _EVAL_109 = _EVAL_36 == 4'h1;
  assign _EVAL_219 = _EVAL_234 | _EVAL_109;
  assign _EVAL_319 = _EVAL_261[7:0];
  assign _EVAL_32 = ~ _EVAL_319;
  assign _EVAL_88 = _EVAL_32[7:2];
  assign _EVAL_292 = _EVAL_152 == 6'h0;
  assign _EVAL_133 = _EVAL_292 == 1'h0;
  assign _EVAL_296 = _EVAL_11 & _EVAL_133;
  assign _EVAL_65 = _EVAL_9 == 3'h0;
  assign _EVAL_184 = _EVAL_2[2:0];
  assign _EVAL_100 = 3'h1 <= _EVAL_184;
  assign _EVAL_154 = _EVAL_30 | _EVAL_5;
  assign _EVAL_254 = _EVAL_154 == 1'h0;
  assign _EVAL_150 = _EVAL_87 == 1'h0;
  assign _EVAL_228 = _EVAL_150 | _EVAL_5;
  assign _EVAL_86 = _EVAL == 3'h1;
  assign _EVAL_289 = ~ _EVAL_304;
  assign _EVAL_103 = _EVAL_125 & _EVAL_289;
  assign _EVAL_224 = ~ _EVAL_159;
  assign _EVAL_274 = _EVAL_4 & _EVAL_224;
  assign _EVAL_90 = _EVAL_274 == 4'h0;
  assign _EVAL_231 = _EVAL_90 | _EVAL_5;
  assign _EVAL_59 = _EVAL_9 <= 3'h2;
  assign _EVAL_70 = _EVAL_208 == 1'h0;
  assign _EVAL_50 = _EVAL_2 == 7'h48;
  assign _EVAL_209 = {{6'd0}, _EVAL_32};
  assign _EVAL_178 = _EVAL_2 == _EVAL_77;
  assign _EVAL_130 = _EVAL_178 | _EVAL_5;
  assign _EVAL_104 = _EVAL_13 == _EVAL_169;
  assign _EVAL_297 = _EVAL_104 | _EVAL_5;
  assign _EVAL_225 = _EVAL_18 <= 4'h8;
  assign _EVAL_207 = _EVAL_225 & _EVAL_117;
  assign _EVAL_176 = _EVAL_207 | _EVAL_5;
  assign _EVAL_139 = _EVAL_176 == 1'h0;
  assign _EVAL_267 = _EVAL_53 == 1'h0;
  assign _EVAL_39 = _EVAL == 3'h4;
  assign _EVAL_107 = _EVAL_11 & _EVAL_39;
  assign _EVAL_294 = _EVAL_194 | _EVAL_120;
  assign _EVAL_134 = _EVAL_259 + 32'h1;
  assign _EVAL_210 = _EVAL_11 & _EVAL_149;
  assign _EVAL_162 = _EVAL_55 == 4'h0;
  assign _EVAL_57 = _EVAL_167 | _EVAL_5;
  assign _EVAL_215 = _EVAL == 3'h2;
  assign _EVAL_316 = _EVAL_11 & _EVAL_215;
  assign _EVAL_266 = _EVAL_10 == 1'h0;
  assign _EVAL_190 = _EVAL_239 | _EVAL_3;
  assign _EVAL_144 = _EVAL_5 == 1'h0;
  assign _EVAL_148 = _EVAL_266 | _EVAL_5;
  assign _EVAL_278 = _EVAL_148 == 1'h0;
  assign _EVAL_170 = _EVAL_54 == 1'h0;
  assign _EVAL_280 = _EVAL_3 == 1'h0;
  assign _EVAL_240 = _EVAL_280 | _EVAL_5;
  assign _EVAL_79 = _EVAL_11 & _EVAL_86;
  assign _EVAL_111 = _EVAL == 3'h0;
  assign _EVAL_204 = _EVAL_55 == 4'h8;
  assign _EVAL_96 = _EVAL_204 & _EVAL_100;
  assign _EVAL_141 = _EVAL_11 & _EVAL_111;
  assign _EVAL_44 = _EVAL_7 >= 4'h2;
  assign _EVAL_160 = _EVAL_44 | _EVAL_5;
  assign _EVAL_108 = _EVAL_36 == 4'h2;
  assign _EVAL_137 = _EVAL_1 == _EVAL_196;
  assign _EVAL_326 = _EVAL_137 | _EVAL_5;
  assign _EVAL_166 = _EVAL_326 == 1'h0;
  assign _EVAL_140 = _EVAL_50 | _EVAL_318;
  assign _EVAL_168 = _EVAL_140 | _EVAL_96;
  assign _EVAL_123 = _EVAL_2 == 7'h20;
  assign _EVAL_189 = _EVAL_168 | _EVAL_123;
  assign _EVAL_101 = _EVAL_189 | _EVAL_162;
  assign _EVAL_98 = _EVAL_219 | _EVAL_108;
  assign _EVAL_324 = _EVAL_36 == 4'h3;
  assign _EVAL_229 = _EVAL_98 | _EVAL_324;
  assign _EVAL_175 = _EVAL_229 | _EVAL_5;
  assign _EVAL_165 = _EVAL_175 == 1'h0;
  assign _EVAL_271 = _EVAL_284 | _EVAL_5;
  assign _EVAL_118 = _EVAL_271 == 1'h0;
  assign _EVAL_295 = _EVAL_12 & _EVAL_209;
  assign _EVAL_127 = _EVAL_295 == 14'h0;
  assign _EVAL_217 = _EVAL <= 3'h6;
  assign _EVAL_73 = _EVAL_27 | _EVAL_5;
  assign _EVAL_180 = _EVAL_13 == 3'h1;
  assign _EVAL_102 = _EVAL_14 & _EVAL_180;
  assign _EVAL_232 = 4'h6 == _EVAL_18;
  assign _EVAL_51 = _EVAL_318 ? _EVAL_232 : 1'h0;
  assign _EVAL_233 = _EVAL_51 | _EVAL_5;
  assign _EVAL_61 = _EVAL_233 == 1'h0;
  assign _EVAL_308 = _EVAL_263 | _EVAL_5;
  assign _EVAL_52 = _EVAL_308 == 1'h0;
  assign _EVAL_275 = _EVAL_152 - 6'h1;
  assign _EVAL_281 = _EVAL_113 == 1'h0;
  assign _EVAL_251 = _EVAL_18 == _EVAL_110;
  assign _EVAL_198 = _EVAL_251 | _EVAL_5;
  assign _EVAL_221 = _EVAL_127 | _EVAL_5;
  assign _EVAL_177 = _EVAL_221 == 1'h0;
  assign _EVAL_45 = _EVAL_13 == 3'h6;
  assign _EVAL_200 = _EVAL_14 & _EVAL_45;
  assign _EVAL_25 = _EVAL_14 & _EVAL_192;
  assign _EVAL_82 = _EVAL_285 | _EVAL_5;
  assign _EVAL_47 = _EVAL_82 == 1'h0;
  assign _EVAL_218 = _EVAL_101 | _EVAL_78;
  assign _EVAL_250 = _EVAL_55 == 4'h2;
  assign _EVAL_161 = _EVAL_218 | _EVAL_250;
  assign _EVAL_174 = _EVAL_55 == 4'h3;
  assign _EVAL_202 = _EVAL_161 | _EVAL_174;
  assign _EVAL_121 = _EVAL_202 | _EVAL_5;
  assign _EVAL_307 = _EVAL_91 == 1'h0;
  assign _EVAL_66 = _EVAL_217 | _EVAL_5;
  assign _EVAL_235 = _EVAL_66 == 1'h0;
  assign _EVAL_313 = _EVAL_0 != 2'h2;
  assign _EVAL_306 = _EVAL_313 | _EVAL_5;
  assign _EVAL_323 = _EVAL_306 == 1'h0;
  assign _EVAL_99 = _EVAL_190 | _EVAL_5;
  assign _EVAL_42 = _EVAL_65 | _EVAL_5;
  assign _EVAL_74 = _EVAL_231 == 1'h0;
  assign _EVAL_155 = _EVAL_13 == 3'h7;
  assign _EVAL_322 = _EVAL_14 & _EVAL_155;
  assign _EVAL_28 = _EVAL_160 == 1'h0;
  assign _EVAL_309 = _EVAL_257 == 1'h0;
  assign _EVAL_269 = _EVAL_0 == _EVAL_312;
  assign _EVAL_273 = _EVAL_269 | _EVAL_5;
  assign _EVAL_220 = _EVAL_273 == 1'h0;
  assign _EVAL_138 = _EVAL_297 == 1'h0;
  assign _EVAL_185 = _EVAL_228 == 1'h0;
  assign _EVAL_122 = _EVAL_73 == 1'h0;
  assign _EVAL_114 = _EVAL_42 == 1'h0;
  assign _EVAL_23 = _EVAL_59 | _EVAL_5;
  assign _EVAL_201 = _EVAL_130 == 1'h0;
  assign _EVAL_92 = _EVAL_57 == 1'h0;
  assign _EVAL_132 = _EVAL_121 == 1'h0;
  assign _EVAL_68 = _EVAL_240 == 1'h0;
  assign _EVAL_241 = _EVAL_198 == 1'h0;
  assign _EVAL_288 = _EVAL_23 == 1'h0;
  assign _EVAL_277 = _EVAL_120 & _EVAL_292;
  assign _EVAL_135 = _EVAL_99 == 1'h0;
  assign _EVAL_71 = _EVAL_11 & _EVAL_46;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_33 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_77 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {3{`RANDOM}};
  _EVAL_89 = _RAND_2[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_105 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_110 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_115 = _RAND_5[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_124 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_147 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_152 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_163 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_169 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_196 = _RAND_11[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_197 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_245 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_259 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_298 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_312 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_16) begin
    if (_EVAL_277) begin
      _EVAL_33 <= _EVAL_17;
    end
    if (_EVAL_222) begin
      _EVAL_77 <= _EVAL_2;
    end
    if (_EVAL_5) begin
      _EVAL_89 <= 73'h0;
    end else begin
      _EVAL_89 <= _EVAL_103;
    end
    if (_EVAL_5) begin
      _EVAL_105 <= 6'h0;
    end else begin
      if (_EVAL_194) begin
        if (_EVAL_182) begin
          if (_EVAL_170) begin
            _EVAL_105 <= _EVAL_88;
          end else begin
            _EVAL_105 <= 6'h0;
          end
        end else begin
          _EVAL_105 <= _EVAL_293;
        end
      end
    end
    if (_EVAL_222) begin
      _EVAL_110 <= _EVAL_18;
    end
    if (_EVAL_222) begin
      _EVAL_115 <= _EVAL_12;
    end
    if (_EVAL_5) begin
      _EVAL_124 <= 6'h0;
    end else begin
      if (_EVAL_194) begin
        if (_EVAL_305) begin
          if (_EVAL_170) begin
            _EVAL_124 <= _EVAL_88;
          end else begin
            _EVAL_124 <= 6'h0;
          end
        end else begin
          _EVAL_124 <= _EVAL_136;
        end
      end
    end
    if (_EVAL_222) begin
      _EVAL_147 <= _EVAL_9;
    end
    if (_EVAL_5) begin
      _EVAL_152 <= 6'h0;
    end else begin
      if (_EVAL_120) begin
        if (_EVAL_292) begin
          if (_EVAL_243) begin
            _EVAL_152 <= _EVAL_181;
          end else begin
            _EVAL_152 <= 6'h0;
          end
        end else begin
          _EVAL_152 <= _EVAL_275;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_163 <= 6'h0;
    end else begin
      if (_EVAL_120) begin
        if (_EVAL_20) begin
          if (_EVAL_243) begin
            _EVAL_163 <= _EVAL_181;
          end else begin
            _EVAL_163 <= 6'h0;
          end
        end else begin
          _EVAL_163 <= _EVAL_287;
        end
      end
    end
    if (_EVAL_222) begin
      _EVAL_169 <= _EVAL_13;
    end
    if (_EVAL_277) begin
      _EVAL_196 <= _EVAL_1;
    end
    if (_EVAL_277) begin
      _EVAL_197 <= _EVAL_7;
    end
    if (_EVAL_277) begin
      _EVAL_245 <= _EVAL_15;
    end
    if (_EVAL_5) begin
      _EVAL_259 <= 32'h0;
    end else begin
      if (_EVAL_294) begin
        _EVAL_259 <= 32'h0;
      end else begin
        _EVAL_259 <= _EVAL_134;
      end
    end
    if (_EVAL_277) begin
      _EVAL_298 <= _EVAL;
    end
    if (_EVAL_277) begin
      _EVAL_312 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(471ba33d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d232913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d398eaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57f7545d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df4c00ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(937068bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b50caba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f651189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2930aba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(708c9fe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d02e68bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee375ff1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5233168)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad8dc383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9348a325)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30621e8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f2e4121)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7da939a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e860007c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d795dc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(646062f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67929e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5563580d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3edcba7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41cf0556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83c61105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98b3f668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d70b7d97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(564d0655)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e5baa13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa0b94c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2019c04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caf05452)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67aa57ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88f53481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(166739c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(976b1268)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3525c5b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dd172f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b12b301)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44fe41e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e777df2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb5fc1d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a53f61b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fbdc3ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d51b018)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb2e49fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(944d44b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dbb9561)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19815436)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87d8e2ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d254b540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b6fe31e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f34954)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a333c51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a56852ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cef74e88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f7a294)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(384eae72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(584d0121)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b532d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53c8ec31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baaec57a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d783e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebc8cb29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1600c2bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fbe1c06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6134c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4b75863)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(302f661f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d21f7cc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c8d6394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c137914d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(701c56fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7c33f10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0fc0687)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f06f559c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4df494b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2efa1692)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f69eff3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(480f3a53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cffee1c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37d7335)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(732f2697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8e653e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80117d38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75418224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac1ef2ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8619de0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14fce006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
