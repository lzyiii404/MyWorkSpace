//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_150_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input  [6:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input  [6:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [24:0] _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [6:0] _EVAL_26;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_43;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_50;
  reg [31:0] _RAND_3;
  reg [24:0] _EVAL_55;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_67;
  reg [31:0] _RAND_5;
  reg  _EVAL_82;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_116;
  reg [31:0] _RAND_7;
  reg  _EVAL_125;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_179;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_224;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_232;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_252;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_298;
  reg [31:0] _RAND_13;
  reg [72:0] _EVAL_308;
  reg [95:0] _RAND_14;
  reg [3:0] _EVAL_315;
  reg [31:0] _RAND_15;
  reg [6:0] _EVAL_323;
  reg [31:0] _RAND_16;
  wire  _EVAL_311;
  wire  _EVAL_299;
  wire [1:0] _EVAL_132;
  wire [1:0] _EVAL_56;
  wire  _EVAL_75;
  wire  _EVAL_233;
  wire  _EVAL_61;
  wire  _EVAL_230;
  wire  _EVAL_133;
  wire  _EVAL_248;
  wire  _EVAL_135;
  wire  _EVAL_181;
  wire  _EVAL_207;
  wire  _EVAL_36;
  wire  _EVAL_282;
  wire  _EVAL_205;
  wire [24:0] _EVAL_326;
  wire [25:0] _EVAL_57;
  wire  _EVAL_115;
  wire  _EVAL_62;
  wire  _EVAL_153;
  wire  _EVAL_296;
  wire  _EVAL_301;
  wire  _EVAL_72;
  wire [3:0] _EVAL_316;
  wire  _EVAL_264;
  wire [2:0] _EVAL_145;
  wire  _EVAL_76;
  wire  _EVAL_168;
  wire  _EVAL_297;
  wire  _EVAL_210;
  wire  _EVAL_49;
  wire  _EVAL_198;
  wire  _EVAL_280;
  wire  _EVAL_226;
  wire  _EVAL_63;
  wire  _EVAL_29;
  wire  _EVAL_107;
  wire  _EVAL_177;
  wire  _EVAL_141;
  wire  _EVAL_262;
  wire  _EVAL_74;
  wire  _EVAL_220;
  wire  _EVAL_175;
  wire  _EVAL_314;
  wire  _EVAL_212;
  wire  _EVAL_184;
  wire  _EVAL_28;
  wire  _EVAL_113;
  wire  _EVAL_152;
  wire [12:0] _EVAL_173;
  wire  _EVAL_186;
  wire [24:0] _EVAL_204;
  wire [25:0] _EVAL_209;
  wire [25:0] _EVAL_165;
  wire [25:0] _EVAL_201;
  wire  _EVAL_257;
  wire [25:0] _EVAL_254;
  wire [25:0] _EVAL_250;
  wire  _EVAL_274;
  wire  _EVAL_247;
  wire  _EVAL_243;
  wire  _EVAL_219;
  wire  _EVAL_35;
  wire  _EVAL_39;
  wire  _EVAL_223;
  wire  _EVAL_304;
  wire  _EVAL_244;
  wire  _EVAL_196;
  wire  _EVAL_24;
  wire  _EVAL_249;
  wire [3:0] _EVAL_89;
  wire  _EVAL_40;
  wire  _EVAL_126;
  wire  _EVAL_193;
  wire  _EVAL_265;
  wire  _EVAL_288;
  wire  _EVAL_42;
  wire  _EVAL_120;
  wire  _EVAL_53;
  wire [3:0] _EVAL_300;
  wire  _EVAL_48;
  wire  _EVAL_279;
  wire  _EVAL_134;
  wire  _EVAL_138;
  wire  _EVAL_70;
  wire  _EVAL_189;
  wire [127:0] _EVAL_237;
  wire [127:0] _EVAL_157;
  wire [72:0] _EVAL_142;
  wire  _EVAL_234;
  wire  _EVAL_216;
  wire  _EVAL_222;
  wire  _EVAL_266;
  wire  _EVAL_229;
  wire  _EVAL_228;
  wire  _EVAL_97;
  wire  _EVAL_172;
  wire  _EVAL_148;
  wire  _EVAL_45;
  wire  _EVAL_136;
  wire [2:0] _EVAL_51;
  wire  _EVAL_290;
  wire  _EVAL_20;
  wire  _EVAL_114;
  wire  _EVAL_65;
  wire  _EVAL_215;
  wire  _EVAL_30;
  wire  _EVAL_161;
  wire  _EVAL_86;
  wire  _EVAL_122;
  wire  _EVAL_276;
  wire  _EVAL_236;
  wire  _EVAL_218;
  wire [5:0] _EVAL_146;
  wire [5:0] _EVAL_149;
  wire [3:0] _EVAL_278;
  wire [3:0] _EVAL_174;
  wire [72:0] _EVAL_199;
  wire  _EVAL_259;
  wire  _EVAL_211;
  wire  _EVAL_103;
  wire  _EVAL_270;
  wire  _EVAL_46;
  wire [127:0] _EVAL_33;
  wire [127:0] _EVAL_267;
  wire [72:0] _EVAL_90;
  wire [72:0] _EVAL_183;
  wire [72:0] _EVAL_128;
  wire [72:0] _EVAL_263;
  wire [72:0] _EVAL_52;
  wire  _EVAL_69;
  wire  _EVAL_214;
  wire  _EVAL_98;
  wire  _EVAL_291;
  wire  _EVAL_41;
  wire  _EVAL_144;
  wire  _EVAL_292;
  wire  _EVAL_318;
  wire  _EVAL_167;
  wire  _EVAL_130;
  wire  _EVAL_150;
  wire  _EVAL_225;
  wire  _EVAL_191;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_112;
  wire  _EVAL_307;
  wire  _EVAL_242;
  wire  _EVAL_221;
  wire  _EVAL_281;
  wire  _EVAL_213;
  wire  _EVAL_241;
  wire [12:0] _EVAL_64;
  wire [5:0] _EVAL_151;
  wire [5:0] _EVAL_71;
  wire [3:0] _EVAL_38;
  wire [3:0] _EVAL_255;
  wire  _EVAL_185;
  wire  _EVAL_235;
  wire  _EVAL_169;
  wire  _EVAL_245;
  wire  _EVAL_124;
  wire  _EVAL_83;
  wire  _EVAL_104;
  wire  _EVAL_246;
  wire  _EVAL_277;
  wire  _EVAL_319;
  wire  _EVAL_143;
  wire  _EVAL_27;
  wire  _EVAL_162;
  wire  _EVAL_85;
  wire  _EVAL_272;
  wire  _EVAL_295;
  wire  _EVAL_129;
  wire [31:0] _EVAL_127;
  wire [3:0] _EVAL_154;
  wire  _EVAL_139;
  wire  _EVAL_190;
  wire [72:0] _EVAL_118;
  wire  _EVAL_59;
  wire  _EVAL_310;
  wire  _EVAL_95;
  wire  _EVAL_159;
  wire  _EVAL_147;
  wire  _EVAL_66;
  wire  _EVAL_155;
  wire  _EVAL_88;
  wire [24:0] _EVAL_92;
  wire [24:0] _EVAL_171;
  wire  _EVAL_325;
  wire  _EVAL_324;
  wire  _EVAL_294;
  wire  _EVAL_111;
  wire  _EVAL_322;
  wire  _EVAL_187;
  wire  _EVAL_268;
  wire  _EVAL_188;
  wire  _EVAL_25;
  wire  _EVAL_289;
  wire  _EVAL_331;
  wire  _EVAL_121;
  wire  _EVAL_275;
  wire  _EVAL_321;
  wire  _EVAL_178;
  wire  _EVAL_117;
  wire  _EVAL_313;
  wire  _EVAL_96;
  wire  _EVAL_239;
  wire  _EVAL_156;
  wire  _EVAL_87;
  wire  _EVAL_269;
  wire  _EVAL_192;
  wire  _EVAL_284;
  wire  _EVAL_105;
  wire  _EVAL_78;
  wire  _EVAL_195;
  wire  _EVAL_197;
  wire  _EVAL_286;
  wire  _EVAL_320;
  wire  _EVAL_100;
  wire  _EVAL_312;
  wire  _EVAL_37;
  wire [3:0] _EVAL_80;
  wire  _EVAL_176;
  wire  _EVAL_160;
  wire  _EVAL_332;
  wire  _EVAL_271;
  wire  _EVAL_253;
  wire  _EVAL_327;
  wire  _EVAL_21;
  wire  _EVAL_106;
  wire  _EVAL_293;
  wire  _EVAL_158;
  wire  _EVAL_260;
  wire  _EVAL_328;
  wire  _EVAL_206;
  wire  _EVAL_273;
  wire  _EVAL_170;
  wire  _EVAL_164;
  wire  _EVAL_203;
  wire  _EVAL_285;
  wire  _EVAL_231;
  wire  _EVAL_60;
  wire [3:0] _EVAL_22;
  wire [3:0] _EVAL_110;
  wire  _EVAL_309;
  wire  _EVAL_317;
  wire  _EVAL_99;
  wire  _EVAL_305;
  wire  _EVAL_238;
  wire  _EVAL_194;
  wire  _EVAL_44;
  wire  _EVAL_261;
  wire  _EVAL_23;
  wire [3:0] _EVAL_108;
  wire  _EVAL_329;
  wire  _EVAL_287;
  wire  _EVAL_227;
  wire  _EVAL_202;
  wire  _EVAL_180;
  wire  _EVAL_163;
  wire  _EVAL_251;
  wire  _EVAL_182;
  wire  _EVAL_109;
  wire  _EVAL_73;
  wire  _EVAL_101;
  wire  _EVAL_137;
  wire  _EVAL_306;
  wire  _EVAL_47;
  wire  _EVAL_166;
  wire  _EVAL_68;
  wire  _EVAL_102;
  wire  _EVAL_217;
  wire  _EVAL_19;
  wire  _EVAL_84;
  wire  _EVAL_140;
  wire  _EVAL_81;
  wire  _EVAL_256;
  wire  _EVAL_91;
  wire  _EVAL_119;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_311 = _EVAL_5 >= 3'h2;
  assign _EVAL_299 = _EVAL_5[0];
  assign _EVAL_132 = 2'h1 << _EVAL_299;
  assign _EVAL_56 = _EVAL_132 | 2'h1;
  assign _EVAL_75 = _EVAL_56[1];
  assign _EVAL_233 = _EVAL_16[1];
  assign _EVAL_61 = _EVAL_233 == 1'h0;
  assign _EVAL_230 = _EVAL_75 & _EVAL_61;
  assign _EVAL_133 = _EVAL_311 | _EVAL_230;
  assign _EVAL_248 = _EVAL_56[0];
  assign _EVAL_135 = _EVAL_16[0];
  assign _EVAL_181 = _EVAL_61 & _EVAL_135;
  assign _EVAL_207 = _EVAL_248 & _EVAL_181;
  assign _EVAL_36 = _EVAL_133 | _EVAL_207;
  assign _EVAL_282 = _EVAL_116 == 4'h0;
  assign _EVAL_205 = _EVAL_13 == _EVAL_26;
  assign _EVAL_326 = _EVAL_16 ^ 25'h1900000;
  assign _EVAL_57 = {1'b0,$signed(_EVAL_326)};
  assign _EVAL_115 = _EVAL_11 <= 2'h2;
  assign _EVAL_62 = _EVAL_115 | _EVAL_8;
  assign _EVAL_153 = _EVAL_62 == 1'h0;
  assign _EVAL_296 = _EVAL_2 == 7'h48;
  assign _EVAL_301 = _EVAL_2 == 7'h40;
  assign _EVAL_72 = _EVAL_296 | _EVAL_301;
  assign _EVAL_316 = _EVAL_2[6:3];
  assign _EVAL_264 = _EVAL_316 == 4'h8;
  assign _EVAL_145 = _EVAL_2[2:0];
  assign _EVAL_76 = 3'h1 <= _EVAL_145;
  assign _EVAL_168 = _EVAL_264 & _EVAL_76;
  assign _EVAL_297 = _EVAL_72 | _EVAL_168;
  assign _EVAL_210 = _EVAL_2 == 7'h20;
  assign _EVAL_49 = _EVAL_297 | _EVAL_210;
  assign _EVAL_198 = _EVAL_316 == 4'h0;
  assign _EVAL_280 = _EVAL_49 | _EVAL_198;
  assign _EVAL_226 = _EVAL_316 == 4'h1;
  assign _EVAL_63 = _EVAL_280 | _EVAL_226;
  assign _EVAL_29 = _EVAL_316 == 4'h2;
  assign _EVAL_107 = _EVAL_63 | _EVAL_29;
  assign _EVAL_177 = _EVAL_316 == 4'h3;
  assign _EVAL_141 = _EVAL_107 | _EVAL_177;
  assign _EVAL_262 = _EVAL_141 | _EVAL_8;
  assign _EVAL_74 = _EVAL_262 == 1'h0;
  assign _EVAL_220 = _EVAL_3 == _EVAL_82;
  assign _EVAL_175 = _EVAL_220 | _EVAL_8;
  assign _EVAL_314 = _EVAL_6 == 3'h1;
  assign _EVAL_212 = _EVAL_9 & _EVAL_314;
  assign _EVAL_184 = _EVAL_308 != 73'h0;
  assign _EVAL_28 = _EVAL_184 == 1'h0;
  assign _EVAL_113 = plusarg_reader_out == 32'h0;
  assign _EVAL_152 = _EVAL_28 | _EVAL_113;
  assign _EVAL_173 = 13'h3f << _EVAL_14;
  assign _EVAL_186 = _EVAL_5 <= 3'h6;
  assign _EVAL_204 = _EVAL_16 ^ 25'h1800000;
  assign _EVAL_209 = {1'b0,$signed(_EVAL_204)};
  assign _EVAL_165 = $signed(_EVAL_209) & $signed(-26'sh8000);
  assign _EVAL_201 = $signed(_EVAL_165);
  assign _EVAL_257 = $signed(_EVAL_201) == $signed(26'sh0);
  assign _EVAL_254 = $signed(_EVAL_57) & $signed(-26'sh2000);
  assign _EVAL_250 = $signed(_EVAL_254);
  assign _EVAL_274 = $signed(_EVAL_250) == $signed(26'sh0);
  assign _EVAL_247 = _EVAL_257 | _EVAL_274;
  assign _EVAL_243 = _EVAL_186 & _EVAL_247;
  assign _EVAL_219 = _EVAL_243 | _EVAL_8;
  assign _EVAL_35 = _EVAL_3 == 1'h0;
  assign _EVAL_39 = _EVAL_35 | _EVAL_1;
  assign _EVAL_223 = _EVAL_39 | _EVAL_8;
  assign _EVAL_304 = _EVAL_223 == 1'h0;
  assign _EVAL_244 = 3'h6 == _EVAL_5;
  assign _EVAL_196 = _EVAL_301 ? _EVAL_244 : 1'h0;
  assign _EVAL_24 = _EVAL_196 | _EVAL_8;
  assign _EVAL_249 = _EVAL_4 <= 3'h4;
  assign _EVAL_89 = _EVAL_13[6:3];
  assign _EVAL_40 = _EVAL_89 == 4'h3;
  assign _EVAL_126 = _EVAL_175 == 1'h0;
  assign _EVAL_193 = _EVAL_4 != 3'h0;
  assign _EVAL_265 = _EVAL_193 | _EVAL_8;
  assign _EVAL_288 = _EVAL_265 == 1'h0;
  assign _EVAL_42 = _EVAL_4 <= 3'h2;
  assign _EVAL_120 = _EVAL_42 | _EVAL_8;
  assign _EVAL_53 = _EVAL_120 == 1'h0;
  assign _EVAL_300 = ~ _EVAL_0;
  assign _EVAL_48 = _EVAL_300 == 4'h0;
  assign _EVAL_279 = _EVAL_48 | _EVAL_8;
  assign _EVAL_134 = _EVAL_279 == 1'h0;
  assign _EVAL_138 = _EVAL_89 == 4'h8;
  assign _EVAL_70 = _EVAL_17 & _EVAL_9;
  assign _EVAL_189 = _EVAL_70 & _EVAL_282;
  assign _EVAL_237 = 128'h1 << _EVAL_2;
  assign _EVAL_157 = _EVAL_189 ? _EVAL_237 : 128'h0;
  assign _EVAL_142 = _EVAL_157[72:0];
  assign _EVAL_234 = _EVAL_142 != 73'h0;
  assign _EVAL_216 = _EVAL_205 | _EVAL_8;
  assign _EVAL_222 = _EVAL_216 == 1'h0;
  assign _EVAL_266 = _EVAL == _EVAL_125;
  assign _EVAL_229 = _EVAL_11 == _EVAL_224;
  assign _EVAL_228 = _EVAL_229 | _EVAL_8;
  assign _EVAL_97 = _EVAL_228 == 1'h0;
  assign _EVAL_172 = _EVAL_232 == 4'h0;
  assign _EVAL_148 = _EVAL_13 == 7'h48;
  assign _EVAL_45 = _EVAL_13 == 7'h40;
  assign _EVAL_136 = _EVAL_148 | _EVAL_45;
  assign _EVAL_51 = _EVAL_13[2:0];
  assign _EVAL_290 = 3'h1 <= _EVAL_51;
  assign _EVAL_20 = _EVAL_138 & _EVAL_290;
  assign _EVAL_114 = _EVAL_136 | _EVAL_20;
  assign _EVAL_65 = _EVAL_13 == 7'h20;
  assign _EVAL_215 = _EVAL_114 | _EVAL_65;
  assign _EVAL_30 = _EVAL_89 == 4'h0;
  assign _EVAL_161 = _EVAL_215 | _EVAL_30;
  assign _EVAL_86 = _EVAL_5 == _EVAL_179;
  assign _EVAL_122 = _EVAL_86 | _EVAL_8;
  assign _EVAL_276 = _EVAL_122 == 1'h0;
  assign _EVAL_236 = _EVAL_67 == 4'h0;
  assign _EVAL_218 = _EVAL_15[0];
  assign _EVAL_146 = _EVAL_173[5:0];
  assign _EVAL_149 = ~ _EVAL_146;
  assign _EVAL_278 = _EVAL_149[5:2];
  assign _EVAL_174 = _EVAL_67 - 4'h1;
  assign _EVAL_199 = _EVAL_308 | _EVAL_142;
  assign _EVAL_259 = _EVAL_12 & _EVAL_10;
  assign _EVAL_211 = _EVAL_259 & _EVAL_172;
  assign _EVAL_103 = _EVAL_15 == 3'h6;
  assign _EVAL_270 = _EVAL_103 == 1'h0;
  assign _EVAL_46 = _EVAL_211 & _EVAL_270;
  assign _EVAL_33 = 128'h1 << _EVAL_13;
  assign _EVAL_267 = _EVAL_46 ? _EVAL_33 : 128'h0;
  assign _EVAL_90 = _EVAL_267[72:0];
  assign _EVAL_183 = ~ _EVAL_90;
  assign _EVAL_128 = _EVAL_199 & _EVAL_183;
  assign _EVAL_263 = _EVAL_142 | _EVAL_308;
  assign _EVAL_52 = _EVAL_263 >> _EVAL_13;
  assign _EVAL_69 = _EVAL_52[0];
  assign _EVAL_214 = _EVAL_135 == 1'h0;
  assign _EVAL_98 = _EVAL_61 & _EVAL_214;
  assign _EVAL_291 = _EVAL_248 & _EVAL_98;
  assign _EVAL_41 = _EVAL_5 <= 3'h2;
  assign _EVAL_144 = _EVAL_41 & _EVAL_274;
  assign _EVAL_292 = _EVAL_144 | _EVAL_8;
  assign _EVAL_318 = _EVAL_292 == 1'h0;
  assign _EVAL_167 = _EVAL_10 & _EVAL_103;
  assign _EVAL_130 = _EVAL_298 < plusarg_reader_out;
  assign _EVAL_150 = _EVAL_152 | _EVAL_130;
  assign _EVAL_225 = _EVAL_150 | _EVAL_8;
  assign _EVAL_191 = _EVAL_2 == _EVAL_323;
  assign _EVAL_302 = _EVAL_191 | _EVAL_8;
  assign _EVAL_303 = _EVAL_302 == 1'h0;
  assign _EVAL_112 = _EVAL_6 == _EVAL_32;
  assign _EVAL_307 = _EVAL_112 | _EVAL_8;
  assign _EVAL_242 = _EVAL_307 == 1'h0;
  assign _EVAL_221 = _EVAL_14 >= 3'h2;
  assign _EVAL_281 = _EVAL_315 == 4'h0;
  assign _EVAL_213 = _EVAL_6[2];
  assign _EVAL_241 = _EVAL_213 == 1'h0;
  assign _EVAL_64 = 13'h3f << _EVAL_5;
  assign _EVAL_151 = _EVAL_64[5:0];
  assign _EVAL_71 = ~ _EVAL_151;
  assign _EVAL_38 = _EVAL_71[5:2];
  assign _EVAL_255 = _EVAL_315 - 4'h1;
  assign _EVAL_185 = _EVAL_142 != _EVAL_90;
  assign _EVAL_235 = _EVAL_234 == 1'h0;
  assign _EVAL_169 = _EVAL_185 | _EVAL_235;
  assign _EVAL_245 = _EVAL_169 | _EVAL_8;
  assign _EVAL_124 = _EVAL_281 == 1'h0;
  assign _EVAL_83 = _EVAL_9 & _EVAL_124;
  assign _EVAL_104 = _EVAL_311 | _EVAL_8;
  assign _EVAL_246 = _EVAL_89 == 4'h1;
  assign _EVAL_277 = _EVAL_161 | _EVAL_246;
  assign _EVAL_319 = _EVAL_89 == 4'h2;
  assign _EVAL_143 = _EVAL_277 | _EVAL_319;
  assign _EVAL_27 = _EVAL_15 == 3'h5;
  assign _EVAL_162 = _EVAL_6 == 3'h2;
  assign _EVAL_85 = _EVAL_4 == 3'h0;
  assign _EVAL_272 = _EVAL_85 | _EVAL_8;
  assign _EVAL_295 = _EVAL_266 | _EVAL_8;
  assign _EVAL_129 = _EVAL_295 == 1'h0;
  assign _EVAL_127 = _EVAL_298 + 32'h1;
  assign _EVAL_154 = _EVAL_232 - 4'h1;
  assign _EVAL_139 = _EVAL_221 | _EVAL_8;
  assign _EVAL_190 = _EVAL_139 == 1'h0;
  assign _EVAL_118 = _EVAL_308 >> _EVAL_2;
  assign _EVAL_59 = _EVAL_118[0];
  assign _EVAL_310 = _EVAL_59 == 1'h0;
  assign _EVAL_95 = _EVAL_310 | _EVAL_8;
  assign _EVAL_159 = _EVAL_95 == 1'h0;
  assign _EVAL_147 = _EVAL_236 == 1'h0;
  assign _EVAL_66 = _EVAL_15 == 3'h2;
  assign _EVAL_155 = _EVAL_7 == 1'h0;
  assign _EVAL_88 = _EVAL_16 == _EVAL_55;
  assign _EVAL_92 = {{19'd0}, _EVAL_71};
  assign _EVAL_171 = _EVAL_16 & _EVAL_92;
  assign _EVAL_325 = _EVAL_104 == 1'h0;
  assign _EVAL_324 = _EVAL_15 <= 3'h6;
  assign _EVAL_294 = _EVAL_324 | _EVAL_8;
  assign _EVAL_111 = _EVAL_294 == 1'h0;
  assign _EVAL_322 = _EVAL_1 == 1'h0;
  assign _EVAL_187 = _EVAL_322 | _EVAL_8;
  assign _EVAL_268 = _EVAL_15 == 3'h4;
  assign _EVAL_188 = _EVAL_10 & _EVAL_268;
  assign _EVAL_25 = _EVAL_6 == 3'h0;
  assign _EVAL_289 = _EVAL_9 & _EVAL_25;
  assign _EVAL_331 = _EVAL_249 | _EVAL_8;
  assign _EVAL_121 = _EVAL_331 == 1'h0;
  assign _EVAL_275 = _EVAL_225 == 1'h0;
  assign _EVAL_321 = _EVAL_10 & _EVAL_66;
  assign _EVAL_178 = _EVAL_14 == _EVAL_50;
  assign _EVAL_117 = _EVAL_178 | _EVAL_8;
  assign _EVAL_313 = _EVAL_117 == 1'h0;
  assign _EVAL_96 = _EVAL_233 & _EVAL_135;
  assign _EVAL_239 = _EVAL_248 & _EVAL_96;
  assign _EVAL_156 = _EVAL_24 == 1'h0;
  assign _EVAL_87 = _EVAL_171 == 25'h0;
  assign _EVAL_269 = _EVAL_6 == 3'h3;
  assign _EVAL_192 = _EVAL_9 & _EVAL_269;
  assign _EVAL_284 = _EVAL_4 <= 3'h3;
  assign _EVAL_105 = _EVAL_284 | _EVAL_8;
  assign _EVAL_78 = _EVAL_105 == 1'h0;
  assign _EVAL_195 = _EVAL_75 & _EVAL_233;
  assign _EVAL_197 = _EVAL_311 | _EVAL_195;
  assign _EVAL_286 = _EVAL_197 | _EVAL_239;
  assign _EVAL_320 = _EVAL_233 & _EVAL_214;
  assign _EVAL_100 = _EVAL_248 & _EVAL_320;
  assign _EVAL_312 = _EVAL_197 | _EVAL_100;
  assign _EVAL_37 = _EVAL_133 | _EVAL_291;
  assign _EVAL_80 = {_EVAL_286,_EVAL_312,_EVAL_36,_EVAL_37};
  assign _EVAL_176 = _EVAL_0 == _EVAL_80;
  assign _EVAL_160 = _EVAL_176 | _EVAL_8;
  assign _EVAL_332 = _EVAL_15 == _EVAL_43;
  assign _EVAL_271 = _EVAL_332 | _EVAL_8;
  assign _EVAL_253 = _EVAL_271 == 1'h0;
  assign _EVAL_327 = _EVAL_70 & _EVAL_281;
  assign _EVAL_21 = _EVAL_11 == 2'h0;
  assign _EVAL_106 = _EVAL_21 | _EVAL_8;
  assign _EVAL_293 = _EVAL_106 == 1'h0;
  assign _EVAL_158 = _EVAL_6 == 3'h7;
  assign _EVAL_260 = _EVAL_70 | _EVAL_259;
  assign _EVAL_328 = _EVAL_35 | _EVAL_8;
  assign _EVAL_206 = _EVAL_328 == 1'h0;
  assign _EVAL_273 = _EVAL_155 | _EVAL_8;
  assign _EVAL_170 = _EVAL_273 == 1'h0;
  assign _EVAL_164 = _EVAL_4 == _EVAL_252;
  assign _EVAL_203 = _EVAL_164 | _EVAL_8;
  assign _EVAL_285 = _EVAL_203 == 1'h0;
  assign _EVAL_231 = _EVAL_6 == 3'h5;
  assign _EVAL_60 = _EVAL_9 & _EVAL_231;
  assign _EVAL_22 = ~ _EVAL_80;
  assign _EVAL_110 = _EVAL_0 & _EVAL_22;
  assign _EVAL_309 = _EVAL_219 == 1'h0;
  assign _EVAL_317 = _EVAL_69 | _EVAL_8;
  assign _EVAL_99 = _EVAL_317 == 1'h0;
  assign _EVAL_305 = _EVAL_88 | _EVAL_8;
  assign _EVAL_238 = _EVAL_305 == 1'h0;
  assign _EVAL_194 = _EVAL_11 != 2'h2;
  assign _EVAL_44 = _EVAL_194 | _EVAL_8;
  assign _EVAL_261 = _EVAL_44 == 1'h0;
  assign _EVAL_23 = _EVAL_160 == 1'h0;
  assign _EVAL_108 = _EVAL_116 - 4'h1;
  assign _EVAL_329 = _EVAL_6 == 3'h4;
  assign _EVAL_287 = _EVAL_9 & _EVAL_329;
  assign _EVAL_227 = _EVAL_6 == 3'h6;
  assign _EVAL_202 = _EVAL_9 & _EVAL_227;
  assign _EVAL_180 = _EVAL_9 & _EVAL_158;
  assign _EVAL_163 = _EVAL_110 == 4'h0;
  assign _EVAL_251 = _EVAL_272 == 1'h0;
  assign _EVAL_182 = _EVAL_15 == 3'h0;
  assign _EVAL_109 = _EVAL_10 & _EVAL_182;
  assign _EVAL_73 = _EVAL_163 | _EVAL_8;
  assign _EVAL_101 = _EVAL_73 == 1'h0;
  assign _EVAL_137 = _EVAL_143 | _EVAL_40;
  assign _EVAL_306 = _EVAL_137 | _EVAL_8;
  assign _EVAL_47 = _EVAL_259 & _EVAL_236;
  assign _EVAL_166 = _EVAL_10 & _EVAL_147;
  assign _EVAL_68 = _EVAL_87 | _EVAL_8;
  assign _EVAL_102 = _EVAL_187 == 1'h0;
  assign _EVAL_217 = _EVAL_15 == 3'h1;
  assign _EVAL_19 = _EVAL_8 == 1'h0;
  assign _EVAL_84 = _EVAL_10 & _EVAL_27;
  assign _EVAL_140 = _EVAL_245 == 1'h0;
  assign _EVAL_81 = _EVAL_10 & _EVAL_217;
  assign _EVAL_256 = _EVAL_9 & _EVAL_162;
  assign _EVAL_91 = _EVAL_68 == 1'h0;
  assign _EVAL_119 = _EVAL_306 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_32 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_43 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_50 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_55 = _RAND_4[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_67 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_82 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_116 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_125 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_179 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_224 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_232 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_252 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_298 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {3{`RANDOM}};
  _EVAL_308 = _RAND_14[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_315 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_323 = _RAND_16[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_18) begin
    if (_EVAL_47) begin
      _EVAL_26 <= _EVAL_13;
    end
    if (_EVAL_327) begin
      _EVAL_32 <= _EVAL_6;
    end
    if (_EVAL_47) begin
      _EVAL_43 <= _EVAL_15;
    end
    if (_EVAL_47) begin
      _EVAL_50 <= _EVAL_14;
    end
    if (_EVAL_327) begin
      _EVAL_55 <= _EVAL_16;
    end
    if (_EVAL_8) begin
      _EVAL_67 <= 4'h0;
    end else begin
      if (_EVAL_259) begin
        if (_EVAL_236) begin
          if (_EVAL_218) begin
            _EVAL_67 <= _EVAL_278;
          end else begin
            _EVAL_67 <= 4'h0;
          end
        end else begin
          _EVAL_67 <= _EVAL_174;
        end
      end
    end
    if (_EVAL_47) begin
      _EVAL_82 <= _EVAL_3;
    end
    if (_EVAL_8) begin
      _EVAL_116 <= 4'h0;
    end else begin
      if (_EVAL_70) begin
        if (_EVAL_282) begin
          if (_EVAL_241) begin
            _EVAL_116 <= _EVAL_38;
          end else begin
            _EVAL_116 <= 4'h0;
          end
        end else begin
          _EVAL_116 <= _EVAL_108;
        end
      end
    end
    if (_EVAL_47) begin
      _EVAL_125 <= _EVAL;
    end
    if (_EVAL_327) begin
      _EVAL_179 <= _EVAL_5;
    end
    if (_EVAL_47) begin
      _EVAL_224 <= _EVAL_11;
    end
    if (_EVAL_8) begin
      _EVAL_232 <= 4'h0;
    end else begin
      if (_EVAL_259) begin
        if (_EVAL_172) begin
          if (_EVAL_218) begin
            _EVAL_232 <= _EVAL_278;
          end else begin
            _EVAL_232 <= 4'h0;
          end
        end else begin
          _EVAL_232 <= _EVAL_154;
        end
      end
    end
    if (_EVAL_327) begin
      _EVAL_252 <= _EVAL_4;
    end
    if (_EVAL_8) begin
      _EVAL_298 <= 32'h0;
    end else begin
      if (_EVAL_260) begin
        _EVAL_298 <= 32'h0;
      end else begin
        _EVAL_298 <= _EVAL_127;
      end
    end
    if (_EVAL_8) begin
      _EVAL_308 <= 73'h0;
    end else begin
      _EVAL_308 <= _EVAL_128;
    end
    if (_EVAL_8) begin
      _EVAL_315 <= 4'h0;
    end else begin
      if (_EVAL_70) begin
        if (_EVAL_281) begin
          if (_EVAL_241) begin
            _EVAL_315 <= _EVAL_38;
          end else begin
            _EVAL_315 <= 4'h0;
          end
        end else begin
          _EVAL_315 <= _EVAL_255;
        end
      end
    end
    if (_EVAL_327) begin
      _EVAL_323 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8f69b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f9d871c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14f7c3d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc6c7724)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8399eafc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ec6ba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ce10529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0a7bd56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b394ea4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45afabf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c5e1544)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84dcab23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87c69517)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(316c6a9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2e792a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(363c4a4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e583ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ed1d4f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6195e102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef0d4179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe347374)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(717bb7d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4520fe4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ef4b42e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9050c223)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4dd3ae3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbd9982f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e0c93c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fa1a46d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa236594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3811d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e7b352)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(255c8928)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82aa08d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5ee59c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a970e4ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de04b1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4e8fd22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9ae5486)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7a088fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e04a3b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd93e6ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e23af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e069e96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77942d8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aef1a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aabf70a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7a949e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277aacec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33d4755c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2314036a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bd7c247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdcd548f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0d1fe6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab33a95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7814ad50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53430c74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(571c6197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cd6d5b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81607f60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fe1948a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d99b011)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8334c61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2b7cc9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57ce9f34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50222b8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a26db1c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(184e47ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbdef0c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2c1a4e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61d428f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0270bc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8976ae3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31bb2e5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52beb5e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5748ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1388490)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4da81b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e52b2365)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a28247d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e34d3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad9bd2ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed80eb91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(959e30aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dde29db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b49967d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b57f4889)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2403d351)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17c45c27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4031c5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97041ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(529c9db1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a22c8506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87a2ff4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e0b31e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
