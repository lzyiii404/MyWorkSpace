//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_61_assert(
  input  [4:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [4:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [1:0] _EVAL_38;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_129;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_133;
  reg [31:0] _RAND_2;
  reg  _EVAL_142;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_161;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_163;
  reg [31:0] _RAND_5;
  reg [31:0] _EVAL_171;
  reg [31:0] _RAND_6;
  reg [5:0] _EVAL_227;
  reg [31:0] _RAND_7;
  reg [31:0] _EVAL_231;
  reg [31:0] _RAND_8;
  reg  _EVAL_265;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_268;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_279;
  reg [31:0] _RAND_11;
  reg [5:0] _EVAL_285;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_311;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_319;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_339;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_344;
  reg [31:0] _RAND_16;
  wire [3:0] _EVAL_114;
  wire  _EVAL_152;
  wire [5:0] _EVAL_146;
  wire [31:0] _EVAL_267;
  wire  _EVAL_175;
  wire  _EVAL_263;
  wire [31:0] _EVAL_109;
  wire [32:0] _EVAL_206;
  wire  _EVAL_182;
  wire [22:0] _EVAL_149;
  wire [7:0] _EVAL_259;
  wire [7:0] _EVAL_232;
  wire [5:0] _EVAL_75;
  wire [31:0] _EVAL_249;
  wire  _EVAL_293;
  wire [31:0] _EVAL_349;
  wire [32:0] _EVAL_120;
  wire [1:0] _EVAL_140;
  wire [1:0] _EVAL_266;
  wire  _EVAL_66;
  wire  _EVAL_200;
  wire  _EVAL_221;
  wire  _EVAL_88;
  wire  _EVAL_78;
  wire  _EVAL_219;
  wire  _EVAL_76;
  wire  _EVAL_145;
  wire  _EVAL_125;
  wire [22:0] _EVAL_42;
  wire [7:0] _EVAL_304;
  wire [7:0] _EVAL_211;
  wire [5:0] _EVAL_72;
  wire [31:0] _EVAL_351;
  wire  _EVAL_168;
  wire  _EVAL_191;
  wire  _EVAL_180;
  wire [31:0] _EVAL_223;
  wire [31:0] _EVAL_210;
  wire  _EVAL_101;
  wire  _EVAL_299;
  wire  _EVAL_106;
  wire  _EVAL_79;
  wire  _EVAL_22;
  wire  _EVAL_203;
  wire [31:0] _EVAL_312;
  wire  _EVAL_243;
  wire  _EVAL_306;
  wire  _EVAL_278;
  wire  _EVAL_283;
  wire  _EVAL_160;
  wire  _EVAL_190;
  wire  _EVAL_233;
  wire  _EVAL_57;
  wire  _EVAL_208;
  wire  _EVAL_63;
  wire  _EVAL_326;
  wire  _EVAL_64;
  wire  _EVAL_49;
  wire  _EVAL_130;
  wire  _EVAL_143;
  wire  _EVAL_287;
  wire  _EVAL_340;
  wire [32:0] _EVAL_241;
  wire [32:0] _EVAL_217;
  wire [32:0] _EVAL_92;
  wire  _EVAL_85;
  wire [31:0] _EVAL_325;
  wire [32:0] _EVAL_33;
  wire [32:0] _EVAL_350;
  wire [32:0] _EVAL_230;
  wire  _EVAL_238;
  wire  _EVAL_103;
  wire [32:0] _EVAL_218;
  wire [32:0] _EVAL_195;
  wire  _EVAL_261;
  wire  _EVAL_357;
  wire [32:0] _EVAL_316;
  wire [32:0] _EVAL_305;
  wire [32:0] _EVAL_167;
  wire  _EVAL_122;
  wire  _EVAL_226;
  wire [31:0] _EVAL_30;
  wire [32:0] _EVAL_136;
  wire [32:0] _EVAL_118;
  wire [32:0] _EVAL_262;
  wire  _EVAL_187;
  wire  _EVAL_225;
  wire [31:0] _EVAL_48;
  wire [32:0] _EVAL_333;
  wire [32:0] _EVAL_84;
  wire [32:0] _EVAL_248;
  wire  _EVAL_173;
  wire  _EVAL_23;
  wire [31:0] _EVAL_300;
  wire [31:0] _EVAL_289;
  wire  _EVAL_215;
  wire [1:0] _EVAL_194;
  wire  _EVAL_213;
  wire  _EVAL_199;
  wire  _EVAL_34;
  wire  _EVAL_197;
  wire  _EVAL_164;
  wire  _EVAL_60;
  wire  _EVAL_205;
  wire  _EVAL_318;
  wire  _EVAL_98;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_86;
  wire  _EVAL_162;
  wire [32:0] _EVAL_341;
  wire [32:0] _EVAL_290;
  wire [32:0] _EVAL_117;
  wire  _EVAL_159;
  wire  _EVAL_354;
  wire  _EVAL_181;
  wire  _EVAL_31;
  wire  _EVAL_70;
  wire  _EVAL_274;
  wire  _EVAL_315;
  wire [31:0] _EVAL_158;
  wire  _EVAL_220;
  wire  _EVAL_235;
  wire  _EVAL_127;
  wire  _EVAL_260;
  wire  _EVAL_59;
  wire  _EVAL_282;
  wire  _EVAL_332;
  wire  _EVAL_54;
  wire [5:0] _EVAL_329;
  wire  _EVAL_358;
  wire  _EVAL_240;
  wire  _EVAL_337;
  wire  _EVAL_153;
  wire  _EVAL_322;
  wire  _EVAL_291;
  wire  _EVAL_273;
  wire  _EVAL_77;
  wire [31:0] _EVAL_176;
  wire  _EVAL_327;
  wire  _EVAL_55;
  wire  _EVAL_275;
  wire  _EVAL_95;
  wire  _EVAL_192;
  wire  _EVAL_124;
  wire [1:0] _EVAL_99;
  wire  _EVAL_147;
  wire  _EVAL_157;
  wire  _EVAL_151;
  wire  _EVAL_336;
  wire  _EVAL_320;
  wire  _EVAL_280;
  wire  _EVAL_113;
  wire  _EVAL_250;
  wire  _EVAL_43;
  wire  _EVAL_111;
  wire  _EVAL_198;
  wire  _EVAL_24;
  wire  _EVAL_328;
  wire  _EVAL_121;
  wire  _EVAL_323;
  wire  _EVAL_154;
  wire  _EVAL_294;
  wire  _EVAL_74;
  wire  _EVAL_28;
  wire  _EVAL_155;
  wire  _EVAL_269;
  wire  _EVAL_355;
  wire  _EVAL_35;
  wire  _EVAL_97;
  wire [31:0] _EVAL_126;
  wire [32:0] _EVAL_338;
  wire [32:0] _EVAL_138;
  wire  _EVAL_132;
  wire  _EVAL_73;
  wire  _EVAL_44;
  wire  _EVAL_255;
  wire  _EVAL_330;
  wire  _EVAL_288;
  wire  _EVAL_62;
  wire  _EVAL_134;
  wire [32:0] _EVAL_68;
  wire  _EVAL_139;
  wire  _EVAL_242;
  wire  _EVAL_239;
  wire  _EVAL_244;
  wire  _EVAL_298;
  wire  _EVAL_183;
  wire  _EVAL_135;
  wire  _EVAL_247;
  wire  _EVAL_228;
  wire  _EVAL_61;
  wire  _EVAL_348;
  wire  _EVAL_144;
  wire  _EVAL_222;
  wire  _EVAL_100;
  wire  _EVAL_331;
  wire  _EVAL_356;
  wire  _EVAL_264;
  wire  _EVAL_204;
  wire  _EVAL_116;
  wire  _EVAL_276;
  wire  _EVAL_303;
  wire  _EVAL_174;
  wire  _EVAL_257;
  wire [3:0] _EVAL_309;
  wire [3:0] _EVAL_131;
  wire [3:0] _EVAL_272;
  wire [31:0] _EVAL_179;
  wire  _EVAL_246;
  wire  _EVAL_150;
  wire  _EVAL_91;
  wire  _EVAL_39;
  wire  _EVAL_189;
  wire  _EVAL_94;
  wire  _EVAL_216;
  wire  _EVAL_156;
  wire  _EVAL_193;
  wire  _EVAL_284;
  wire  _EVAL_110;
  wire  _EVAL_295;
  wire  _EVAL_82;
  wire  _EVAL_128;
  wire  _EVAL_148;
  wire  _EVAL_251;
  wire  _EVAL_245;
  wire  _EVAL_286;
  wire  _EVAL_196;
  wire  _EVAL_352;
  wire  _EVAL_32;
  wire  _EVAL_292;
  wire  _EVAL_141;
  wire [31:0] _EVAL_342;
  wire [31:0] _EVAL_90;
  wire  _EVAL_80;
  wire  _EVAL_308;
  wire  _EVAL_310;
  wire  _EVAL_335;
  wire  _EVAL_45;
  wire [31:0] _EVAL_65;
  wire  _EVAL_29;
  wire  _EVAL_50;
  wire  _EVAL_119;
  wire  _EVAL_277;
  wire  _EVAL_108;
  wire  _EVAL_178;
  wire  _EVAL_102;
  wire  _EVAL_67;
  wire  _EVAL_170;
  wire  _EVAL_186;
  wire  _EVAL_256;
  wire [5:0] _EVAL_234;
  wire  _EVAL_201;
  wire  _EVAL_253;
  wire  _EVAL_20;
  wire  _EVAL_81;
  wire  _EVAL_346;
  wire  _EVAL_207;
  wire  _EVAL_137;
  wire  _EVAL_297;
  wire  _EVAL_296;
  wire  _EVAL_115;
  wire  _EVAL_302;
  wire  _EVAL_112;
  wire  _EVAL_87;
  wire  _EVAL_36;
  wire  _EVAL_301;
  wire  _EVAL_40;
  wire  _EVAL_51;
  wire  _EVAL_123;
  wire  _EVAL_93;
  wire  _EVAL_314;
  wire  _EVAL_229;
  wire  _EVAL_209;
  wire  _EVAL_317;
  wire  _EVAL_89;
  wire  _EVAL_105;
  wire  _EVAL_270;
  wire  _EVAL_25;
  wire  _EVAL_172;
  wire [5:0] _EVAL_347;
  wire  _EVAL_224;
  wire  _EVAL_96;
  wire  _EVAL_324;
  wire  _EVAL_258;
  wire  _EVAL_236;
  wire  _EVAL_353;
  wire  _EVAL_345;
  wire  _EVAL_58;
  wire  _EVAL_56;
  wire  _EVAL_53;
  wire  _EVAL_166;
  wire  _EVAL_19;
  wire  _EVAL_71;
  wire  _EVAL_313;
  wire  _EVAL_202;
  wire  _EVAL_254;
  wire  _EVAL_52;
  wire  _EVAL_271;
  wire  _EVAL_46;
  wire  _EVAL_26;
  wire  _EVAL_321;
  wire [31:0] _EVAL_169;
  wire  _EVAL_307;
  wire  _EVAL_185;
  wire  _EVAL_184;
  wire  _EVAL_165;
  wire  _EVAL_237;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_114 = ~ _EVAL_10;
  assign _EVAL_152 = _EVAL_114 == 4'h0;
  assign _EVAL_146 = _EVAL_227 - 6'h1;
  assign _EVAL_267 = _EVAL_17 ^ 32'h80000000;
  assign _EVAL_175 = _EVAL_16 == _EVAL_265;
  assign _EVAL_263 = _EVAL_2[0];
  assign _EVAL_109 = _EVAL_17 ^ 32'h2000000;
  assign _EVAL_206 = {1'b0,$signed(_EVAL_109)};
  assign _EVAL_182 = _EVAL_8[0];
  assign _EVAL_149 = 23'hff << _EVAL_18;
  assign _EVAL_259 = _EVAL_149[7:0];
  assign _EVAL_232 = ~ _EVAL_259;
  assign _EVAL_75 = _EVAL_232[7:2];
  assign _EVAL_249 = _EVAL_17 ^ 32'h3000;
  assign _EVAL_293 = _EVAL_4 != 2'h2;
  assign _EVAL_349 = _EVAL_17 ^ 32'h40000000;
  assign _EVAL_120 = {1'b0,$signed(_EVAL_349)};
  assign _EVAL_140 = 2'h1 << _EVAL_263;
  assign _EVAL_266 = _EVAL_140 | 2'h1;
  assign _EVAL_66 = _EVAL_266[0];
  assign _EVAL_200 = _EVAL_17[1];
  assign _EVAL_221 = _EVAL_200 == 1'h0;
  assign _EVAL_88 = _EVAL_17[0];
  assign _EVAL_78 = _EVAL_88 == 1'h0;
  assign _EVAL_219 = _EVAL_221 & _EVAL_78;
  assign _EVAL_76 = _EVAL_66 & _EVAL_219;
  assign _EVAL_145 = _EVAL_7[2];
  assign _EVAL_125 = _EVAL_145 == 1'h0;
  assign _EVAL_42 = 23'hff << _EVAL_2;
  assign _EVAL_304 = _EVAL_42[7:0];
  assign _EVAL_211 = ~ _EVAL_304;
  assign _EVAL_72 = _EVAL_211[7:2];
  assign _EVAL_351 = {{24'd0}, _EVAL_211};
  assign _EVAL_168 = _EVAL_11 & _EVAL_1;
  assign _EVAL_191 = _EVAL_227 == 6'h0;
  assign _EVAL_180 = _EVAL_168 & _EVAL_191;
  assign _EVAL_223 = 32'h1 << _EVAL_5;
  assign _EVAL_210 = _EVAL_180 ? _EVAL_223 : 32'h0;
  assign _EVAL_101 = _EVAL_210 != 32'h0;
  assign _EVAL_299 = _EVAL_15 == 1'h0;
  assign _EVAL_106 = _EVAL_231 != 32'h0;
  assign _EVAL_79 = _EVAL_106 == 1'h0;
  assign _EVAL_22 = _EVAL_3 == 3'h0;
  assign _EVAL_203 = _EVAL_22 | _EVAL_12;
  assign _EVAL_312 = _EVAL_231 >> _EVAL_5;
  assign _EVAL_243 = _EVAL_312[0];
  assign _EVAL_306 = _EVAL_243 == 1'h0;
  assign _EVAL_278 = _EVAL_306 | _EVAL_12;
  assign _EVAL_283 = _EVAL_278 == 1'h0;
  assign _EVAL_160 = _EVAL_14 & _EVAL_0;
  assign _EVAL_190 = _EVAL_268 == 6'h0;
  assign _EVAL_233 = _EVAL_160 & _EVAL_190;
  assign _EVAL_57 = _EVAL_8 == 3'h6;
  assign _EVAL_208 = _EVAL_57 == 1'h0;
  assign _EVAL_63 = _EVAL_233 & _EVAL_208;
  assign _EVAL_326 = _EVAL_4 == _EVAL_38;
  assign _EVAL_64 = _EVAL_326 | _EVAL_12;
  assign _EVAL_49 = _EVAL_64 == 1'h0;
  assign _EVAL_130 = _EVAL_8 == 3'h5;
  assign _EVAL_143 = _EVAL_0 & _EVAL_130;
  assign _EVAL_287 = _EVAL_13 == 1'h0;
  assign _EVAL_340 = _EVAL_3 == _EVAL_279;
  assign _EVAL_241 = {1'b0,$signed(_EVAL_249)};
  assign _EVAL_217 = $signed(_EVAL_241) & $signed(-33'sh1000);
  assign _EVAL_92 = $signed(_EVAL_217);
  assign _EVAL_85 = $signed(_EVAL_92) == $signed(33'sh0);
  assign _EVAL_325 = _EVAL_17 ^ 32'hc000000;
  assign _EVAL_33 = {1'b0,$signed(_EVAL_325)};
  assign _EVAL_350 = $signed(_EVAL_33) & $signed(-33'sh4000000);
  assign _EVAL_230 = $signed(_EVAL_350);
  assign _EVAL_238 = $signed(_EVAL_230) == $signed(33'sh0);
  assign _EVAL_103 = _EVAL_85 | _EVAL_238;
  assign _EVAL_218 = $signed(_EVAL_206) & $signed(-33'sh10000);
  assign _EVAL_195 = $signed(_EVAL_218);
  assign _EVAL_261 = $signed(_EVAL_195) == $signed(33'sh0);
  assign _EVAL_357 = _EVAL_103 | _EVAL_261;
  assign _EVAL_316 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_305 = $signed(_EVAL_316) & $signed(-33'sh5000);
  assign _EVAL_167 = $signed(_EVAL_305);
  assign _EVAL_122 = $signed(_EVAL_167) == $signed(33'sh0);
  assign _EVAL_226 = _EVAL_357 | _EVAL_122;
  assign _EVAL_30 = _EVAL_17 ^ 32'h1800000;
  assign _EVAL_136 = {1'b0,$signed(_EVAL_30)};
  assign _EVAL_118 = $signed(_EVAL_136) & $signed(-33'sh8000);
  assign _EVAL_262 = $signed(_EVAL_118);
  assign _EVAL_187 = $signed(_EVAL_262) == $signed(33'sh0);
  assign _EVAL_225 = _EVAL_226 | _EVAL_187;
  assign _EVAL_48 = _EVAL_17 ^ 32'h1900000;
  assign _EVAL_333 = {1'b0,$signed(_EVAL_48)};
  assign _EVAL_84 = $signed(_EVAL_333) & $signed(-33'sh2000);
  assign _EVAL_248 = $signed(_EVAL_84);
  assign _EVAL_173 = $signed(_EVAL_248) == $signed(33'sh0);
  assign _EVAL_23 = _EVAL_225 | _EVAL_173;
  assign _EVAL_300 = 32'h1 << _EVAL;
  assign _EVAL_289 = _EVAL_63 ? _EVAL_300 : 32'h0;
  assign _EVAL_215 = _EVAL_210 != _EVAL_289;
  assign _EVAL_194 = _EVAL[4:3];
  assign _EVAL_213 = _EVAL_194 == 2'h0;
  assign _EVAL_199 = _EVAL_194 == 2'h1;
  assign _EVAL_34 = _EVAL_213 | _EVAL_199;
  assign _EVAL_197 = _EVAL_194 == 2'h2;
  assign _EVAL_164 = _EVAL_34 | _EVAL_197;
  assign _EVAL_60 = _EVAL_194 == 2'h3;
  assign _EVAL_205 = _EVAL_164 | _EVAL_60;
  assign _EVAL_318 = _EVAL_205 | _EVAL_12;
  assign _EVAL_98 = _EVAL_318 == 1'h0;
  assign _EVAL_104 = $signed(_EVAL_120) & $signed(-33'sh2000);
  assign _EVAL_86 = $signed(_EVAL_104);
  assign _EVAL_162 = $signed(_EVAL_86) == $signed(33'sh0);
  assign _EVAL_341 = {1'b0,$signed(_EVAL_267)};
  assign _EVAL_290 = $signed(_EVAL_341) & $signed(-33'sh20000);
  assign _EVAL_117 = $signed(_EVAL_290);
  assign _EVAL_159 = $signed(_EVAL_117) == $signed(33'sh0);
  assign _EVAL_354 = _EVAL_162 | _EVAL_159;
  assign _EVAL_181 = _EVAL_354 | _EVAL_238;
  assign _EVAL_31 = _EVAL_18 >= 4'h2;
  assign _EVAL_70 = _EVAL_31 | _EVAL_12;
  assign _EVAL_274 = _EVAL_7 == _EVAL_339;
  assign _EVAL_315 = _EVAL_2 <= 4'h6;
  assign _EVAL_158 = _EVAL_231 | _EVAL_210;
  assign _EVAL_220 = _EVAL_7 == 3'h1;
  assign _EVAL_235 = _EVAL_2 >= 4'h2;
  assign _EVAL_127 = _EVAL_235 | _EVAL_12;
  assign _EVAL_260 = _EVAL_127 == 1'h0;
  assign _EVAL_59 = _EVAL_16 == 1'h0;
  assign _EVAL_282 = _EVAL_59 | _EVAL_15;
  assign _EVAL_332 = _EVAL_282 | _EVAL_12;
  assign _EVAL_54 = _EVAL_133 == 6'h0;
  assign _EVAL_329 = _EVAL_133 - 6'h1;
  assign _EVAL_358 = _EVAL_18 == _EVAL_129;
  assign _EVAL_240 = _EVAL_358 | _EVAL_12;
  assign _EVAL_337 = _EVAL_7 == 3'h4;
  assign _EVAL_153 = _EVAL_1 & _EVAL_337;
  assign _EVAL_322 = _EVAL_101 == 1'h0;
  assign _EVAL_291 = _EVAL_215 | _EVAL_322;
  assign _EVAL_273 = _EVAL_291 | _EVAL_12;
  assign _EVAL_77 = _EVAL_168 | _EVAL_160;
  assign _EVAL_176 = _EVAL_171 + 32'h1;
  assign _EVAL_327 = _EVAL_285 == 6'h0;
  assign _EVAL_55 = _EVAL_327 == 1'h0;
  assign _EVAL_275 = _EVAL_340 | _EVAL_12;
  assign _EVAL_95 = _EVAL_274 | _EVAL_12;
  assign _EVAL_192 = _EVAL_95 == 1'h0;
  assign _EVAL_124 = _EVAL_293 | _EVAL_12;
  assign _EVAL_99 = _EVAL_5[4:3];
  assign _EVAL_147 = _EVAL_99 == 2'h0;
  assign _EVAL_157 = _EVAL_3 != 3'h0;
  assign _EVAL_151 = _EVAL_2 == _EVAL_163;
  assign _EVAL_336 = _EVAL_240 == 1'h0;
  assign _EVAL_320 = _EVAL_7 == 3'h7;
  assign _EVAL_280 = _EVAL_8 == 3'h0;
  assign _EVAL_113 = _EVAL_0 & _EVAL_280;
  assign _EVAL_250 = _EVAL_160 & _EVAL_327;
  assign _EVAL_43 = _EVAL_2 <= 4'h2;
  assign _EVAL_111 = _EVAL_200 & _EVAL_78;
  assign _EVAL_198 = plusarg_reader_out == 32'h0;
  assign _EVAL_24 = _EVAL_3 <= 3'h2;
  assign _EVAL_328 = _EVAL_24 | _EVAL_12;
  assign _EVAL_121 = _EVAL_4 <= 2'h2;
  assign _EVAL_323 = _EVAL_2 <= 4'h8;
  assign _EVAL_154 = _EVAL_323 & _EVAL_85;
  assign _EVAL_294 = _EVAL_181 | _EVAL_261;
  assign _EVAL_74 = _EVAL_294 | _EVAL_122;
  assign _EVAL_28 = _EVAL_59 | _EVAL_12;
  assign _EVAL_155 = _EVAL_299 | _EVAL_12;
  assign _EVAL_269 = _EVAL_155 == 1'h0;
  assign _EVAL_355 = _EVAL_12 == 1'h0;
  assign _EVAL_35 = _EVAL_200 & _EVAL_88;
  assign _EVAL_97 = _EVAL_66 & _EVAL_35;
  assign _EVAL_126 = _EVAL_17 ^ 32'h20000000;
  assign _EVAL_338 = {1'b0,$signed(_EVAL_126)};
  assign _EVAL_138 = $signed(_EVAL_338) & $signed(-33'sh2000);
  assign _EVAL_132 = _EVAL_99 == 2'h1;
  assign _EVAL_73 = _EVAL_147 | _EVAL_132;
  assign _EVAL_44 = _EVAL_99 == 2'h2;
  assign _EVAL_255 = _EVAL_73 | _EVAL_44;
  assign _EVAL_330 = _EVAL_99 == 2'h3;
  assign _EVAL_288 = _EVAL_255 | _EVAL_330;
  assign _EVAL_62 = _EVAL_288 | _EVAL_12;
  assign _EVAL_134 = _EVAL_62 == 1'h0;
  assign _EVAL_68 = $signed(_EVAL_138);
  assign _EVAL_139 = $signed(_EVAL_68) == $signed(33'sh0);
  assign _EVAL_242 = _EVAL_275 == 1'h0;
  assign _EVAL_239 = _EVAL_23 | _EVAL_139;
  assign _EVAL_244 = _EVAL_74 | _EVAL_187;
  assign _EVAL_298 = _EVAL_8 == 3'h2;
  assign _EVAL_183 = _EVAL_0 & _EVAL_298;
  assign _EVAL_135 = _EVAL_266[1];
  assign _EVAL_247 = _EVAL_135 & _EVAL_221;
  assign _EVAL_228 = _EVAL_235 | _EVAL_247;
  assign _EVAL_61 = _EVAL_221 & _EVAL_88;
  assign _EVAL_348 = _EVAL_66 & _EVAL_61;
  assign _EVAL_144 = _EVAL_228 | _EVAL_348;
  assign _EVAL_222 = _EVAL_3 <= 3'h3;
  assign _EVAL_100 = _EVAL_222 | _EVAL_12;
  assign _EVAL_331 = _EVAL_100 == 1'h0;
  assign _EVAL_356 = _EVAL_152 | _EVAL_12;
  assign _EVAL_264 = _EVAL_356 == 1'h0;
  assign _EVAL_204 = _EVAL_135 & _EVAL_200;
  assign _EVAL_116 = _EVAL_235 | _EVAL_204;
  assign _EVAL_276 = _EVAL_116 | _EVAL_97;
  assign _EVAL_303 = _EVAL_66 & _EVAL_111;
  assign _EVAL_174 = _EVAL_116 | _EVAL_303;
  assign _EVAL_257 = _EVAL_228 | _EVAL_76;
  assign _EVAL_309 = {_EVAL_276,_EVAL_174,_EVAL_144,_EVAL_257};
  assign _EVAL_131 = ~ _EVAL_309;
  assign _EVAL_272 = _EVAL_10 & _EVAL_131;
  assign _EVAL_179 = _EVAL_17 & _EVAL_351;
  assign _EVAL_246 = _EVAL_179 == 32'h0;
  assign _EVAL_150 = _EVAL_8 <= 3'h6;
  assign _EVAL_91 = _EVAL_150 | _EVAL_12;
  assign _EVAL_39 = _EVAL_3 <= 3'h4;
  assign _EVAL_189 = _EVAL_39 | _EVAL_12;
  assign _EVAL_94 = _EVAL_189 == 1'h0;
  assign _EVAL_216 = _EVAL_1 & _EVAL_220;
  assign _EVAL_156 = _EVAL_1 & _EVAL_320;
  assign _EVAL_193 = _EVAL_8 == _EVAL_344;
  assign _EVAL_284 = _EVAL_193 | _EVAL_12;
  assign _EVAL_110 = _EVAL_244 | _EVAL_173;
  assign _EVAL_295 = _EVAL_110 | _EVAL_139;
  assign _EVAL_82 = _EVAL_315 & _EVAL_295;
  assign _EVAL_128 = _EVAL_82 | _EVAL_154;
  assign _EVAL_148 = _EVAL_128 | _EVAL_12;
  assign _EVAL_251 = _EVAL_148 == 1'h0;
  assign _EVAL_245 = _EVAL_287 | _EVAL_12;
  assign _EVAL_286 = _EVAL == _EVAL_161;
  assign _EVAL_196 = _EVAL_286 | _EVAL_12;
  assign _EVAL_352 = _EVAL_272 == 4'h0;
  assign _EVAL_32 = _EVAL_352 | _EVAL_12;
  assign _EVAL_292 = _EVAL_7 == 3'h2;
  assign _EVAL_141 = _EVAL_1 & _EVAL_292;
  assign _EVAL_342 = _EVAL_210 | _EVAL_231;
  assign _EVAL_90 = _EVAL_342 >> _EVAL;
  assign _EVAL_80 = _EVAL_90[0];
  assign _EVAL_308 = _EVAL_8 == 3'h1;
  assign _EVAL_310 = _EVAL_28 == 1'h0;
  assign _EVAL_335 = _EVAL_17 == _EVAL_311;
  assign _EVAL_45 = _EVAL_328 == 1'h0;
  assign _EVAL_65 = ~ _EVAL_289;
  assign _EVAL_29 = _EVAL_5 == _EVAL_319;
  assign _EVAL_50 = _EVAL_29 | _EVAL_12;
  assign _EVAL_119 = _EVAL_50 == 1'h0;
  assign _EVAL_277 = _EVAL_4 == 2'h0;
  assign _EVAL_108 = _EVAL_277 | _EVAL_12;
  assign _EVAL_178 = _EVAL_108 == 1'h0;
  assign _EVAL_102 = _EVAL_80 | _EVAL_12;
  assign _EVAL_67 = _EVAL_332 == 1'h0;
  assign _EVAL_170 = _EVAL_43 & _EVAL_239;
  assign _EVAL_186 = _EVAL_170 | _EVAL_12;
  assign _EVAL_256 = _EVAL_246 | _EVAL_12;
  assign _EVAL_234 = _EVAL_285 - 6'h1;
  assign _EVAL_201 = _EVAL_168 & _EVAL_54;
  assign _EVAL_253 = _EVAL_196 == 1'h0;
  assign _EVAL_20 = _EVAL_121 | _EVAL_12;
  assign _EVAL_81 = _EVAL_10 == _EVAL_309;
  assign _EVAL_346 = _EVAL_81 | _EVAL_12;
  assign _EVAL_207 = _EVAL_346 == 1'h0;
  assign _EVAL_137 = _EVAL_7 == 3'h5;
  assign _EVAL_297 = _EVAL_1 & _EVAL_137;
  assign _EVAL_296 = _EVAL_7 == 3'h0;
  assign _EVAL_115 = _EVAL_154 | _EVAL_12;
  assign _EVAL_302 = _EVAL_79 | _EVAL_198;
  assign _EVAL_112 = _EVAL_171 < plusarg_reader_out;
  assign _EVAL_87 = _EVAL_302 | _EVAL_112;
  assign _EVAL_36 = _EVAL_87 | _EVAL_12;
  assign _EVAL_301 = _EVAL_54 == 1'h0;
  assign _EVAL_40 = _EVAL_7 == 3'h6;
  assign _EVAL_51 = _EVAL_32 == 1'h0;
  assign _EVAL_123 = _EVAL_315 & _EVAL_159;
  assign _EVAL_93 = _EVAL_123 | _EVAL_12;
  assign _EVAL_314 = _EVAL_175 | _EVAL_12;
  assign _EVAL_229 = _EVAL_124 == 1'h0;
  assign _EVAL_209 = _EVAL_335 | _EVAL_12;
  assign _EVAL_317 = _EVAL_209 == 1'h0;
  assign _EVAL_89 = _EVAL_8 == 3'h4;
  assign _EVAL_105 = _EVAL_9 == _EVAL_142;
  assign _EVAL_270 = _EVAL_105 | _EVAL_12;
  assign _EVAL_25 = _EVAL_270 == 1'h0;
  assign _EVAL_172 = _EVAL_284 == 1'h0;
  assign _EVAL_347 = _EVAL_268 - 6'h1;
  assign _EVAL_224 = _EVAL_203 == 1'h0;
  assign _EVAL_96 = _EVAL_36 == 1'h0;
  assign _EVAL_324 = _EVAL_91 == 1'h0;
  assign _EVAL_258 = _EVAL_1 & _EVAL_296;
  assign _EVAL_236 = _EVAL_93 == 1'h0;
  assign _EVAL_353 = _EVAL_314 == 1'h0;
  assign _EVAL_345 = _EVAL_273 == 1'h0;
  assign _EVAL_58 = _EVAL_0 & _EVAL_89;
  assign _EVAL_56 = _EVAL_0 & _EVAL_308;
  assign _EVAL_53 = _EVAL_151 | _EVAL_12;
  assign _EVAL_166 = _EVAL_53 == 1'h0;
  assign _EVAL_19 = _EVAL_102 == 1'h0;
  assign _EVAL_71 = _EVAL_186 == 1'h0;
  assign _EVAL_313 = _EVAL_157 | _EVAL_12;
  assign _EVAL_202 = _EVAL_313 == 1'h0;
  assign _EVAL_254 = _EVAL_1 & _EVAL_301;
  assign _EVAL_52 = _EVAL_7 == 3'h3;
  assign _EVAL_271 = _EVAL_1 & _EVAL_40;
  assign _EVAL_46 = _EVAL_245 == 1'h0;
  assign _EVAL_26 = _EVAL_115 == 1'h0;
  assign _EVAL_321 = _EVAL_0 & _EVAL_57;
  assign _EVAL_169 = _EVAL_158 & _EVAL_65;
  assign _EVAL_307 = _EVAL_256 == 1'h0;
  assign _EVAL_185 = _EVAL_0 & _EVAL_55;
  assign _EVAL_184 = _EVAL_20 == 1'h0;
  assign _EVAL_165 = _EVAL_70 == 1'h0;
  assign _EVAL_237 = _EVAL_1 & _EVAL_52;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_38 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_129 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_133 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_142 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_161 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_163 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_171 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_227 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_231 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_265 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_268 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_279 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_285 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_311 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_319 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_339 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_344 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_6) begin
    if (_EVAL_250) begin
      _EVAL_38 <= _EVAL_4;
    end
    if (_EVAL_250) begin
      _EVAL_129 <= _EVAL_18;
    end
    if (_EVAL_12) begin
      _EVAL_133 <= 6'h0;
    end else begin
      if (_EVAL_168) begin
        if (_EVAL_54) begin
          if (_EVAL_125) begin
            _EVAL_133 <= _EVAL_72;
          end else begin
            _EVAL_133 <= 6'h0;
          end
        end else begin
          _EVAL_133 <= _EVAL_329;
        end
      end
    end
    if (_EVAL_250) begin
      _EVAL_142 <= _EVAL_9;
    end
    if (_EVAL_250) begin
      _EVAL_161 <= _EVAL;
    end
    if (_EVAL_201) begin
      _EVAL_163 <= _EVAL_2;
    end
    if (_EVAL_12) begin
      _EVAL_171 <= 32'h0;
    end else begin
      if (_EVAL_77) begin
        _EVAL_171 <= 32'h0;
      end else begin
        _EVAL_171 <= _EVAL_176;
      end
    end
    if (_EVAL_12) begin
      _EVAL_227 <= 6'h0;
    end else begin
      if (_EVAL_168) begin
        if (_EVAL_191) begin
          if (_EVAL_125) begin
            _EVAL_227 <= _EVAL_72;
          end else begin
            _EVAL_227 <= 6'h0;
          end
        end else begin
          _EVAL_227 <= _EVAL_146;
        end
      end
    end
    if (_EVAL_12) begin
      _EVAL_231 <= 32'h0;
    end else begin
      _EVAL_231 <= _EVAL_169;
    end
    if (_EVAL_250) begin
      _EVAL_265 <= _EVAL_16;
    end
    if (_EVAL_12) begin
      _EVAL_268 <= 6'h0;
    end else begin
      if (_EVAL_160) begin
        if (_EVAL_190) begin
          if (_EVAL_182) begin
            _EVAL_268 <= _EVAL_75;
          end else begin
            _EVAL_268 <= 6'h0;
          end
        end else begin
          _EVAL_268 <= _EVAL_347;
        end
      end
    end
    if (_EVAL_201) begin
      _EVAL_279 <= _EVAL_3;
    end
    if (_EVAL_12) begin
      _EVAL_285 <= 6'h0;
    end else begin
      if (_EVAL_160) begin
        if (_EVAL_327) begin
          if (_EVAL_182) begin
            _EVAL_285 <= _EVAL_75;
          end else begin
            _EVAL_285 <= 6'h0;
          end
        end else begin
          _EVAL_285 <= _EVAL_234;
        end
      end
    end
    if (_EVAL_201) begin
      _EVAL_311 <= _EVAL_17;
    end
    if (_EVAL_201) begin
      _EVAL_319 <= _EVAL_5;
    end
    if (_EVAL_201) begin
      _EVAL_339 <= _EVAL_7;
    end
    if (_EVAL_250) begin
      _EVAL_344 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a07ddc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cc3dac1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cbf7e08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91ae9c7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_336) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e537a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca4edcc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbbfff61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c82a4c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9ad9ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96dd48ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_336) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c76f185e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(229b0c80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c74c9db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6252)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b295cf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(882be9f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca760424)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_310) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8276e1d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a9fb2f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(555a970c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1163ea4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bca2acc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4189e15b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e81f9356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5099e0a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd3ad708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e1eaf1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c751c757)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(638a3502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29c308f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73f3abab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17b0779e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e106e86b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ee129e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(710e38d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a875fc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2909259)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cffecb78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb16259e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e241b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba6bc78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(764b4eb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1ff4741)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4244f337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f31e343a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dce4d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28056808)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18ebc176)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(359ab8c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(410ab672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4e56bb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf578a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d289a95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b91e7f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ca5c8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8a9b1b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaa62b06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_310) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d24f969)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e78e161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e90adc9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d690eb30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb5ccae0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28903174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ca9bec5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d147e796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea6f07ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9f0886)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(587c6f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4f77a4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f8ca505)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(251b337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c863c7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b900f016)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62eb8917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf074481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c3a475c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4467bc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83291e2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3668dfd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd5cfd33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c26aab02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea1fbb54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2f4c4a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b54e4fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2423657)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64b2e731)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88132a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4416a49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
