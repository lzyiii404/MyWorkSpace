//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_20(
  input  [3:0]  _EVAL,
  output [10:0] _EVAL_0,
  output [31:0] _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  output [7:0]  _EVAL_4,
  output [1:0]  _EVAL_5,
  output        _EVAL_6,
  output [2:0]  _EVAL_7,
  output        _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [7:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  output [3:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  output [3:0]  _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  input  [30:0] _EVAL_22,
  input         _EVAL_23,
  input  [10:0] _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  output        _EVAL_27,
  output [10:0] _EVAL_28,
  input         _EVAL_29,
  input  [31:0] _EVAL_30,
  input  [31:0] _EVAL_31,
  output [10:0] _EVAL_32,
  input         _EVAL_33,
  output        _EVAL_34,
  output [30:0] _EVAL_35,
  output [3:0]  _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  input  [1:0]  _EVAL_39,
  output        _EVAL_40,
  output [3:0]  _EVAL_41,
  input  [3:0]  _EVAL_42,
  input  [10:0] _EVAL_43,
  output        _EVAL_44,
  input         _EVAL_45,
  output [3:0]  _EVAL_46,
  input  [1:0]  _EVAL_47,
  output        _EVAL_48,
  output [1:0]  _EVAL_49,
  output [1:0]  _EVAL_50,
  input  [3:0]  _EVAL_51,
  output [30:0] _EVAL_52,
  output        _EVAL_53,
  output [3:0]  _EVAL_54,
  output [31:0] _EVAL_55,
  output [7:0]  _EVAL_56,
  input  [10:0] _EVAL_57,
  input  [3:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  output [2:0]  _EVAL_60,
  input  [7:0]  _EVAL_61,
  input  [2:0]  _EVAL_62,
  output [3:0]  _EVAL_63,
  output [2:0]  _EVAL_64,
  input         _EVAL_65,
  output        _EVAL_66,
  input  [3:0]  _EVAL_67,
  input  [2:0]  _EVAL_68,
  input  [1:0]  _EVAL_69,
  output [3:0]  _EVAL_70,
  input  [2:0]  _EVAL_71,
  output [1:0]  _EVAL_72,
  input  [10:0] _EVAL_73,
  input  [30:0] _EVAL_74,
  output        _EVAL_75,
  input         _EVAL_76,
  input         _EVAL_77,
  output [2:0]  _EVAL_78,
  input  [3:0]  _EVAL_79,
  input  [1:0]  _EVAL_80,
  input         _EVAL_81,
  output [10:0] _EVAL_82
);
  wire [10:0] Queue_5__EVAL;
  wire  Queue_5__EVAL_0;
  wire [31:0] Queue_5__EVAL_1;
  wire [1:0] Queue_5__EVAL_2;
  wire  Queue_5__EVAL_3;
  wire  Queue_5__EVAL_4;
  wire  Queue_5__EVAL_5;
  wire  Queue_5__EVAL_6;
  wire [31:0] Queue_5__EVAL_7;
  wire  Queue_5__EVAL_8;
  wire [3:0] Queue_5__EVAL_9;
  wire [1:0] Queue_5__EVAL_10;
  wire  Queue_5__EVAL_11;
  wire [10:0] Queue_5__EVAL_12;
  wire [3:0] Queue_5__EVAL_13;
  wire  Queue_5__EVAL_14;
  wire [10:0] Queue_2__EVAL;
  wire  Queue_2__EVAL_0;
  wire [31:0] Queue_2__EVAL_1;
  wire [1:0] Queue_2__EVAL_2;
  wire  Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire  Queue_2__EVAL_5;
  wire  Queue_2__EVAL_6;
  wire [31:0] Queue_2__EVAL_7;
  wire  Queue_2__EVAL_8;
  wire [3:0] Queue_2__EVAL_9;
  wire [1:0] Queue_2__EVAL_10;
  wire  Queue_2__EVAL_11;
  wire [10:0] Queue_2__EVAL_12;
  wire [3:0] Queue_2__EVAL_13;
  wire  Queue_2__EVAL_14;
  wire [10:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire [31:0] Queue_1__EVAL_1;
  wire [1:0] Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire [31:0] Queue_1__EVAL_7;
  wire  Queue_1__EVAL_8;
  wire [3:0] Queue_1__EVAL_9;
  wire [1:0] Queue_1__EVAL_10;
  wire  Queue_1__EVAL_11;
  wire [10:0] Queue_1__EVAL_12;
  wire [3:0] Queue_1__EVAL_13;
  wire  Queue_1__EVAL_14;
  wire [10:0] Queue_4__EVAL;
  wire  Queue_4__EVAL_0;
  wire [31:0] Queue_4__EVAL_1;
  wire [1:0] Queue_4__EVAL_2;
  wire  Queue_4__EVAL_3;
  wire  Queue_4__EVAL_4;
  wire  Queue_4__EVAL_5;
  wire  Queue_4__EVAL_6;
  wire [31:0] Queue_4__EVAL_7;
  wire  Queue_4__EVAL_8;
  wire [3:0] Queue_4__EVAL_9;
  wire [1:0] Queue_4__EVAL_10;
  wire  Queue_4__EVAL_11;
  wire [10:0] Queue_4__EVAL_12;
  wire [3:0] Queue_4__EVAL_13;
  wire  Queue_4__EVAL_14;
  wire [10:0] Queue_7__EVAL;
  wire  Queue_7__EVAL_0;
  wire [31:0] Queue_7__EVAL_1;
  wire [1:0] Queue_7__EVAL_2;
  wire  Queue_7__EVAL_3;
  wire  Queue_7__EVAL_4;
  wire  Queue_7__EVAL_5;
  wire  Queue_7__EVAL_6;
  wire [31:0] Queue_7__EVAL_7;
  wire  Queue_7__EVAL_8;
  wire [3:0] Queue_7__EVAL_9;
  wire [1:0] Queue_7__EVAL_10;
  wire  Queue_7__EVAL_11;
  wire [10:0] Queue_7__EVAL_12;
  wire [3:0] Queue_7__EVAL_13;
  wire  Queue_7__EVAL_14;
  wire [10:0] Queue_6__EVAL;
  wire  Queue_6__EVAL_0;
  wire [31:0] Queue_6__EVAL_1;
  wire [1:0] Queue_6__EVAL_2;
  wire  Queue_6__EVAL_3;
  wire  Queue_6__EVAL_4;
  wire  Queue_6__EVAL_5;
  wire  Queue_6__EVAL_6;
  wire [31:0] Queue_6__EVAL_7;
  wire  Queue_6__EVAL_8;
  wire [3:0] Queue_6__EVAL_9;
  wire [1:0] Queue_6__EVAL_10;
  wire  Queue_6__EVAL_11;
  wire [10:0] Queue_6__EVAL_12;
  wire [3:0] Queue_6__EVAL_13;
  wire  Queue_6__EVAL_14;
  wire [10:0] Queue_3__EVAL;
  wire  Queue_3__EVAL_0;
  wire [31:0] Queue_3__EVAL_1;
  wire [1:0] Queue_3__EVAL_2;
  wire  Queue_3__EVAL_3;
  wire  Queue_3__EVAL_4;
  wire  Queue_3__EVAL_5;
  wire  Queue_3__EVAL_6;
  wire [31:0] Queue_3__EVAL_7;
  wire  Queue_3__EVAL_8;
  wire [3:0] Queue_3__EVAL_9;
  wire [1:0] Queue_3__EVAL_10;
  wire  Queue_3__EVAL_11;
  wire [10:0] Queue_3__EVAL_12;
  wire [3:0] Queue_3__EVAL_13;
  wire  Queue_3__EVAL_14;
  wire [10:0] Queue__EVAL;
  wire  Queue__EVAL_0;
  wire [31:0] Queue__EVAL_1;
  wire [1:0] Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire [31:0] Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire [3:0] Queue__EVAL_9;
  wire [1:0] Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire [10:0] Queue__EVAL_12;
  wire [3:0] Queue__EVAL_13;
  wire  Queue__EVAL_14;
  reg [4:0] _EVAL_201;
  reg [31:0] _RAND_0;
  reg [4:0] _EVAL_263;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_302;
  reg [31:0] _RAND_2;
  reg [4:0] _EVAL_305;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_347;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_348;
  reg [31:0] _RAND_5;
  reg  _EVAL_364;
  reg [31:0] _RAND_6;
  reg [4:0] _EVAL_407;
  reg [31:0] _RAND_7;
  reg [4:0] _EVAL_431;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_451;
  reg [31:0] _RAND_9;
  wire [31:0] _EVAL_375;
  wire [31:0] _EVAL_261;
  wire [31:0] _EVAL_253;
  wire [31:0] _EVAL_352;
  wire [31:0] _EVAL_96;
  wire [31:0] _EVAL_455;
  wire [31:0] _EVAL_137;
  wire [31:0] _EVAL_125;
  wire [31:0] _EVAL_435;
  wire [31:0] _EVAL_121;
  wire [31:0] _EVAL_424;
  wire [31:0] _EVAL_133;
  wire [31:0] _EVAL_427;
  wire [31:0] _EVAL_262;
  wire [31:0] _EVAL_141;
  wire [31:0] _EVAL_324;
  wire [31:0] _EVAL_353;
  wire [31:0] _EVAL_443;
  wire [31:0] _EVAL_393;
  wire [15:0] _EVAL_94;
  wire  _EVAL_145;
  wire  _EVAL_377;
  wire  _EVAL_110;
  wire  _EVAL_441;
  wire  _EVAL_350;
  wire  _EVAL_317;
  wire  _EVAL_360;
  wire  _EVAL_139;
  wire  _EVAL_135;
  wire  _EVAL_105;
  wire  _EVAL_430;
  wire  _EVAL_390;
  wire  _EVAL_276;
  wire  _EVAL_99;
  wire  _EVAL_374;
  wire  _EVAL_178;
  wire  _EVAL_298;
  wire  _EVAL_97;
  wire  _EVAL_362;
  wire  _EVAL_299;
  wire  _EVAL_90;
  wire  _EVAL_208;
  wire  _EVAL_337;
  wire  _EVAL_397;
  wire  _EVAL_164;
  wire  _EVAL_416;
  wire  _EVAL_207;
  wire [4:0] _EVAL_402;
  wire [4:0] _EVAL_93;
  wire [15:0] _EVAL_138;
  wire  _EVAL_351;
  wire  _EVAL_391;
  wire  _EVAL_192;
  wire  _EVAL_368;
  wire  _EVAL_366;
  wire  _EVAL_274;
  wire  _EVAL_232;
  wire  _EVAL_161;
  wire  _EVAL_421;
  wire  _EVAL_149;
  wire  _EVAL_383;
  wire  _EVAL_84;
  wire  _EVAL_381;
  wire  _EVAL_411;
  wire  _EVAL_220;
  wire  _EVAL_156;
  wire  _EVAL_289;
  wire  _EVAL_426;
  wire  _EVAL_296;
  wire  _EVAL_420;
  wire  _EVAL_425;
  wire  _EVAL_211;
  wire  _EVAL_365;
  wire  _EVAL_268;
  wire  _EVAL_338;
  wire  _EVAL_242;
  wire  _EVAL_331;
  wire [4:0] _EVAL_131;
  wire [4:0] _EVAL_184;
  wire  _EVAL_234;
  wire [31:0] _EVAL_256;
  wire [31:0] _EVAL_114;
  wire  _EVAL_303;
  wire  _EVAL_323;
  wire  _EVAL_342;
  wire  _EVAL_444;
  wire  _EVAL_270;
  wire  _EVAL_180;
  wire  _EVAL_422;
  wire  _EVAL_372;
  wire [4:0] _EVAL_226;
  wire [4:0] _EVAL_91;
  wire  _EVAL_206;
  wire  _EVAL_132;
  wire  _EVAL_328;
  wire [4:0] _EVAL_450;
  wire [4:0] _EVAL_209;
  wire  _EVAL_442;
  wire [4:0] _EVAL_129;
  wire [4:0] _EVAL_388;
  wire  _EVAL_314;
  wire  _EVAL_147;
  wire  _EVAL_439;
  wire [4:0] _EVAL_406;
  wire [4:0] _EVAL_225;
  wire  _EVAL_310;
  wire  _EVAL_446;
  wire  _EVAL_290;
  wire  _EVAL_230;
  wire [4:0] _EVAL_130;
  wire [4:0] _EVAL_239;
  wire  _EVAL_171;
  wire  _EVAL_126;
  wire  _EVAL_238;
  wire [4:0] _EVAL_85;
  wire [4:0] _EVAL_399;
  wire  _EVAL_152;
  wire  _EVAL_437;
  wire [4:0] _EVAL_370;
  wire [4:0] _EVAL_200;
  wire  _EVAL_240;
  wire  _EVAL_387;
  wire  _EVAL_186;
  wire [4:0] _EVAL_144;
  wire [4:0] _EVAL_326;
  wire  _EVAL_396;
  wire  _EVAL_354;
  wire  _EVAL_282;
  wire  _EVAL_334;
  wire [4:0] _EVAL_409;
  wire [4:0] _EVAL_359;
  wire  _EVAL_449;
  wire  _EVAL_166;
  wire  _EVAL_107;
  wire [4:0] _EVAL_321;
  wire [4:0] _EVAL_394;
  wire  _EVAL_101;
  wire  _EVAL_143;
  wire  _EVAL_349;
  wire  _EVAL_384;
  wire [4:0] _EVAL_122;
  wire [4:0] _EVAL_241;
  wire  _EVAL_332;
  wire  _EVAL_408;
  wire  _EVAL_357;
  wire [4:0] _EVAL_254;
  wire [4:0] _EVAL_404;
  wire  _EVAL_313;
  wire  _EVAL_188;
  wire  _EVAL_116;
  wire  _EVAL_300;
  wire [4:0] _EVAL_369;
  wire [4:0] _EVAL_403;
  wire  _EVAL_223;
  wire  _EVAL_410;
  wire  _EVAL_340;
  wire [4:0] _EVAL_136;
  wire [4:0] _EVAL_320;
  wire  _EVAL_285;
  wire [15:0] _EVAL_280;
  wire [16:0] _EVAL_378;
  wire [15:0] _EVAL_284;
  wire [15:0] _EVAL_355;
  wire [17:0] _EVAL_405;
  wire [15:0] _EVAL_89;
  wire [15:0] _EVAL_198;
  wire [19:0] _EVAL_273;
  wire [15:0] _EVAL_356;
  wire [15:0] _EVAL_423;
  wire [23:0] _EVAL_127;
  wire [15:0] _EVAL_189;
  wire [15:0] _EVAL_215;
  wire [16:0] _EVAL_336;
  wire [16:0] _EVAL_214;
  wire [16:0] _EVAL_327;
  wire [16:0] _EVAL_271;
  wire  _EVAL_237;
  wire [15:0] _EVAL_119;
  wire [15:0] _EVAL_429;
  wire [15:0] _EVAL_386;
  wire [7:0] _EVAL_217;
  wire [7:0] _EVAL_150;
  wire [7:0] _EVAL_447;
  wire [3:0] _EVAL_176;
  wire [3:0] _EVAL_218;
  wire [3:0] _EVAL_181;
  wire [1:0] _EVAL_177;
  wire  _EVAL_438;
  wire [3:0] _EVAL_109;
  wire [3:0] _EVAL_168;
  wire [3:0] _EVAL_295;
  wire [3:0] _EVAL_115;
  wire [3:0] _EVAL_108;
  wire [3:0] _EVAL_293;
  wire [3:0] _EVAL_245;
  wire [10:0] _EVAL_255;
  wire [10:0] _EVAL_452;
  wire [10:0] _EVAL_316;
  wire [10:0] _EVAL_222;
  wire [10:0] _EVAL_249;
  wire [10:0] _EVAL_281;
  wire [10:0] _EVAL_124;
  wire  _EVAL_371;
  wire  _EVAL_160;
  wire  _EVAL_92;
  wire  _EVAL_202;
  wire  _EVAL_229;
  wire [1:0] _EVAL_221;
  wire [1:0] _EVAL_413;
  wire  _EVAL_395;
  wire [4:0] _EVAL_236;
  wire [4:0] _EVAL_278;
  wire [10:0] _EVAL_419;
  wire [10:0] _EVAL_260;
  wire [10:0] _EVAL_345;
  wire [10:0] _EVAL_190;
  wire [10:0] _EVAL_418;
  wire [10:0] _EVAL_247;
  wire [10:0] _EVAL_227;
  wire [10:0] _EVAL_311;
  wire [10:0] _EVAL_159;
  wire [10:0] _EVAL_155;
  wire [10:0] _EVAL_257;
  wire [10:0] _EVAL_194;
  wire [10:0] _EVAL_318;
  wire [10:0] _EVAL_179;
  wire [3:0] _EVAL_283;
  wire [3:0] _EVAL_172;
  wire [3:0] _EVAL_264;
  wire [3:0] _EVAL_219;
  wire [3:0] _EVAL_306;
  wire [3:0] _EVAL_197;
  wire [3:0] _EVAL_251;
  wire [3:0] _EVAL_297;
  wire [3:0] _EVAL_205;
  wire [3:0] _EVAL_191;
  wire [3:0] _EVAL_100;
  wire [3:0] _EVAL_210;
  wire [1:0] _EVAL_286;
  wire [1:0] _EVAL_432;
  wire [1:0] _EVAL_165;
  wire [1:0] _EVAL_330;
  wire [1:0] _EVAL_275;
  wire [1:0] _EVAL_106;
  wire [1:0] _EVAL_319;
  wire [1:0] _EVAL_346;
  wire [1:0] _EVAL_380;
  wire [1:0] _EVAL_183;
  wire [1:0] _EVAL_454;
  wire [1:0] _EVAL_233;
  wire [1:0] _EVAL_134;
  wire [1:0] _EVAL_162;
  wire [1:0] _EVAL_307;
  wire [1:0] _EVAL_98;
  wire [1:0] _EVAL_412;
  wire [1:0] _EVAL_367;
  wire [31:0] _EVAL_175;
  wire [1:0] _EVAL_140;
  wire [1:0] _EVAL_301;
  wire [1:0] _EVAL_158;
  wire  _EVAL_203;
  wire [10:0] _EVAL_102;
  wire [3:0] _EVAL_228;
  wire [3:0] _EVAL_287;
  wire [3:0] _EVAL_248;
  wire [1:0] _EVAL_434;
  SiFive__EVAL_19 Queue_5 (
    ._EVAL(Queue_5__EVAL),
    ._EVAL_0(Queue_5__EVAL_0),
    ._EVAL_1(Queue_5__EVAL_1),
    ._EVAL_2(Queue_5__EVAL_2),
    ._EVAL_3(Queue_5__EVAL_3),
    ._EVAL_4(Queue_5__EVAL_4),
    ._EVAL_5(Queue_5__EVAL_5),
    ._EVAL_6(Queue_5__EVAL_6),
    ._EVAL_7(Queue_5__EVAL_7),
    ._EVAL_8(Queue_5__EVAL_8),
    ._EVAL_9(Queue_5__EVAL_9),
    ._EVAL_10(Queue_5__EVAL_10),
    ._EVAL_11(Queue_5__EVAL_11),
    ._EVAL_12(Queue_5__EVAL_12),
    ._EVAL_13(Queue_5__EVAL_13),
    ._EVAL_14(Queue_5__EVAL_14)
  );
  SiFive__EVAL_19 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6),
    ._EVAL_7(Queue_2__EVAL_7),
    ._EVAL_8(Queue_2__EVAL_8),
    ._EVAL_9(Queue_2__EVAL_9),
    ._EVAL_10(Queue_2__EVAL_10),
    ._EVAL_11(Queue_2__EVAL_11),
    ._EVAL_12(Queue_2__EVAL_12),
    ._EVAL_13(Queue_2__EVAL_13),
    ._EVAL_14(Queue_2__EVAL_14)
  );
  SiFive__EVAL_19 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14)
  );
  SiFive__EVAL_19 Queue_4 (
    ._EVAL(Queue_4__EVAL),
    ._EVAL_0(Queue_4__EVAL_0),
    ._EVAL_1(Queue_4__EVAL_1),
    ._EVAL_2(Queue_4__EVAL_2),
    ._EVAL_3(Queue_4__EVAL_3),
    ._EVAL_4(Queue_4__EVAL_4),
    ._EVAL_5(Queue_4__EVAL_5),
    ._EVAL_6(Queue_4__EVAL_6),
    ._EVAL_7(Queue_4__EVAL_7),
    ._EVAL_8(Queue_4__EVAL_8),
    ._EVAL_9(Queue_4__EVAL_9),
    ._EVAL_10(Queue_4__EVAL_10),
    ._EVAL_11(Queue_4__EVAL_11),
    ._EVAL_12(Queue_4__EVAL_12),
    ._EVAL_13(Queue_4__EVAL_13),
    ._EVAL_14(Queue_4__EVAL_14)
  );
  SiFive__EVAL_19 Queue_7 (
    ._EVAL(Queue_7__EVAL),
    ._EVAL_0(Queue_7__EVAL_0),
    ._EVAL_1(Queue_7__EVAL_1),
    ._EVAL_2(Queue_7__EVAL_2),
    ._EVAL_3(Queue_7__EVAL_3),
    ._EVAL_4(Queue_7__EVAL_4),
    ._EVAL_5(Queue_7__EVAL_5),
    ._EVAL_6(Queue_7__EVAL_6),
    ._EVAL_7(Queue_7__EVAL_7),
    ._EVAL_8(Queue_7__EVAL_8),
    ._EVAL_9(Queue_7__EVAL_9),
    ._EVAL_10(Queue_7__EVAL_10),
    ._EVAL_11(Queue_7__EVAL_11),
    ._EVAL_12(Queue_7__EVAL_12),
    ._EVAL_13(Queue_7__EVAL_13),
    ._EVAL_14(Queue_7__EVAL_14)
  );
  SiFive__EVAL_19 Queue_6 (
    ._EVAL(Queue_6__EVAL),
    ._EVAL_0(Queue_6__EVAL_0),
    ._EVAL_1(Queue_6__EVAL_1),
    ._EVAL_2(Queue_6__EVAL_2),
    ._EVAL_3(Queue_6__EVAL_3),
    ._EVAL_4(Queue_6__EVAL_4),
    ._EVAL_5(Queue_6__EVAL_5),
    ._EVAL_6(Queue_6__EVAL_6),
    ._EVAL_7(Queue_6__EVAL_7),
    ._EVAL_8(Queue_6__EVAL_8),
    ._EVAL_9(Queue_6__EVAL_9),
    ._EVAL_10(Queue_6__EVAL_10),
    ._EVAL_11(Queue_6__EVAL_11),
    ._EVAL_12(Queue_6__EVAL_12),
    ._EVAL_13(Queue_6__EVAL_13),
    ._EVAL_14(Queue_6__EVAL_14)
  );
  SiFive__EVAL_19 Queue_3 (
    ._EVAL(Queue_3__EVAL),
    ._EVAL_0(Queue_3__EVAL_0),
    ._EVAL_1(Queue_3__EVAL_1),
    ._EVAL_2(Queue_3__EVAL_2),
    ._EVAL_3(Queue_3__EVAL_3),
    ._EVAL_4(Queue_3__EVAL_4),
    ._EVAL_5(Queue_3__EVAL_5),
    ._EVAL_6(Queue_3__EVAL_6),
    ._EVAL_7(Queue_3__EVAL_7),
    ._EVAL_8(Queue_3__EVAL_8),
    ._EVAL_9(Queue_3__EVAL_9),
    ._EVAL_10(Queue_3__EVAL_10),
    ._EVAL_11(Queue_3__EVAL_11),
    ._EVAL_12(Queue_3__EVAL_12),
    ._EVAL_13(Queue_3__EVAL_13),
    ._EVAL_14(Queue_3__EVAL_14)
  );
  SiFive__EVAL_19 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14)
  );
  assign _EVAL_375 = Queue_7__EVAL_1;
  assign _EVAL_261 = Queue_6__EVAL_1;
  assign _EVAL_253 = Queue_5__EVAL_1;
  assign _EVAL_352 = Queue_4__EVAL_1;
  assign _EVAL_96 = Queue_3__EVAL_1;
  assign _EVAL_455 = Queue_2__EVAL_1;
  assign _EVAL_137 = Queue_1__EVAL_1;
  assign _EVAL_125 = Queue__EVAL_1;
  assign _EVAL_435 = 4'h1 == _EVAL_451 ? _EVAL_137 : _EVAL_125;
  assign _EVAL_121 = 4'h2 == _EVAL_451 ? _EVAL_455 : _EVAL_435;
  assign _EVAL_424 = 4'h3 == _EVAL_451 ? _EVAL_96 : _EVAL_121;
  assign _EVAL_133 = 4'h4 == _EVAL_451 ? _EVAL_352 : _EVAL_424;
  assign _EVAL_427 = 4'h5 == _EVAL_451 ? _EVAL_253 : _EVAL_133;
  assign _EVAL_262 = 4'h6 == _EVAL_451 ? _EVAL_261 : _EVAL_427;
  assign _EVAL_141 = 4'h7 == _EVAL_451 ? _EVAL_375 : _EVAL_262;
  assign _EVAL_324 = 4'h8 == _EVAL_451 ? 32'h0 : _EVAL_141;
  assign _EVAL_353 = 4'h9 == _EVAL_451 ? 32'h0 : _EVAL_324;
  assign _EVAL_443 = 4'ha == _EVAL_451 ? 32'h0 : _EVAL_353;
  assign _EVAL_393 = 4'hb == _EVAL_451 ? 32'h0 : _EVAL_443;
  assign _EVAL_94 = 16'h1 << _EVAL_58;
  assign _EVAL_145 = _EVAL_94[0];
  assign _EVAL_377 = Queue_7__EVAL_4;
  assign _EVAL_110 = Queue_6__EVAL_4;
  assign _EVAL_441 = Queue_5__EVAL_4;
  assign _EVAL_350 = Queue_4__EVAL_4;
  assign _EVAL_317 = Queue_3__EVAL_4;
  assign _EVAL_360 = Queue_2__EVAL_4;
  assign _EVAL_139 = Queue_1__EVAL_4;
  assign _EVAL_135 = Queue__EVAL_4;
  assign _EVAL_105 = 4'h1 == _EVAL_58 ? _EVAL_139 : _EVAL_135;
  assign _EVAL_430 = 4'h2 == _EVAL_58 ? _EVAL_360 : _EVAL_105;
  assign _EVAL_390 = 4'h3 == _EVAL_58 ? _EVAL_317 : _EVAL_430;
  assign _EVAL_276 = 4'h4 == _EVAL_58 ? _EVAL_350 : _EVAL_390;
  assign _EVAL_99 = 4'h5 == _EVAL_58 ? _EVAL_441 : _EVAL_276;
  assign _EVAL_374 = 4'h6 == _EVAL_58 ? _EVAL_110 : _EVAL_99;
  assign _EVAL_178 = 4'h7 == _EVAL_58 ? _EVAL_377 : _EVAL_374;
  assign _EVAL_298 = 4'h8 == _EVAL_58 ? 1'h0 : _EVAL_178;
  assign _EVAL_97 = 4'h9 == _EVAL_58 ? 1'h0 : _EVAL_298;
  assign _EVAL_362 = 4'ha == _EVAL_58 ? 1'h0 : _EVAL_97;
  assign _EVAL_299 = 4'hb == _EVAL_58 ? 1'h0 : _EVAL_362;
  assign _EVAL_90 = 4'hc == _EVAL_58 ? 1'h0 : _EVAL_299;
  assign _EVAL_208 = 4'hd == _EVAL_58 ? 1'h0 : _EVAL_90;
  assign _EVAL_337 = 4'he == _EVAL_58 ? 1'h0 : _EVAL_208;
  assign _EVAL_397 = 4'hf == _EVAL_58 ? 1'h0 : _EVAL_337;
  assign _EVAL_164 = _EVAL_397 & _EVAL_23;
  assign _EVAL_416 = _EVAL_145 & _EVAL_164;
  assign _EVAL_207 = _EVAL_416 & _EVAL_45;
  assign _EVAL_402 = {{4'd0}, _EVAL_207};
  assign _EVAL_93 = _EVAL_263 + _EVAL_402;
  assign _EVAL_138 = 16'h1 << _EVAL_451;
  assign _EVAL_351 = _EVAL_138[0];
  assign _EVAL_391 = _EVAL_25 & _EVAL_364;
  assign _EVAL_192 = _EVAL_351 & _EVAL_391;
  assign _EVAL_368 = Queue_7__EVAL_5;
  assign _EVAL_366 = Queue_6__EVAL_5;
  assign _EVAL_274 = Queue_5__EVAL_5;
  assign _EVAL_232 = Queue_4__EVAL_5;
  assign _EVAL_161 = Queue_3__EVAL_5;
  assign _EVAL_421 = Queue_2__EVAL_5;
  assign _EVAL_149 = Queue_1__EVAL_5;
  assign _EVAL_383 = Queue__EVAL_5;
  assign _EVAL_84 = 4'h1 == _EVAL_451 ? _EVAL_149 : _EVAL_383;
  assign _EVAL_381 = 4'h2 == _EVAL_451 ? _EVAL_421 : _EVAL_84;
  assign _EVAL_411 = 4'h3 == _EVAL_451 ? _EVAL_161 : _EVAL_381;
  assign _EVAL_220 = 4'h4 == _EVAL_451 ? _EVAL_232 : _EVAL_411;
  assign _EVAL_156 = 4'h5 == _EVAL_451 ? _EVAL_274 : _EVAL_220;
  assign _EVAL_289 = 4'h6 == _EVAL_451 ? _EVAL_366 : _EVAL_156;
  assign _EVAL_426 = 4'h7 == _EVAL_451 ? _EVAL_368 : _EVAL_289;
  assign _EVAL_296 = 4'h8 == _EVAL_451 ? 1'h0 : _EVAL_426;
  assign _EVAL_420 = 4'h9 == _EVAL_451 ? 1'h0 : _EVAL_296;
  assign _EVAL_425 = 4'ha == _EVAL_451 ? 1'h0 : _EVAL_420;
  assign _EVAL_211 = 4'hb == _EVAL_451 ? 1'h0 : _EVAL_425;
  assign _EVAL_365 = 4'hc == _EVAL_451 ? 1'h0 : _EVAL_211;
  assign _EVAL_268 = 4'hd == _EVAL_451 ? 1'h0 : _EVAL_365;
  assign _EVAL_338 = 4'he == _EVAL_451 ? 1'h0 : _EVAL_268;
  assign _EVAL_242 = 4'hf == _EVAL_451 ? 1'h0 : _EVAL_338;
  assign _EVAL_331 = _EVAL_192 & _EVAL_242;
  assign _EVAL_131 = {{4'd0}, _EVAL_331};
  assign _EVAL_184 = _EVAL_93 - _EVAL_131;
  assign _EVAL_234 = _EVAL_184 != 5'h0;
  assign _EVAL_256 = 4'hc == _EVAL_451 ? 32'h0 : _EVAL_393;
  assign _EVAL_114 = 4'hd == _EVAL_451 ? 32'h0 : _EVAL_256;
  assign _EVAL_303 = _EVAL_94[4];
  assign _EVAL_323 = _EVAL_303 & _EVAL_164;
  assign _EVAL_342 = _EVAL_94[6];
  assign _EVAL_444 = _EVAL_342 & _EVAL_164;
  assign _EVAL_270 = _EVAL_444 & _EVAL_45;
  assign _EVAL_180 = _EVAL_94[7];
  assign _EVAL_422 = _EVAL_180 & _EVAL_164;
  assign _EVAL_372 = _EVAL_422 & _EVAL_45;
  assign _EVAL_226 = {{4'd0}, _EVAL_372};
  assign _EVAL_91 = _EVAL_347 + _EVAL_226;
  assign _EVAL_206 = _EVAL_138[7];
  assign _EVAL_132 = _EVAL_206 & _EVAL_391;
  assign _EVAL_328 = _EVAL_132 & _EVAL_242;
  assign _EVAL_450 = {{4'd0}, _EVAL_328};
  assign _EVAL_209 = _EVAL_91 - _EVAL_450;
  assign _EVAL_442 = _EVAL_209 != 5'h0;
  assign _EVAL_129 = {{4'd0}, _EVAL_270};
  assign _EVAL_388 = _EVAL_201 + _EVAL_129;
  assign _EVAL_314 = _EVAL_138[6];
  assign _EVAL_147 = _EVAL_314 & _EVAL_391;
  assign _EVAL_439 = _EVAL_147 & _EVAL_242;
  assign _EVAL_406 = {{4'd0}, _EVAL_439};
  assign _EVAL_225 = _EVAL_388 - _EVAL_406;
  assign _EVAL_310 = _EVAL_225 != 5'h0;
  assign _EVAL_446 = _EVAL_94[5];
  assign _EVAL_290 = _EVAL_446 & _EVAL_164;
  assign _EVAL_230 = _EVAL_290 & _EVAL_45;
  assign _EVAL_130 = {{4'd0}, _EVAL_230};
  assign _EVAL_239 = _EVAL_407 + _EVAL_130;
  assign _EVAL_171 = _EVAL_138[5];
  assign _EVAL_126 = _EVAL_171 & _EVAL_391;
  assign _EVAL_238 = _EVAL_126 & _EVAL_242;
  assign _EVAL_85 = {{4'd0}, _EVAL_238};
  assign _EVAL_399 = _EVAL_239 - _EVAL_85;
  assign _EVAL_152 = _EVAL_399 != 5'h0;
  assign _EVAL_437 = _EVAL_323 & _EVAL_45;
  assign _EVAL_370 = {{4'd0}, _EVAL_437};
  assign _EVAL_200 = _EVAL_305 + _EVAL_370;
  assign _EVAL_240 = _EVAL_138[4];
  assign _EVAL_387 = _EVAL_240 & _EVAL_391;
  assign _EVAL_186 = _EVAL_387 & _EVAL_242;
  assign _EVAL_144 = {{4'd0}, _EVAL_186};
  assign _EVAL_326 = _EVAL_200 - _EVAL_144;
  assign _EVAL_396 = _EVAL_326 != 5'h0;
  assign _EVAL_354 = _EVAL_94[3];
  assign _EVAL_282 = _EVAL_354 & _EVAL_164;
  assign _EVAL_334 = _EVAL_282 & _EVAL_45;
  assign _EVAL_409 = {{4'd0}, _EVAL_334};
  assign _EVAL_359 = _EVAL_348 + _EVAL_409;
  assign _EVAL_449 = _EVAL_138[3];
  assign _EVAL_166 = _EVAL_449 & _EVAL_391;
  assign _EVAL_107 = _EVAL_166 & _EVAL_242;
  assign _EVAL_321 = {{4'd0}, _EVAL_107};
  assign _EVAL_394 = _EVAL_359 - _EVAL_321;
  assign _EVAL_101 = _EVAL_394 != 5'h0;
  assign _EVAL_143 = _EVAL_94[2];
  assign _EVAL_349 = _EVAL_143 & _EVAL_164;
  assign _EVAL_384 = _EVAL_349 & _EVAL_45;
  assign _EVAL_122 = {{4'd0}, _EVAL_384};
  assign _EVAL_241 = _EVAL_302 + _EVAL_122;
  assign _EVAL_332 = _EVAL_138[2];
  assign _EVAL_408 = _EVAL_332 & _EVAL_391;
  assign _EVAL_357 = _EVAL_408 & _EVAL_242;
  assign _EVAL_254 = {{4'd0}, _EVAL_357};
  assign _EVAL_404 = _EVAL_241 - _EVAL_254;
  assign _EVAL_313 = _EVAL_404 != 5'h0;
  assign _EVAL_188 = _EVAL_94[1];
  assign _EVAL_116 = _EVAL_188 & _EVAL_164;
  assign _EVAL_300 = _EVAL_116 & _EVAL_45;
  assign _EVAL_369 = {{4'd0}, _EVAL_300};
  assign _EVAL_403 = _EVAL_431 + _EVAL_369;
  assign _EVAL_223 = _EVAL_138[1];
  assign _EVAL_410 = _EVAL_223 & _EVAL_391;
  assign _EVAL_340 = _EVAL_410 & _EVAL_242;
  assign _EVAL_136 = {{4'd0}, _EVAL_340};
  assign _EVAL_320 = _EVAL_403 - _EVAL_136;
  assign _EVAL_285 = _EVAL_320 != 5'h0;
  assign _EVAL_280 = {8'h0,_EVAL_442,_EVAL_310,_EVAL_152,_EVAL_396,_EVAL_101,_EVAL_313,_EVAL_285,_EVAL_234};
  assign _EVAL_378 = {_EVAL_280, 1'h0};
  assign _EVAL_284 = _EVAL_378[15:0];
  assign _EVAL_355 = _EVAL_280 | _EVAL_284;
  assign _EVAL_405 = {_EVAL_355, 2'h0};
  assign _EVAL_89 = _EVAL_405[15:0];
  assign _EVAL_198 = _EVAL_355 | _EVAL_89;
  assign _EVAL_273 = {_EVAL_198, 4'h0};
  assign _EVAL_356 = _EVAL_273[15:0];
  assign _EVAL_423 = _EVAL_198 | _EVAL_356;
  assign _EVAL_127 = {_EVAL_423, 8'h0};
  assign _EVAL_189 = _EVAL_127[15:0];
  assign _EVAL_215 = _EVAL_423 | _EVAL_189;
  assign _EVAL_336 = {{1'd0}, _EVAL_280};
  assign _EVAL_214 = {_EVAL_215, 1'h0};
  assign _EVAL_327 = ~ _EVAL_214;
  assign _EVAL_271 = _EVAL_336 & _EVAL_327;
  assign _EVAL_237 = _EVAL_271[16];
  assign _EVAL_119 = {{15'd0}, _EVAL_237};
  assign _EVAL_429 = _EVAL_271[15:0];
  assign _EVAL_386 = _EVAL_119 | _EVAL_429;
  assign _EVAL_217 = _EVAL_386[15:8];
  assign _EVAL_150 = _EVAL_386[7:0];
  assign _EVAL_447 = _EVAL_217 | _EVAL_150;
  assign _EVAL_176 = _EVAL_447[7:4];
  assign _EVAL_218 = _EVAL_447[3:0];
  assign _EVAL_181 = _EVAL_176 | _EVAL_218;
  assign _EVAL_177 = _EVAL_181[3:2];
  assign _EVAL_438 = _EVAL_364 == 1'h0;
  assign _EVAL_109 = Queue_3__EVAL_13;
  assign _EVAL_168 = Queue_2__EVAL_13;
  assign _EVAL_295 = Queue_1__EVAL_13;
  assign _EVAL_115 = Queue__EVAL_13;
  assign _EVAL_108 = 4'h1 == _EVAL_451 ? _EVAL_295 : _EVAL_115;
  assign _EVAL_293 = 4'h2 == _EVAL_451 ? _EVAL_168 : _EVAL_108;
  assign _EVAL_245 = 4'h3 == _EVAL_451 ? _EVAL_109 : _EVAL_293;
  assign _EVAL_255 = Queue_3__EVAL;
  assign _EVAL_452 = Queue_2__EVAL;
  assign _EVAL_316 = Queue_1__EVAL;
  assign _EVAL_222 = Queue__EVAL;
  assign _EVAL_249 = 4'h1 == _EVAL_451 ? _EVAL_316 : _EVAL_222;
  assign _EVAL_281 = 4'h2 == _EVAL_451 ? _EVAL_452 : _EVAL_249;
  assign _EVAL_124 = 4'h3 == _EVAL_451 ? _EVAL_255 : _EVAL_281;
  assign _EVAL_371 = _EVAL_391 & _EVAL_242;
  assign _EVAL_160 = _EVAL_438 | _EVAL_371;
  assign _EVAL_92 = _EVAL_217 != 8'h0;
  assign _EVAL_202 = _EVAL_176 != 4'h0;
  assign _EVAL_229 = _EVAL_177 != 2'h0;
  assign _EVAL_221 = _EVAL_181[1:0];
  assign _EVAL_413 = _EVAL_177 | _EVAL_221;
  assign _EVAL_395 = _EVAL_413[1];
  assign _EVAL_236 = {_EVAL_237,_EVAL_92,_EVAL_202,_EVAL_229,_EVAL_395};
  assign _EVAL_278 = _EVAL_160 ? _EVAL_236 : {{1'd0}, _EVAL_451};
  assign _EVAL_419 = Queue_7__EVAL;
  assign _EVAL_260 = Queue_6__EVAL;
  assign _EVAL_345 = Queue_5__EVAL;
  assign _EVAL_190 = Queue_4__EVAL;
  assign _EVAL_418 = 4'h4 == _EVAL_451 ? _EVAL_190 : _EVAL_124;
  assign _EVAL_247 = 4'h5 == _EVAL_451 ? _EVAL_345 : _EVAL_418;
  assign _EVAL_227 = 4'h6 == _EVAL_451 ? _EVAL_260 : _EVAL_247;
  assign _EVAL_311 = 4'h7 == _EVAL_451 ? _EVAL_419 : _EVAL_227;
  assign _EVAL_159 = 4'h8 == _EVAL_451 ? 11'h0 : _EVAL_311;
  assign _EVAL_155 = 4'h9 == _EVAL_451 ? 11'h0 : _EVAL_159;
  assign _EVAL_257 = 4'ha == _EVAL_451 ? 11'h0 : _EVAL_155;
  assign _EVAL_194 = 4'hb == _EVAL_451 ? 11'h0 : _EVAL_257;
  assign _EVAL_318 = 4'hc == _EVAL_451 ? 11'h0 : _EVAL_194;
  assign _EVAL_179 = 4'hd == _EVAL_451 ? 11'h0 : _EVAL_318;
  assign _EVAL_283 = Queue_7__EVAL_13;
  assign _EVAL_172 = Queue_6__EVAL_13;
  assign _EVAL_264 = Queue_5__EVAL_13;
  assign _EVAL_219 = Queue_4__EVAL_13;
  assign _EVAL_306 = 4'h4 == _EVAL_451 ? _EVAL_219 : _EVAL_245;
  assign _EVAL_197 = 4'h5 == _EVAL_451 ? _EVAL_264 : _EVAL_306;
  assign _EVAL_251 = 4'h6 == _EVAL_451 ? _EVAL_172 : _EVAL_197;
  assign _EVAL_297 = 4'h7 == _EVAL_451 ? _EVAL_283 : _EVAL_251;
  assign _EVAL_205 = 4'h8 == _EVAL_451 ? 4'h0 : _EVAL_297;
  assign _EVAL_191 = 4'h9 == _EVAL_451 ? 4'h0 : _EVAL_205;
  assign _EVAL_100 = 4'ha == _EVAL_451 ? 4'h0 : _EVAL_191;
  assign _EVAL_210 = 4'hb == _EVAL_451 ? 4'h0 : _EVAL_100;
  assign _EVAL_286 = Queue_4__EVAL_10;
  assign _EVAL_432 = Queue_7__EVAL_10;
  assign _EVAL_165 = Queue_6__EVAL_10;
  assign _EVAL_330 = Queue_5__EVAL_10;
  assign _EVAL_275 = Queue_3__EVAL_10;
  assign _EVAL_106 = Queue_2__EVAL_10;
  assign _EVAL_319 = Queue_1__EVAL_10;
  assign _EVAL_346 = Queue__EVAL_10;
  assign _EVAL_380 = 4'h1 == _EVAL_451 ? _EVAL_319 : _EVAL_346;
  assign _EVAL_183 = 4'h2 == _EVAL_451 ? _EVAL_106 : _EVAL_380;
  assign _EVAL_454 = 4'h3 == _EVAL_451 ? _EVAL_275 : _EVAL_183;
  assign _EVAL_233 = 4'h4 == _EVAL_451 ? _EVAL_286 : _EVAL_454;
  assign _EVAL_134 = 4'h5 == _EVAL_451 ? _EVAL_330 : _EVAL_233;
  assign _EVAL_162 = 4'h6 == _EVAL_451 ? _EVAL_165 : _EVAL_134;
  assign _EVAL_307 = 4'h7 == _EVAL_451 ? _EVAL_432 : _EVAL_162;
  assign _EVAL_98 = 4'h8 == _EVAL_451 ? 2'h0 : _EVAL_307;
  assign _EVAL_412 = 4'h9 == _EVAL_451 ? 2'h0 : _EVAL_98;
  assign _EVAL_367 = 4'ha == _EVAL_451 ? 2'h0 : _EVAL_412;
  assign _EVAL_175 = 4'he == _EVAL_451 ? 32'h0 : _EVAL_114;
  assign _EVAL_140 = 4'hb == _EVAL_451 ? 2'h0 : _EVAL_367;
  assign _EVAL_301 = 4'hc == _EVAL_451 ? 2'h0 : _EVAL_140;
  assign _EVAL_158 = 4'hd == _EVAL_451 ? 2'h0 : _EVAL_301;
  assign _EVAL_203 = _EVAL_280 != 16'h0;
  assign _EVAL_102 = 4'he == _EVAL_451 ? 11'h0 : _EVAL_179;
  assign _EVAL_228 = 4'hc == _EVAL_451 ? 4'h0 : _EVAL_210;
  assign _EVAL_287 = 4'hd == _EVAL_451 ? 4'h0 : _EVAL_228;
  assign _EVAL_248 = 4'he == _EVAL_451 ? 4'h0 : _EVAL_287;
  assign _EVAL_434 = 4'he == _EVAL_451 ? 2'h0 : _EVAL_158;
  assign Queue_4__EVAL_7 = _EVAL_31;
  assign Queue_2__EVAL_8 = _EVAL_3;
  assign _EVAL_4 = _EVAL_10;
  assign Queue_4__EVAL_8 = _EVAL_3;
  assign Queue_7__EVAL_6 = _EVAL_180 & _EVAL_23;
  assign Queue_2__EVAL_9 = _EVAL_58;
  assign Queue_7__EVAL_2 = _EVAL_39;
  assign Queue_5__EVAL_6 = _EVAL_446 & _EVAL_23;
  assign _EVAL_0 = 4'hf == _EVAL_451 ? 11'h0 : _EVAL_102;
  assign _EVAL_53 = _EVAL_65;
  assign Queue_7__EVAL_8 = _EVAL_3;
  assign Queue_3__EVAL_12 = _EVAL_73;
  assign Queue__EVAL_3 = _EVAL_45;
  assign Queue_6__EVAL_8 = _EVAL_3;
  assign Queue_6__EVAL_12 = _EVAL_73;
  assign Queue_2__EVAL_6 = _EVAL_143 & _EVAL_23;
  assign Queue_1__EVAL_8 = _EVAL_3;
  assign Queue_6__EVAL_2 = _EVAL_39;
  assign Queue_2__EVAL_2 = _EVAL_39;
  assign Queue_6__EVAL_0 = _EVAL_314 & _EVAL_391;
  assign _EVAL_54 = _EVAL_67;
  assign _EVAL_50 = _EVAL_69;
  assign _EVAL_52 = _EVAL_22;
  assign Queue_2__EVAL_12 = _EVAL_73;
  assign Queue_6__EVAL_7 = _EVAL_31;
  assign _EVAL_28 = _EVAL_43;
  assign _EVAL_2 = _EVAL_26;
  assign _EVAL_36 = _EVAL_11;
  assign _EVAL_6 = _EVAL_364;
  assign _EVAL_32 = _EVAL_24;
  assign Queue_4__EVAL_2 = _EVAL_39;
  assign Queue_7__EVAL_3 = _EVAL_45;
  assign _EVAL_5 = _EVAL_47;
  assign Queue_5__EVAL_7 = _EVAL_31;
  assign _EVAL_70 = _EVAL_17;
  assign Queue_5__EVAL_2 = _EVAL_39;
  assign _EVAL_41 = 4'hf == _EVAL_451 ? 4'h0 : _EVAL_248;
  assign Queue_3__EVAL_6 = _EVAL_354 & _EVAL_23;
  assign Queue_7__EVAL_9 = _EVAL_58;
  assign Queue_4__EVAL_9 = _EVAL_58;
  assign Queue_4__EVAL_11 = _EVAL_76;
  assign _EVAL_7 = _EVAL_71;
  assign _EVAL_1 = _EVAL_30;
  assign _EVAL_44 = 4'hf == _EVAL_58 ? 1'h0 : _EVAL_337;
  assign _EVAL_75 = _EVAL_16;
  assign Queue_1__EVAL_9 = _EVAL_58;
  assign Queue_3__EVAL_0 = _EVAL_449 & _EVAL_391;
  assign Queue_4__EVAL_12 = _EVAL_73;
  assign Queue_5__EVAL_8 = _EVAL_3;
  assign _EVAL_14 = _EVAL_51;
  assign Queue__EVAL_12 = _EVAL_73;
  assign Queue_2__EVAL_11 = _EVAL_76;
  assign Queue_4__EVAL_3 = _EVAL_45;
  assign Queue_3__EVAL_3 = _EVAL_45;
  assign Queue_6__EVAL_6 = _EVAL_342 & _EVAL_23;
  assign Queue_4__EVAL_6 = _EVAL_303 & _EVAL_23;
  assign Queue_3__EVAL_2 = _EVAL_39;
  assign Queue_6__EVAL_3 = _EVAL_45;
  assign Queue__EVAL_2 = _EVAL_39;
  assign Queue_1__EVAL_11 = _EVAL_76;
  assign _EVAL_82 = _EVAL_57;
  assign Queue__EVAL_9 = _EVAL_58;
  assign _EVAL_60 = _EVAL_62;
  assign _EVAL_20 = _EVAL_15;
  assign Queue_7__EVAL_7 = _EVAL_31;
  assign Queue_6__EVAL_11 = _EVAL_76;
  assign _EVAL_40 = 4'hf == _EVAL_451 ? 1'h0 : _EVAL_338;
  assign Queue_1__EVAL_0 = _EVAL_223 & _EVAL_391;
  assign Queue_5__EVAL_9 = _EVAL_58;
  assign Queue_6__EVAL_9 = _EVAL_58;
  assign Queue_1__EVAL_7 = _EVAL_31;
  assign _EVAL_38 = _EVAL_12;
  assign Queue_5__EVAL_11 = _EVAL_76;
  assign _EVAL_8 = _EVAL_81;
  assign _EVAL_49 = _EVAL_80;
  assign _EVAL_59 = _EVAL;
  assign Queue__EVAL_0 = _EVAL_351 & _EVAL_391;
  assign _EVAL_66 = _EVAL_29;
  assign Queue__EVAL_8 = _EVAL_3;
  assign Queue_2__EVAL_3 = _EVAL_45;
  assign Queue_5__EVAL_3 = _EVAL_45;
  assign _EVAL_72 = 4'hf == _EVAL_451 ? 2'h0 : _EVAL_434;
  assign Queue__EVAL_11 = _EVAL_76;
  assign Queue_3__EVAL_9 = _EVAL_58;
  assign _EVAL_55 = 4'hf == _EVAL_451 ? 32'h0 : _EVAL_175;
  assign Queue_1__EVAL_3 = _EVAL_45;
  assign _EVAL_27 = _EVAL_33;
  assign Queue__EVAL_6 = _EVAL_145 & _EVAL_23;
  assign _EVAL_37 = _EVAL_19;
  assign Queue_3__EVAL_7 = _EVAL_31;
  assign Queue_5__EVAL_12 = _EVAL_73;
  assign Queue_3__EVAL_8 = _EVAL_3;
  assign _EVAL_48 = _EVAL_21;
  assign _EVAL_64 = _EVAL_9;
  assign Queue_2__EVAL_7 = _EVAL_31;
  assign _EVAL_56 = _EVAL_61;
  assign _EVAL_78 = _EVAL_68;
  assign _EVAL_18 = _EVAL_79;
  assign Queue_3__EVAL_11 = _EVAL_76;
  assign _EVAL_46 = _EVAL_13;
  assign Queue_1__EVAL_6 = _EVAL_188 & _EVAL_23;
  assign Queue_7__EVAL_11 = _EVAL_76;
  assign Queue_7__EVAL_12 = _EVAL_73;
  assign _EVAL_35 = _EVAL_74;
  assign Queue_7__EVAL_0 = _EVAL_206 & _EVAL_391;
  assign Queue_4__EVAL_0 = _EVAL_240 & _EVAL_391;
  assign Queue_2__EVAL_0 = _EVAL_332 & _EVAL_391;
  assign Queue__EVAL_7 = _EVAL_31;
  assign Queue_1__EVAL_12 = _EVAL_73;
  assign Queue_5__EVAL_0 = _EVAL_171 & _EVAL_391;
  assign _EVAL_34 = _EVAL_77;
  assign _EVAL_63 = _EVAL_42;
  assign Queue_1__EVAL_2 = _EVAL_39;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_201 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_263 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_302 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_305 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_347 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_348 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_364 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_407 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_431 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_451 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_76) begin
      _EVAL_201 <= 5'h0;
    end else begin
      _EVAL_201 <= _EVAL_225;
    end
    if (_EVAL_76) begin
      _EVAL_263 <= 5'h0;
    end else begin
      _EVAL_263 <= _EVAL_184;
    end
    if (_EVAL_76) begin
      _EVAL_302 <= 5'h0;
    end else begin
      _EVAL_302 <= _EVAL_404;
    end
    if (_EVAL_76) begin
      _EVAL_305 <= 5'h0;
    end else begin
      _EVAL_305 <= _EVAL_326;
    end
    if (_EVAL_76) begin
      _EVAL_347 <= 5'h0;
    end else begin
      _EVAL_347 <= _EVAL_209;
    end
    if (_EVAL_76) begin
      _EVAL_348 <= 5'h0;
    end else begin
      _EVAL_348 <= _EVAL_394;
    end
    if (_EVAL_76) begin
      _EVAL_364 <= 1'h0;
    end else begin
      if (_EVAL_160) begin
        _EVAL_364 <= _EVAL_203;
      end
    end
    if (_EVAL_76) begin
      _EVAL_407 <= 5'h0;
    end else begin
      _EVAL_407 <= _EVAL_399;
    end
    if (_EVAL_76) begin
      _EVAL_431 <= 5'h0;
    end else begin
      _EVAL_431 <= _EVAL_320;
    end
    _EVAL_451 <= _EVAL_278[3:0];
  end
endmodule
