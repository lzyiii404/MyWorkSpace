//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_250_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input  [24:0] _EVAL_3,
  input  [7:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [7:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_39;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_92;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_115;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_153;
  reg [31:0] _RAND_3;
  reg [7:0] _EVAL_156;
  reg [31:0] _RAND_4;
  reg [31:0] _EVAL_181;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_201;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_223;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_227;
  reg [31:0] _RAND_8;
  reg [24:0] _EVAL_230;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_241;
  reg [31:0] _RAND_10;
  reg [7:0] _EVAL_266;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_281;
  reg [31:0] _RAND_12;
  reg [135:0] _EVAL_301;
  reg [159:0] _RAND_13;
  wire  _EVAL_233;
  wire [4:0] _EVAL_276;
  wire  _EVAL_206;
  wire [24:0] _EVAL_22;
  wire [25:0] _EVAL_297;
  wire [25:0] _EVAL_46;
  wire [2:0] _EVAL_205;
  wire [25:0] _EVAL_106;
  wire  _EVAL_200;
  wire  _EVAL_255;
  wire  _EVAL_175;
  wire  _EVAL_254;
  wire  _EVAL_277;
  wire  _EVAL_237;
  wire  _EVAL_17;
  wire  _EVAL_167;
  wire [4:0] _EVAL_26;
  wire  _EVAL_179;
  wire  _EVAL_134;
  wire [1:0] _EVAL_129;
  wire [1:0] _EVAL_32;
  wire  _EVAL_78;
  wire  _EVAL_303;
  wire  _EVAL_216;
  wire  _EVAL_114;
  wire  _EVAL_79;
  wire  _EVAL_256;
  wire  _EVAL_23;
  wire  _EVAL_66;
  wire [255:0] _EVAL_75;
  wire [255:0] _EVAL_211;
  wire [135:0] _EVAL_183;
  wire [135:0] _EVAL_300;
  wire  _EVAL_267;
  wire  _EVAL_251;
  wire  _EVAL_70;
  wire  _EVAL_212;
  wire  _EVAL_52;
  wire  _EVAL_15;
  wire [255:0] _EVAL_18;
  wire [255:0] _EVAL_187;
  wire [135:0] _EVAL_27;
  wire [135:0] _EVAL_264;
  wire [135:0] _EVAL_172;
  wire  _EVAL_118;
  wire  _EVAL_173;
  wire  _EVAL_109;
  wire  _EVAL_126;
  wire  _EVAL_108;
  wire  _EVAL_76;
  wire  _EVAL_294;
  wire  _EVAL_272;
  wire  _EVAL_143;
  wire  _EVAL_215;
  wire  _EVAL_157;
  wire  _EVAL_219;
  wire  _EVAL_38;
  wire  _EVAL_99;
  wire  _EVAL_213;
  wire  _EVAL_304;
  wire  _EVAL_51;
  wire  _EVAL_194;
  wire  _EVAL_105;
  wire  _EVAL_121;
  wire  _EVAL_204;
  wire  _EVAL_16;
  wire  _EVAL_77;
  wire [12:0] _EVAL_226;
  wire [5:0] _EVAL_25;
  wire [5:0] _EVAL_148;
  wire [3:0] _EVAL_189;
  wire [3:0] _EVAL_142;
  wire  _EVAL_130;
  wire  _EVAL_90;
  wire  _EVAL_265;
  wire  _EVAL_138;
  wire  _EVAL_73;
  wire  _EVAL_147;
  wire  _EVAL_299;
  wire  _EVAL_69;
  wire [135:0] _EVAL_29;
  wire  _EVAL_222;
  wire  _EVAL_199;
  wire  _EVAL_152;
  wire  _EVAL_31;
  wire  _EVAL_101;
  wire  _EVAL_214;
  wire  _EVAL_195;
  wire  _EVAL_269;
  wire  _EVAL_136;
  wire  _EVAL_43;
  wire  _EVAL_244;
  wire  _EVAL_182;
  wire  _EVAL_111;
  wire  _EVAL_74;
  wire  _EVAL_224;
  wire  _EVAL_278;
  wire  _EVAL_135;
  wire  _EVAL_61;
  wire [3:0] _EVAL_280;
  wire  _EVAL_252;
  wire  _EVAL_170;
  wire [3:0] _EVAL_287;
  wire  _EVAL_56;
  wire  _EVAL_117;
  wire  _EVAL_58;
  wire  _EVAL_178;
  wire [2:0] _EVAL_41;
  wire  _EVAL_273;
  wire  _EVAL_84;
  wire  _EVAL_235;
  wire  _EVAL_293;
  wire  _EVAL_295;
  wire  _EVAL_98;
  wire  _EVAL_275;
  wire  _EVAL_296;
  wire  _EVAL_85;
  wire  _EVAL_112;
  wire  _EVAL_232;
  wire  _EVAL_144;
  wire  _EVAL_80;
  wire  _EVAL_124;
  wire  _EVAL_229;
  wire  _EVAL_190;
  wire  _EVAL_250;
  wire  _EVAL_208;
  wire [3:0] _EVAL_174;
  wire  _EVAL_193;
  wire  _EVAL_171;
  wire  _EVAL_47;
  wire  _EVAL_63;
  wire [31:0] _EVAL_72;
  wire [135:0] _EVAL_128;
  wire [135:0] _EVAL_95;
  wire  _EVAL_261;
  wire  _EVAL_21;
  wire  _EVAL_59;
  wire  _EVAL_139;
  wire  _EVAL_209;
  wire  _EVAL_28;
  wire  _EVAL_288;
  wire  _EVAL_197;
  wire [3:0] _EVAL_104;
  wire  _EVAL_91;
  wire  _EVAL_253;
  wire  _EVAL_202;
  wire  _EVAL_113;
  wire  _EVAL_225;
  wire  _EVAL_48;
  wire  _EVAL_176;
  wire [3:0] _EVAL_50;
  wire [3:0] _EVAL_68;
  wire  _EVAL_107;
  wire  _EVAL_158;
  wire  _EVAL_282;
  wire  _EVAL_218;
  wire  _EVAL_236;
  wire  _EVAL_247;
  wire  _EVAL_274;
  wire  _EVAL_164;
  wire  _EVAL_65;
  wire  _EVAL_151;
  wire  _EVAL_86;
  wire  _EVAL_119;
  wire  _EVAL_150;
  wire  _EVAL_145;
  wire  _EVAL_163;
  wire  _EVAL_246;
  wire  _EVAL_166;
  wire [12:0] _EVAL_283;
  wire [5:0] _EVAL_198;
  wire [5:0] _EVAL_184;
  wire [3:0] _EVAL_291;
  wire  _EVAL_160;
  wire  _EVAL_165;
  wire  _EVAL_97;
  wire  _EVAL_238;
  wire  _EVAL_243;
  wire  _EVAL_83;
  wire  _EVAL_185;
  wire [24:0] _EVAL_55;
  wire [24:0] _EVAL_240;
  wire  _EVAL_257;
  wire  _EVAL_54;
  wire  _EVAL_123;
  wire  _EVAL_44;
  wire  _EVAL_140;
  wire  _EVAL_188;
  wire  _EVAL_149;
  wire  _EVAL_290;
  wire  _EVAL_220;
  wire  _EVAL_289;
  wire  _EVAL_60;
  wire  _EVAL_34;
  wire  _EVAL_207;
  wire  _EVAL_62;
  wire  _EVAL_96;
  wire  _EVAL_53;
  wire  _EVAL_67;
  wire  _EVAL_103;
  wire  _EVAL_42;
  wire  _EVAL_191;
  wire  _EVAL_137;
  wire [3:0] _EVAL_217;
  wire  _EVAL_125;
  wire  _EVAL_93;
  wire  _EVAL_180;
  wire  _EVAL_177;
  wire  _EVAL_49;
  wire  _EVAL_19;
  wire  _EVAL_120;
  wire  _EVAL_196;
  wire  _EVAL_258;
  wire  _EVAL_245;
  wire  _EVAL_57;
  wire  _EVAL_186;
  wire  _EVAL_110;
  wire  _EVAL_221;
  wire  _EVAL_81;
  wire  _EVAL_284;
  wire  _EVAL_155;
  wire  _EVAL_89;
  wire  _EVAL_20;
  wire  _EVAL_162;
  wire  _EVAL_231;
  wire  _EVAL_203;
  wire  _EVAL_285;
  wire  _EVAL_141;
  wire  _EVAL_279;
  wire  _EVAL_260;
  wire  _EVAL_154;
  wire  _EVAL_228;
  wire  _EVAL_146;
  wire  _EVAL_292;
  wire  _EVAL_263;
  wire  _EVAL_159;
  wire  _EVAL_210;
  wire  _EVAL_33;
  wire  _EVAL_192;
  wire  _EVAL_100;
  wire  _EVAL_286;
  wire  _EVAL_37;
  wire  _EVAL_122;
  wire  _EVAL_259;
  wire  _EVAL_116;
  wire  _EVAL_40;
  wire  _EVAL_169;
  wire  _EVAL_24;
  wire  _EVAL_64;
  wire  _EVAL_35;
  wire  _EVAL_102;
  wire  _EVAL_30;
  wire  _EVAL_302;
  wire  _EVAL_87;
  wire  _EVAL_239;
  wire  _EVAL_36;
  wire  _EVAL_248;
  wire  _EVAL_45;
  wire  _EVAL_132;
  wire  _EVAL_94;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_233 = _EVAL_8 == 1'h0;
  assign _EVAL_276 = _EVAL_9[7:3];
  assign _EVAL_206 = _EVAL_276 == 5'h3;
  assign _EVAL_22 = _EVAL_3 ^ 25'h1900000;
  assign _EVAL_297 = {1'b0,$signed(_EVAL_22)};
  assign _EVAL_46 = $signed(_EVAL_297) & $signed(-26'sh2000);
  assign _EVAL_205 = _EVAL_4[2:0];
  assign _EVAL_106 = $signed(_EVAL_46);
  assign _EVAL_200 = _EVAL_4 == 8'h40;
  assign _EVAL_255 = 3'h6 == _EVAL_11;
  assign _EVAL_175 = _EVAL_200 ? _EVAL_255 : 1'h0;
  assign _EVAL_254 = _EVAL_4 == 8'h80;
  assign _EVAL_277 = _EVAL_254 ? _EVAL_255 : 1'h0;
  assign _EVAL_237 = _EVAL_175 | _EVAL_277;
  assign _EVAL_17 = _EVAL_237 | _EVAL_1;
  assign _EVAL_167 = _EVAL_17 == 1'h0;
  assign _EVAL_26 = _EVAL_4[7:3];
  assign _EVAL_179 = _EVAL_26 == 5'h1;
  assign _EVAL_134 = _EVAL_11[0];
  assign _EVAL_129 = 2'h1 << _EVAL_134;
  assign _EVAL_32 = _EVAL_129 | 2'h1;
  assign _EVAL_78 = _EVAL_32[0];
  assign _EVAL_303 = _EVAL_3[1];
  assign _EVAL_216 = _EVAL_3[0];
  assign _EVAL_114 = _EVAL_303 & _EVAL_216;
  assign _EVAL_79 = _EVAL_78 & _EVAL_114;
  assign _EVAL_256 = _EVAL & _EVAL_6;
  assign _EVAL_23 = _EVAL_227 == 4'h0;
  assign _EVAL_66 = _EVAL_256 & _EVAL_23;
  assign _EVAL_75 = 256'h1 << _EVAL_4;
  assign _EVAL_211 = _EVAL_66 ? _EVAL_75 : 256'h0;
  assign _EVAL_183 = _EVAL_211[135:0];
  assign _EVAL_300 = _EVAL_301 | _EVAL_183;
  assign _EVAL_267 = _EVAL_5 & _EVAL_13;
  assign _EVAL_251 = _EVAL_241 == 4'h0;
  assign _EVAL_70 = _EVAL_267 & _EVAL_251;
  assign _EVAL_212 = _EVAL_0 == 3'h6;
  assign _EVAL_52 = _EVAL_212 == 1'h0;
  assign _EVAL_15 = _EVAL_70 & _EVAL_52;
  assign _EVAL_18 = 256'h1 << _EVAL_9;
  assign _EVAL_187 = _EVAL_15 ? _EVAL_18 : 256'h0;
  assign _EVAL_27 = _EVAL_187[135:0];
  assign _EVAL_264 = ~ _EVAL_27;
  assign _EVAL_172 = _EVAL_300 & _EVAL_264;
  assign _EVAL_118 = _EVAL_4 == 8'h48;
  assign _EVAL_173 = _EVAL_118 | _EVAL_200;
  assign _EVAL_109 = _EVAL_26 == 5'h8;
  assign _EVAL_126 = 3'h1 <= _EVAL_205;
  assign _EVAL_108 = _EVAL_109 & _EVAL_126;
  assign _EVAL_76 = _EVAL_173 | _EVAL_108;
  assign _EVAL_294 = _EVAL_4 == 8'h20;
  assign _EVAL_272 = _EVAL_76 | _EVAL_294;
  assign _EVAL_143 = _EVAL_26 == 5'h0;
  assign _EVAL_215 = _EVAL_272 | _EVAL_143;
  assign _EVAL_157 = _EVAL_215 | _EVAL_179;
  assign _EVAL_219 = _EVAL_26 == 5'h2;
  assign _EVAL_38 = _EVAL_157 | _EVAL_219;
  assign _EVAL_99 = _EVAL_26 == 5'h3;
  assign _EVAL_213 = _EVAL_38 | _EVAL_99;
  assign _EVAL_304 = _EVAL_213 | _EVAL_254;
  assign _EVAL_51 = _EVAL_26 == 5'h10;
  assign _EVAL_194 = _EVAL_51 & _EVAL_126;
  assign _EVAL_105 = _EVAL_304 | _EVAL_194;
  assign _EVAL_121 = _EVAL_105 | _EVAL_1;
  assign _EVAL_204 = _EVAL_121 == 1'h0;
  assign _EVAL_16 = _EVAL_7[2];
  assign _EVAL_77 = _EVAL_16 == 1'h0;
  assign _EVAL_226 = 13'h3f << _EVAL_11;
  assign _EVAL_25 = _EVAL_226[5:0];
  assign _EVAL_148 = ~ _EVAL_25;
  assign _EVAL_189 = _EVAL_148[5:2];
  assign _EVAL_142 = _EVAL_227 - 4'h1;
  assign _EVAL_130 = _EVAL_11 == _EVAL_223;
  assign _EVAL_90 = _EVAL_7 == 3'h6;
  assign _EVAL_265 = _EVAL_6 & _EVAL_90;
  assign _EVAL_138 = _EVAL_183 != _EVAL_27;
  assign _EVAL_73 = _EVAL_183 != 136'h0;
  assign _EVAL_147 = _EVAL_73 == 1'h0;
  assign _EVAL_299 = _EVAL_138 | _EVAL_147;
  assign _EVAL_69 = _EVAL_256 | _EVAL_267;
  assign _EVAL_29 = _EVAL_301 >> _EVAL_4;
  assign _EVAL_222 = _EVAL_11 >= 3'h2;
  assign _EVAL_199 = _EVAL_32[1];
  assign _EVAL_152 = _EVAL_199 & _EVAL_303;
  assign _EVAL_31 = _EVAL_222 | _EVAL_152;
  assign _EVAL_101 = _EVAL_31 | _EVAL_79;
  assign _EVAL_214 = _EVAL_216 == 1'h0;
  assign _EVAL_195 = _EVAL_303 & _EVAL_214;
  assign _EVAL_269 = _EVAL_78 & _EVAL_195;
  assign _EVAL_136 = _EVAL_31 | _EVAL_269;
  assign _EVAL_43 = _EVAL_303 == 1'h0;
  assign _EVAL_244 = _EVAL_199 & _EVAL_43;
  assign _EVAL_182 = _EVAL_222 | _EVAL_244;
  assign _EVAL_111 = _EVAL_43 & _EVAL_216;
  assign _EVAL_74 = _EVAL_78 & _EVAL_111;
  assign _EVAL_224 = _EVAL_182 | _EVAL_74;
  assign _EVAL_278 = _EVAL_43 & _EVAL_214;
  assign _EVAL_135 = _EVAL_78 & _EVAL_278;
  assign _EVAL_61 = _EVAL_182 | _EVAL_135;
  assign _EVAL_280 = {_EVAL_101,_EVAL_136,_EVAL_224,_EVAL_61};
  assign _EVAL_252 = _EVAL_2 == _EVAL_280;
  assign _EVAL_170 = _EVAL_252 | _EVAL_1;
  assign _EVAL_287 = _EVAL_153 - 4'h1;
  assign _EVAL_56 = _EVAL_9 == 8'h48;
  assign _EVAL_117 = _EVAL_9 == 8'h40;
  assign _EVAL_58 = _EVAL_56 | _EVAL_117;
  assign _EVAL_178 = _EVAL_276 == 5'h8;
  assign _EVAL_41 = _EVAL_9[2:0];
  assign _EVAL_273 = 3'h1 <= _EVAL_41;
  assign _EVAL_84 = _EVAL_178 & _EVAL_273;
  assign _EVAL_235 = _EVAL_58 | _EVAL_84;
  assign _EVAL_293 = _EVAL_9 == 8'h20;
  assign _EVAL_295 = _EVAL_235 | _EVAL_293;
  assign _EVAL_98 = _EVAL_276 == 5'h0;
  assign _EVAL_275 = _EVAL_295 | _EVAL_98;
  assign _EVAL_296 = _EVAL_276 == 5'h1;
  assign _EVAL_85 = _EVAL_275 | _EVAL_296;
  assign _EVAL_112 = _EVAL_276 == 5'h2;
  assign _EVAL_232 = _EVAL_85 | _EVAL_112;
  assign _EVAL_144 = _EVAL_232 | _EVAL_206;
  assign _EVAL_80 = _EVAL_9 == 8'h80;
  assign _EVAL_124 = _EVAL_144 | _EVAL_80;
  assign _EVAL_229 = _EVAL_276 == 5'h10;
  assign _EVAL_190 = _EVAL_229 & _EVAL_273;
  assign _EVAL_250 = _EVAL_124 | _EVAL_190;
  assign _EVAL_208 = _EVAL_250 | _EVAL_1;
  assign _EVAL_174 = ~ _EVAL_2;
  assign _EVAL_193 = _EVAL_174 == 4'h0;
  assign _EVAL_171 = _EVAL_193 | _EVAL_1;
  assign _EVAL_47 = _EVAL_171 == 1'h0;
  assign _EVAL_63 = _EVAL_233 | _EVAL_1;
  assign _EVAL_72 = _EVAL_181 + 32'h1;
  assign _EVAL_128 = _EVAL_183 | _EVAL_301;
  assign _EVAL_95 = _EVAL_128 >> _EVAL_9;
  assign _EVAL_261 = _EVAL_95[0];
  assign _EVAL_21 = _EVAL_261 | _EVAL_1;
  assign _EVAL_59 = _EVAL_153 == 4'h0;
  assign _EVAL_139 = _EVAL_267 & _EVAL_59;
  assign _EVAL_209 = _EVAL_7 == 3'h4;
  assign _EVAL_28 = _EVAL_6 & _EVAL_209;
  assign _EVAL_288 = _EVAL_12 == _EVAL_201;
  assign _EVAL_197 = _EVAL_115 == 4'h0;
  assign _EVAL_104 = _EVAL_115 - 4'h1;
  assign _EVAL_91 = _EVAL_301 != 136'h0;
  assign _EVAL_253 = _EVAL_91 == 1'h0;
  assign _EVAL_202 = _EVAL_10 == _EVAL_281;
  assign _EVAL_113 = _EVAL_202 | _EVAL_1;
  assign _EVAL_225 = _EVAL_113 == 1'h0;
  assign _EVAL_48 = _EVAL_0 == _EVAL_92;
  assign _EVAL_176 = _EVAL_7 == 3'h3;
  assign _EVAL_50 = ~ _EVAL_280;
  assign _EVAL_68 = _EVAL_2 & _EVAL_50;
  assign _EVAL_107 = _EVAL_68 == 4'h0;
  assign _EVAL_158 = _EVAL_107 | _EVAL_1;
  assign _EVAL_282 = _EVAL_11 <= 3'h6;
  assign _EVAL_218 = _EVAL_10 >= 3'h2;
  assign _EVAL_236 = _EVAL_218 | _EVAL_1;
  assign _EVAL_247 = _EVAL_4 == _EVAL_266;
  assign _EVAL_274 = _EVAL_29[0];
  assign _EVAL_164 = _EVAL_274 == 1'h0;
  assign _EVAL_65 = _EVAL_164 | _EVAL_1;
  assign _EVAL_151 = _EVAL_65 == 1'h0;
  assign _EVAL_86 = _EVAL_3 == _EVAL_230;
  assign _EVAL_119 = _EVAL_86 | _EVAL_1;
  assign _EVAL_150 = _EVAL_299 | _EVAL_1;
  assign _EVAL_145 = _EVAL_150 == 1'h0;
  assign _EVAL_163 = _EVAL_13 & _EVAL_212;
  assign _EVAL_246 = _EVAL_0 == 3'h5;
  assign _EVAL_166 = _EVAL_0[0];
  assign _EVAL_283 = 13'h3f << _EVAL_10;
  assign _EVAL_198 = _EVAL_283[5:0];
  assign _EVAL_184 = ~ _EVAL_198;
  assign _EVAL_291 = _EVAL_184[5:2];
  assign _EVAL_160 = _EVAL_0 == 3'h4;
  assign _EVAL_165 = _EVAL_119 == 1'h0;
  assign _EVAL_97 = _EVAL_170 == 1'h0;
  assign _EVAL_238 = _EVAL_48 | _EVAL_1;
  assign _EVAL_243 = _EVAL_238 == 1'h0;
  assign _EVAL_83 = plusarg_reader_out == 32'h0;
  assign _EVAL_185 = _EVAL_253 | _EVAL_83;
  assign _EVAL_55 = {{19'd0}, _EVAL_148};
  assign _EVAL_240 = _EVAL_3 & _EVAL_55;
  assign _EVAL_257 = _EVAL_240 == 25'h0;
  assign _EVAL_54 = _EVAL_257 | _EVAL_1;
  assign _EVAL_123 = _EVAL_54 == 1'h0;
  assign _EVAL_44 = _EVAL_12 <= 3'h2;
  assign _EVAL_140 = _EVAL_44 | _EVAL_1;
  assign _EVAL_188 = _EVAL_140 == 1'h0;
  assign _EVAL_149 = $signed(_EVAL_106) == $signed(26'sh0);
  assign _EVAL_290 = _EVAL_11 <= 3'h2;
  assign _EVAL_220 = _EVAL_290 & _EVAL_149;
  assign _EVAL_289 = _EVAL_220 | _EVAL_1;
  assign _EVAL_60 = _EVAL_289 == 1'h0;
  assign _EVAL_34 = _EVAL_0 <= 3'h6;
  assign _EVAL_207 = _EVAL_1 == 1'h0;
  assign _EVAL_62 = _EVAL_6 & _EVAL_176;
  assign _EVAL_96 = _EVAL_0 == 3'h2;
  assign _EVAL_53 = _EVAL_13 & _EVAL_96;
  assign _EVAL_67 = _EVAL_247 | _EVAL_1;
  assign _EVAL_103 = _EVAL_67 == 1'h0;
  assign _EVAL_42 = _EVAL_12 == 3'h0;
  assign _EVAL_191 = _EVAL_42 | _EVAL_1;
  assign _EVAL_137 = _EVAL_191 == 1'h0;
  assign _EVAL_217 = _EVAL_241 - 4'h1;
  assign _EVAL_125 = _EVAL_181 < plusarg_reader_out;
  assign _EVAL_93 = _EVAL_130 | _EVAL_1;
  assign _EVAL_180 = _EVAL_222 | _EVAL_1;
  assign _EVAL_177 = _EVAL_180 == 1'h0;
  assign _EVAL_49 = _EVAL_288 | _EVAL_1;
  assign _EVAL_19 = _EVAL_49 == 1'h0;
  assign _EVAL_120 = _EVAL_21 == 1'h0;
  assign _EVAL_196 = _EVAL_7 == 3'h7;
  assign _EVAL_258 = _EVAL_6 & _EVAL_196;
  assign _EVAL_245 = _EVAL_0 == 3'h0;
  assign _EVAL_57 = _EVAL_12 <= 3'h4;
  assign _EVAL_186 = _EVAL_57 | _EVAL_1;
  assign _EVAL_110 = _EVAL_7 == _EVAL_39;
  assign _EVAL_221 = _EVAL_110 | _EVAL_1;
  assign _EVAL_81 = _EVAL_9 == _EVAL_156;
  assign _EVAL_284 = _EVAL_256 & _EVAL_197;
  assign _EVAL_155 = _EVAL_197 == 1'h0;
  assign _EVAL_89 = _EVAL_6 & _EVAL_155;
  assign _EVAL_20 = _EVAL_59 == 1'h0;
  assign _EVAL_162 = _EVAL_282 & _EVAL_149;
  assign _EVAL_231 = _EVAL_162 | _EVAL_1;
  assign _EVAL_203 = _EVAL_231 == 1'h0;
  assign _EVAL_285 = _EVAL_7 == 3'h1;
  assign _EVAL_141 = _EVAL_185 | _EVAL_125;
  assign _EVAL_279 = _EVAL_141 | _EVAL_1;
  assign _EVAL_260 = _EVAL_279 == 1'h0;
  assign _EVAL_154 = _EVAL_12 <= 3'h3;
  assign _EVAL_228 = _EVAL_154 | _EVAL_1;
  assign _EVAL_146 = _EVAL_0 == 3'h1;
  assign _EVAL_292 = _EVAL_13 & _EVAL_146;
  assign _EVAL_263 = _EVAL_34 | _EVAL_1;
  assign _EVAL_159 = _EVAL_6 & _EVAL_285;
  assign _EVAL_210 = _EVAL_208 == 1'h0;
  assign _EVAL_33 = _EVAL_13 & _EVAL_160;
  assign _EVAL_192 = _EVAL_7 == 3'h5;
  assign _EVAL_100 = _EVAL_6 & _EVAL_192;
  assign _EVAL_286 = _EVAL_7 == 3'h0;
  assign _EVAL_37 = _EVAL_6 & _EVAL_286;
  assign _EVAL_122 = _EVAL_236 == 1'h0;
  assign _EVAL_259 = _EVAL_13 & _EVAL_20;
  assign _EVAL_116 = _EVAL_12 != 3'h0;
  assign _EVAL_40 = _EVAL_7 == 3'h2;
  assign _EVAL_169 = _EVAL_116 | _EVAL_1;
  assign _EVAL_24 = _EVAL_13 & _EVAL_245;
  assign _EVAL_64 = _EVAL_158 == 1'h0;
  assign _EVAL_35 = _EVAL_228 == 1'h0;
  assign _EVAL_102 = _EVAL_186 == 1'h0;
  assign _EVAL_30 = _EVAL_93 == 1'h0;
  assign _EVAL_302 = _EVAL_13 & _EVAL_246;
  assign _EVAL_87 = _EVAL_169 == 1'h0;
  assign _EVAL_239 = _EVAL_263 == 1'h0;
  assign _EVAL_36 = _EVAL_63 == 1'h0;
  assign _EVAL_248 = _EVAL_81 | _EVAL_1;
  assign _EVAL_45 = _EVAL_248 == 1'h0;
  assign _EVAL_132 = _EVAL_6 & _EVAL_40;
  assign _EVAL_94 = _EVAL_221 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_39 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_92 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_115 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_153 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_156 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_181 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_201 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_223 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_227 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_230 = _RAND_9[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_241 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_266 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_281 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {5{`RANDOM}};
  _EVAL_301 = _RAND_13[135:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL_284) begin
      _EVAL_39 <= _EVAL_7;
    end
    if (_EVAL_139) begin
      _EVAL_92 <= _EVAL_0;
    end
    if (_EVAL_1) begin
      _EVAL_115 <= 4'h0;
    end else begin
      if (_EVAL_256) begin
        if (_EVAL_197) begin
          if (_EVAL_77) begin
            _EVAL_115 <= _EVAL_189;
          end else begin
            _EVAL_115 <= 4'h0;
          end
        end else begin
          _EVAL_115 <= _EVAL_104;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_153 <= 4'h0;
    end else begin
      if (_EVAL_267) begin
        if (_EVAL_59) begin
          if (_EVAL_166) begin
            _EVAL_153 <= _EVAL_291;
          end else begin
            _EVAL_153 <= 4'h0;
          end
        end else begin
          _EVAL_153 <= _EVAL_287;
        end
      end
    end
    if (_EVAL_139) begin
      _EVAL_156 <= _EVAL_9;
    end
    if (_EVAL_1) begin
      _EVAL_181 <= 32'h0;
    end else begin
      if (_EVAL_69) begin
        _EVAL_181 <= 32'h0;
      end else begin
        _EVAL_181 <= _EVAL_72;
      end
    end
    if (_EVAL_284) begin
      _EVAL_201 <= _EVAL_12;
    end
    if (_EVAL_284) begin
      _EVAL_223 <= _EVAL_11;
    end
    if (_EVAL_1) begin
      _EVAL_227 <= 4'h0;
    end else begin
      if (_EVAL_256) begin
        if (_EVAL_23) begin
          if (_EVAL_77) begin
            _EVAL_227 <= _EVAL_189;
          end else begin
            _EVAL_227 <= 4'h0;
          end
        end else begin
          _EVAL_227 <= _EVAL_142;
        end
      end
    end
    if (_EVAL_284) begin
      _EVAL_230 <= _EVAL_3;
    end
    if (_EVAL_1) begin
      _EVAL_241 <= 4'h0;
    end else begin
      if (_EVAL_267) begin
        if (_EVAL_251) begin
          if (_EVAL_166) begin
            _EVAL_241 <= _EVAL_291;
          end else begin
            _EVAL_241 <= 4'h0;
          end
        end else begin
          _EVAL_241 <= _EVAL_217;
        end
      end
    end
    if (_EVAL_284) begin
      _EVAL_266 <= _EVAL_4;
    end
    if (_EVAL_139) begin
      _EVAL_281 <= _EVAL_10;
    end
    if (_EVAL_1) begin
      _EVAL_301 <= 136'h0;
    end else begin
      _EVAL_301 <= _EVAL_172;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc3352a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f7e5e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb310e2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8842479)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f747e6e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dc63c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb611bfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c90b3f7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41d58e9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b9f3759)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55bc9d3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c70ab4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8efea4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed73bdec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42b363b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e61e560e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c50c85f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(610de59f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba472dbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc170e74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a92aec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d63973a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(849bb17e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb4624e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(978cbb4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ed0bdd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d120246)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9188d231)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8f1801c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daaee3d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cca05e7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbc13e6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97f4d334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed4350f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea96da71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69f1d6b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbfa0bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daf60fed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90fbebe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5785be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f337c358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f69ee573)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e803eda7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25c15ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4b900b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ec2f8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4669aab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7739ae8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd1e3962)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46be1adb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a575dca7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b566539)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d27fbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7408e68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a575a11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c79ec80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(242c57d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a9dc2ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c407f737)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77b7e18e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeea9afa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79e4456d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6d193ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2752e770)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15afe35b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33158d8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c249764)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(146bdd98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2deb6aed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c5df710)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d7c42ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab9abba5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
