//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_213(
  input         _EVAL,
  input         _EVAL_0,
  input  [3:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  input  [7:0]  _EVAL_7,
  output [1:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  output [31:0] _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [11:0] _EVAL_16,
  output [3:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output [1:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  input  [11:0] _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  output [7:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [8:0]  _EVAL_32,
  output        _EVAL_33,
  input  [31:0] _EVAL_34,
  output [2:0]  _EVAL_35,
  input  [31:0] _EVAL_36,
  output        _EVAL_37,
  output [31:0] _EVAL_38,
  input         _EVAL_39,
  output        _EVAL_40,
  input         _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  output [2:0]  _EVAL_44,
  input  [9:0]  _EVAL_45,
  output [31:0] _EVAL_46,
  output        _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49,
  input         _EVAL_50,
  input  [11:0] _EVAL_51
);
  wire  sb2tlOpt__EVAL;
  wire  sb2tlOpt__EVAL_0;
  wire [7:0] sb2tlOpt__EVAL_1;
  wire  sb2tlOpt__EVAL_2;
  wire  sb2tlOpt__EVAL_3;
  wire  sb2tlOpt__EVAL_4;
  wire [2:0] sb2tlOpt__EVAL_5;
  wire  sb2tlOpt__EVAL_6;
  wire  sb2tlOpt__EVAL_7;
  wire  sb2tlOpt__EVAL_8;
  wire  sb2tlOpt__EVAL_9;
  wire [31:0] sb2tlOpt__EVAL_10;
  wire  sb2tlOpt__EVAL_11;
  wire  sb2tlOpt__EVAL_12;
  wire [3:0] sb2tlOpt__EVAL_13;
  wire [2:0] sb2tlOpt__EVAL_14;
  wire  sb2tlOpt__EVAL_15;
  wire  sb2tlOpt__EVAL_16;
  wire  sb2tlOpt__EVAL_17;
  wire  sb2tlOpt__EVAL_18;
  wire [7:0] sb2tlOpt__EVAL_19;
  wire  sb2tlOpt__EVAL_20;
  wire [127:0] sb2tlOpt__EVAL_21;
  wire  sb2tlOpt__EVAL_22;
  wire [2:0] sb2tlOpt__EVAL_23;
  wire  sb2tlOpt__EVAL_24;
  wire  sb2tlOpt__EVAL_25;
  wire  sb2tlOpt__EVAL_26;
  wire [7:0] sb2tlOpt__EVAL_27;
  wire [127:0] sb2tlOpt__EVAL_28;
  reg  _EVAL_54;
  reg [31:0] _RAND_0;
  reg [7:0] _EVAL_56;
  reg [31:0] _RAND_1;
  reg [7:0] _EVAL_72;
  reg [31:0] _RAND_2;
  reg [7:0] _EVAL_75;
  reg [31:0] _RAND_3;
  reg [7:0] _EVAL_92;
  reg [31:0] _RAND_4;
  reg [7:0] _EVAL_130;
  reg [31:0] _RAND_5;
  reg [7:0] _EVAL_174;
  reg [31:0] _RAND_6;
  reg [7:0] _EVAL_182;
  reg [31:0] _RAND_7;
  reg  _EVAL_212;
  reg [31:0] _RAND_8;
  reg [7:0] _EVAL_229;
  reg [31:0] _RAND_9;
  reg [7:0] _EVAL_254;
  reg [31:0] _RAND_10;
  reg [7:0] _EVAL_277;
  reg [31:0] _RAND_11;
  reg  _EVAL_284;
  reg [31:0] _RAND_12;
  reg [7:0] _EVAL_329;
  reg [31:0] _RAND_13;
  reg [7:0] _EVAL_438;
  reg [31:0] _RAND_14;
  reg [7:0] _EVAL_446;
  reg [31:0] _RAND_15;
  reg [7:0] _EVAL_532;
  reg [31:0] _RAND_16;
  reg  _EVAL_593;
  reg [31:0] _RAND_17;
  reg [7:0] _EVAL_606;
  reg [31:0] _RAND_18;
  reg  _EVAL_616;
  reg [31:0] _RAND_19;
  reg [23:0] _EVAL_623;
  reg [31:0] _RAND_20;
  reg  _EVAL_634;
  reg [31:0] _RAND_21;
  reg [7:0] _EVAL_658;
  reg [31:0] _RAND_22;
  reg [7:0] _EVAL_732;
  reg [31:0] _RAND_23;
  reg  _EVAL_734;
  reg [31:0] _RAND_24;
  reg [7:0] _EVAL_737;
  reg [31:0] _RAND_25;
  reg [7:0] _EVAL_739;
  reg [31:0] _RAND_26;
  reg [7:0] _EVAL_751;
  reg [31:0] _RAND_27;
  reg [7:0] _EVAL_804;
  reg [31:0] _RAND_28;
  reg [1:0] _EVAL_838;
  reg [31:0] _RAND_29;
  reg [7:0] _EVAL_846;
  reg [31:0] _RAND_30;
  reg [7:0] _EVAL_858;
  reg [31:0] _RAND_31;
  reg  _EVAL_861;
  reg [31:0] _RAND_32;
  reg [7:0] _EVAL_864;
  reg [31:0] _RAND_33;
  reg [7:0] _EVAL_881;
  reg [31:0] _RAND_34;
  reg [7:0] _EVAL_915;
  reg [31:0] _RAND_35;
  reg [31:0] _EVAL_916;
  reg [31:0] _RAND_36;
  reg [7:0] _EVAL_961;
  reg [31:0] _RAND_37;
  reg [7:0] _EVAL_1001;
  reg [31:0] _RAND_38;
  reg [7:0] _EVAL_1019;
  reg [31:0] _RAND_39;
  reg [7:0] _EVAL_1040;
  reg [31:0] _RAND_40;
  reg [7:0] _EVAL_1055;
  reg [31:0] _RAND_41;
  reg  _EVAL_1065;
  reg [31:0] _RAND_42;
  reg [7:0] _EVAL_1100;
  reg [31:0] _RAND_43;
  reg [7:0] _EVAL_1132;
  reg [31:0] _RAND_44;
  reg [7:0] _EVAL_1134;
  reg [31:0] _RAND_45;
  reg [11:0] _EVAL_1135;
  reg [31:0] _RAND_46;
  reg [15:0] _EVAL_1137;
  reg [31:0] _RAND_47;
  reg [7:0] _EVAL_1154;
  reg [31:0] _RAND_48;
  reg [7:0] _EVAL_1200;
  reg [31:0] _RAND_49;
  reg [7:0] _EVAL_1207;
  reg [31:0] _RAND_50;
  reg [7:0] _EVAL_1250;
  reg [31:0] _RAND_51;
  reg [2:0] _EVAL_1263;
  reg [31:0] _RAND_52;
  reg [7:0] _EVAL_1264;
  reg [31:0] _RAND_53;
  reg [7:0] _EVAL_1349;
  reg [31:0] _RAND_54;
  reg [7:0] _EVAL_1350;
  reg [31:0] _RAND_55;
  reg [7:0] _EVAL_1370;
  reg [31:0] _RAND_56;
  reg [7:0] _EVAL_1383;
  reg [31:0] _RAND_57;
  reg [7:0] _EVAL_1402;
  reg [31:0] _RAND_58;
  reg [7:0] _EVAL_1447;
  reg [31:0] _RAND_59;
  reg [7:0] _EVAL_1469;
  reg [31:0] _RAND_60;
  reg [7:0] _EVAL_1499;
  reg [31:0] _RAND_61;
  reg [7:0] _EVAL_1508;
  reg [31:0] _RAND_62;
  reg [7:0] _EVAL_1516;
  reg [31:0] _RAND_63;
  reg [7:0] _EVAL_1562;
  reg [31:0] _RAND_64;
  reg [7:0] _EVAL_1572;
  reg [31:0] _RAND_65;
  reg [7:0] _EVAL_1595;
  reg [31:0] _RAND_66;
  reg [7:0] _EVAL_1599;
  reg [31:0] _RAND_67;
  reg [7:0] _EVAL_1646;
  reg [31:0] _RAND_68;
  reg [7:0] _EVAL_1649;
  reg [31:0] _RAND_69;
  reg [7:0] _EVAL_1652;
  reg [31:0] _RAND_70;
  reg [7:0] _EVAL_1694;
  reg [31:0] _RAND_71;
  reg [7:0] _EVAL_1716;
  reg [31:0] _RAND_72;
  reg [7:0] _EVAL_1768;
  reg [31:0] _RAND_73;
  reg [7:0] _EVAL_1785;
  reg [31:0] _RAND_74;
  reg  _EVAL_1803;
  reg [31:0] _RAND_75;
  reg  _EVAL_1829;
  reg [31:0] _RAND_76;
  reg [7:0] _EVAL_1859;
  reg [31:0] _RAND_77;
  reg [31:0] _EVAL_1866;
  reg [31:0] _RAND_78;
  reg [7:0] _EVAL_1869;
  reg [31:0] _RAND_79;
  reg [7:0] _EVAL_1916;
  reg [31:0] _RAND_80;
  reg [7:0] _EVAL_1943;
  reg [31:0] _RAND_81;
  reg  _EVAL_1951;
  reg [31:0] _RAND_82;
  reg [7:0] _EVAL_1991;
  reg [31:0] _RAND_83;
  reg [7:0] _EVAL_2000;
  reg [31:0] _RAND_84;
  reg [7:0] _EVAL_2026;
  reg [31:0] _RAND_85;
  reg  _EVAL_2054;
  reg [31:0] _RAND_86;
  reg [7:0] _EVAL_2057;
  reg [31:0] _RAND_87;
  reg [7:0] _EVAL_2058;
  reg [31:0] _RAND_88;
  reg [7:0] _EVAL_2082;
  reg [31:0] _RAND_89;
  reg [7:0] _EVAL_2097;
  reg [31:0] _RAND_90;
  reg  _EVAL_2117;
  reg [31:0] _RAND_91;
  reg [7:0] _EVAL_2154;
  reg [31:0] _RAND_92;
  reg [7:0] _EVAL_2165;
  reg [31:0] _RAND_93;
  reg [2:0] _EVAL_2167;
  reg [31:0] _RAND_94;
  reg [31:0] _EVAL_2220;
  reg [31:0] _RAND_95;
  wire  _EVAL_1129;
  wire  _EVAL_2174;
  wire [7:0] _EVAL_642;
  wire  _EVAL_1252;
  wire [7:0] _EVAL_1528;
  wire  _EVAL_416;
  wire [7:0] _EVAL_1543;
  wire  _EVAL_1139;
  wire [7:0] _EVAL_1743;
  wire [31:0] _EVAL_1582;
  wire  _EVAL_1048;
  wire  _EVAL_644;
  wire [9:0] _EVAL_145;
  wire  _EVAL_181;
  wire  _EVAL_219;
  wire  _EVAL_1000;
  wire  _EVAL_1908;
  wire  _EVAL_1774;
  wire  _EVAL_1405;
  wire  _EVAL_1054;
  wire  _EVAL_1573;
  wire  _EVAL_1853;
  wire [8:0] _EVAL_390;
  wire [511:0] _EVAL_631;
  wire [9:0] _EVAL_643;
  wire  _EVAL_502;
  wire  _EVAL_1760;
  wire  _EVAL_1604;
  wire [7:0] _EVAL_1076;
  wire  _EVAL_1928;
  wire [7:0] _EVAL_1567;
  wire  _EVAL_2187;
  wire [7:0] _EVAL_1668;
  wire  _EVAL_1292;
  wire [7:0] _EVAL_1707;
  wire [31:0] _EVAL_332;
  wire [7:0] _EVAL_1017;
  wire  _EVAL_1486;
  wire [31:0] _EVAL_1500;
  wire  _EVAL_1492;
  wire  _EVAL_681;
  wire  _EVAL_1503;
  wire  _EVAL_2076;
  wire [6:0] _EVAL_177;
  wire  _EVAL_583;
  wire  _EVAL_171;
  wire  _EVAL_540;
  wire  _EVAL_594;
  wire  _EVAL_1878;
  wire  _EVAL_1632;
  wire [5:0] _EVAL_433;
  wire [63:0] _EVAL_1421;
  wire  _EVAL_610;
  wire  _EVAL_376;
  wire [6:0] _EVAL_2056;
  wire  _EVAL_680;
  wire  _EVAL_581;
  wire [7:0] _EVAL_2136;
  wire  _EVAL_1964;
  wire  _EVAL_139;
  wire  _EVAL_1971;
  wire  _EVAL_1858;
  wire [7:0] _EVAL_142;
  wire  _EVAL_1992;
  wire  _EVAL_749;
  wire [7:0] _EVAL_573;
  wire  _EVAL_1387;
  wire  _EVAL_1691;
  wire  _EVAL_1961;
  wire  _EVAL_646;
  wire  _EVAL_1686;
  wire [7:0] _EVAL_366;
  wire  _EVAL_234;
  wire  _EVAL_1145;
  wire  _EVAL_1459;
  wire [7:0] _EVAL_55;
  wire  _EVAL_729;
  wire [3:0] _EVAL_1323;
  wire [2:0] _EVAL_1537;
  wire [23:0] _EVAL_106;
  wire [7:0] _EVAL_1563;
  wire  _EVAL_758;
  wire  _EVAL_886;
  wire  _EVAL_57;
  wire  _EVAL_1020;
  wire  _EVAL_1319;
  wire [7:0] _EVAL_1753;
  wire  _EVAL_1638;
  wire  _EVAL_857;
  wire [127:0] _EVAL_2029;
  wire  _EVAL_531;
  wire  _EVAL_1009;
  wire  _EVAL_714;
  wire  _EVAL_1093;
  wire  _EVAL_568;
  wire  _EVAL_1556;
  wire  _EVAL_451;
  wire  _EVAL_214;
  wire  _EVAL_1732;
  wire  _EVAL_305;
  wire  _EVAL_1303;
  wire  _EVAL_1376;
  wire  _EVAL_1580;
  wire  _EVAL_633;
  wire  _EVAL_2178;
  wire  _EVAL_1311;
  wire  _EVAL_603;
  wire  _EVAL_1782;
  wire  _EVAL_1501;
  wire  _EVAL_1078;
  wire  _EVAL_1780;
  wire  _EVAL_518;
  wire  _EVAL_109;
  wire  _EVAL_721;
  wire  _EVAL_1737;
  wire  _EVAL_987;
  wire  _EVAL_205;
  wire  _EVAL_1274;
  wire  _EVAL_1085;
  wire  _EVAL_153;
  wire  _EVAL_750;
  wire  _EVAL_1299;
  wire  _EVAL_1607;
  wire  _EVAL_224;
  wire  _EVAL_1209;
  wire  _EVAL_420;
  wire  _EVAL_900;
  wire  _EVAL_1615;
  wire  _EVAL_924;
  wire  _EVAL_350;
  wire  _EVAL_2148;
  wire  _EVAL_505;
  wire  _EVAL_374;
  wire  _EVAL_1590;
  wire  _EVAL_2031;
  wire  _EVAL_1424;
  wire  _EVAL_1312;
  wire  _EVAL_1830;
  wire  _EVAL_715;
  wire  _EVAL_1736;
  wire  _EVAL_752;
  wire  _EVAL_1331;
  wire  _EVAL_1745;
  wire  _EVAL_560;
  wire  _EVAL_753;
  wire  _EVAL_779;
  wire  _EVAL_1086;
  wire  _EVAL_127;
  wire  _EVAL_1709;
  wire  _EVAL_1119;
  wire  _EVAL_1966;
  wire  _EVAL_529;
  wire  _EVAL_165;
  wire  _EVAL_901;
  wire  _EVAL_1931;
  wire  _EVAL_1090;
  wire  _EVAL_2051;
  wire  _EVAL_189;
  wire  _EVAL_1449;
  wire  _EVAL_173;
  wire  _EVAL_827;
  wire  _EVAL_1841;
  wire  _EVAL_869;
  wire  _EVAL_2150;
  wire  _EVAL_462;
  wire  _EVAL_862;
  wire  _EVAL_2125;
  wire  _EVAL_67;
  wire  _EVAL_395;
  wire  _EVAL_2006;
  wire  _EVAL_1059;
  wire  _EVAL_612;
  wire  _EVAL_447;
  wire  _EVAL_950;
  wire  _EVAL_1050;
  wire  _EVAL_382;
  wire  _EVAL_1381;
  wire  _EVAL_159;
  wire  _EVAL_1464;
  wire  _EVAL_266;
  wire  _EVAL_2104;
  wire  _EVAL_1175;
  wire  _EVAL_1844;
  wire  _EVAL_453;
  wire  _EVAL_255;
  wire  _EVAL_268;
  wire  _EVAL_823;
  wire  _EVAL_1696;
  wire  _EVAL_2126;
  wire  _EVAL_1114;
  wire  _EVAL_883;
  wire  _EVAL_1628;
  wire  _EVAL_818;
  wire  _EVAL_140;
  wire  _EVAL_2215;
  wire  _EVAL_1494;
  wire  _EVAL_1470;
  wire  _EVAL_415;
  wire  _EVAL_381;
  wire  _EVAL_1483;
  wire  _EVAL_1335;
  wire  _EVAL_771;
  wire  _EVAL_193;
  wire  _EVAL_1245;
  wire  _EVAL_885;
  wire  _EVAL_1744;
  wire  _EVAL_516;
  wire  _EVAL_1270;
  wire  _EVAL_547;
  wire  _EVAL_1392;
  wire  _EVAL_1226;
  wire  _EVAL_621;
  wire  _EVAL_261;
  wire  _EVAL_1008;
  wire  _EVAL_148;
  wire  _EVAL_934;
  wire  _EVAL_1036;
  wire  _EVAL_1549;
  wire  _EVAL_2169;
  wire  _EVAL_114;
  wire  _EVAL_2111;
  wire  _EVAL_742;
  wire  _EVAL_364;
  wire  _EVAL_655;
  wire  _EVAL_772;
  wire  _EVAL_1979;
  wire  _EVAL_1968;
  wire  _EVAL_64;
  wire  _EVAL_2101;
  wire  _EVAL_2106;
  wire  _EVAL_370;
  wire  _EVAL_1986;
  wire [7:0] _EVAL_1888;
  wire  _EVAL_1246;
  wire  _EVAL_614;
  wire  _EVAL_129;
  wire  _EVAL_507;
  wire  _EVAL_168;
  wire  _EVAL_1824;
  wire  _EVAL_1286;
  wire  _EVAL_410;
  wire  _EVAL_299;
  wire  _EVAL_538;
  wire  _EVAL_2235;
  wire  _EVAL_2137;
  wire  _EVAL_1545;
  wire  _EVAL_339;
  wire [31:0] _EVAL_545;
  wire [31:0] _EVAL_1799;
  wire [31:0] _EVAL_1141;
  wire [31:0] _EVAL_1658;
  wire [31:0] _EVAL_1635;
  wire [31:0] _EVAL_1302;
  wire [31:0] _EVAL_905;
  wire [31:0] _EVAL_478;
  wire [31:0] _EVAL_2234;
  wire [31:0] _EVAL_2182;
  wire [31:0] _EVAL_222;
  wire [31:0] _EVAL_460;
  wire [31:0] _EVAL_1810;
  wire [31:0] _EVAL_490;
  wire [31:0] _EVAL_1704;
  wire [31:0] _EVAL_2181;
  wire [31:0] _EVAL_794;
  wire [31:0] _EVAL_1398;
  wire [31:0] _EVAL_1356;
  wire [31:0] _EVAL_741;
  wire [31:0] _EVAL_495;
  wire [31:0] _EVAL_1253;
  wire [31:0] _EVAL_228;
  wire [31:0] _EVAL_443;
  wire [31:0] _EVAL_248;
  wire [31:0] _EVAL_1360;
  wire [31:0] _EVAL_757;
  wire [31:0] _EVAL_1131;
  wire [31:0] _EVAL_795;
  wire [31:0] _EVAL_1860;
  wire [31:0] _EVAL_1359;
  wire [31:0] _EVAL_1577;
  wire [31:0] _EVAL_1345;
  wire [31:0] _EVAL_110;
  wire [31:0] _EVAL_1451;
  wire [31:0] _EVAL_904;
  wire [31:0] _EVAL_353;
  wire [31:0] _EVAL_196;
  wire [31:0] _EVAL_716;
  wire [31:0] _EVAL_1419;
  wire  _EVAL_637;
  wire  _EVAL_1900;
  wire  _EVAL_627;
  wire  _EVAL_1366;
  wire  _EVAL_1608;
  wire  _EVAL_880;
  wire  _EVAL_1096;
  wire  _EVAL_295;
  wire  _EVAL_994;
  wire [7:0] _EVAL_2060;
  wire  _EVAL_423;
  wire  _EVAL_328;
  wire  _EVAL_2095;
  wire  _EVAL_2017;
  wire  _EVAL_1798;
  wire  _EVAL_986;
  wire  _EVAL_1845;
  wire [9:0] _EVAL_190;
  wire  _EVAL_1188;
  wire  _EVAL_2080;
  wire  _EVAL_272;
  wire  _EVAL_665;
  wire  _EVAL_1831;
  wire  _EVAL_539;
  wire  _EVAL_731;
  wire  _EVAL_1104;
  wire  _EVAL_1304;
  wire [7:0] _EVAL_1827;
  wire  _EVAL_619;
  wire  _EVAL_556;
  wire  _EVAL_820;
  wire  _EVAL_1880;
  wire  _EVAL_107;
  wire  _EVAL_1558;
  wire  _EVAL_647;
  wire  _EVAL_1654;
  wire  _EVAL_544;
  wire  _EVAL_1680;
  wire  _EVAL_2030;
  wire  _EVAL_1720;
  wire  _EVAL_2102;
  wire  _EVAL_1570;
  wire  _EVAL_971;
  wire  _EVAL_1742;
  wire  _EVAL_233;
  wire  _EVAL_2190;
  wire  _EVAL_418;
  wire  _EVAL_1400;
  wire  _EVAL_1721;
  wire  _EVAL_1532;
  wire  _EVAL_1053;
  wire  _EVAL_1229;
  wire  _EVAL_2088;
  wire  _EVAL_2092;
  wire  _EVAL_113;
  wire  _EVAL_1551;
  wire  _EVAL_166;
  wire  _EVAL_1975;
  wire  _EVAL_727;
  wire  _EVAL_1163;
  wire  _EVAL_1317;
  wire  _EVAL_569;
  wire  _EVAL_2205;
  wire  _EVAL_1192;
  wire  _EVAL_360;
  wire  _EVAL_1038;
  wire  _EVAL_1296;
  wire  _EVAL_333;
  wire  _EVAL_719;
  wire  _EVAL_1133;
  wire  _EVAL_914;
  wire  _EVAL_736;
  wire  _EVAL_958;
  wire  _EVAL_1524;
  wire  _EVAL_204;
  wire  _EVAL_1171;
  wire  _EVAL_1490;
  wire  _EVAL_1756;
  wire  _EVAL_1698;
  wire  _EVAL_884;
  wire  _EVAL_408;
  wire  _EVAL_1083;
  wire  _EVAL_1636;
  wire  _EVAL_1136;
  wire  _EVAL_236;
  wire  _EVAL_133;
  wire  _EVAL_483;
  wire  _EVAL_1947;
  wire  _EVAL_2153;
  wire  _EVAL_620;
  wire  _EVAL_1318;
  wire  _EVAL_1201;
  wire  _EVAL_559;
  wire  _EVAL_1708;
  wire  _EVAL_1914;
  wire  _EVAL_1593;
  wire  _EVAL_1752;
  wire  _EVAL_2195;
  wire  _EVAL_1004;
  wire  _EVAL_440;
  wire  _EVAL_669;
  wire  _EVAL_1237;
  wire  _EVAL_879;
  wire  _EVAL_303;
  wire  _EVAL_1242;
  wire  _EVAL_1903;
  wire  _EVAL_330;
  wire  _EVAL_686;
  wire  _EVAL_104;
  wire  _EVAL_334;
  wire  _EVAL_191;
  wire  _EVAL_101;
  wire  _EVAL_384;
  wire  _EVAL_221;
  wire  _EVAL_1003;
  wire  _EVAL_660;
  wire  _EVAL_264;
  wire  _EVAL_957;
  wire  _EVAL_2068;
  wire  _EVAL_519;
  wire  _EVAL_639;
  wire  _EVAL_469;
  wire  _EVAL_361;
  wire  _EVAL_760;
  wire  _EVAL_403;
  wire  _EVAL_164;
  wire  _EVAL_1322;
  wire [31:0] _EVAL_1965;
  wire [7:0] _EVAL_1925;
  wire  _EVAL_898;
  wire  _EVAL_2147;
  wire  _EVAL_61;
  wire  _EVAL_1254;
  wire  _EVAL_1838;
  wire  _EVAL_1473;
  wire  _EVAL_2236;
  wire  _EVAL_1885;
  wire  _EVAL_1244;
  wire  _EVAL_1854;
  wire  _EVAL_1193;
  wire  _EVAL_1094;
  wire  _EVAL_1771;
  wire  _EVAL_548;
  wire  _EVAL_1512;
  wire  _EVAL_918;
  wire  _EVAL_237;
  wire  _EVAL_1051;
  wire  _EVAL_195;
  wire  _EVAL_455;
  wire  _EVAL_2210;
  wire  _EVAL_1630;
  wire  _EVAL_508;
  wire  _EVAL_1491;
  wire  _EVAL_803;
  wire  _EVAL_2161;
  wire  _EVAL_789;
  wire  _EVAL_1592;
  wire  _EVAL_2233;
  wire  _EVAL_1057;
  wire  _EVAL_435;
  wire  _EVAL_2116;
  wire  _EVAL_244;
  wire  _EVAL_1791;
  wire  _EVAL_2086;
  wire  _EVAL_1993;
  wire  _EVAL_439;
  wire  _EVAL_1458;
  wire  _EVAL_2192;
  wire  _EVAL_570;
  wire  _EVAL_461;
  wire  _EVAL_590;
  wire  _EVAL_1662;
  wire  _EVAL_1548;
  wire  _EVAL_836;
  wire  _EVAL_553;
  wire  _EVAL_692;
  wire  _EVAL_988;
  wire  _EVAL_1308;
  wire  _EVAL_1535;
  wire  _EVAL_702;
  wire  _EVAL_970;
  wire  _EVAL_1103;
  wire  _EVAL_200;
  wire  _EVAL_1982;
  wire  _EVAL_436;
  wire  _EVAL_1305;
  wire  _EVAL_1750;
  wire  _EVAL_1079;
  wire  _EVAL_1932;
  wire  _EVAL_1071;
  wire  _EVAL_442;
  wire  _EVAL_1962;
  wire  _EVAL_401;
  wire  _EVAL_1879;
  wire  _EVAL_1062;
  wire  _EVAL_136;
  wire  _EVAL_1872;
  wire  _EVAL_1773;
  wire  _EVAL_1239;
  wire  _EVAL_94;
  wire  _EVAL_1998;
  wire  _EVAL_1769;
  wire  _EVAL_96;
  wire  _EVAL_1157;
  wire  _EVAL_1893;
  wire  _EVAL_1044;
  wire  _EVAL_2093;
  wire  _EVAL_865;
  wire  _EVAL_517;
  wire  _EVAL_693;
  wire  _EVAL_2127;
  wire  _EVAL_833;
  wire  _EVAL_1772;
  wire  _EVAL_2094;
  wire  _EVAL_270;
  wire  _EVAL_1765;
  wire  _EVAL_320;
  wire  _EVAL_839;
  wire  _EVAL_1610;
  wire  _EVAL_1677;
  wire  _EVAL_1836;
  wire  _EVAL_1277;
  wire  _EVAL_2044;
  wire  _EVAL_1637;
  wire  _EVAL_756;
  wire  _EVAL_790;
  wire  _EVAL_530;
  wire  _EVAL_1598;
  wire  _EVAL_380;
  wire  _EVAL_144;
  wire  _EVAL_1820;
  wire  _EVAL_695;
  wire  _EVAL_1243;
  wire  _EVAL_1840;
  wire  _EVAL_1722;
  wire  _EVAL_504;
  wire  _EVAL_372;
  wire  _EVAL_247;
  wire  _EVAL_319;
  wire  _EVAL_2087;
  wire  _EVAL_743;
  wire  _EVAL_1480;
  wire  _EVAL_85;
  wire  _EVAL_1138;
  wire  _EVAL_2069;
  wire  _EVAL_53;
  wire  _EVAL_728;
  wire  _EVAL_2012;
  wire  _EVAL_1276;
  wire  _EVAL_1225;
  wire  _EVAL_740;
  wire  _EVAL_1374;
  wire  _EVAL_2202;
  wire  _EVAL_1927;
  wire  _EVAL_1889;
  wire  _EVAL_1334;
  wire  _EVAL_2225;
  wire  _EVAL_141;
  wire  _EVAL_437;
  wire  _EVAL_936;
  wire  _EVAL_1396;
  wire  _EVAL_1174;
  wire  _EVAL_1960;
  wire  _EVAL_407;
  wire  _EVAL_859;
  wire  _EVAL_773;
  wire  _EVAL_1361;
  wire  _EVAL_175;
  wire  _EVAL_1222;
  wire  _EVAL_2185;
  wire  _EVAL_1847;
  wire  _EVAL_1391;
  wire  _EVAL_953;
  wire  _EVAL_2146;
  wire [31:0] _EVAL_726;
  wire  _EVAL_1327;
  wire  _EVAL_471;
  wire  _EVAL_2004;
  wire  _EVAL_137;
  wire  _EVAL_1538;
  wire  _EVAL_1815;
  wire  _EVAL_801;
  wire  _EVAL_558;
  wire  _EVAL_985;
  wire  _EVAL_1959;
  wire  _EVAL_256;
  wire  _EVAL_1169;
  wire  _EVAL_1301;
  wire  _EVAL_2110;
  wire  _EVAL_774;
  wire [2:0] _EVAL_2081;
  wire [15:0] _EVAL_1644;
  wire [15:0] _EVAL_2238;
  wire [4:0] _EVAL_345;
  wire [31:0] _EVAL_882;
  wire [31:0] _EVAL_1800;
  wire  _EVAL_172;
  wire  _EVAL_2011;
  wire [31:0] _EVAL_445;
  wire [3:0] _EVAL_1121;
  wire  _EVAL_1702;
  wire  _EVAL_778;
  wire  _EVAL_126;
  wire  _EVAL_1843;
  wire  _EVAL_989;
  wire  _EVAL_1484;
  wire  _EVAL_979;
  wire  _EVAL_349;
  wire  _EVAL_1153;
  wire  _EVAL_767;
  wire  _EVAL_452;
  wire  _EVAL_1988;
  wire  _EVAL_465;
  wire [7:0] _EVAL_1352;
  wire  _EVAL_1429;
  wire  _EVAL_1251;
  wire  _EVAL_1198;
  wire  _EVAL_1703;
  wire [7:0] _EVAL_1755;
  wire  _EVAL_2224;
  wire  _EVAL_311;
  wire  _EVAL_766;
  wire  _EVAL_1160;
  wire  _EVAL_73;
  wire  _EVAL_321;
  wire  _EVAL_105;
  wire  _EVAL_273;
  wire  _EVAL_847;
  wire  _EVAL_199;
  wire  _EVAL_485;
  wire  _EVAL_962;
  wire  _EVAL_1266;
  wire  _EVAL_630;
  wire  _EVAL_920;
  wire  _EVAL_1554;
  wire  _EVAL_336;
  wire  _EVAL_2197;
  wire  _EVAL_1766;
  wire  _EVAL_1404;
  wire  _EVAL_1997;
  wire  _EVAL_894;
  wire  _EVAL_1813;
  wire  _EVAL_656;
  wire  _EVAL_351;
  wire  _EVAL_1987;
  wire  _EVAL_1534;
  wire  _EVAL_554;
  wire  _EVAL_59;
  wire  _EVAL_1435;
  wire  _EVAL_1147;
  wire  _EVAL_2079;
  wire  _EVAL_323;
  wire  _EVAL_770;
  wire  _EVAL_2114;
  wire  _EVAL_1890;
  wire [9:0] _EVAL_975;
  wire  _EVAL_589;
  wire  _EVAL_527;
  wire  _EVAL_855;
  wire  _EVAL_1973;
  wire  _EVAL_1958;
  wire [7:0] _EVAL_562;
  wire  _EVAL_1711;
  wire  _EVAL_385;
  wire  _EVAL_835;
  wire  _EVAL_598;
  wire  _EVAL_260;
  wire  _EVAL_1985;
  wire  _EVAL_278;
  wire  _EVAL_487;
  wire  _EVAL_685;
  wire  _EVAL_1594;
  wire  _EVAL_1641;
  wire  _EVAL_1671;
  wire  _EVAL_60;
  wire  _EVAL_1241;
  wire  _EVAL_688;
  wire  _EVAL_1452;
  wire  _EVAL_1542;
  wire  _EVAL_322;
  wire  _EVAL_2075;
  wire  _EVAL_1485;
  wire  _EVAL_1441;
  wire [127:0] _EVAL_1422;
  wire [7:0] _EVAL_1616;
  wire [127:0] _EVAL_817;
  wire  _EVAL_1047;
  wire  _EVAL_357;
  wire  _EVAL_291;
  wire  _EVAL_783;
  wire  _EVAL_1493;
  wire  _EVAL_2067;
  wire  _EVAL_1627;
  wire  _EVAL_240;
  wire  _EVAL_840;
  wire  _EVAL_1210;
  wire  _EVAL_1969;
  wire  _EVAL_281;
  wire  _EVAL_1864;
  wire  _EVAL_480;
  wire  _EVAL_422;
  wire  _EVAL_1462;
  wire  _EVAL_1386;
  wire  _EVAL_63;
  wire  _EVAL_1415;
  wire  _EVAL_1609;
  wire  _EVAL_162;
  wire [2:0] _EVAL_1511;
  wire  _EVAL_841;
  wire  _EVAL_155;
  wire [2:0] _EVAL_1436;
  wire  _EVAL_1082;
  wire  _EVAL_2157;
  wire  _EVAL_285;
  wire  _EVAL_923;
  wire  _EVAL_1589;
  wire  _EVAL_796;
  wire [7:0] _EVAL_1205;
  wire  _EVAL_513;
  wire  _EVAL_1984;
  wire  _EVAL_135;
  wire  _EVAL_1357;
  wire  _EVAL_1414;
  wire  _EVAL_475;
  wire  _EVAL_648;
  wire  _EVAL_88;
  wire  _EVAL_555;
  wire  _EVAL_895;
  wire  _EVAL_2222;
  wire  _EVAL_1098;
  wire  _EVAL_1920;
  wire  _EVAL_1184;
  wire  _EVAL_1942;
  wire  _EVAL_1606;
  wire  _EVAL_371;
  wire  _EVAL_1430;
  wire  _EVAL_95;
  wire  _EVAL_722;
  wire [31:0] _EVAL_124;
  wire  _EVAL_1066;
  wire  _EVAL_1833;
  wire  _EVAL_1806;
  wire  _EVAL_628;
  wire  _EVAL_528;
  wire  _EVAL_131;
  wire  _EVAL_697;
  wire  _EVAL_1316;
  wire  _EVAL_2109;
  wire  _EVAL_1996;
  wire  _EVAL_169;
  wire  _EVAL_217;
  wire  _EVAL_1540;
  wire [15:0] _EVAL_744;
  wire  _EVAL_1465;
  wire  _EVAL_1977;
  wire  _EVAL_701;
  wire  _EVAL_1818;
  wire  _EVAL_1101;
  wire  _EVAL_324;
  wire  _EVAL_943;
  wire [31:0] _EVAL_1466;
  wire [31:0] _EVAL_352;
  wire [31:0] _EVAL_1074;
  wire [31:0] _EVAL_492;
  wire [31:0] _EVAL_1362;
  wire [31:0] _EVAL_1240;
  wire [31:0] _EVAL_152;
  wire [31:0] _EVAL_123;
  wire [31:0] _EVAL_1221;
  wire [31:0] _EVAL_1874;
  wire [31:0] _EVAL_2073;
  wire [31:0] _EVAL_409;
  wire [31:0] _EVAL_1740;
  wire [31:0] _EVAL_2219;
  wire [31:0] _EVAL_1695;
  wire  _EVAL_811;
  wire  _EVAL_2204;
  wire [16:0] _EVAL_1125;
  wire [20:0] _EVAL_899;
  wire  _EVAL_2113;
  wire  _EVAL_1428;
  wire  _EVAL_1822;
  wire  _EVAL_1902;
  wire  _EVAL_1789;
  wire  _EVAL_1227;
  wire  _EVAL_1216;
  wire  _EVAL_2194;
  wire  _EVAL_2036;
  wire  _EVAL_1794;
  wire  _EVAL_444;
  wire  _EVAL_1282;
  wire  _EVAL_1413;
  wire  _EVAL_1238;
  wire  _EVAL_1306;
  wire  _EVAL_1790;
  wire  _EVAL_458;
  wire  _EVAL_122;
  wire [31:0] _EVAL_657;
  wire [31:0] _EVAL_1173;
  wire [31:0] _EVAL_2133;
  wire [31:0] _EVAL_501;
  wire  _EVAL_710;
  wire  _EVAL_251;
  wire  _EVAL_822;
  wire  _EVAL_1807;
  wire  _EVAL_611;
  wire  _EVAL_208;
  wire  _EVAL_808;
  wire  _EVAL_1107;
  wire  _EVAL_2152;
  wire  _EVAL_777;
  wire  _EVAL_782;
  wire  _EVAL_1021;
  wire  _EVAL_2230;
  wire  _EVAL_860;
  wire  _EVAL_62;
  wire  _EVAL_1579;
  wire  _EVAL_2015;
  wire  _EVAL_666;
  wire  _EVAL_347;
  wire  _EVAL_1690;
  wire  _EVAL_1022;
  wire  _EVAL_1427;
  wire  _EVAL_709;
  wire  _EVAL_1995;
  wire  _EVAL_1337;
  wire  _EVAL_1310;
  wire  _EVAL_1793;
  wire  _EVAL_1081;
  wire  _EVAL_2218;
  wire  _EVAL_2020;
  wire  _EVAL_1394;
  wire  _EVAL_1069;
  wire  _EVAL_1401;
  wire  _EVAL_577;
  wire  _EVAL_1518;
  wire  _EVAL_856;
  wire  _EVAL_306;
  wire  _EVAL_622;
  wire  _EVAL_1926;
  wire  _EVAL_467;
  wire  _EVAL_1230;
  wire  _EVAL_1314;
  wire  _EVAL_375;
  wire  _EVAL_1821;
  wire  _EVAL_1111;
  wire  _EVAL_1180;
  wire  _EVAL_117;
  wire  _EVAL_1089;
  wire  _EVAL_2108;
  wire  _EVAL_1271;
  wire  _EVAL_1648;
  wire  _EVAL_2201;
  wire  _EVAL_1187;
  wire  _EVAL_1176;
  wire  _EVAL_312;
  wire  _EVAL_872;
  wire  _EVAL_434;
  wire  _EVAL_1935;
  wire  _EVAL_1850;
  wire  _EVAL_2191;
  wire  _EVAL_143;
  wire  _EVAL_1034;
  wire  _EVAL_1906;
  wire  _EVAL_866;
  wire  _EVAL_1583;
  wire  _EVAL_1273;
  wire  _EVAL_776;
  wire  _EVAL_1565;
  wire  _EVAL_1049;
  wire  _EVAL_1425;
  wire  _EVAL_557;
  wire  _EVAL_781;
  wire  _EVAL_1197;
  wire  _EVAL_2021;
  wire  _EVAL_274;
  wire  _EVAL_1105;
  wire  _EVAL_503;
  wire  _EVAL_1479;
  wire  _EVAL_826;
  wire  _EVAL_2160;
  wire  _EVAL_69;
  wire  _EVAL_1923;
  wire  _EVAL_1569;
  wire  _EVAL_1095;
  wire  _EVAL_1112;
  wire  _EVAL_2130;
  wire  _EVAL_1326;
  wire  _EVAL_207;
  wire  _EVAL_1329;
  wire  _EVAL_356;
  wire  _EVAL_1602;
  wire  _EVAL_383;
  wire  _EVAL_1898;
  wire  _EVAL_2200;
  wire  _EVAL_2041;
  wire  _EVAL_2071;
  wire  _EVAL_1976;
  wire  _EVAL_1832;
  wire  _EVAL_1432;
  wire  _EVAL_472;
  wire  _EVAL_1851;
  wire  _EVAL_887;
  wire [7:0] _EVAL_868;
  wire  _EVAL_1234;
  wire [2:0] _EVAL_1297;
  wire  _EVAL_68;
  wire  _EVAL_785;
  wire [28:0] _EVAL_1495;
  wire [31:0] _EVAL_1710;
  wire [31:0] _EVAL_1320;
  wire [31:0] _EVAL_98;
  wire [31:0] _EVAL_1295;
  wire [31:0] _EVAL_896;
  wire [31:0] _EVAL_809;
  wire [31:0] _EVAL_1461;
  wire [31:0] _EVAL_763;
  wire [31:0] _EVAL_1052;
  wire [31:0] _EVAL_968;
  wire [31:0] _EVAL_300;
  wire [31:0] _EVAL_2177;
  wire [31:0] _EVAL_1980;
  wire [31:0] _EVAL_600;
  wire [31:0] _EVAL_1664;
  wire [2:0] _EVAL_1892;
  wire  _EVAL_1571;
  wire  _EVAL_1517;
  wire  _EVAL_2019;
  wire [11:0] _EVAL_1509;
  wire  _EVAL_1371;
  wire  _EVAL_567;
  wire  _EVAL_115;
  wire  _EVAL_245;
  wire [2:0] _EVAL_1377;
  wire  _EVAL_290;
  wire  _EVAL_118;
  wire  _EVAL_498;
  wire  _EVAL_388;
  wire  _EVAL_1037;
  wire  _EVAL_929;
  wire  _EVAL_2214;
  wire  _EVAL_1219;
  wire  _EVAL_1092;
  wire [31:0] _EVAL_1379;
  wire  _EVAL_1113;
  wire  _EVAL_1189;
  wire [1:0] _EVAL_1487;
  wire  _EVAL_1970;
  wire  _EVAL_1603;
  wire  _EVAL_377;
  wire [2:0] _EVAL_738;
  wire  _EVAL_470;
  wire  _EVAL_157;
  wire  _EVAL_906;
  wire  _EVAL_1454;
  wire  _EVAL_179;
  wire  _EVAL_1406;
  wire [2:0] _EVAL_431;
  wire  _EVAL_1247;
  wire  _EVAL_511;
  wire  _EVAL_1596;
  wire  _EVAL_1010;
  wire  _EVAL_1856;
  wire  _EVAL_194;
  wire  _EVAL_315;
  wire  _EVAL_1717;
  wire  _EVAL_1805;
  wire  _EVAL_1936;
  wire  _EVAL_1045;
  wire [21:0] _EVAL_959;
  wire [22:0] _EVAL_1862;
  wire  _EVAL_1185;
  wire  _EVAL_1639;
  wire  _EVAL_1029;
  wire  _EVAL_2038;
  wire  _EVAL_699;
  wire [31:0] _EVAL_662;
  wire  _EVAL_810;
  wire  _EVAL_65;
  wire  _EVAL_2025;
  wire  _EVAL_663;
  wire  _EVAL_1618;
  wire [127:0] _EVAL_1861;
  wire [31:0] _EVAL_928;
  wire  _EVAL_307;
  wire  _EVAL_1777;
  wire  _EVAL_209;
  wire  _EVAL_2014;
  wire  _EVAL_1678;
  wire  _EVAL_877;
  wire  _EVAL_1622;
  wire  _EVAL_596;
  wire  _EVAL_1870;
  wire  _EVAL_2032;
  wire  _EVAL_1725;
  wire  _EVAL_108;
  wire  _EVAL_450;
  wire  _EVAL_1612;
  wire  _EVAL_1990;
  wire  _EVAL_533;
  wire  _EVAL_981;
  wire  _EVAL_1520;
  wire  _EVAL_399;
  wire  _EVAL_907;
  wire  _EVAL_1474;
  wire  _EVAL_1808;
  wire  _EVAL_1324;
  wire  _EVAL_363;
  wire  _EVAL_1685;
  wire  _EVAL_1631;
  wire  _EVAL_613;
  wire  _EVAL_635;
  wire [31:0] _EVAL_1478;
  wire  _EVAL_935;
  wire  _EVAL_1560;
  wire  _EVAL_786;
  wire  _EVAL_386;
  wire  _EVAL_1642;
  wire  _EVAL_1194;
  wire  _EVAL_1541;
  wire  _EVAL_1749;
  wire  _EVAL_670;
  wire  _EVAL_500;
  wire  _EVAL_706;
  wire  _EVAL_1747;
  wire  _EVAL_1633;
  wire  _EVAL_1191;
  wire  _EVAL_232;
  wire  _EVAL_1199;
  wire  _EVAL_1344;
  wire  _EVAL_298;
  wire [11:0] _EVAL_225;
  wire  _EVAL_1269;
  wire  _EVAL_1460;
  wire  _EVAL_1877;
  wire  _EVAL_1940;
  wire  _EVAL_712;
  wire  _EVAL_464;
  wire  _EVAL_2212;
  wire  _EVAL_1307;
  wire [1:0] _EVAL_1056;
  wire [15:0] _EVAL_79;
  wire [31:0] _EVAL_625;
  wire [31:0] _EVAL_1776;
  wire [31:0] _EVAL_459;
  wire [31:0] _EVAL_1911;
  wire [31:0] _EVAL_1795;
  wire [31:0] _EVAL_66;
  wire [31:0] _EVAL_393;
  wire [15:0] _EVAL_482;
  wire  _EVAL_718;
  wire  _EVAL_848;
  wire  _EVAL_845;
  wire  _EVAL_521;
  wire  _EVAL_151;
  wire  _EVAL_941;
  wire  _EVAL_454;
  wire  _EVAL_1547;
  wire  _EVAL_1873;
  wire  _EVAL_1471;
  wire  _EVAL_404;
  wire  _EVAL_515;
  wire  _EVAL_2199;
  wire  _EVAL_77;
  wire  _EVAL_192;
  wire  _EVAL_1918;
  wire  _EVAL_1564;
  wire  _EVAL_1536;
  wire  _EVAL_523;
  wire  _EVAL_210;
  wire  _EVAL_2096;
  wire  _EVAL_933;
  wire  _EVAL_1917;
  wire [2:0] _EVAL_1754;
  wire [2:0] _EVAL_1482;
  wire  _EVAL_925;
  wire  _EVAL_1656;
  wire [13:0] _EVAL_1731;
  wire [23:0] _EVAL_1006;
  wire  _EVAL_2229;
  wire  _EVAL_80;
  wire  _EVAL_588;
  wire  _EVAL_969;
  wire  _EVAL_1294;
  wire  _EVAL_1012;
  wire  _EVAL_908;
  wire  _EVAL_522;
  wire  _EVAL_359;
  wire  _EVAL_1108;
  wire  _EVAL_463;
  wire  _EVAL_1952;
  wire  _EVAL_955;
  wire  _EVAL_2134;
  wire  _EVAL_1697;
  wire  _EVAL_875;
  wire  _EVAL_2226;
  wire  _EVAL_2001;
  wire  _EVAL_1751;
  wire  _EVAL_2216;
  wire  _EVAL_591;
  wire  _EVAL_1275;
  wire  _EVAL_391;
  wire  _EVAL_2170;
  wire  _EVAL_313;
  wire  _EVAL_805;
  wire  _EVAL_1218;
  wire  _EVAL_253;
  wire  _EVAL_82;
  wire  _EVAL_843;
  wire  _EVAL_1339;
  wire  _EVAL_1456;
  wire  _EVAL_1688;
  wire  _EVAL_1403;
  wire  _EVAL_990;
  wire  _EVAL_1313;
  wire [31:0] _EVAL_373;
  wire [28:0] _EVAL_1533;
  wire [31:0] _EVAL_1881;
  wire [31:0] _EVAL_636;
  wire [31:0] _EVAL_100;
  wire [13:0] _EVAL_156;
  wire  _EVAL_1115;
  wire  _EVAL_1158;
  wire  _EVAL_279;
  wire [23:0] _EVAL_331;
  wire  _EVAL_2048;
  wire [127:0] _EVAL_457;
  wire [31:0] _EVAL_632;
  wire  _EVAL_1826;
  wire  _EVAL_1912;
  wire  _EVAL_703;
  wire  _EVAL_1353;
  wire  _EVAL_103;
  wire  _EVAL_1060;
  wire  _EVAL_814;
  wire  _EVAL_784;
  wire  _EVAL_671;
  wire  _EVAL_52;
  wire  _EVAL_1523;
  wire  _EVAL_1183;
  wire  _EVAL_1787;
  wire  _EVAL_149;
  wire  _EVAL_543;
  wire  _EVAL_2034;
  wire  _EVAL_2047;
  wire  _EVAL_211;
  wire  _EVAL_185;
  wire  _EVAL_2138;
  wire  _EVAL_1797;
  wire  _EVAL_2144;
  wire  _EVAL_2166;
  wire  _EVAL_1433;
  wire  _EVAL_1762;
  wire [127:0] _EVAL_1653;
  wire  _EVAL_1279;
  wire [31:0] _EVAL_1665;
  wire [31:0] _EVAL_705;
  wire  _EVAL_112;
  wire  _EVAL_1522;
  wire  _EVAL_1215;
  wire  _EVAL_362;
  wire  _EVAL_724;
  wire [15:0] _EVAL_1863;
  wire  _EVAL_912;
  wire [2:0] _EVAL_867;
  wire  _EVAL_761;
  wire  _EVAL_1938;
  wire  _EVAL_2228;
  wire  _EVAL_678;
  wire  _EVAL_690;
  wire  _EVAL_74;
  wire [31:0] _EVAL_318;
  wire  _EVAL_1196;
  wire  _EVAL_1643;
  wire  _EVAL_1232;
  wire  _EVAL_2139;
  wire  _EVAL_694;
  wire  _EVAL_1939;
  wire  _EVAL_449;
  wire [31:0] _EVAL_1439;
  SiFive__EVAL_210 sb2tlOpt (
    ._EVAL(sb2tlOpt__EVAL),
    ._EVAL_0(sb2tlOpt__EVAL_0),
    ._EVAL_1(sb2tlOpt__EVAL_1),
    ._EVAL_2(sb2tlOpt__EVAL_2),
    ._EVAL_3(sb2tlOpt__EVAL_3),
    ._EVAL_4(sb2tlOpt__EVAL_4),
    ._EVAL_5(sb2tlOpt__EVAL_5),
    ._EVAL_6(sb2tlOpt__EVAL_6),
    ._EVAL_7(sb2tlOpt__EVAL_7),
    ._EVAL_8(sb2tlOpt__EVAL_8),
    ._EVAL_9(sb2tlOpt__EVAL_9),
    ._EVAL_10(sb2tlOpt__EVAL_10),
    ._EVAL_11(sb2tlOpt__EVAL_11),
    ._EVAL_12(sb2tlOpt__EVAL_12),
    ._EVAL_13(sb2tlOpt__EVAL_13),
    ._EVAL_14(sb2tlOpt__EVAL_14),
    ._EVAL_15(sb2tlOpt__EVAL_15),
    ._EVAL_16(sb2tlOpt__EVAL_16),
    ._EVAL_17(sb2tlOpt__EVAL_17),
    ._EVAL_18(sb2tlOpt__EVAL_18),
    ._EVAL_19(sb2tlOpt__EVAL_19),
    ._EVAL_20(sb2tlOpt__EVAL_20),
    ._EVAL_21(sb2tlOpt__EVAL_21),
    ._EVAL_22(sb2tlOpt__EVAL_22),
    ._EVAL_23(sb2tlOpt__EVAL_23),
    ._EVAL_24(sb2tlOpt__EVAL_24),
    ._EVAL_25(sb2tlOpt__EVAL_25),
    ._EVAL_26(sb2tlOpt__EVAL_26),
    ._EVAL_27(sb2tlOpt__EVAL_27),
    ._EVAL_28(sb2tlOpt__EVAL_28)
  );
  assign _EVAL_1129 = _EVAL_1137[3];
  assign _EVAL_2174 = _EVAL_1[3];
  assign _EVAL_642 = _EVAL_2174 ? 8'hff : 8'h0;
  assign _EVAL_1252 = _EVAL_1[2];
  assign _EVAL_1528 = _EVAL_1252 ? 8'hff : 8'h0;
  assign _EVAL_416 = _EVAL_1[1];
  assign _EVAL_1543 = _EVAL_416 ? 8'hff : 8'h0;
  assign _EVAL_1139 = _EVAL_1[0];
  assign _EVAL_1743 = _EVAL_1139 ? 8'hff : 8'h0;
  assign _EVAL_1582 = {_EVAL_642,_EVAL_1528,_EVAL_1543,_EVAL_1743};
  assign _EVAL_1048 = _EVAL_28 & _EVAL_48;
  assign _EVAL_644 = _EVAL_3 == 3'h4;
  assign _EVAL_145 = _EVAL_23[11:2];
  assign _EVAL_181 = _EVAL_145[9];
  assign _EVAL_219 = _EVAL_145[7];
  assign _EVAL_1000 = _EVAL_145[6];
  assign _EVAL_1908 = _EVAL_145[5];
  assign _EVAL_1774 = _EVAL_145[4];
  assign _EVAL_1405 = _EVAL_145[3];
  assign _EVAL_1054 = _EVAL_145[2];
  assign _EVAL_1573 = _EVAL_145[1];
  assign _EVAL_1853 = _EVAL_145[0];
  assign _EVAL_390 = {_EVAL_181,_EVAL_219,_EVAL_1000,_EVAL_1908,_EVAL_1774,_EVAL_1405,_EVAL_1054,_EVAL_1573,_EVAL_1853};
  assign _EVAL_631 = 512'h1 << _EVAL_390;
  assign _EVAL_643 = _EVAL_145 & 10'h100;
  assign _EVAL_502 = _EVAL_643 == 10'h0;
  assign _EVAL_1760 = _EVAL_631[221];
  assign _EVAL_1604 = _EVAL_14[3];
  assign _EVAL_1076 = _EVAL_1604 ? 8'hff : 8'h0;
  assign _EVAL_1928 = _EVAL_14[2];
  assign _EVAL_1567 = _EVAL_1928 ? 8'hff : 8'h0;
  assign _EVAL_2187 = _EVAL_14[1];
  assign _EVAL_1668 = _EVAL_2187 ? 8'hff : 8'h0;
  assign _EVAL_1292 = _EVAL_14[0];
  assign _EVAL_1707 = _EVAL_1292 ? 8'hff : 8'h0;
  assign _EVAL_332 = {_EVAL_1076,_EVAL_1567,_EVAL_1668,_EVAL_1707};
  assign _EVAL_1017 = _EVAL_332[31:24];
  assign _EVAL_1486 = _EVAL_631[208];
  assign _EVAL_1500 = {_EVAL_1040,_EVAL_1768,_EVAL_1562,_EVAL_438};
  assign _EVAL_1492 = _EVAL_13 & _EVAL_18;
  assign _EVAL_681 = _EVAL_9 == 3'h4;
  assign _EVAL_1503 = _EVAL_681 == 1'h0;
  assign _EVAL_2076 = _EVAL_1492 & _EVAL_1503;
  assign _EVAL_177 = _EVAL_32[8:2];
  assign _EVAL_583 = _EVAL_177[5];
  assign _EVAL_171 = _EVAL_177[4];
  assign _EVAL_540 = _EVAL_177[3];
  assign _EVAL_594 = _EVAL_177[2];
  assign _EVAL_1878 = _EVAL_177[1];
  assign _EVAL_1632 = _EVAL_177[0];
  assign _EVAL_433 = {_EVAL_583,_EVAL_171,_EVAL_540,_EVAL_594,_EVAL_1878,_EVAL_1632};
  assign _EVAL_1421 = 64'h1 << _EVAL_433;
  assign _EVAL_610 = _EVAL_1421[33];
  assign _EVAL_376 = _EVAL_2076 & _EVAL_610;
  assign _EVAL_2056 = _EVAL_177 & 7'h40;
  assign _EVAL_680 = _EVAL_2056 == 7'h0;
  assign _EVAL_581 = _EVAL_376 & _EVAL_680;
  assign _EVAL_2136 = _EVAL_1582[31:24];
  assign _EVAL_1964 = _EVAL_2136 == 8'hff;
  assign _EVAL_139 = _EVAL_581 & _EVAL_1964;
  assign _EVAL_1971 = _EVAL_838 == 2'h0;
  assign _EVAL_1858 = _EVAL_139 & _EVAL_1971;
  assign _EVAL_142 = _EVAL_34[31:24];
  assign _EVAL_1992 = _EVAL_644 == 1'h0;
  assign _EVAL_749 = _EVAL_1048 & _EVAL_1992;
  assign _EVAL_573 = _EVAL_332[23:16];
  assign _EVAL_1387 = _EVAL_573 == 8'hff;
  assign _EVAL_1691 = 6'h20 == _EVAL_433;
  assign _EVAL_1961 = _EVAL_1421[43];
  assign _EVAL_646 = _EVAL_2076 & _EVAL_1961;
  assign _EVAL_1686 = _EVAL_646 & _EVAL_680;
  assign _EVAL_366 = _EVAL_1582[23:16];
  assign _EVAL_234 = _EVAL_366 == 8'hff;
  assign _EVAL_1145 = _EVAL_1686 & _EVAL_234;
  assign _EVAL_1459 = _EVAL_1145 & _EVAL_1971;
  assign _EVAL_55 = _EVAL_34[23:16];
  assign _EVAL_729 = sb2tlOpt__EVAL_14 != 3'h0;
  assign _EVAL_1323 = {1'h0,_EVAL_284,_EVAL_212,_EVAL_1803};
  assign _EVAL_1537 = _EVAL_1323[2:0];
  assign _EVAL_106 = {1'h0,_EVAL_734,_EVAL_729,_EVAL_1951,_EVAL_2167,_EVAL_1829,_EVAL_2117,_EVAL_1537,12'h407};
  assign _EVAL_1563 = _EVAL_332[7:0];
  assign _EVAL_758 = _EVAL_1563 == 8'hff;
  assign _EVAL_886 = _EVAL_631[212];
  assign _EVAL_57 = _EVAL_631[218];
  assign _EVAL_1020 = _EVAL_749 & _EVAL_57;
  assign _EVAL_1319 = _EVAL_1020 & _EVAL_502;
  assign _EVAL_1753 = _EVAL_332[15:8];
  assign _EVAL_1638 = _EVAL_1753 == 8'hff;
  assign _EVAL_857 = _EVAL_1319 & _EVAL_1638;
  assign _EVAL_2029 = {96'h0,_EVAL_34};
  assign _EVAL_531 = _EVAL_1421[47];
  assign _EVAL_1009 = _EVAL_2076 & _EVAL_531;
  assign _EVAL_714 = _EVAL_1009 & _EVAL_680;
  assign _EVAL_1093 = _EVAL_714 & _EVAL_234;
  assign _EVAL_568 = _EVAL_1421[57];
  assign _EVAL_1556 = _EVAL_2076 & _EVAL_568;
  assign _EVAL_451 = _EVAL_1556 & _EVAL_680;
  assign _EVAL_214 = _EVAL_1582 == 32'hffffffff;
  assign _EVAL_1732 = _EVAL_451 & _EVAL_214;
  assign _EVAL_305 = _EVAL_1732 & _EVAL_729;
  assign _EVAL_1303 = _EVAL_1492 & _EVAL_681;
  assign _EVAL_1376 = _EVAL_1421[60];
  assign _EVAL_1580 = _EVAL_1303 & _EVAL_1376;
  assign _EVAL_633 = _EVAL_1580 & _EVAL_680;
  assign _EVAL_2178 = _EVAL_1582 != 32'h0;
  assign _EVAL_1311 = _EVAL_633 & _EVAL_2178;
  assign _EVAL_603 = _EVAL_2076 & _EVAL_1376;
  assign _EVAL_1782 = _EVAL_603 & _EVAL_680;
  assign _EVAL_1501 = _EVAL_1782 & _EVAL_214;
  assign _EVAL_1078 = _EVAL_1311 | _EVAL_1501;
  assign _EVAL_1780 = _EVAL_1078 & _EVAL_729;
  assign _EVAL_518 = 6'h21 == _EVAL_433;
  assign _EVAL_109 = 6'h22 == _EVAL_433;
  assign _EVAL_721 = 6'h23 == _EVAL_433;
  assign _EVAL_1737 = 6'h24 == _EVAL_433;
  assign _EVAL_987 = 6'h25 == _EVAL_433;
  assign _EVAL_205 = 6'h26 == _EVAL_433;
  assign _EVAL_1274 = 6'h27 == _EVAL_433;
  assign _EVAL_1085 = 6'h28 == _EVAL_433;
  assign _EVAL_153 = 6'h29 == _EVAL_433;
  assign _EVAL_750 = 6'h2a == _EVAL_433;
  assign _EVAL_1299 = 6'h2b == _EVAL_433;
  assign _EVAL_1607 = 6'h2c == _EVAL_433;
  assign _EVAL_224 = 6'h2d == _EVAL_433;
  assign _EVAL_1209 = 6'h2e == _EVAL_433;
  assign _EVAL_420 = 6'h2f == _EVAL_433;
  assign _EVAL_900 = 6'h38 == _EVAL_433;
  assign _EVAL_1615 = 6'h39 == _EVAL_433;
  assign _EVAL_924 = 6'h3c == _EVAL_433;
  assign _EVAL_350 = _EVAL_924 ? _EVAL_680 : 1'h1;
  assign _EVAL_2148 = _EVAL_1615 ? _EVAL_680 : _EVAL_350;
  assign _EVAL_505 = _EVAL_900 ? _EVAL_680 : _EVAL_2148;
  assign _EVAL_374 = _EVAL_420 ? _EVAL_680 : _EVAL_505;
  assign _EVAL_1590 = _EVAL_1209 ? _EVAL_680 : _EVAL_374;
  assign _EVAL_2031 = _EVAL_224 ? _EVAL_680 : _EVAL_1590;
  assign _EVAL_1424 = _EVAL_1607 ? _EVAL_680 : _EVAL_2031;
  assign _EVAL_1312 = _EVAL_1299 ? _EVAL_680 : _EVAL_1424;
  assign _EVAL_1830 = _EVAL_750 ? _EVAL_680 : _EVAL_1312;
  assign _EVAL_715 = _EVAL_153 ? _EVAL_680 : _EVAL_1830;
  assign _EVAL_1736 = _EVAL_1085 ? _EVAL_680 : _EVAL_715;
  assign _EVAL_752 = _EVAL_1274 ? _EVAL_680 : _EVAL_1736;
  assign _EVAL_1331 = _EVAL_205 ? _EVAL_680 : _EVAL_752;
  assign _EVAL_1745 = _EVAL_987 ? _EVAL_680 : _EVAL_1331;
  assign _EVAL_560 = _EVAL_1737 ? _EVAL_680 : _EVAL_1745;
  assign _EVAL_753 = _EVAL_721 ? _EVAL_680 : _EVAL_560;
  assign _EVAL_779 = _EVAL_109 ? _EVAL_680 : _EVAL_753;
  assign _EVAL_1086 = _EVAL_518 ? _EVAL_680 : _EVAL_779;
  assign _EVAL_127 = _EVAL_1691 ? _EVAL_680 : _EVAL_1086;
  assign _EVAL_1709 = _EVAL_1582[20];
  assign _EVAL_1119 = 9'hce == _EVAL_390;
  assign _EVAL_1966 = 9'hcf == _EVAL_390;
  assign _EVAL_529 = 9'hd0 == _EVAL_390;
  assign _EVAL_165 = 9'hd1 == _EVAL_390;
  assign _EVAL_901 = 9'hd2 == _EVAL_390;
  assign _EVAL_1931 = 9'hd3 == _EVAL_390;
  assign _EVAL_1090 = 9'hd4 == _EVAL_390;
  assign _EVAL_2051 = 9'hd5 == _EVAL_390;
  assign _EVAL_189 = 9'hd6 == _EVAL_390;
  assign _EVAL_1449 = 9'hd7 == _EVAL_390;
  assign _EVAL_173 = 9'hd8 == _EVAL_390;
  assign _EVAL_827 = 9'hd9 == _EVAL_390;
  assign _EVAL_1841 = 9'hda == _EVAL_390;
  assign _EVAL_869 = 9'hdb == _EVAL_390;
  assign _EVAL_2150 = 9'hdc == _EVAL_390;
  assign _EVAL_462 = 9'hdd == _EVAL_390;
  assign _EVAL_862 = 9'hde == _EVAL_390;
  assign _EVAL_2125 = 9'hdf == _EVAL_390;
  assign _EVAL_67 = 9'he0 == _EVAL_390;
  assign _EVAL_395 = 9'h100 == _EVAL_390;
  assign _EVAL_2006 = 9'h101 == _EVAL_390;
  assign _EVAL_1059 = 9'h102 == _EVAL_390;
  assign _EVAL_612 = 9'h103 == _EVAL_390;
  assign _EVAL_447 = 9'h104 == _EVAL_390;
  assign _EVAL_950 = 9'h105 == _EVAL_390;
  assign _EVAL_1050 = 9'h106 == _EVAL_390;
  assign _EVAL_382 = 9'h107 == _EVAL_390;
  assign _EVAL_1381 = 9'h108 == _EVAL_390;
  assign _EVAL_159 = 9'h109 == _EVAL_390;
  assign _EVAL_1464 = 9'h10a == _EVAL_390;
  assign _EVAL_266 = 9'h10b == _EVAL_390;
  assign _EVAL_2104 = 9'h10c == _EVAL_390;
  assign _EVAL_1175 = 9'h10d == _EVAL_390;
  assign _EVAL_1844 = 9'h10e == _EVAL_390;
  assign _EVAL_453 = 9'h10f == _EVAL_390;
  assign _EVAL_255 = 9'h110 == _EVAL_390;
  assign _EVAL_268 = 9'h111 == _EVAL_390;
  assign _EVAL_823 = 9'h112 == _EVAL_390;
  assign _EVAL_1696 = 9'h113 == _EVAL_390;
  assign _EVAL_2126 = 9'h114 == _EVAL_390;
  assign _EVAL_1114 = _EVAL_2126 ? _EVAL_502 : 1'h1;
  assign _EVAL_883 = _EVAL_1696 ? _EVAL_502 : _EVAL_1114;
  assign _EVAL_1628 = _EVAL_823 ? _EVAL_502 : _EVAL_883;
  assign _EVAL_818 = _EVAL_268 ? _EVAL_502 : _EVAL_1628;
  assign _EVAL_140 = _EVAL_255 ? _EVAL_502 : _EVAL_818;
  assign _EVAL_2215 = _EVAL_453 ? _EVAL_502 : _EVAL_140;
  assign _EVAL_1494 = _EVAL_1844 ? _EVAL_502 : _EVAL_2215;
  assign _EVAL_1470 = _EVAL_1175 ? _EVAL_502 : _EVAL_1494;
  assign _EVAL_415 = _EVAL_2104 ? _EVAL_502 : _EVAL_1470;
  assign _EVAL_381 = _EVAL_266 ? _EVAL_502 : _EVAL_415;
  assign _EVAL_1483 = _EVAL_1464 ? _EVAL_502 : _EVAL_381;
  assign _EVAL_1335 = _EVAL_159 ? _EVAL_502 : _EVAL_1483;
  assign _EVAL_771 = _EVAL_1381 ? _EVAL_502 : _EVAL_1335;
  assign _EVAL_193 = _EVAL_382 ? _EVAL_502 : _EVAL_771;
  assign _EVAL_1245 = _EVAL_1050 ? _EVAL_502 : _EVAL_193;
  assign _EVAL_885 = _EVAL_950 ? _EVAL_502 : _EVAL_1245;
  assign _EVAL_1744 = _EVAL_447 ? _EVAL_502 : _EVAL_885;
  assign _EVAL_516 = _EVAL_612 ? _EVAL_502 : _EVAL_1744;
  assign _EVAL_1270 = _EVAL_1059 ? _EVAL_502 : _EVAL_516;
  assign _EVAL_547 = _EVAL_2006 ? _EVAL_502 : _EVAL_1270;
  assign _EVAL_1392 = _EVAL_395 ? _EVAL_502 : _EVAL_547;
  assign _EVAL_1226 = _EVAL_67 ? _EVAL_502 : _EVAL_1392;
  assign _EVAL_621 = _EVAL_2125 ? _EVAL_502 : _EVAL_1226;
  assign _EVAL_261 = _EVAL_862 ? _EVAL_502 : _EVAL_621;
  assign _EVAL_1008 = _EVAL_462 ? _EVAL_502 : _EVAL_261;
  assign _EVAL_148 = _EVAL_2150 ? _EVAL_502 : _EVAL_1008;
  assign _EVAL_934 = _EVAL_869 ? _EVAL_502 : _EVAL_148;
  assign _EVAL_1036 = _EVAL_1841 ? _EVAL_502 : _EVAL_934;
  assign _EVAL_1549 = _EVAL_827 ? _EVAL_502 : _EVAL_1036;
  assign _EVAL_2169 = _EVAL_173 ? _EVAL_502 : _EVAL_1549;
  assign _EVAL_114 = _EVAL_1449 ? _EVAL_502 : _EVAL_2169;
  assign _EVAL_2111 = _EVAL_189 ? _EVAL_502 : _EVAL_114;
  assign _EVAL_742 = _EVAL_2051 ? _EVAL_502 : _EVAL_2111;
  assign _EVAL_364 = _EVAL_1090 ? _EVAL_502 : _EVAL_742;
  assign _EVAL_655 = _EVAL_1931 ? _EVAL_502 : _EVAL_364;
  assign _EVAL_772 = _EVAL_901 ? _EVAL_502 : _EVAL_655;
  assign _EVAL_1979 = _EVAL_165 ? _EVAL_502 : _EVAL_772;
  assign _EVAL_1968 = _EVAL_529 ? _EVAL_502 : _EVAL_1979;
  assign _EVAL_64 = _EVAL_1966 ? _EVAL_502 : _EVAL_1968;
  assign _EVAL_2101 = _EVAL_1119 ? _EVAL_502 : _EVAL_64;
  assign _EVAL_2106 = _EVAL_1421[36];
  assign _EVAL_370 = _EVAL_2076 & _EVAL_2106;
  assign _EVAL_1986 = _EVAL_370 & _EVAL_680;
  assign _EVAL_1888 = _EVAL_1582[15:8];
  assign _EVAL_1246 = _EVAL_1888 == 8'hff;
  assign _EVAL_614 = _EVAL_1986 & _EVAL_1246;
  assign _EVAL_129 = _EVAL_631[67];
  assign _EVAL_507 = _EVAL_1421[40];
  assign _EVAL_168 = _EVAL_2076 & _EVAL_507;
  assign _EVAL_1824 = _EVAL_168 & _EVAL_680;
  assign _EVAL_1286 = _EVAL_1824 & _EVAL_234;
  assign _EVAL_410 = _EVAL_1286 & _EVAL_1971;
  assign _EVAL_299 = _EVAL_1421[22];
  assign _EVAL_538 = _EVAL_1732 & _EVAL_1951;
  assign _EVAL_2235 = _EVAL_1311 & _EVAL_2117;
  assign _EVAL_2137 = _EVAL_538 | _EVAL_2235;
  assign _EVAL_1545 = _EVAL_1501 | _EVAL_2137;
  assign _EVAL_339 = _EVAL_366 != 8'h0;
  assign _EVAL_545 = {_EVAL_1649,_EVAL_1055,_EVAL_1264,_EVAL_130};
  assign _EVAL_1799 = {_EVAL_2058,_EVAL_229,_EVAL_858,_EVAL_1859};
  assign _EVAL_1141 = {_EVAL_1370,_EVAL_658,_EVAL_739,_EVAL_92};
  assign _EVAL_1658 = {_EVAL_2057,_EVAL_2154,_EVAL_1599,_EVAL_2165};
  assign _EVAL_1635 = {_EVAL_1785,_EVAL_1200,_EVAL_961,_EVAL_1447};
  assign _EVAL_1302 = {_EVAL_915,_EVAL_1646,_EVAL_1869,_EVAL_1652};
  assign _EVAL_905 = {_EVAL_732,_EVAL_1694,_EVAL_72,_EVAL_182};
  assign _EVAL_478 = {_EVAL_1100,_EVAL_174,_EVAL_1943,_EVAL_329};
  assign _EVAL_2234 = {_EVAL_804,_EVAL_881,_EVAL_532,_EVAL_846};
  assign _EVAL_2182 = _EVAL_2126 ? 32'h100073 : 32'h0;
  assign _EVAL_222 = _EVAL_1696 ? 32'h10002623 : _EVAL_2182;
  assign _EVAL_460 = _EVAL_823 ? 32'h7b200073 : _EVAL_222;
  assign _EVAL_1810 = _EVAL_268 ? 32'h7b202473 : _EVAL_460;
  assign _EVAL_490 = _EVAL_255 ? 32'h10802423 : _EVAL_1810;
  assign _EVAL_1704 = _EVAL_453 ? 32'hf1402473 : _EVAL_490;
  assign _EVAL_2181 = _EVAL_1844 ? 32'h30000067 : _EVAL_1704;
  assign _EVAL_794 = _EVAL_1175 ? 32'h10002223 : _EVAL_2181;
  assign _EVAL_1398 = _EVAL_2104 ? 32'h7b202473 : _EVAL_794;
  assign _EVAL_1356 = _EVAL_266 ? 32'h40863 : _EVAL_1398;
  assign _EVAL_741 = _EVAL_1464 ? 32'h147413 : _EVAL_1356;
  assign _EVAL_495 = _EVAL_159 ? 32'hfe0408e3 : _EVAL_741;
  assign _EVAL_1253 = _EVAL_1381 ? 32'h347413 : _EVAL_495;
  assign _EVAL_228 = _EVAL_382 ? 32'h40044403 : _EVAL_1253;
  assign _EVAL_443 = _EVAL_1050 ? 32'h10802023 : _EVAL_228;
  assign _EVAL_248 = _EVAL_950 ? 32'hf1402473 : _EVAL_443;
  assign _EVAL_1360 = _EVAL_447 ? 32'h7b241073 : _EVAL_248;
  assign _EVAL_757 = _EVAL_612 ? 32'hff0000f : _EVAL_1360;
  assign _EVAL_1131 = _EVAL_1059 ? 32'h440006f : _EVAL_757;
  assign _EVAL_795 = _EVAL_2006 ? 32'h380006f : _EVAL_1131;
  assign _EVAL_1860 = _EVAL_395 ? 32'hc0006f : _EVAL_795;
  assign _EVAL_1359 = _EVAL_67 ? _EVAL_2234 : _EVAL_1860;
  assign _EVAL_1577 = _EVAL_2125 ? _EVAL_1500 : _EVAL_1359;
  assign _EVAL_1345 = _EVAL_862 ? _EVAL_478 : _EVAL_1577;
  assign _EVAL_110 = _EVAL_462 ? _EVAL_905 : _EVAL_1345;
  assign _EVAL_1451 = _EVAL_2150 ? _EVAL_1302 : _EVAL_110;
  assign _EVAL_904 = _EVAL_869 ? _EVAL_1635 : _EVAL_1451;
  assign _EVAL_353 = _EVAL_1841 ? _EVAL_1658 : _EVAL_904;
  assign _EVAL_196 = _EVAL_827 ? _EVAL_1141 : _EVAL_353;
  assign _EVAL_716 = _EVAL_173 ? _EVAL_1799 : _EVAL_196;
  assign _EVAL_1419 = _EVAL_1449 ? _EVAL_545 : _EVAL_716;
  assign _EVAL_637 = _EVAL_631[211];
  assign _EVAL_1900 = _EVAL_1421[4];
  assign _EVAL_627 = _EVAL_2076 & _EVAL_1900;
  assign _EVAL_1366 = _EVAL_627 & _EVAL_680;
  assign _EVAL_1608 = _EVAL_1366 & _EVAL_1246;
  assign _EVAL_880 = _EVAL_1421[34];
  assign _EVAL_1096 = _EVAL_2076 & _EVAL_880;
  assign _EVAL_295 = _EVAL_1096 & _EVAL_680;
  assign _EVAL_994 = _EVAL_295 & _EVAL_1246;
  assign _EVAL_2060 = _EVAL_34[15:8];
  assign _EVAL_423 = _EVAL_2076 & _EVAL_299;
  assign _EVAL_328 = _EVAL_423 & _EVAL_680;
  assign _EVAL_2095 = _EVAL_631[219];
  assign _EVAL_2017 = _EVAL_749 & _EVAL_2095;
  assign _EVAL_1798 = _EVAL_2017 & _EVAL_502;
  assign _EVAL_986 = _EVAL_1798 & _EVAL_1387;
  assign _EVAL_1845 = _EVAL_631[66];
  assign _EVAL_190 = _EVAL_332[9:0];
  assign _EVAL_1188 = _EVAL_631[217];
  assign _EVAL_2080 = _EVAL_1421[46];
  assign _EVAL_272 = _EVAL_2076 & _EVAL_2080;
  assign _EVAL_665 = _EVAL_272 & _EVAL_680;
  assign _EVAL_1831 = _EVAL_665 & _EVAL_1246;
  assign _EVAL_539 = _EVAL_1831 & _EVAL_1971;
  assign _EVAL_731 = _EVAL_1421[32];
  assign _EVAL_1104 = _EVAL_2076 & _EVAL_731;
  assign _EVAL_1304 = _EVAL_1104 & _EVAL_680;
  assign _EVAL_1827 = _EVAL_1582[7:0];
  assign _EVAL_619 = _EVAL_1827 == 8'hff;
  assign _EVAL_556 = _EVAL_1304 & _EVAL_619;
  assign _EVAL_820 = _EVAL_1303 & _EVAL_731;
  assign _EVAL_1880 = _EVAL_820 & _EVAL_680;
  assign _EVAL_107 = _EVAL_1827 != 8'h0;
  assign _EVAL_1558 = _EVAL_1880 & _EVAL_107;
  assign _EVAL_647 = _EVAL_556 | _EVAL_1558;
  assign _EVAL_1654 = _EVAL_1304 & _EVAL_1246;
  assign _EVAL_544 = _EVAL_1888 != 8'h0;
  assign _EVAL_1680 = _EVAL_1880 & _EVAL_544;
  assign _EVAL_2030 = _EVAL_1654 | _EVAL_1680;
  assign _EVAL_1720 = _EVAL_647 | _EVAL_2030;
  assign _EVAL_2102 = _EVAL_1304 & _EVAL_234;
  assign _EVAL_1570 = _EVAL_1880 & _EVAL_339;
  assign _EVAL_971 = _EVAL_2102 | _EVAL_1570;
  assign _EVAL_1742 = _EVAL_1720 | _EVAL_971;
  assign _EVAL_233 = _EVAL_1304 & _EVAL_1964;
  assign _EVAL_2190 = _EVAL_2136 != 8'h0;
  assign _EVAL_418 = _EVAL_1880 & _EVAL_2190;
  assign _EVAL_1400 = _EVAL_233 | _EVAL_418;
  assign _EVAL_1721 = _EVAL_1742 | _EVAL_1400;
  assign _EVAL_1532 = _EVAL_581 & _EVAL_619;
  assign _EVAL_1053 = _EVAL_1303 & _EVAL_610;
  assign _EVAL_1229 = _EVAL_1053 & _EVAL_680;
  assign _EVAL_2088 = _EVAL_1229 & _EVAL_107;
  assign _EVAL_2092 = _EVAL_1532 | _EVAL_2088;
  assign _EVAL_113 = _EVAL_1721 | _EVAL_2092;
  assign _EVAL_1551 = _EVAL_581 & _EVAL_1246;
  assign _EVAL_166 = _EVAL_1229 & _EVAL_544;
  assign _EVAL_1975 = _EVAL_1551 | _EVAL_166;
  assign _EVAL_727 = _EVAL_113 | _EVAL_1975;
  assign _EVAL_1163 = _EVAL_581 & _EVAL_234;
  assign _EVAL_1317 = _EVAL_1229 & _EVAL_339;
  assign _EVAL_569 = _EVAL_1163 | _EVAL_1317;
  assign _EVAL_2205 = _EVAL_727 | _EVAL_569;
  assign _EVAL_1192 = _EVAL_1229 & _EVAL_2190;
  assign _EVAL_360 = _EVAL_139 | _EVAL_1192;
  assign _EVAL_1038 = _EVAL_2205 | _EVAL_360;
  assign _EVAL_1296 = _EVAL_295 & _EVAL_619;
  assign _EVAL_333 = _EVAL_1303 & _EVAL_880;
  assign _EVAL_719 = _EVAL_333 & _EVAL_680;
  assign _EVAL_1133 = _EVAL_719 & _EVAL_107;
  assign _EVAL_914 = _EVAL_1296 | _EVAL_1133;
  assign _EVAL_736 = _EVAL_1038 | _EVAL_914;
  assign _EVAL_958 = _EVAL_719 & _EVAL_544;
  assign _EVAL_1524 = _EVAL_994 | _EVAL_958;
  assign _EVAL_204 = _EVAL_736 | _EVAL_1524;
  assign _EVAL_1171 = _EVAL_295 & _EVAL_234;
  assign _EVAL_1490 = _EVAL_719 & _EVAL_339;
  assign _EVAL_1756 = _EVAL_1171 | _EVAL_1490;
  assign _EVAL_1698 = _EVAL_204 | _EVAL_1756;
  assign _EVAL_884 = _EVAL_295 & _EVAL_1964;
  assign _EVAL_408 = _EVAL_719 & _EVAL_2190;
  assign _EVAL_1083 = _EVAL_884 | _EVAL_408;
  assign _EVAL_1636 = _EVAL_1698 | _EVAL_1083;
  assign _EVAL_1136 = _EVAL_1421[35];
  assign _EVAL_236 = _EVAL_2076 & _EVAL_1136;
  assign _EVAL_133 = _EVAL_236 & _EVAL_680;
  assign _EVAL_483 = _EVAL_133 & _EVAL_619;
  assign _EVAL_1947 = _EVAL_1303 & _EVAL_1136;
  assign _EVAL_2153 = _EVAL_1947 & _EVAL_680;
  assign _EVAL_620 = _EVAL_2153 & _EVAL_107;
  assign _EVAL_1318 = _EVAL_483 | _EVAL_620;
  assign _EVAL_1201 = _EVAL_1636 | _EVAL_1318;
  assign _EVAL_559 = _EVAL_133 & _EVAL_1246;
  assign _EVAL_1708 = _EVAL_2153 & _EVAL_544;
  assign _EVAL_1914 = _EVAL_559 | _EVAL_1708;
  assign _EVAL_1593 = _EVAL_1201 | _EVAL_1914;
  assign _EVAL_1752 = _EVAL_133 & _EVAL_234;
  assign _EVAL_2195 = _EVAL_2153 & _EVAL_339;
  assign _EVAL_1004 = _EVAL_1752 | _EVAL_2195;
  assign _EVAL_440 = _EVAL_1593 | _EVAL_1004;
  assign _EVAL_669 = _EVAL_133 & _EVAL_1964;
  assign _EVAL_1237 = _EVAL_2153 & _EVAL_2190;
  assign _EVAL_879 = _EVAL_669 | _EVAL_1237;
  assign _EVAL_303 = _EVAL_440 | _EVAL_879;
  assign _EVAL_1242 = _EVAL_1986 & _EVAL_619;
  assign _EVAL_1903 = _EVAL_1303 & _EVAL_2106;
  assign _EVAL_330 = _EVAL_1903 & _EVAL_680;
  assign _EVAL_686 = _EVAL_330 & _EVAL_107;
  assign _EVAL_104 = _EVAL_1242 | _EVAL_686;
  assign _EVAL_334 = _EVAL_303 | _EVAL_104;
  assign _EVAL_191 = _EVAL_330 & _EVAL_544;
  assign _EVAL_101 = _EVAL_614 | _EVAL_191;
  assign _EVAL_384 = _EVAL_334 | _EVAL_101;
  assign _EVAL_221 = _EVAL_1986 & _EVAL_234;
  assign _EVAL_1003 = _EVAL_330 & _EVAL_339;
  assign _EVAL_660 = _EVAL_221 | _EVAL_1003;
  assign _EVAL_264 = _EVAL_384 | _EVAL_660;
  assign _EVAL_957 = _EVAL_1986 & _EVAL_1964;
  assign _EVAL_2068 = _EVAL_330 & _EVAL_2190;
  assign _EVAL_519 = _EVAL_957 | _EVAL_2068;
  assign _EVAL_639 = _EVAL_264 | _EVAL_519;
  assign _EVAL_469 = _EVAL_631[214];
  assign _EVAL_361 = _EVAL_1421[23];
  assign _EVAL_760 = _EVAL_2076 & _EVAL_361;
  assign _EVAL_403 = _EVAL_760 & _EVAL_680;
  assign _EVAL_164 = _EVAL_403 & _EVAL_214;
  assign _EVAL_1322 = _EVAL_164 & _EVAL_1971;
  assign _EVAL_1965 = _EVAL_164 ? _EVAL_34 : 32'h0;
  assign _EVAL_1925 = _EVAL_1965[31:24];
  assign _EVAL_898 = _EVAL_1925 == 8'h0;
  assign _EVAL_2147 = _EVAL_1322 & _EVAL_898;
  assign _EVAL_61 = _EVAL_1263 == 3'h0;
  assign _EVAL_1254 = _EVAL_2147 & _EVAL_61;
  assign _EVAL_1838 = _EVAL_1366 & _EVAL_619;
  assign _EVAL_1473 = _EVAL_1303 & _EVAL_1900;
  assign _EVAL_2236 = _EVAL_1473 & _EVAL_680;
  assign _EVAL_1885 = _EVAL_2236 & _EVAL_107;
  assign _EVAL_1244 = _EVAL_1838 | _EVAL_1885;
  assign _EVAL_1854 = _EVAL_1135[0];
  assign _EVAL_1193 = _EVAL_1244 & _EVAL_1854;
  assign _EVAL_1094 = _EVAL_1137[0];
  assign _EVAL_1771 = _EVAL_647 & _EVAL_1094;
  assign _EVAL_548 = _EVAL_1137[1];
  assign _EVAL_1512 = _EVAL_2092 & _EVAL_548;
  assign _EVAL_918 = _EVAL_1771 | _EVAL_1512;
  assign _EVAL_237 = _EVAL_1137[2];
  assign _EVAL_1051 = _EVAL_914 & _EVAL_237;
  assign _EVAL_195 = _EVAL_918 | _EVAL_1051;
  assign _EVAL_455 = _EVAL_1318 & _EVAL_1129;
  assign _EVAL_2210 = _EVAL_195 | _EVAL_455;
  assign _EVAL_1630 = _EVAL_1137[4];
  assign _EVAL_508 = _EVAL_104 & _EVAL_1630;
  assign _EVAL_1491 = _EVAL_2210 | _EVAL_508;
  assign _EVAL_803 = _EVAL_1421[37];
  assign _EVAL_2161 = _EVAL_2076 & _EVAL_803;
  assign _EVAL_789 = _EVAL_2161 & _EVAL_680;
  assign _EVAL_1592 = _EVAL_789 & _EVAL_619;
  assign _EVAL_2233 = _EVAL_1303 & _EVAL_803;
  assign _EVAL_1057 = _EVAL_2233 & _EVAL_680;
  assign _EVAL_435 = _EVAL_1057 & _EVAL_107;
  assign _EVAL_2116 = _EVAL_1592 | _EVAL_435;
  assign _EVAL_244 = _EVAL_1137[5];
  assign _EVAL_1791 = _EVAL_2116 & _EVAL_244;
  assign _EVAL_2086 = _EVAL_1491 | _EVAL_1791;
  assign _EVAL_1993 = _EVAL_1421[38];
  assign _EVAL_439 = _EVAL_2076 & _EVAL_1993;
  assign _EVAL_1458 = _EVAL_439 & _EVAL_680;
  assign _EVAL_2192 = _EVAL_1458 & _EVAL_619;
  assign _EVAL_570 = _EVAL_1303 & _EVAL_1993;
  assign _EVAL_461 = _EVAL_570 & _EVAL_680;
  assign _EVAL_590 = _EVAL_461 & _EVAL_107;
  assign _EVAL_1662 = _EVAL_2192 | _EVAL_590;
  assign _EVAL_1548 = _EVAL_1137[6];
  assign _EVAL_836 = _EVAL_1662 & _EVAL_1548;
  assign _EVAL_553 = _EVAL_2086 | _EVAL_836;
  assign _EVAL_692 = _EVAL_1421[39];
  assign _EVAL_988 = _EVAL_2076 & _EVAL_692;
  assign _EVAL_1308 = _EVAL_988 & _EVAL_680;
  assign _EVAL_1535 = _EVAL_1308 & _EVAL_619;
  assign _EVAL_702 = _EVAL_1303 & _EVAL_692;
  assign _EVAL_970 = _EVAL_702 & _EVAL_680;
  assign _EVAL_1103 = _EVAL_970 & _EVAL_107;
  assign _EVAL_200 = _EVAL_1535 | _EVAL_1103;
  assign _EVAL_1982 = _EVAL_1137[7];
  assign _EVAL_436 = _EVAL_200 & _EVAL_1982;
  assign _EVAL_1305 = _EVAL_553 | _EVAL_436;
  assign _EVAL_1750 = _EVAL_1824 & _EVAL_619;
  assign _EVAL_1079 = _EVAL_1303 & _EVAL_507;
  assign _EVAL_1932 = _EVAL_1079 & _EVAL_680;
  assign _EVAL_1071 = _EVAL_1932 & _EVAL_107;
  assign _EVAL_442 = _EVAL_1750 | _EVAL_1071;
  assign _EVAL_1962 = _EVAL_1137[8];
  assign _EVAL_401 = _EVAL_442 & _EVAL_1962;
  assign _EVAL_1879 = _EVAL_1305 | _EVAL_401;
  assign _EVAL_1062 = _EVAL_1421[41];
  assign _EVAL_136 = _EVAL_2076 & _EVAL_1062;
  assign _EVAL_1872 = _EVAL_136 & _EVAL_680;
  assign _EVAL_1773 = _EVAL_1872 & _EVAL_619;
  assign _EVAL_1239 = _EVAL_1303 & _EVAL_1062;
  assign _EVAL_94 = _EVAL_1239 & _EVAL_680;
  assign _EVAL_1998 = _EVAL_94 & _EVAL_107;
  assign _EVAL_1769 = _EVAL_1773 | _EVAL_1998;
  assign _EVAL_96 = _EVAL_1137[9];
  assign _EVAL_1157 = _EVAL_1769 & _EVAL_96;
  assign _EVAL_1893 = _EVAL_1879 | _EVAL_1157;
  assign _EVAL_1044 = _EVAL_1421[42];
  assign _EVAL_2093 = _EVAL_2076 & _EVAL_1044;
  assign _EVAL_865 = _EVAL_2093 & _EVAL_680;
  assign _EVAL_517 = _EVAL_865 & _EVAL_619;
  assign _EVAL_693 = _EVAL_1303 & _EVAL_1044;
  assign _EVAL_2127 = _EVAL_693 & _EVAL_680;
  assign _EVAL_833 = _EVAL_2127 & _EVAL_107;
  assign _EVAL_1772 = _EVAL_517 | _EVAL_833;
  assign _EVAL_2094 = _EVAL_1137[10];
  assign _EVAL_270 = _EVAL_1772 & _EVAL_2094;
  assign _EVAL_1765 = _EVAL_1893 | _EVAL_270;
  assign _EVAL_320 = _EVAL_1686 & _EVAL_619;
  assign _EVAL_839 = _EVAL_1303 & _EVAL_1961;
  assign _EVAL_1610 = _EVAL_839 & _EVAL_680;
  assign _EVAL_1677 = _EVAL_1610 & _EVAL_107;
  assign _EVAL_1836 = _EVAL_320 | _EVAL_1677;
  assign _EVAL_1277 = _EVAL_1137[11];
  assign _EVAL_2044 = _EVAL_1836 & _EVAL_1277;
  assign _EVAL_1637 = _EVAL_1765 | _EVAL_2044;
  assign _EVAL_756 = _EVAL_1421[44];
  assign _EVAL_790 = _EVAL_2076 & _EVAL_756;
  assign _EVAL_530 = _EVAL_790 & _EVAL_680;
  assign _EVAL_1598 = _EVAL_530 & _EVAL_619;
  assign _EVAL_380 = _EVAL_1303 & _EVAL_756;
  assign _EVAL_144 = _EVAL_380 & _EVAL_680;
  assign _EVAL_1820 = _EVAL_144 & _EVAL_107;
  assign _EVAL_695 = _EVAL_1598 | _EVAL_1820;
  assign _EVAL_1243 = _EVAL_1137[12];
  assign _EVAL_1840 = _EVAL_695 & _EVAL_1243;
  assign _EVAL_1722 = _EVAL_1637 | _EVAL_1840;
  assign _EVAL_504 = _EVAL_1421[45];
  assign _EVAL_372 = _EVAL_2076 & _EVAL_504;
  assign _EVAL_247 = _EVAL_372 & _EVAL_680;
  assign _EVAL_319 = _EVAL_247 & _EVAL_619;
  assign _EVAL_2087 = _EVAL_1303 & _EVAL_504;
  assign _EVAL_743 = _EVAL_2087 & _EVAL_680;
  assign _EVAL_1480 = _EVAL_743 & _EVAL_107;
  assign _EVAL_85 = _EVAL_319 | _EVAL_1480;
  assign _EVAL_1138 = _EVAL_1137[13];
  assign _EVAL_2069 = _EVAL_85 & _EVAL_1138;
  assign _EVAL_53 = _EVAL_1722 | _EVAL_2069;
  assign _EVAL_728 = _EVAL_665 & _EVAL_619;
  assign _EVAL_2012 = _EVAL_1303 & _EVAL_2080;
  assign _EVAL_1276 = _EVAL_2012 & _EVAL_680;
  assign _EVAL_1225 = _EVAL_1276 & _EVAL_107;
  assign _EVAL_740 = _EVAL_728 | _EVAL_1225;
  assign _EVAL_1374 = _EVAL_1137[14];
  assign _EVAL_2202 = _EVAL_740 & _EVAL_1374;
  assign _EVAL_1927 = _EVAL_53 | _EVAL_2202;
  assign _EVAL_1889 = _EVAL_714 & _EVAL_619;
  assign _EVAL_1334 = _EVAL_1303 & _EVAL_531;
  assign _EVAL_2225 = _EVAL_1334 & _EVAL_680;
  assign _EVAL_141 = _EVAL_2225 & _EVAL_107;
  assign _EVAL_437 = _EVAL_1889 | _EVAL_141;
  assign _EVAL_936 = _EVAL_1137[15];
  assign _EVAL_1396 = _EVAL_437 & _EVAL_936;
  assign _EVAL_1174 = _EVAL_1927 | _EVAL_1396;
  assign _EVAL_1960 = _EVAL_1193 | _EVAL_1174;
  assign _EVAL_407 = _EVAL_1154 == 8'h0;
  assign _EVAL_859 = _EVAL_1960 & _EVAL_407;
  assign _EVAL_773 = _EVAL_859 & _EVAL_61;
  assign _EVAL_1361 = _EVAL_1254 | _EVAL_773;
  assign _EVAL_175 = _EVAL_1017 == 8'hff;
  assign _EVAL_1222 = _EVAL_1824 & _EVAL_1964;
  assign _EVAL_2185 = _EVAL_1222 & _EVAL_1971;
  assign _EVAL_1847 = _EVAL_461 & _EVAL_2190;
  assign _EVAL_1391 = _EVAL_631[209];
  assign _EVAL_953 = _EVAL_665 & _EVAL_234;
  assign _EVAL_2146 = _EVAL_953 & _EVAL_1971;
  assign _EVAL_726 = {_EVAL_1154,_EVAL_623};
  assign _EVAL_1327 = _EVAL_726[18];
  assign _EVAL_471 = _EVAL_616 == 1'h0;
  assign _EVAL_2004 = _EVAL_1501 & _EVAL_471;
  assign _EVAL_137 = _EVAL_734 == 1'h0;
  assign _EVAL_1538 = _EVAL_2004 & _EVAL_137;
  assign _EVAL_1815 = _EVAL_1537 == 3'h0;
  assign _EVAL_801 = _EVAL_1538 & _EVAL_1815;
  assign _EVAL_558 = _EVAL_749 & _EVAL_637;
  assign _EVAL_985 = _EVAL_558 & _EVAL_502;
  assign _EVAL_1959 = _EVAL_985 & _EVAL_175;
  assign _EVAL_256 = _EVAL_1308 & _EVAL_1964;
  assign _EVAL_1169 = _EVAL_2137 & _EVAL_471;
  assign _EVAL_1301 = _EVAL_1169 & _EVAL_137;
  assign _EVAL_2110 = _EVAL_256 & _EVAL_1971;
  assign _EVAL_774 = _EVAL_726[16];
  assign _EVAL_2081 = _EVAL_726[22:20];
  assign _EVAL_1644 = _EVAL_726[15:0];
  assign _EVAL_2238 = _EVAL_1644 & 16'h1f;
  assign _EVAL_345 = _EVAL_2238[4:0];
  assign _EVAL_882 = {17'h7000,_EVAL_2081,_EVAL_345,7'h3};
  assign _EVAL_1800 = {7'h1c,_EVAL_345,5'h0,_EVAL_2081,5'h0,7'h23};
  assign _EVAL_172 = _EVAL_631[222];
  assign _EVAL_2011 = _EVAL_2167 == 3'h4;
  assign _EVAL_445 = _EVAL_1732 ? _EVAL_34 : _EVAL_916;
  assign _EVAL_1121 = _EVAL_445[3:0];
  assign _EVAL_1702 = _EVAL_1121 != 4'h0;
  assign _EVAL_778 = _EVAL_2011 & _EVAL_1702;
  assign _EVAL_126 = _EVAL_1732 & _EVAL_1815;
  assign _EVAL_1843 = _EVAL_749 & _EVAL_129;
  assign _EVAL_989 = _EVAL_1421[56];
  assign _EVAL_1484 = _EVAL_2076 & _EVAL_989;
  assign _EVAL_979 = _EVAL_1484 & _EVAL_680;
  assign _EVAL_349 = _EVAL_1582[22];
  assign _EVAL_1153 = _EVAL_979 & _EVAL_349;
  assign _EVAL_767 = _EVAL_749 & _EVAL_1188;
  assign _EVAL_452 = _EVAL_767 & _EVAL_502;
  assign _EVAL_1988 = _EVAL_452 & _EVAL_1387;
  assign _EVAL_465 = _EVAL_517 & _EVAL_1971;
  assign _EVAL_1352 = _EVAL_34[7:0];
  assign _EVAL_1429 = _EVAL_631[215];
  assign _EVAL_1251 = _EVAL_749 & _EVAL_1429;
  assign _EVAL_1198 = _EVAL_1251 & _EVAL_502;
  assign _EVAL_1703 = _EVAL_1198 & _EVAL_175;
  assign _EVAL_1755 = _EVAL_36[31:24];
  assign _EVAL_2224 = _EVAL_838 == 2'h1;
  assign _EVAL_311 = _EVAL_2056 == 7'h40;
  assign _EVAL_766 = _EVAL_2236 & _EVAL_544;
  assign _EVAL_1160 = _EVAL_1608 | _EVAL_766;
  assign _EVAL_73 = _EVAL_726[17];
  assign _EVAL_321 = _EVAL_73 == 1'h0;
  assign _EVAL_105 = _EVAL_1644 >= 16'h1000;
  assign _EVAL_273 = _EVAL_1644 <= 16'h101f;
  assign _EVAL_847 = _EVAL_105 & _EVAL_273;
  assign _EVAL_199 = _EVAL_321 | _EVAL_847;
  assign _EVAL_485 = _EVAL_199 ? 1'h0 : 1'h1;
  assign _EVAL_962 = _EVAL_407 ? _EVAL_485 : 1'h1;
  assign _EVAL_1266 = ~ _EVAL_1065;
  assign _EVAL_630 = _EVAL_199 ? _EVAL_1266 : 1'h0;
  assign _EVAL_920 = _EVAL_407 ? _EVAL_630 : 1'h0;
  assign _EVAL_1554 = _EVAL_962 ? 1'h0 : _EVAL_920;
  assign _EVAL_336 = _EVAL_2224 ? _EVAL_1554 : 1'h0;
  assign _EVAL_2197 = _EVAL_1971 ? 1'h0 : _EVAL_336;
  assign _EVAL_1766 = _EVAL_714 & _EVAL_1964;
  assign _EVAL_1404 = _EVAL_1766 & _EVAL_1971;
  assign _EVAL_1997 = _EVAL_2167 == 3'h3;
  assign _EVAL_894 = _EVAL_1997 | _EVAL_2011;
  assign _EVAL_1813 = _EVAL_2167 > 3'h4;
  assign _EVAL_656 = _EVAL_894 | _EVAL_1813;
  assign _EVAL_351 = _EVAL_1545 & _EVAL_656;
  assign _EVAL_1987 = _EVAL_631[220];
  assign _EVAL_1534 = _EVAL_631[224];
  assign _EVAL_554 = _EVAL_749 & _EVAL_1534;
  assign _EVAL_59 = _EVAL_554 & _EVAL_502;
  assign _EVAL_1435 = _EVAL_59 & _EVAL_175;
  assign _EVAL_1147 = _EVAL_2167 == 3'h2;
  assign _EVAL_2079 = _EVAL_631[65];
  assign _EVAL_323 = _EVAL_749 & _EVAL_1845;
  assign _EVAL_770 = _EVAL_323 & _EVAL_502;
  assign _EVAL_2114 = _EVAL_190 == 10'h3ff;
  assign _EVAL_1890 = _EVAL_770 & _EVAL_2114;
  assign _EVAL_975 = _EVAL_36[9:0];
  assign _EVAL_589 = _EVAL_975 == 10'h0;
  assign _EVAL_527 = _EVAL_42 & _EVAL_0;
  assign _EVAL_855 = _EVAL_527 & _EVAL_19;
  assign _EVAL_1973 = _EVAL_247 & _EVAL_234;
  assign _EVAL_1958 = _EVAL_1973 & _EVAL_1971;
  assign _EVAL_562 = _EVAL_36[15:8];
  assign _EVAL_1711 = _EVAL_865 & _EVAL_1246;
  assign _EVAL_385 = _EVAL_1711 & _EVAL_1971;
  assign _EVAL_835 = _EVAL_639 | _EVAL_2116;
  assign _EVAL_598 = _EVAL_789 & _EVAL_1246;
  assign _EVAL_260 = _EVAL_1057 & _EVAL_544;
  assign _EVAL_1985 = _EVAL_598 | _EVAL_260;
  assign _EVAL_278 = _EVAL_835 | _EVAL_1985;
  assign _EVAL_487 = _EVAL_789 & _EVAL_234;
  assign _EVAL_685 = _EVAL_1057 & _EVAL_339;
  assign _EVAL_1594 = _EVAL_487 | _EVAL_685;
  assign _EVAL_1641 = _EVAL_278 | _EVAL_1594;
  assign _EVAL_1671 = _EVAL_789 & _EVAL_1964;
  assign _EVAL_60 = _EVAL_1057 & _EVAL_2190;
  assign _EVAL_1241 = _EVAL_1671 | _EVAL_60;
  assign _EVAL_688 = _EVAL_1641 | _EVAL_1241;
  assign _EVAL_1452 = _EVAL_688 | _EVAL_1662;
  assign _EVAL_1542 = _EVAL_1458 & _EVAL_1246;
  assign _EVAL_322 = _EVAL_461 & _EVAL_544;
  assign _EVAL_2075 = _EVAL_1542 | _EVAL_322;
  assign _EVAL_1485 = _EVAL_1452 | _EVAL_2075;
  assign _EVAL_1441 = _EVAL_643 == 10'h100;
  assign _EVAL_1422 = {64'h0,32'h0,_EVAL_916};
  assign _EVAL_1616 = 8'h1 << _EVAL_2167;
  assign _EVAL_817 = {{120'd0}, _EVAL_1616};
  assign _EVAL_1047 = _EVAL_59 & _EVAL_1387;
  assign _EVAL_357 = _EVAL_749 & _EVAL_469;
  assign _EVAL_291 = _EVAL_357 & _EVAL_502;
  assign _EVAL_783 = _EVAL_291 & _EVAL_758;
  assign _EVAL_1493 = _EVAL_749 & _EVAL_1486;
  assign _EVAL_2067 = _EVAL_1493 & _EVAL_502;
  assign _EVAL_1627 = _EVAL_2067 & _EVAL_175;
  assign _EVAL_240 = _EVAL_957 & _EVAL_1971;
  assign _EVAL_840 = _EVAL_1198 & _EVAL_1638;
  assign _EVAL_1210 = _EVAL_631[213];
  assign _EVAL_1969 = _EVAL_749 & _EVAL_1210;
  assign _EVAL_281 = _EVAL_1969 & _EVAL_502;
  assign _EVAL_1864 = _EVAL_281 & _EVAL_175;
  assign _EVAL_480 = _EVAL_1654 & _EVAL_1971;
  assign _EVAL_422 = 6'h16 == _EVAL_433;
  assign _EVAL_1462 = 6'h17 == _EVAL_433;
  assign _EVAL_1386 = 6'h18 == _EVAL_433;
  assign _EVAL_63 = _EVAL_1386 ? _EVAL_680 : _EVAL_127;
  assign _EVAL_1415 = _EVAL_1462 ? _EVAL_680 : _EVAL_63;
  assign _EVAL_1609 = _EVAL_422 ? _EVAL_680 : _EVAL_1415;
  assign _EVAL_162 = _EVAL_556 & _EVAL_1971;
  assign _EVAL_1511 = _EVAL_1582[19:17];
  assign _EVAL_841 = _EVAL_1511 == 3'h7;
  assign _EVAL_155 = _EVAL_979 & _EVAL_841;
  assign _EVAL_1436 = _EVAL_34[19:17];
  assign _EVAL_1082 = _EVAL_631[216];
  assign _EVAL_2157 = _EVAL_749 & _EVAL_1082;
  assign _EVAL_285 = _EVAL_2157 & _EVAL_502;
  assign _EVAL_923 = _EVAL_285 & _EVAL_1638;
  assign _EVAL_1589 = _EVAL_1824 & _EVAL_1246;
  assign _EVAL_796 = _EVAL_1589 & _EVAL_1971;
  assign _EVAL_1205 = _EVAL_36[7:0];
  assign _EVAL_513 = _EVAL_749 & _EVAL_1987;
  assign _EVAL_1984 = _EVAL_513 & _EVAL_502;
  assign _EVAL_135 = _EVAL_1984 & _EVAL_758;
  assign _EVAL_1357 = _EVAL_1798 & _EVAL_758;
  assign _EVAL_1414 = _EVAL_320 & _EVAL_1971;
  assign _EVAL_475 = _EVAL_749 & _EVAL_886;
  assign _EVAL_648 = _EVAL_475 & _EVAL_502;
  assign _EVAL_88 = _EVAL_648 & _EVAL_175;
  assign _EVAL_555 = _EVAL_838 == 2'h2;
  assign _EVAL_895 = _EVAL_1843 & _EVAL_502;
  assign _EVAL_2222 = _EVAL_895 & _EVAL_2114;
  assign _EVAL_1098 = _EVAL_898 == 1'h0;
  assign _EVAL_1920 = _EVAL_1322 & _EVAL_1098;
  assign _EVAL_1184 = _EVAL_1960 & _EVAL_962;
  assign _EVAL_1942 = _EVAL_1920 ? 1'h1 : _EVAL_1184;
  assign _EVAL_1606 = _EVAL_2102 & _EVAL_1971;
  assign _EVAL_371 = _EVAL_530 & _EVAL_1964;
  assign _EVAL_1430 = _EVAL_144 & _EVAL_2190;
  assign _EVAL_95 = _EVAL_371 | _EVAL_1430;
  assign _EVAL_722 = _EVAL_994 & _EVAL_1971;
  assign _EVAL_124 = {_EVAL_1350,_EVAL_1508,_EVAL_56,_EVAL_1469};
  assign _EVAL_1066 = _EVAL_2225 & _EVAL_2190;
  assign _EVAL_1833 = _EVAL_1766 | _EVAL_1066;
  assign _EVAL_1806 = _EVAL_656 == 1'h0;
  assign _EVAL_628 = sb2tlOpt__EVAL_7 == 1'h0;
  assign _EVAL_528 = sb2tlOpt__EVAL_25 & _EVAL_628;
  assign _EVAL_131 = _EVAL_126 & _EVAL_471;
  assign _EVAL_697 = _EVAL_131 & _EVAL_137;
  assign _EVAL_1316 = _EVAL_1984 & _EVAL_1387;
  assign _EVAL_2109 = _EVAL_865 & _EVAL_234;
  assign _EVAL_1996 = _EVAL_34[22];
  assign _EVAL_169 = _EVAL_1153 & _EVAL_1996;
  assign _EVAL_217 = _EVAL_45 == 10'h0;
  assign _EVAL_1540 = _EVAL_855 & _EVAL_217;
  assign _EVAL_744 = _EVAL_1582[31:16];
  assign _EVAL_1465 = _EVAL_1458 & _EVAL_234;
  assign _EVAL_1977 = _EVAL_461 & _EVAL_339;
  assign _EVAL_701 = _EVAL_1465 | _EVAL_1977;
  assign _EVAL_1818 = _EVAL_1485 | _EVAL_701;
  assign _EVAL_1101 = _EVAL_1458 & _EVAL_1964;
  assign _EVAL_324 = _EVAL_1101 | _EVAL_1847;
  assign _EVAL_943 = _EVAL_1818 | _EVAL_324;
  assign _EVAL_1466 = {_EVAL_1595,_EVAL_1572,_EVAL_1516,_EVAL_2000};
  assign _EVAL_352 = {_EVAL_1001,_EVAL_1402,_EVAL_277,_EVAL_75};
  assign _EVAL_1074 = {_EVAL_1716,_EVAL_2026,_EVAL_606,_EVAL_751};
  assign _EVAL_492 = {_EVAL_446,_EVAL_254,_EVAL_1991,_EVAL_1916};
  assign _EVAL_1362 = {_EVAL_1132,_EVAL_2082,_EVAL_1349,_EVAL_1250};
  assign _EVAL_1240 = {_EVAL_1499,_EVAL_1207,_EVAL_1134,_EVAL_737};
  assign _EVAL_152 = _EVAL_189 ? _EVAL_1240 : _EVAL_1419;
  assign _EVAL_123 = _EVAL_2051 ? _EVAL_1362 : _EVAL_152;
  assign _EVAL_1221 = _EVAL_1090 ? _EVAL_492 : _EVAL_123;
  assign _EVAL_1874 = _EVAL_1931 ? _EVAL_124 : _EVAL_1221;
  assign _EVAL_2073 = _EVAL_901 ? _EVAL_1074 : _EVAL_1874;
  assign _EVAL_409 = _EVAL_165 ? _EVAL_352 : _EVAL_2073;
  assign _EVAL_1740 = _EVAL_529 ? _EVAL_1466 : _EVAL_409;
  assign _EVAL_2219 = _EVAL_1966 ? _EVAL_1866 : _EVAL_1740;
  assign _EVAL_1695 = _EVAL_1119 ? _EVAL_2220 : _EVAL_2219;
  assign _EVAL_811 = _EVAL_54 == 1'h0;
  assign _EVAL_2204 = _EVAL_1065 == 1'h0;
  assign _EVAL_1125 = {_EVAL_811,1'h0,1'h0,1'h0,1'h0,_EVAL_2204,_EVAL_2204,_EVAL_1065,_EVAL_1065,8'ha2};
  assign _EVAL_899 = {1'h0,_EVAL_861,_EVAL_861,_EVAL_811,_EVAL_1125};
  assign _EVAL_2113 = _EVAL_445[0];
  assign _EVAL_1428 = _EVAL_985 & _EVAL_758;
  assign _EVAL_1822 = _EVAL_1610 & _EVAL_339;
  assign _EVAL_1902 = _EVAL_1421[24];
  assign _EVAL_1789 = _EVAL_631[210];
  assign _EVAL_1227 = _EVAL_749 & _EVAL_1789;
  assign _EVAL_1216 = _EVAL_1227 & _EVAL_502;
  assign _EVAL_2194 = _EVAL_1216 & _EVAL_175;
  assign _EVAL_2036 = _EVAL_884 & _EVAL_1971;
  assign _EVAL_1794 = _EVAL_1101 & _EVAL_1971;
  assign _EVAL_444 = _EVAL_530 & _EVAL_1246;
  assign _EVAL_1282 = _EVAL_1598 & _EVAL_1971;
  assign _EVAL_1413 = _EVAL_1932 & _EVAL_544;
  assign _EVAL_1238 = _EVAL_1589 | _EVAL_1413;
  assign _EVAL_1306 = 9'h41 == _EVAL_390;
  assign _EVAL_1790 = 9'h42 == _EVAL_390;
  assign _EVAL_458 = 9'h43 == _EVAL_390;
  assign _EVAL_122 = 9'hc0 == _EVAL_390;
  assign _EVAL_657 = _EVAL_122 ? 32'h380006f : _EVAL_1695;
  assign _EVAL_1173 = _EVAL_458 ? 32'h0 : _EVAL_657;
  assign _EVAL_2133 = _EVAL_1790 ? 32'h0 : _EVAL_1173;
  assign _EVAL_501 = _EVAL_1306 ? 32'h0 : _EVAL_2133;
  assign _EVAL_710 = _EVAL_1361 ? 1'h0 : _EVAL_1942;
  assign _EVAL_251 = _EVAL_2076 & _EVAL_1902;
  assign _EVAL_822 = _EVAL_251 & _EVAL_680;
  assign _EVAL_1807 = _EVAL_943 | _EVAL_200;
  assign _EVAL_611 = _EVAL_1308 & _EVAL_1246;
  assign _EVAL_208 = _EVAL_970 & _EVAL_544;
  assign _EVAL_808 = _EVAL_611 | _EVAL_208;
  assign _EVAL_1107 = _EVAL_1807 | _EVAL_808;
  assign _EVAL_2152 = _EVAL_1308 & _EVAL_234;
  assign _EVAL_777 = _EVAL_970 & _EVAL_339;
  assign _EVAL_782 = _EVAL_2152 | _EVAL_777;
  assign _EVAL_1021 = _EVAL_1107 | _EVAL_782;
  assign _EVAL_2230 = _EVAL_970 & _EVAL_2190;
  assign _EVAL_860 = _EVAL_256 | _EVAL_2230;
  assign _EVAL_62 = _EVAL_1021 | _EVAL_860;
  assign _EVAL_1579 = _EVAL_62 | _EVAL_442;
  assign _EVAL_2015 = _EVAL_1579 | _EVAL_1238;
  assign _EVAL_666 = _EVAL_1932 & _EVAL_339;
  assign _EVAL_347 = _EVAL_1286 | _EVAL_666;
  assign _EVAL_1690 = _EVAL_2015 | _EVAL_347;
  assign _EVAL_1022 = _EVAL_1932 & _EVAL_2190;
  assign _EVAL_1427 = _EVAL_1222 | _EVAL_1022;
  assign _EVAL_709 = _EVAL_1690 | _EVAL_1427;
  assign _EVAL_1995 = _EVAL_709 | _EVAL_1769;
  assign _EVAL_1337 = _EVAL_1872 & _EVAL_1246;
  assign _EVAL_1310 = _EVAL_94 & _EVAL_544;
  assign _EVAL_1793 = _EVAL_1337 | _EVAL_1310;
  assign _EVAL_1081 = _EVAL_1995 | _EVAL_1793;
  assign _EVAL_2218 = _EVAL_1872 & _EVAL_234;
  assign _EVAL_2020 = _EVAL_94 & _EVAL_339;
  assign _EVAL_1394 = _EVAL_2218 | _EVAL_2020;
  assign _EVAL_1069 = _EVAL_1081 | _EVAL_1394;
  assign _EVAL_1401 = _EVAL_1872 & _EVAL_1964;
  assign _EVAL_577 = _EVAL_94 & _EVAL_2190;
  assign _EVAL_1518 = _EVAL_1401 | _EVAL_577;
  assign _EVAL_856 = _EVAL_1069 | _EVAL_1518;
  assign _EVAL_306 = _EVAL_856 | _EVAL_1772;
  assign _EVAL_622 = _EVAL_2127 & _EVAL_544;
  assign _EVAL_1926 = _EVAL_1711 | _EVAL_622;
  assign _EVAL_467 = _EVAL_306 | _EVAL_1926;
  assign _EVAL_1230 = _EVAL_2127 & _EVAL_339;
  assign _EVAL_1314 = _EVAL_2109 | _EVAL_1230;
  assign _EVAL_375 = _EVAL_467 | _EVAL_1314;
  assign _EVAL_1821 = _EVAL_865 & _EVAL_1964;
  assign _EVAL_1111 = _EVAL_2127 & _EVAL_2190;
  assign _EVAL_1180 = _EVAL_1821 | _EVAL_1111;
  assign _EVAL_117 = _EVAL_375 | _EVAL_1180;
  assign _EVAL_1089 = _EVAL_117 | _EVAL_1836;
  assign _EVAL_2108 = _EVAL_1686 & _EVAL_1246;
  assign _EVAL_1271 = _EVAL_1610 & _EVAL_544;
  assign _EVAL_1648 = _EVAL_2108 | _EVAL_1271;
  assign _EVAL_2201 = _EVAL_1089 | _EVAL_1648;
  assign _EVAL_1187 = _EVAL_1145 | _EVAL_1822;
  assign _EVAL_1176 = _EVAL_2201 | _EVAL_1187;
  assign _EVAL_312 = _EVAL_1686 & _EVAL_1964;
  assign _EVAL_872 = _EVAL_1610 & _EVAL_2190;
  assign _EVAL_434 = _EVAL_312 | _EVAL_872;
  assign _EVAL_1935 = _EVAL_1176 | _EVAL_434;
  assign _EVAL_1850 = _EVAL_1935 | _EVAL_695;
  assign _EVAL_2191 = _EVAL_144 & _EVAL_544;
  assign _EVAL_143 = _EVAL_444 | _EVAL_2191;
  assign _EVAL_1034 = _EVAL_1850 | _EVAL_143;
  assign _EVAL_1906 = _EVAL_530 & _EVAL_234;
  assign _EVAL_866 = _EVAL_144 & _EVAL_339;
  assign _EVAL_1583 = _EVAL_1906 | _EVAL_866;
  assign _EVAL_1273 = _EVAL_1034 | _EVAL_1583;
  assign _EVAL_776 = _EVAL_1273 | _EVAL_95;
  assign _EVAL_1565 = _EVAL_776 | _EVAL_85;
  assign _EVAL_1049 = _EVAL_247 & _EVAL_1246;
  assign _EVAL_1425 = _EVAL_743 & _EVAL_544;
  assign _EVAL_557 = _EVAL_1049 | _EVAL_1425;
  assign _EVAL_781 = _EVAL_1565 | _EVAL_557;
  assign _EVAL_1197 = _EVAL_743 & _EVAL_339;
  assign _EVAL_2021 = _EVAL_1973 | _EVAL_1197;
  assign _EVAL_274 = _EVAL_781 | _EVAL_2021;
  assign _EVAL_1105 = _EVAL_247 & _EVAL_1964;
  assign _EVAL_503 = _EVAL_743 & _EVAL_2190;
  assign _EVAL_1479 = _EVAL_1105 | _EVAL_503;
  assign _EVAL_826 = _EVAL_274 | _EVAL_1479;
  assign _EVAL_2160 = _EVAL_826 | _EVAL_740;
  assign _EVAL_69 = _EVAL_1276 & _EVAL_544;
  assign _EVAL_1923 = _EVAL_1831 | _EVAL_69;
  assign _EVAL_1569 = _EVAL_2160 | _EVAL_1923;
  assign _EVAL_1095 = _EVAL_1276 & _EVAL_339;
  assign _EVAL_1112 = _EVAL_953 | _EVAL_1095;
  assign _EVAL_2130 = _EVAL_1569 | _EVAL_1112;
  assign _EVAL_1326 = _EVAL_665 & _EVAL_1964;
  assign _EVAL_207 = _EVAL_1276 & _EVAL_2190;
  assign _EVAL_1329 = _EVAL_1326 | _EVAL_207;
  assign _EVAL_356 = _EVAL_2130 | _EVAL_1329;
  assign _EVAL_1602 = _EVAL_356 | _EVAL_437;
  assign _EVAL_383 = _EVAL_1216 & _EVAL_1638;
  assign _EVAL_1898 = _EVAL_2054 == 1'h0;
  assign _EVAL_2200 = _EVAL_631[64];
  assign _EVAL_2041 = _EVAL_749 & _EVAL_2200;
  assign _EVAL_2071 = _EVAL_2041 & _EVAL_502;
  assign _EVAL_1976 = _EVAL_2071 & _EVAL_2114;
  assign _EVAL_1832 = _EVAL_1898 & _EVAL_1976;
  assign _EVAL_1432 = _EVAL_1832 & _EVAL_589;
  assign _EVAL_472 = _EVAL_1366 & _EVAL_1964;
  assign _EVAL_1851 = _EVAL_472 & _EVAL_1971;
  assign _EVAL_887 = _EVAL_281 & _EVAL_1387;
  assign _EVAL_868 = _EVAL_36[23:16];
  assign _EVAL_1234 = _EVAL_487 & _EVAL_1971;
  assign _EVAL_1297 = _EVAL_34[14:12];
  assign _EVAL_68 = _EVAL_1297[0];
  assign _EVAL_785 = _EVAL_2236 & _EVAL_2190;
  assign _EVAL_1495 = {{5'd0}, _EVAL_106};
  assign _EVAL_1710 = {3'h1,_EVAL_1495};
  assign _EVAL_1320 = {_EVAL_864,_EVAL_1019,_EVAL_1383,_EVAL_2097};
  assign _EVAL_98 = _EVAL_924 ? _EVAL_1320 : 32'h0;
  assign _EVAL_1295 = _EVAL_1615 ? _EVAL_916 : _EVAL_98;
  assign _EVAL_896 = _EVAL_900 ? _EVAL_1710 : _EVAL_1295;
  assign _EVAL_809 = _EVAL_420 ? _EVAL_1500 : _EVAL_896;
  assign _EVAL_1461 = _EVAL_1209 ? _EVAL_478 : _EVAL_809;
  assign _EVAL_763 = _EVAL_224 ? _EVAL_905 : _EVAL_1461;
  assign _EVAL_1052 = _EVAL_1607 ? _EVAL_1302 : _EVAL_763;
  assign _EVAL_968 = _EVAL_1299 ? _EVAL_1635 : _EVAL_1052;
  assign _EVAL_300 = _EVAL_750 ? _EVAL_1658 : _EVAL_968;
  assign _EVAL_2177 = _EVAL_153 ? _EVAL_1141 : _EVAL_300;
  assign _EVAL_1980 = _EVAL_1085 ? _EVAL_1799 : _EVAL_2177;
  assign _EVAL_600 = _EVAL_1274 ? _EVAL_545 : _EVAL_1980;
  assign _EVAL_1664 = _EVAL_205 ? _EVAL_1240 : _EVAL_600;
  assign _EVAL_1892 = _EVAL_1582[10:8];
  assign _EVAL_1571 = _EVAL_1892 == 3'h7;
  assign _EVAL_1517 = _EVAL_1582[15];
  assign _EVAL_2019 = _EVAL_34[0];
  assign _EVAL_1509 = {{11'd0}, _EVAL_2019};
  assign _EVAL_1371 = _EVAL_1984 & _EVAL_175;
  assign _EVAL_567 = _EVAL_1319 & _EVAL_175;
  assign _EVAL_115 = _EVAL_1821 & _EVAL_1971;
  assign _EVAL_245 = _EVAL_801 & _EVAL_1806;
  assign _EVAL_1377 = _EVAL_34[10:8];
  assign _EVAL_290 = _EVAL_611 & _EVAL_1971;
  assign _EVAL_118 = sb2tlOpt__EVAL_15 | sb2tlOpt__EVAL_9;
  assign _EVAL_498 = _EVAL_631[223];
  assign _EVAL_388 = _EVAL_749 & _EVAL_498;
  assign _EVAL_1037 = _EVAL_388 & _EVAL_502;
  assign _EVAL_929 = _EVAL_1037 & _EVAL_1387;
  assign _EVAL_2214 = _EVAL_1093 & _EVAL_1971;
  assign _EVAL_1219 = _EVAL_744 == 16'hffff;
  assign _EVAL_1092 = _EVAL_822 & _EVAL_1219;
  assign _EVAL_1379 = _EVAL_987 ? _EVAL_1362 : _EVAL_1664;
  assign _EVAL_1113 = _EVAL_2167 == 3'h1;
  assign _EVAL_1189 = _EVAL_1113 & _EVAL_2113;
  assign _EVAL_1487 = _EVAL_445[1:0];
  assign _EVAL_1970 = _EVAL_1487 != 2'h0;
  assign _EVAL_1603 = _EVAL_1147 & _EVAL_1970;
  assign _EVAL_377 = _EVAL_1189 | _EVAL_1603;
  assign _EVAL_738 = _EVAL_445[2:0];
  assign _EVAL_470 = _EVAL_738 != 3'h0;
  assign _EVAL_157 = _EVAL_1997 & _EVAL_470;
  assign _EVAL_906 = _EVAL_377 | _EVAL_157;
  assign _EVAL_1454 = _EVAL_906 | _EVAL_778;
  assign _EVAL_179 = _EVAL_1454 == 1'h0;
  assign _EVAL_1406 = _EVAL_2067 & _EVAL_1638;
  assign _EVAL_431 = _EVAL_1582[14:12];
  assign _EVAL_1247 = _EVAL_431 == 3'h7;
  assign _EVAL_511 = _EVAL_979 & _EVAL_1247;
  assign _EVAL_1596 = _EVAL_511 & _EVAL_68;
  assign _EVAL_1010 = _EVAL_483 & _EVAL_1971;
  assign _EVAL_1856 = _EVAL_221 & _EVAL_1971;
  assign _EVAL_194 = _EVAL_749 & _EVAL_1391;
  assign _EVAL_315 = _EVAL_194 & _EVAL_502;
  assign _EVAL_1717 = _EVAL_315 & _EVAL_1638;
  assign _EVAL_1805 = _EVAL_1465 & _EVAL_1971;
  assign _EVAL_1936 = _EVAL_281 & _EVAL_1638;
  assign _EVAL_1045 = _EVAL_598 & _EVAL_1971;
  assign _EVAL_959 = {{1'd0}, _EVAL_899};
  assign _EVAL_1862 = {1'h0,_EVAL_959};
  assign _EVAL_1185 = _EVAL_34[20];
  assign _EVAL_1639 = _EVAL_2192 & _EVAL_1971;
  assign _EVAL_1029 = _EVAL_118 & sb2tlOpt__EVAL_8;
  assign _EVAL_2038 = _EVAL_714 & _EVAL_1246;
  assign _EVAL_699 = _EVAL_2038 & _EVAL_1971;
  assign _EVAL_662 = {{31'd0}, _EVAL_1065};
  assign _EVAL_810 = _EVAL_371 & _EVAL_1971;
  assign _EVAL_65 = _EVAL_2218 & _EVAL_1971;
  assign _EVAL_2025 = _EVAL_1049 & _EVAL_1971;
  assign _EVAL_663 = _EVAL_1671 & _EVAL_1971;
  assign _EVAL_1618 = _EVAL_118 & _EVAL_1829;
  assign _EVAL_1861 = _EVAL_1422 + _EVAL_817;
  assign _EVAL_928 = _EVAL_1861[31:0];
  assign _EVAL_307 = _EVAL_319 & _EVAL_1971;
  assign _EVAL_1777 = _EVAL_749 & _EVAL_172;
  assign _EVAL_209 = _EVAL_1777 & _EVAL_502;
  assign _EVAL_2014 = _EVAL_209 & _EVAL_1638;
  assign _EVAL_1678 = _EVAL_749 & _EVAL_1760;
  assign _EVAL_877 = _EVAL_1678 & _EVAL_502;
  assign _EVAL_1622 = _EVAL_877 & _EVAL_758;
  assign _EVAL_596 = _EVAL_233 & _EVAL_1971;
  assign _EVAL_1870 = _EVAL_1582[0];
  assign _EVAL_2032 = _EVAL_979 & _EVAL_1517;
  assign _EVAL_1725 = _EVAL_527 & _EVAL_31;
  assign _EVAL_108 = _EVAL_648 & _EVAL_758;
  assign _EVAL_450 = _EVAL_1242 & _EVAL_1971;
  assign _EVAL_1612 = _EVAL_1366 & _EVAL_234;
  assign _EVAL_1990 = _EVAL_1612 & _EVAL_1971;
  assign _EVAL_533 = sb2tlOpt__EVAL_6 == 1'h0;
  assign _EVAL_981 = _EVAL_209 & _EVAL_758;
  assign _EVAL_1520 = 6'h0 == _EVAL_433;
  assign _EVAL_399 = 6'h4 == _EVAL_433;
  assign _EVAL_907 = 6'h11 == _EVAL_433;
  assign _EVAL_1474 = 6'h12 == _EVAL_433;
  assign _EVAL_1808 = 6'h13 == _EVAL_433;
  assign _EVAL_1324 = _EVAL_1808 ? _EVAL_680 : _EVAL_1609;
  assign _EVAL_363 = _EVAL_1474 ? _EVAL_680 : _EVAL_1324;
  assign _EVAL_1685 = _EVAL_907 ? _EVAL_680 : _EVAL_363;
  assign _EVAL_1631 = _EVAL_399 ? _EVAL_680 : _EVAL_1685;
  assign _EVAL_613 = _EVAL_1520 ? _EVAL_311 : _EVAL_1631;
  assign _EVAL_635 = _EVAL_1551 & _EVAL_1971;
  assign _EVAL_1478 = _EVAL_1737 ? _EVAL_492 : _EVAL_1379;
  assign _EVAL_935 = _EVAL_555 ? _EVAL_2222 : 1'h0;
  assign _EVAL_1560 = _EVAL_2224 ? 1'h0 : _EVAL_935;
  assign _EVAL_786 = _EVAL_315 & _EVAL_758;
  assign _EVAL_386 = _EVAL_444 & _EVAL_1971;
  assign _EVAL_1642 = ~ _EVAL_1971;
  assign _EVAL_1194 = _EVAL_164 & _EVAL_1642;
  assign _EVAL_1541 = _EVAL_59 & _EVAL_758;
  assign _EVAL_1749 = _EVAL_1838 & _EVAL_1971;
  assign _EVAL_670 = _EVAL_315 & _EVAL_175;
  assign _EVAL_500 = _EVAL_614 & _EVAL_1971;
  assign _EVAL_706 = _EVAL_2225 & _EVAL_544;
  assign _EVAL_1747 = _EVAL_2038 | _EVAL_706;
  assign _EVAL_1633 = _EVAL_1602 | _EVAL_1747;
  assign _EVAL_1191 = _EVAL_2225 & _EVAL_339;
  assign _EVAL_232 = _EVAL_1093 | _EVAL_1191;
  assign _EVAL_1199 = _EVAL_1633 | _EVAL_232;
  assign _EVAL_1344 = _EVAL_1199 | _EVAL_1833;
  assign _EVAL_298 = _EVAL_1344 & _EVAL_1642;
  assign _EVAL_225 = _EVAL_1509 & 12'h1;
  assign _EVAL_1269 = _EVAL_1545 & _EVAL_1454;
  assign _EVAL_1460 = _EVAL_1198 & _EVAL_758;
  assign _EVAL_1877 = _EVAL_1535 & _EVAL_1971;
  assign _EVAL_1940 = _EVAL_1608 & _EVAL_1971;
  assign _EVAL_712 = _EVAL_877 & _EVAL_175;
  assign _EVAL_464 = _EVAL_749 & _EVAL_2079;
  assign _EVAL_2212 = _EVAL_464 & _EVAL_502;
  assign _EVAL_1307 = _EVAL_2224 ? _EVAL_962 : 1'h0;
  assign _EVAL_1056 = {1'h0,_EVAL_1854};
  assign _EVAL_79 = {{14'd0}, _EVAL_1056};
  assign _EVAL_625 = {_EVAL_1137,_EVAL_79};
  assign _EVAL_1776 = _EVAL_721 ? _EVAL_124 : _EVAL_1478;
  assign _EVAL_459 = _EVAL_109 ? _EVAL_1074 : _EVAL_1776;
  assign _EVAL_1911 = _EVAL_518 ? _EVAL_352 : _EVAL_459;
  assign _EVAL_1795 = _EVAL_1691 ? _EVAL_1466 : _EVAL_1911;
  assign _EVAL_66 = _EVAL_1386 ? _EVAL_625 : _EVAL_1795;
  assign _EVAL_393 = _EVAL_1462 ? _EVAL_726 : _EVAL_66;
  assign _EVAL_482 = _EVAL_34[31:16];
  assign _EVAL_718 = _EVAL_1216 & _EVAL_758;
  assign _EVAL_848 = _EVAL_1296 & _EVAL_1971;
  assign _EVAL_845 = _EVAL_1773 & _EVAL_1971;
  assign _EVAL_521 = _EVAL_209 & _EVAL_175;
  assign _EVAL_151 = _EVAL_1326 & _EVAL_1971;
  assign _EVAL_941 = _EVAL_593 & _EVAL_2204;
  assign _EVAL_454 = _EVAL_30 | _EVAL_941;
  assign _EVAL_1547 = _EVAL_634 & _EVAL_454;
  assign _EVAL_1873 = _EVAL_328 & _EVAL_1571;
  assign _EVAL_1471 = _EVAL_1873 & _EVAL_1642;
  assign _EVAL_404 = _EVAL_822 & _EVAL_1870;
  assign _EVAL_515 = _EVAL_404 & _EVAL_1642;
  assign _EVAL_2199 = _EVAL_1471 | _EVAL_515;
  assign _EVAL_77 = _EVAL_404 & _EVAL_1971;
  assign _EVAL_192 = _EVAL_1244 | _EVAL_1160;
  assign _EVAL_1918 = _EVAL_2236 & _EVAL_339;
  assign _EVAL_1564 = _EVAL_1612 | _EVAL_1918;
  assign _EVAL_1536 = _EVAL_192 | _EVAL_1564;
  assign _EVAL_523 = _EVAL_472 | _EVAL_785;
  assign _EVAL_210 = _EVAL_1536 | _EVAL_523;
  assign _EVAL_2096 = _EVAL_210 & _EVAL_1642;
  assign _EVAL_933 = _EVAL_452 & _EVAL_1638;
  assign _EVAL_1917 = _EVAL_1337 & _EVAL_1971;
  assign _EVAL_1754 = ~ _EVAL_1377;
  assign _EVAL_1482 = _EVAL_1263 & _EVAL_1754;
  assign _EVAL_925 = _EVAL_1297[1];
  assign _EVAL_1656 = _EVAL_838 != 2'h0;
  assign _EVAL_1731 = {1'h0,_EVAL_1656,1'h0,_EVAL_1263,8'h1};
  assign _EVAL_1006 = {{10'd0}, _EVAL_1731};
  assign _EVAL_2229 = _EVAL_34[16];
  assign _EVAL_80 = _EVAL_1798 & _EVAL_1638;
  assign _EVAL_588 = _EVAL_1582[16];
  assign _EVAL_969 = _EVAL_979 & _EVAL_588;
  assign _EVAL_1294 = _EVAL_1163 & _EVAL_1971;
  assign _EVAL_1012 = _EVAL_1092 & _EVAL_1642;
  assign _EVAL_908 = _EVAL_2199 | _EVAL_1012;
  assign _EVAL_522 = _EVAL_908 | _EVAL_1194;
  assign _EVAL_359 = _EVAL_522 | _EVAL_2096;
  assign _EVAL_1108 = _EVAL_359 | _EVAL_298;
  assign _EVAL_463 = _EVAL_1971 ? 1'h0 : _EVAL_1560;
  assign _EVAL_1952 = _EVAL_1971 ? _EVAL_710 : _EVAL_1307;
  assign _EVAL_955 = _EVAL_1873 & _EVAL_1971;
  assign _EVAL_2134 = _EVAL_1798 & _EVAL_175;
  assign _EVAL_1697 = _EVAL_312 & _EVAL_1971;
  assign _EVAL_875 = _EVAL_2212 & _EVAL_2114;
  assign _EVAL_2226 = _EVAL_1906 & _EVAL_1971;
  assign _EVAL_2001 = 9'h40 == _EVAL_390;
  assign _EVAL_1751 = _EVAL_122 ? _EVAL_502 : _EVAL_2101;
  assign _EVAL_2216 = _EVAL_458 ? _EVAL_502 : _EVAL_1751;
  assign _EVAL_591 = _EVAL_1790 ? _EVAL_502 : _EVAL_2216;
  assign _EVAL_1275 = _EVAL_1306 ? _EVAL_502 : _EVAL_591;
  assign _EVAL_391 = _EVAL_2001 ? _EVAL_502 : _EVAL_1275;
  assign _EVAL_2170 = _EVAL_985 & _EVAL_1638;
  assign _EVAL_313 = _EVAL_669 & _EVAL_1971;
  assign _EVAL_805 = _EVAL_285 & _EVAL_175;
  assign _EVAL_1218 = _EVAL_648 & _EVAL_1638;
  assign _EVAL_253 = _EVAL_1092 & _EVAL_1971;
  assign _EVAL_82 = _EVAL_1297[2];
  assign _EVAL_843 = _EVAL_511 & _EVAL_82;
  assign _EVAL_1339 = sb2tlOpt__EVAL_11 & _EVAL_533;
  assign _EVAL_1456 = _EVAL_1339 | _EVAL_528;
  assign _EVAL_1688 = _EVAL_452 & _EVAL_758;
  assign _EVAL_1403 = _EVAL_1725 & _EVAL_217;
  assign _EVAL_990 = _EVAL_1171 & _EVAL_1971;
  assign _EVAL_1313 = _EVAL_662 != 32'h0;
  assign _EVAL_373 = {{31'd0}, _EVAL_1313};
  assign _EVAL_1533 = {5'h10,_EVAL_1006};
  assign _EVAL_1881 = _EVAL_422 ? {{3'd0}, _EVAL_1533} : _EVAL_393;
  assign _EVAL_636 = _EVAL_1808 ? _EVAL_373 : _EVAL_1881;
  assign _EVAL_100 = _EVAL_1474 ? 32'h111380 : _EVAL_636;
  assign _EVAL_156 = {_EVAL_51,_EVAL_12};
  assign _EVAL_1115 = _EVAL_1037 & _EVAL_175;
  assign _EVAL_1158 = _EVAL_281 & _EVAL_758;
  assign _EVAL_279 = _EVAL_59 & _EVAL_1638;
  assign _EVAL_331 = _EVAL_1965[23:0];
  assign _EVAL_2048 = _EVAL_2067 & _EVAL_1387;
  assign _EVAL_457 = {64'h0,32'h0,_EVAL_864,_EVAL_1019,_EVAL_1383,_EVAL_2097};
  assign _EVAL_632 = _EVAL_907 ? {{9'd0}, _EVAL_1862} : _EVAL_100;
  assign _EVAL_1826 = _EVAL_1105 & _EVAL_1971;
  assign _EVAL_1912 = _EVAL_2108 & _EVAL_1971;
  assign _EVAL_703 = ~ _EVAL_11;
  assign _EVAL_1353 = _EVAL_285 & _EVAL_1387;
  assign _EVAL_103 = _EVAL_285 & _EVAL_758;
  assign _EVAL_1060 = _EVAL_1592 & _EVAL_1971;
  assign _EVAL_814 = _EVAL_1752 & _EVAL_1971;
  assign _EVAL_784 = _EVAL_985 & _EVAL_1387;
  assign _EVAL_671 = _EVAL_877 & _EVAL_1387;
  assign _EVAL_52 = _EVAL_920 ? 1'h0 : 1'h1;
  assign _EVAL_1523 = _EVAL_962 ? 1'h0 : _EVAL_52;
  assign _EVAL_1183 = _EVAL_2224 ? _EVAL_1523 : 1'h0;
  assign _EVAL_1787 = _EVAL_1971 ? 1'h0 : _EVAL_1183;
  assign _EVAL_149 = _EVAL_1319 & _EVAL_1387;
  assign _EVAL_543 = _EVAL_209 & _EVAL_1387;
  assign _EVAL_2034 = _EVAL_1037 & _EVAL_1638;
  assign _EVAL_2047 = _EVAL_1542 & _EVAL_1971;
  assign _EVAL_211 = _EVAL_1401 & _EVAL_1971;
  assign _EVAL_185 = 9'h0 == _EVAL_390;
  assign _EVAL_2138 = _EVAL_728 & _EVAL_1971;
  assign _EVAL_1797 = _EVAL_291 & _EVAL_175;
  assign _EVAL_2144 = _EVAL_1216 & _EVAL_1387;
  assign _EVAL_2166 = _EVAL_2109 & _EVAL_1971;
  assign _EVAL_1433 = _EVAL_2067 & _EVAL_758;
  assign _EVAL_1762 = _EVAL_34[15];
  assign _EVAL_1653 = {64'h0,32'h0,_EVAL_34};
  assign _EVAL_1279 = _EVAL_1301 & _EVAL_1815;
  assign _EVAL_1665 = _EVAL_399 ? _EVAL_2234 : _EVAL_632;
  assign _EVAL_705 = _EVAL_1520 ? _EVAL_662 : _EVAL_1665;
  assign _EVAL_112 = _EVAL_877 & _EVAL_1638;
  assign _EVAL_1522 = _EVAL_1198 & _EVAL_1387;
  assign _EVAL_1215 = _EVAL_2152 & _EVAL_1971;
  assign _EVAL_362 = _EVAL_291 & _EVAL_1638;
  assign _EVAL_724 = _EVAL_1750 & _EVAL_1971;
  assign _EVAL_1863 = {8'h0,6'h0,_EVAL_54,_EVAL_2054};
  assign _EVAL_912 = _EVAL_1984 & _EVAL_1638;
  assign _EVAL_867 = {_EVAL_4,_EVAL_6};
  assign _EVAL_761 = _EVAL_559 & _EVAL_1971;
  assign _EVAL_1938 = _EVAL_979 & _EVAL_1709;
  assign _EVAL_2228 = _EVAL_511 & _EVAL_925;
  assign _EVAL_678 = _EVAL_648 & _EVAL_1387;
  assign _EVAL_690 = _EVAL_1279 & _EVAL_1806;
  assign _EVAL_74 = _EVAL_1532 & _EVAL_1971;
  assign _EVAL_318 = _EVAL_2001 ? 32'h0 : _EVAL_501;
  assign _EVAL_1196 = _EVAL_185 ? _EVAL_1441 : _EVAL_391;
  assign _EVAL_1643 = _EVAL_291 & _EVAL_1387;
  assign _EVAL_1232 = _EVAL_1889 & _EVAL_1971;
  assign _EVAL_2139 = _EVAL_1319 & _EVAL_758;
  assign _EVAL_694 = _EVAL_452 & _EVAL_175;
  assign _EVAL_1939 = _EVAL_315 & _EVAL_1387;
  assign _EVAL_449 = _EVAL_1037 & _EVAL_758;
  assign _EVAL_1439 = _EVAL_185 ? {{16'd0}, _EVAL_1863} : _EVAL_318;
  assign _EVAL_38 = _EVAL_613 ? _EVAL_705 : 32'h0;
  assign _EVAL_26 = _EVAL_13;
  assign _EVAL_17 = sb2tlOpt__EVAL_13;
  assign _EVAL_42 = 1'h1;
  assign _EVAL_47 = _EVAL_48;
  assign _EVAL_33 = sb2tlOpt__EVAL_26;
  assign sb2tlOpt__EVAL_5 = _EVAL_2167;
  assign _EVAL_29 = sb2tlOpt__EVAL_27;
  assign _EVAL_8 = _EVAL_156[1:0];
  assign sb2tlOpt__EVAL_17 = _EVAL_11;
  assign sb2tlOpt__EVAL_20 = _EVAL_30;
  assign sb2tlOpt__EVAL_4 = _EVAL_5;
  assign sb2tlOpt__EVAL_11 = _EVAL_245 & _EVAL_179;
  assign _EVAL_35 = {{2'd0}, _EVAL_681};
  assign _EVAL_46 = _EVAL_1196 ? _EVAL_1439 : 32'h0;
  assign sb2tlOpt__EVAL_16 = _EVAL_39;
  assign sb2tlOpt__EVAL_18 = _EVAL;
  assign sb2tlOpt__EVAL = _EVAL_50;
  assign _EVAL_44 = {{2'd0}, _EVAL_644};
  assign sb2tlOpt__EVAL_1 = _EVAL_7;
  assign _EVAL_22 = sb2tlOpt__EVAL_23;
  assign _EVAL_40 = _EVAL_28;
  assign sb2tlOpt__EVAL_24 = _EVAL_27;
  assign sb2tlOpt__EVAL_28 = sb2tlOpt__EVAL_25 ? _EVAL_2029 : _EVAL_1422;
  assign _EVAL_37 = sb2tlOpt__EVAL_2;
  assign _EVAL_49 = _EVAL_593;
  assign _EVAL_20 = _EVAL_867[1:0];
  assign sb2tlOpt__EVAL_21 = sb2tlOpt__EVAL_11 ? _EVAL_1653 : _EVAL_457;
  assign sb2tlOpt__EVAL_25 = _EVAL_690 & _EVAL_179;
  assign _EVAL_16 = _EVAL_156[13:2];
  assign _EVAL_25 = _EVAL_867[2];
  assign _EVAL_10 = sb2tlOpt__EVAL_10;
  assign _EVAL_24 = _EVAL_18;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_54 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_56 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_72 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_75 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_92 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_130 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_174 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_182 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_212 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_229 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_254 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_277 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_284 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_329 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_438 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_446 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_532 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_593 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_606 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_616 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_623 = _RAND_20[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_634 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_658 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_732 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_734 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_737 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_739 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_751 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_804 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_838 = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_846 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_858 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_861 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_864 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_881 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_915 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_916 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_961 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_1001 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_1019 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_1040 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_1055 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_1065 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_1100 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_1132 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_1134 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_1135 = _RAND_46[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_1137 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_1154 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_1200 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1207 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1250 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1263 = _RAND_52[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1264 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1349 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1350 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1370 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1383 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1402 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1447 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1469 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1499 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1508 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1516 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1562 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1572 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1595 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1599 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1646 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1649 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1652 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1694 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1716 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1768 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1785 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1803 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1829 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1859 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1866 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1869 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1916 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1943 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1951 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1991 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_2000 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_2026 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_2054 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_2057 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_2058 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_2082 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_2097 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_2117 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_2154 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_2165 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_2167 = _RAND_94[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_2220 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_703) begin
      _EVAL_54 <= 1'h0;
    end else begin
      if (_EVAL_1403) begin
        _EVAL_54 <= 1'h1;
      end else begin
        if (_EVAL_1890) begin
          if (_EVAL_589) begin
            _EVAL_54 <= 1'h0;
          end else begin
            if (_EVAL_30) begin
              _EVAL_54 <= 1'h0;
            end
          end
        end else begin
          if (_EVAL_30) begin
            _EVAL_54 <= 1'h0;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_56 <= 8'h0;
    end else begin
      if (_EVAL_2170) begin
        _EVAL_56 <= _EVAL_562;
      end else begin
        if (_EVAL_761) begin
          if (_EVAL_559) begin
            _EVAL_56 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_72 <= 8'h0;
    end else begin
      if (_EVAL_112) begin
        _EVAL_72 <= _EVAL_562;
      end else begin
        if (_EVAL_2025) begin
          if (_EVAL_1049) begin
            _EVAL_72 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_75 <= 8'h0;
    end else begin
      if (_EVAL_786) begin
        _EVAL_75 <= _EVAL_1205;
      end else begin
        if (_EVAL_74) begin
          if (_EVAL_1532) begin
            _EVAL_75 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_92 <= 8'h0;
    end else begin
      if (_EVAL_1688) begin
        _EVAL_92 <= _EVAL_1205;
      end else begin
        if (_EVAL_845) begin
          if (_EVAL_1773) begin
            _EVAL_92 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_130 <= 8'h0;
    end else begin
      if (_EVAL_1460) begin
        _EVAL_130 <= _EVAL_1205;
      end else begin
        if (_EVAL_1877) begin
          if (_EVAL_1535) begin
            _EVAL_130 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_174 <= 8'h0;
    end else begin
      if (_EVAL_543) begin
        _EVAL_174 <= _EVAL_868;
      end else begin
        if (_EVAL_2146) begin
          if (_EVAL_953) begin
            _EVAL_174 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_182 <= 8'h0;
    end else begin
      if (_EVAL_1622) begin
        _EVAL_182 <= _EVAL_1205;
      end else begin
        if (_EVAL_307) begin
          if (_EVAL_319) begin
            _EVAL_182 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_212 <= 1'h0;
    end else begin
      if (_EVAL_2228) begin
        _EVAL_212 <= 1'h0;
      end else begin
        if (_EVAL_1456) begin
          _EVAL_212 <= 1'h1;
        end else begin
          if (_EVAL_1269) begin
            _EVAL_212 <= 1'h1;
          end else begin
            if (_EVAL_351) begin
              _EVAL_212 <= 1'h0;
            end else begin
              if (_EVAL_1029) begin
                _EVAL_212 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_229 <= 8'h0;
    end else begin
      if (_EVAL_1353) begin
        _EVAL_229 <= _EVAL_868;
      end else begin
        if (_EVAL_410) begin
          if (_EVAL_1286) begin
            _EVAL_229 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_254 <= 8'h0;
    end else begin
      if (_EVAL_678) begin
        _EVAL_254 <= _EVAL_868;
      end else begin
        if (_EVAL_1856) begin
          if (_EVAL_221) begin
            _EVAL_254 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_277 <= 8'h0;
    end else begin
      if (_EVAL_1717) begin
        _EVAL_277 <= _EVAL_562;
      end else begin
        if (_EVAL_635) begin
          if (_EVAL_1551) begin
            _EVAL_277 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_284 <= 1'h0;
    end else begin
      if (_EVAL_843) begin
        _EVAL_284 <= 1'h0;
      end else begin
        if (_EVAL_1456) begin
          _EVAL_284 <= 1'h0;
        end else begin
          if (_EVAL_1269) begin
            _EVAL_284 <= 1'h0;
          end else begin
            if (_EVAL_351) begin
              _EVAL_284 <= 1'h1;
            end else begin
              if (_EVAL_1029) begin
                _EVAL_284 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_329 <= 8'h0;
    end else begin
      if (_EVAL_981) begin
        _EVAL_329 <= _EVAL_1205;
      end else begin
        if (_EVAL_2138) begin
          if (_EVAL_728) begin
            _EVAL_329 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_438 <= 8'h0;
    end else begin
      if (_EVAL_449) begin
        _EVAL_438 <= _EVAL_1205;
      end else begin
        if (_EVAL_1232) begin
          if (_EVAL_1889) begin
            _EVAL_438 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_446 <= 8'h0;
    end else begin
      if (_EVAL_88) begin
        _EVAL_446 <= _EVAL_1755;
      end else begin
        if (_EVAL_240) begin
          if (_EVAL_957) begin
            _EVAL_446 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_532 <= 8'h0;
    end else begin
      if (_EVAL_279) begin
        _EVAL_532 <= _EVAL_562;
      end else begin
        if (_EVAL_1940) begin
          if (_EVAL_1608) begin
            _EVAL_532 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_593 <= 1'h0;
    end else begin
      _EVAL_593 <= _EVAL_1547;
    end
    if (_EVAL_703) begin
      _EVAL_606 <= 8'h0;
    end else begin
      if (_EVAL_383) begin
        _EVAL_606 <= _EVAL_562;
      end else begin
        if (_EVAL_722) begin
          if (_EVAL_994) begin
            _EVAL_606 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_616 <= _EVAL_729;
    end
    if (_EVAL_703) begin
      _EVAL_623 <= 24'h0;
    end else begin
      if (_EVAL_1322) begin
        _EVAL_623 <= _EVAL_331;
      end
    end
    if (_EVAL_703) begin
      _EVAL_634 <= 1'h0;
    end else begin
      if (_EVAL_527) begin
        _EVAL_634 <= _EVAL_43;
      end
    end
    if (_EVAL_703) begin
      _EVAL_658 <= 8'h0;
    end else begin
      if (_EVAL_1988) begin
        _EVAL_658 <= _EVAL_868;
      end else begin
        if (_EVAL_65) begin
          if (_EVAL_2218) begin
            _EVAL_658 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_732 <= 8'h0;
    end else begin
      if (_EVAL_712) begin
        _EVAL_732 <= _EVAL_1755;
      end else begin
        if (_EVAL_1826) begin
          if (_EVAL_1105) begin
            _EVAL_732 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_734 <= 1'h0;
    end else begin
      if (_EVAL_169) begin
        _EVAL_734 <= 1'h0;
      end else begin
        if (_EVAL_305) begin
          _EVAL_734 <= 1'h1;
        end else begin
          if (_EVAL_1780) begin
            _EVAL_734 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_737 <= 8'h0;
    end else begin
      if (_EVAL_783) begin
        _EVAL_737 <= _EVAL_1205;
      end else begin
        if (_EVAL_1639) begin
          if (_EVAL_2192) begin
            _EVAL_737 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_739 <= 8'h0;
    end else begin
      if (_EVAL_933) begin
        _EVAL_739 <= _EVAL_562;
      end else begin
        if (_EVAL_1917) begin
          if (_EVAL_1337) begin
            _EVAL_739 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_751 <= 8'h0;
    end else begin
      if (_EVAL_718) begin
        _EVAL_751 <= _EVAL_1205;
      end else begin
        if (_EVAL_848) begin
          if (_EVAL_1296) begin
            _EVAL_751 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_804 <= 8'h0;
    end else begin
      if (_EVAL_1435) begin
        _EVAL_804 <= _EVAL_1755;
      end else begin
        if (_EVAL_1851) begin
          if (_EVAL_472) begin
            _EVAL_804 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_838 <= 2'h0;
    end else begin
      if (_EVAL_1971) begin
        if (_EVAL_1361) begin
          _EVAL_838 <= 2'h1;
        end
      end else begin
        if (_EVAL_2224) begin
          if (_EVAL_962) begin
            _EVAL_838 <= 2'h0;
          end else begin
            if (_EVAL_920) begin
              _EVAL_838 <= 2'h0;
            end else begin
              _EVAL_838 <= 2'h2;
            end
          end
        end else begin
          if (_EVAL_555) begin
            if (_EVAL_2222) begin
              _EVAL_838 <= 2'h0;
            end else begin
              if (_EVAL_1432) begin
                _EVAL_838 <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_846 <= 8'h0;
    end else begin
      if (_EVAL_1541) begin
        _EVAL_846 <= _EVAL_1205;
      end else begin
        if (_EVAL_1749) begin
          if (_EVAL_1838) begin
            _EVAL_846 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_858 <= 8'h0;
    end else begin
      if (_EVAL_923) begin
        _EVAL_858 <= _EVAL_562;
      end else begin
        if (_EVAL_796) begin
          if (_EVAL_1589) begin
            _EVAL_858 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_861 <= 1'h0;
    end else begin
      if (_EVAL_30) begin
        _EVAL_861 <= 1'h1;
      end else begin
        if (_EVAL_1540) begin
          _EVAL_861 <= 1'h0;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_864 <= 8'h0;
    end else begin
      if (_EVAL_801) begin
        _EVAL_864 <= _EVAL_142;
      end else begin
        if (sb2tlOpt__EVAL_22) begin
          _EVAL_864 <= sb2tlOpt__EVAL_19;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_881 <= 8'h0;
    end else begin
      if (_EVAL_1047) begin
        _EVAL_881 <= _EVAL_868;
      end else begin
        if (_EVAL_1990) begin
          if (_EVAL_1612) begin
            _EVAL_881 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_915 <= 8'h0;
    end else begin
      if (_EVAL_1371) begin
        _EVAL_915 <= _EVAL_1755;
      end else begin
        if (_EVAL_810) begin
          if (_EVAL_371) begin
            _EVAL_915 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_916 <= 32'h0;
    end else begin
      if (_EVAL_697) begin
        _EVAL_916 <= _EVAL_34;
      end else begin
        if (_EVAL_1618) begin
          _EVAL_916 <= _EVAL_928;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_961 <= 8'h0;
    end else begin
      if (_EVAL_80) begin
        _EVAL_961 <= _EVAL_562;
      end else begin
        if (_EVAL_1912) begin
          if (_EVAL_2108) begin
            _EVAL_961 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1001 <= 8'h0;
    end else begin
      if (_EVAL_670) begin
        _EVAL_1001 <= _EVAL_1755;
      end else begin
        if (_EVAL_1858) begin
          if (_EVAL_139) begin
            _EVAL_1001 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1019 <= 8'h0;
    end else begin
      if (_EVAL_801) begin
        _EVAL_1019 <= _EVAL_55;
      end else begin
        if (sb2tlOpt__EVAL_0) begin
          _EVAL_1019 <= sb2tlOpt__EVAL_19;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1040 <= 8'h0;
    end else begin
      if (_EVAL_1115) begin
        _EVAL_1040 <= _EVAL_1755;
      end else begin
        if (_EVAL_1404) begin
          if (_EVAL_1766) begin
            _EVAL_1040 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1055 <= 8'h0;
    end else begin
      if (_EVAL_1522) begin
        _EVAL_1055 <= _EVAL_868;
      end else begin
        if (_EVAL_1215) begin
          if (_EVAL_2152) begin
            _EVAL_1055 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1065 <= 1'h0;
    end else begin
      if (_EVAL_30) begin
        _EVAL_1065 <= 1'h0;
      end else begin
        if (_EVAL_1976) begin
          if (_EVAL_589) begin
            _EVAL_1065 <= 1'h1;
          end
        end else begin
          if (_EVAL_1890) begin
            if (_EVAL_589) begin
              _EVAL_1065 <= 1'h0;
            end
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1100 <= 8'h0;
    end else begin
      if (_EVAL_521) begin
        _EVAL_1100 <= _EVAL_1755;
      end else begin
        if (_EVAL_151) begin
          if (_EVAL_1326) begin
            _EVAL_1100 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1132 <= 8'h0;
    end else begin
      if (_EVAL_1864) begin
        _EVAL_1132 <= _EVAL_1755;
      end else begin
        if (_EVAL_663) begin
          if (_EVAL_1671) begin
            _EVAL_1132 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1134 <= 8'h0;
    end else begin
      if (_EVAL_362) begin
        _EVAL_1134 <= _EVAL_562;
      end else begin
        if (_EVAL_2047) begin
          if (_EVAL_1542) begin
            _EVAL_1134 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1135 <= 12'h0;
    end else begin
      if (_EVAL_77) begin
        _EVAL_1135 <= _EVAL_225;
      end
    end
    if (_EVAL_703) begin
      _EVAL_1137 <= 16'h0;
    end else begin
      if (_EVAL_253) begin
        _EVAL_1137 <= _EVAL_482;
      end
    end
    if (_EVAL_703) begin
      _EVAL_1154 <= 8'h0;
    end else begin
      if (_EVAL_1322) begin
        _EVAL_1154 <= _EVAL_1925;
      end
    end
    if (_EVAL_703) begin
      _EVAL_1200 <= 8'h0;
    end else begin
      if (_EVAL_986) begin
        _EVAL_1200 <= _EVAL_868;
      end else begin
        if (_EVAL_1459) begin
          if (_EVAL_1145) begin
            _EVAL_1200 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1207 <= 8'h0;
    end else begin
      if (_EVAL_1643) begin
        _EVAL_1207 <= _EVAL_868;
      end else begin
        if (_EVAL_1805) begin
          if (_EVAL_1465) begin
            _EVAL_1207 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1250 <= 8'h0;
    end else begin
      if (_EVAL_1158) begin
        _EVAL_1250 <= _EVAL_1205;
      end else begin
        if (_EVAL_1060) begin
          if (_EVAL_1592) begin
            _EVAL_1250 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1263 <= 3'h0;
    end else begin
      if (_EVAL_1108) begin
        _EVAL_1263 <= 3'h1;
      end else begin
        if (_EVAL_463) begin
          _EVAL_1263 <= 3'h3;
        end else begin
          if (_EVAL_1952) begin
            _EVAL_1263 <= 3'h2;
          end else begin
            if (_EVAL_2197) begin
              _EVAL_1263 <= 3'h4;
            end else begin
              if (_EVAL_955) begin
                _EVAL_1263 <= _EVAL_1482;
              end
            end
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1264 <= 8'h0;
    end else begin
      if (_EVAL_840) begin
        _EVAL_1264 <= _EVAL_562;
      end else begin
        if (_EVAL_290) begin
          if (_EVAL_611) begin
            _EVAL_1264 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1349 <= 8'h0;
    end else begin
      if (_EVAL_1936) begin
        _EVAL_1349 <= _EVAL_562;
      end else begin
        if (_EVAL_1045) begin
          if (_EVAL_598) begin
            _EVAL_1349 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1350 <= 8'h0;
    end else begin
      if (_EVAL_1959) begin
        _EVAL_1350 <= _EVAL_1755;
      end else begin
        if (_EVAL_313) begin
          if (_EVAL_669) begin
            _EVAL_1350 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1370 <= 8'h0;
    end else begin
      if (_EVAL_694) begin
        _EVAL_1370 <= _EVAL_1755;
      end else begin
        if (_EVAL_211) begin
          if (_EVAL_1401) begin
            _EVAL_1370 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1383 <= 8'h0;
    end else begin
      if (_EVAL_801) begin
        _EVAL_1383 <= _EVAL_2060;
      end else begin
        if (sb2tlOpt__EVAL_3) begin
          _EVAL_1383 <= sb2tlOpt__EVAL_19;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1402 <= 8'h0;
    end else begin
      if (_EVAL_1939) begin
        _EVAL_1402 <= _EVAL_868;
      end else begin
        if (_EVAL_1294) begin
          if (_EVAL_1163) begin
            _EVAL_1402 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1447 <= 8'h0;
    end else begin
      if (_EVAL_1357) begin
        _EVAL_1447 <= _EVAL_1205;
      end else begin
        if (_EVAL_1414) begin
          if (_EVAL_320) begin
            _EVAL_1447 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1469 <= 8'h0;
    end else begin
      if (_EVAL_1428) begin
        _EVAL_1469 <= _EVAL_1205;
      end else begin
        if (_EVAL_1010) begin
          if (_EVAL_483) begin
            _EVAL_1469 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1499 <= 8'h0;
    end else begin
      if (_EVAL_1797) begin
        _EVAL_1499 <= _EVAL_1755;
      end else begin
        if (_EVAL_1794) begin
          if (_EVAL_1101) begin
            _EVAL_1499 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1508 <= 8'h0;
    end else begin
      if (_EVAL_784) begin
        _EVAL_1508 <= _EVAL_868;
      end else begin
        if (_EVAL_814) begin
          if (_EVAL_1752) begin
            _EVAL_1508 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1516 <= 8'h0;
    end else begin
      if (_EVAL_1406) begin
        _EVAL_1516 <= _EVAL_562;
      end else begin
        if (_EVAL_480) begin
          if (_EVAL_1654) begin
            _EVAL_1516 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1562 <= 8'h0;
    end else begin
      if (_EVAL_2034) begin
        _EVAL_1562 <= _EVAL_562;
      end else begin
        if (_EVAL_699) begin
          if (_EVAL_2038) begin
            _EVAL_1562 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1572 <= 8'h0;
    end else begin
      if (_EVAL_2048) begin
        _EVAL_1572 <= _EVAL_868;
      end else begin
        if (_EVAL_1606) begin
          if (_EVAL_2102) begin
            _EVAL_1572 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1595 <= 8'h0;
    end else begin
      if (_EVAL_1627) begin
        _EVAL_1595 <= _EVAL_1755;
      end else begin
        if (_EVAL_596) begin
          if (_EVAL_233) begin
            _EVAL_1595 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1599 <= 8'h0;
    end else begin
      if (_EVAL_857) begin
        _EVAL_1599 <= _EVAL_562;
      end else begin
        if (_EVAL_385) begin
          if (_EVAL_1711) begin
            _EVAL_1599 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1646 <= 8'h0;
    end else begin
      if (_EVAL_1316) begin
        _EVAL_1646 <= _EVAL_868;
      end else begin
        if (_EVAL_2226) begin
          if (_EVAL_1906) begin
            _EVAL_1646 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1649 <= 8'h0;
    end else begin
      if (_EVAL_1703) begin
        _EVAL_1649 <= _EVAL_1755;
      end else begin
        if (_EVAL_2110) begin
          if (_EVAL_256) begin
            _EVAL_1649 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1652 <= 8'h0;
    end else begin
      if (_EVAL_135) begin
        _EVAL_1652 <= _EVAL_1205;
      end else begin
        if (_EVAL_1282) begin
          if (_EVAL_1598) begin
            _EVAL_1652 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1694 <= 8'h0;
    end else begin
      if (_EVAL_671) begin
        _EVAL_1694 <= _EVAL_868;
      end else begin
        if (_EVAL_1958) begin
          if (_EVAL_1973) begin
            _EVAL_1694 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1716 <= 8'h0;
    end else begin
      if (_EVAL_2194) begin
        _EVAL_1716 <= _EVAL_1755;
      end else begin
        if (_EVAL_2036) begin
          if (_EVAL_884) begin
            _EVAL_1716 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1768 <= 8'h0;
    end else begin
      if (_EVAL_929) begin
        _EVAL_1768 <= _EVAL_868;
      end else begin
        if (_EVAL_2214) begin
          if (_EVAL_1093) begin
            _EVAL_1768 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1785 <= 8'h0;
    end else begin
      if (_EVAL_2134) begin
        _EVAL_1785 <= _EVAL_1755;
      end else begin
        if (_EVAL_1697) begin
          if (_EVAL_312) begin
            _EVAL_1785 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1803 <= 1'h0;
    end else begin
      if (_EVAL_1596) begin
        _EVAL_1803 <= 1'h0;
      end else begin
        if (_EVAL_1456) begin
          _EVAL_1803 <= 1'h0;
        end else begin
          if (_EVAL_1269) begin
            _EVAL_1803 <= 1'h1;
          end else begin
            if (_EVAL_351) begin
              _EVAL_1803 <= 1'h0;
            end else begin
              if (_EVAL_1029) begin
                _EVAL_1803 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1829 <= 1'h0;
    end else begin
      if (_EVAL_969) begin
        _EVAL_1829 <= _EVAL_2229;
      end
    end
    if (_EVAL_703) begin
      _EVAL_1859 <= 8'h0;
    end else begin
      if (_EVAL_103) begin
        _EVAL_1859 <= _EVAL_1205;
      end else begin
        if (_EVAL_724) begin
          if (_EVAL_1750) begin
            _EVAL_1859 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_1787) begin
      if (_EVAL_1327) begin
        _EVAL_1866 <= 32'h13;
      end else begin
        _EVAL_1866 <= 32'h100073;
      end
    end
    if (_EVAL_703) begin
      _EVAL_1869 <= 8'h0;
    end else begin
      if (_EVAL_912) begin
        _EVAL_1869 <= _EVAL_562;
      end else begin
        if (_EVAL_386) begin
          if (_EVAL_444) begin
            _EVAL_1869 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1916 <= 8'h0;
    end else begin
      if (_EVAL_108) begin
        _EVAL_1916 <= _EVAL_1205;
      end else begin
        if (_EVAL_450) begin
          if (_EVAL_1242) begin
            _EVAL_1916 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1943 <= 8'h0;
    end else begin
      if (_EVAL_2014) begin
        _EVAL_1943 <= _EVAL_562;
      end else begin
        if (_EVAL_539) begin
          if (_EVAL_1831) begin
            _EVAL_1943 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_1951 <= 1'h0;
    end else begin
      if (_EVAL_1938) begin
        _EVAL_1951 <= _EVAL_1185;
      end
    end
    if (_EVAL_703) begin
      _EVAL_1991 <= 8'h0;
    end else begin
      if (_EVAL_1218) begin
        _EVAL_1991 <= _EVAL_562;
      end else begin
        if (_EVAL_500) begin
          if (_EVAL_614) begin
            _EVAL_1991 <= _EVAL_2060;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2000 <= 8'h0;
    end else begin
      if (_EVAL_1433) begin
        _EVAL_2000 <= _EVAL_1205;
      end else begin
        if (_EVAL_162) begin
          if (_EVAL_556) begin
            _EVAL_2000 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2026 <= 8'h0;
    end else begin
      if (_EVAL_2144) begin
        _EVAL_2026 <= _EVAL_868;
      end else begin
        if (_EVAL_990) begin
          if (_EVAL_1171) begin
            _EVAL_2026 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2054 <= 1'h0;
    end else begin
      if (_EVAL_1787) begin
        _EVAL_2054 <= 1'h1;
      end else begin
        if (_EVAL_875) begin
          _EVAL_2054 <= 1'h0;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2057 <= 8'h0;
    end else begin
      if (_EVAL_567) begin
        _EVAL_2057 <= _EVAL_1755;
      end else begin
        if (_EVAL_115) begin
          if (_EVAL_1821) begin
            _EVAL_2057 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2058 <= 8'h0;
    end else begin
      if (_EVAL_805) begin
        _EVAL_2058 <= _EVAL_1755;
      end else begin
        if (_EVAL_2185) begin
          if (_EVAL_1222) begin
            _EVAL_2058 <= _EVAL_142;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2082 <= 8'h0;
    end else begin
      if (_EVAL_887) begin
        _EVAL_2082 <= _EVAL_868;
      end else begin
        if (_EVAL_1234) begin
          if (_EVAL_487) begin
            _EVAL_2082 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2097 <= 8'h0;
    end else begin
      if (_EVAL_801) begin
        _EVAL_2097 <= _EVAL_1352;
      end else begin
        if (sb2tlOpt__EVAL_12) begin
          _EVAL_2097 <= sb2tlOpt__EVAL_19;
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2117 <= 1'h0;
    end else begin
      if (_EVAL_2032) begin
        _EVAL_2117 <= _EVAL_1762;
      end
    end
    if (_EVAL_703) begin
      _EVAL_2154 <= 8'h0;
    end else begin
      if (_EVAL_149) begin
        _EVAL_2154 <= _EVAL_868;
      end else begin
        if (_EVAL_2166) begin
          if (_EVAL_2109) begin
            _EVAL_2154 <= _EVAL_55;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2165 <= 8'h0;
    end else begin
      if (_EVAL_2139) begin
        _EVAL_2165 <= _EVAL_1205;
      end else begin
        if (_EVAL_465) begin
          if (_EVAL_517) begin
            _EVAL_2165 <= _EVAL_1352;
          end
        end
      end
    end
    if (_EVAL_703) begin
      _EVAL_2167 <= 3'h0;
    end else begin
      if (_EVAL_155) begin
        _EVAL_2167 <= _EVAL_1436;
      end
    end
    if (_EVAL_1787) begin
      if (_EVAL_73) begin
        if (_EVAL_774) begin
          _EVAL_2220 <= _EVAL_882;
        end else begin
          _EVAL_2220 <= _EVAL_1800;
        end
      end else begin
        _EVAL_2220 <= 32'h13;
      end
    end
  end
endmodule
