//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_255(
  input         _EVAL,
  input         _EVAL_0,
  input  [63:0] _EVAL_1,
  output [2:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [7:0]  _EVAL_7,
  output        _EVAL_8,
  output [2:0]  _EVAL_9,
  output [7:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  output        _EVAL_12,
  output [2:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  output [3:0]  _EVAL_15,
  output        _EVAL_16,
  input  [2:0]  _EVAL_17,
  output [31:0] _EVAL_18,
  output [63:0] _EVAL_19
);
  reg [2:0] _EVAL_22 [0:3];
  reg [31:0] _RAND_0;
  wire [2:0] _EVAL_22__EVAL_23_data;
  wire [1:0] _EVAL_22__EVAL_23_addr;
  wire [2:0] _EVAL_22__EVAL_24_data;
  wire [1:0] _EVAL_22__EVAL_24_addr;
  wire  _EVAL_22__EVAL_24_mask;
  wire  _EVAL_22__EVAL_24_en;
  reg [63:0] _EVAL_25 [0:3];
  reg [63:0] _RAND_1;
  wire [63:0] _EVAL_25__EVAL_26_data;
  wire [1:0] _EVAL_25__EVAL_26_addr;
  wire [63:0] _EVAL_25__EVAL_27_data;
  wire [1:0] _EVAL_25__EVAL_27_addr;
  wire  _EVAL_25__EVAL_27_mask;
  wire  _EVAL_25__EVAL_27_en;
  reg [2:0] _EVAL_31 [0:3];
  reg [31:0] _RAND_2;
  wire [2:0] _EVAL_31__EVAL_32_data;
  wire [1:0] _EVAL_31__EVAL_32_addr;
  wire [2:0] _EVAL_31__EVAL_33_data;
  wire [1:0] _EVAL_31__EVAL_33_addr;
  wire  _EVAL_31__EVAL_33_mask;
  wire  _EVAL_31__EVAL_33_en;
  reg  _EVAL_35 [0:3];
  reg [31:0] _RAND_3;
  wire  _EVAL_35__EVAL_36_data;
  wire [1:0] _EVAL_35__EVAL_36_addr;
  wire  _EVAL_35__EVAL_37_data;
  wire [1:0] _EVAL_35__EVAL_37_addr;
  wire  _EVAL_35__EVAL_37_mask;
  wire  _EVAL_35__EVAL_37_en;
  reg [3:0] _EVAL_38 [0:3];
  reg [31:0] _RAND_4;
  wire [3:0] _EVAL_38__EVAL_39_data;
  wire [1:0] _EVAL_38__EVAL_39_addr;
  wire [3:0] _EVAL_38__EVAL_40_data;
  wire [1:0] _EVAL_38__EVAL_40_addr;
  wire  _EVAL_38__EVAL_40_mask;
  wire  _EVAL_38__EVAL_40_en;
  reg [31:0] _EVAL_48 [0:3];
  reg [31:0] _RAND_5;
  wire [31:0] _EVAL_48__EVAL_49_data;
  wire [1:0] _EVAL_48__EVAL_49_addr;
  wire [31:0] _EVAL_48__EVAL_50_data;
  wire [1:0] _EVAL_48__EVAL_50_addr;
  wire  _EVAL_48__EVAL_50_mask;
  wire  _EVAL_48__EVAL_50_en;
  reg [2:0] _EVAL_51 [0:3];
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_51__EVAL_52_data;
  wire [1:0] _EVAL_51__EVAL_52_addr;
  wire [2:0] _EVAL_51__EVAL_53_data;
  wire [1:0] _EVAL_51__EVAL_53_addr;
  wire  _EVAL_51__EVAL_53_mask;
  wire  _EVAL_51__EVAL_53_en;
  reg [7:0] _EVAL_62 [0:3];
  reg [31:0] _RAND_7;
  wire [7:0] _EVAL_62__EVAL_63_data;
  wire [1:0] _EVAL_62__EVAL_63_addr;
  wire [7:0] _EVAL_62__EVAL_64_data;
  wire [1:0] _EVAL_62__EVAL_64_addr;
  wire  _EVAL_62__EVAL_64_mask;
  wire  _EVAL_62__EVAL_64_en;
  reg [1:0] _EVAL_30;
  reg [31:0] _RAND_8;
  reg  _EVAL_44;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_56;
  reg [31:0] _RAND_10;
  wire [1:0] _EVAL_43;
  wire  _EVAL_46;
  wire  _EVAL_60;
  wire  _EVAL_41;
  wire  _EVAL_55;
  wire  _EVAL_59;
  wire  _EVAL_42;
  wire  _EVAL_28;
  wire  _EVAL_47;
  wire  _EVAL_57;
  wire  _EVAL_21;
  wire  _EVAL_20;
  wire [1:0] _EVAL_58;
  assign _EVAL_22__EVAL_23_addr = _EVAL_30;
  assign _EVAL_22__EVAL_23_data = _EVAL_22[_EVAL_22__EVAL_23_addr];
  assign _EVAL_22__EVAL_24_data = _EVAL_17;
  assign _EVAL_22__EVAL_24_addr = _EVAL_56;
  assign _EVAL_22__EVAL_24_mask = 1'h1;
  assign _EVAL_22__EVAL_24_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_25__EVAL_26_addr = _EVAL_30;
  assign _EVAL_25__EVAL_26_data = _EVAL_25[_EVAL_25__EVAL_26_addr];
  assign _EVAL_25__EVAL_27_data = _EVAL_1;
  assign _EVAL_25__EVAL_27_addr = _EVAL_56;
  assign _EVAL_25__EVAL_27_mask = 1'h1;
  assign _EVAL_25__EVAL_27_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_31__EVAL_32_addr = _EVAL_30;
  assign _EVAL_31__EVAL_32_data = _EVAL_31[_EVAL_31__EVAL_32_addr];
  assign _EVAL_31__EVAL_33_data = _EVAL_11;
  assign _EVAL_31__EVAL_33_addr = _EVAL_56;
  assign _EVAL_31__EVAL_33_mask = 1'h1;
  assign _EVAL_31__EVAL_33_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_35__EVAL_36_addr = _EVAL_30;
  assign _EVAL_35__EVAL_36_data = _EVAL_35[_EVAL_35__EVAL_36_addr];
  assign _EVAL_35__EVAL_37_data = 1'h0;
  assign _EVAL_35__EVAL_37_addr = _EVAL_56;
  assign _EVAL_35__EVAL_37_mask = 1'h1;
  assign _EVAL_35__EVAL_37_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_38__EVAL_39_addr = _EVAL_30;
  assign _EVAL_38__EVAL_39_data = _EVAL_38[_EVAL_38__EVAL_39_addr];
  assign _EVAL_38__EVAL_40_data = _EVAL_3;
  assign _EVAL_38__EVAL_40_addr = _EVAL_56;
  assign _EVAL_38__EVAL_40_mask = 1'h1;
  assign _EVAL_38__EVAL_40_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_48__EVAL_49_addr = _EVAL_30;
  assign _EVAL_48__EVAL_49_data = _EVAL_48[_EVAL_48__EVAL_49_addr];
  assign _EVAL_48__EVAL_50_data = _EVAL_14;
  assign _EVAL_48__EVAL_50_addr = _EVAL_56;
  assign _EVAL_48__EVAL_50_mask = 1'h1;
  assign _EVAL_48__EVAL_50_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_51__EVAL_52_addr = _EVAL_30;
  assign _EVAL_51__EVAL_52_data = _EVAL_51[_EVAL_51__EVAL_52_addr];
  assign _EVAL_51__EVAL_53_data = _EVAL_5;
  assign _EVAL_51__EVAL_53_addr = _EVAL_56;
  assign _EVAL_51__EVAL_53_mask = 1'h1;
  assign _EVAL_51__EVAL_53_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_62__EVAL_63_addr = _EVAL_30;
  assign _EVAL_62__EVAL_63_data = _EVAL_62[_EVAL_62__EVAL_63_addr];
  assign _EVAL_62__EVAL_64_data = _EVAL_7;
  assign _EVAL_62__EVAL_64_addr = _EVAL_56;
  assign _EVAL_62__EVAL_64_mask = 1'h1;
  assign _EVAL_62__EVAL_64_en = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_43 = _EVAL_56 + 2'h1;
  assign _EVAL_46 = _EVAL_8 & _EVAL;
  assign _EVAL_60 = _EVAL_4 ? 1'h0 : _EVAL_46;
  assign _EVAL_41 = _EVAL_56 == _EVAL_30;
  assign _EVAL_55 = _EVAL_44 == 1'h0;
  assign _EVAL_59 = _EVAL_41 & _EVAL_55;
  assign _EVAL_42 = _EVAL_59 ? _EVAL_60 : _EVAL_46;
  assign _EVAL_28 = _EVAL_59 == 1'h0;
  assign _EVAL_47 = _EVAL_4 & _EVAL_16;
  assign _EVAL_57 = _EVAL_41 & _EVAL_44;
  assign _EVAL_21 = _EVAL_59 ? 1'h0 : _EVAL_47;
  assign _EVAL_20 = _EVAL_42 != _EVAL_21;
  assign _EVAL_58 = _EVAL_30 + 2'h1;
  assign _EVAL_15 = _EVAL_59 ? _EVAL_3 : _EVAL_38__EVAL_39_data;
  assign _EVAL_10 = _EVAL_59 ? _EVAL_7 : _EVAL_62__EVAL_63_data;
  assign _EVAL_19 = _EVAL_59 ? _EVAL_1 : _EVAL_25__EVAL_26_data;
  assign _EVAL_12 = _EVAL_59 ? 1'h0 : _EVAL_35__EVAL_36_data;
  assign _EVAL_8 = _EVAL_57 == 1'h0;
  assign _EVAL_2 = _EVAL_59 ? _EVAL_17 : _EVAL_22__EVAL_23_data;
  assign _EVAL_9 = _EVAL_59 ? _EVAL_11 : _EVAL_31__EVAL_32_data;
  assign _EVAL_13 = _EVAL_59 ? _EVAL_5 : _EVAL_51__EVAL_52_data;
  assign _EVAL_16 = _EVAL ? 1'h1 : _EVAL_28;
  assign _EVAL_18 = _EVAL_59 ? _EVAL_14 : _EVAL_48__EVAL_49_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_22[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_25[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_31[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_35[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_38[initvar] = _RAND_4[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_48[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_51[initvar] = _RAND_6[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_62[initvar] = _RAND_7[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_30 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_44 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_56 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if(_EVAL_22__EVAL_24_en & _EVAL_22__EVAL_24_mask) begin
      _EVAL_22[_EVAL_22__EVAL_24_addr] <= _EVAL_22__EVAL_24_data;
    end
    if(_EVAL_25__EVAL_27_en & _EVAL_25__EVAL_27_mask) begin
      _EVAL_25[_EVAL_25__EVAL_27_addr] <= _EVAL_25__EVAL_27_data;
    end
    if(_EVAL_31__EVAL_33_en & _EVAL_31__EVAL_33_mask) begin
      _EVAL_31[_EVAL_31__EVAL_33_addr] <= _EVAL_31__EVAL_33_data;
    end
    if(_EVAL_35__EVAL_37_en & _EVAL_35__EVAL_37_mask) begin
      _EVAL_35[_EVAL_35__EVAL_37_addr] <= _EVAL_35__EVAL_37_data;
    end
    if(_EVAL_38__EVAL_40_en & _EVAL_38__EVAL_40_mask) begin
      _EVAL_38[_EVAL_38__EVAL_40_addr] <= _EVAL_38__EVAL_40_data;
    end
    if(_EVAL_48__EVAL_50_en & _EVAL_48__EVAL_50_mask) begin
      _EVAL_48[_EVAL_48__EVAL_50_addr] <= _EVAL_48__EVAL_50_data;
    end
    if(_EVAL_51__EVAL_53_en & _EVAL_51__EVAL_53_mask) begin
      _EVAL_51[_EVAL_51__EVAL_53_addr] <= _EVAL_51__EVAL_53_data;
    end
    if(_EVAL_62__EVAL_64_en & _EVAL_62__EVAL_64_mask) begin
      _EVAL_62[_EVAL_62__EVAL_64_addr] <= _EVAL_62__EVAL_64_data;
    end
    if (_EVAL_6) begin
      _EVAL_30 <= 2'h0;
    end else begin
      if (_EVAL_21) begin
        _EVAL_30 <= _EVAL_58;
      end
    end
    if (_EVAL_6) begin
      _EVAL_44 <= 1'h0;
    end else begin
      if (_EVAL_20) begin
        if (_EVAL_59) begin
          if (_EVAL_4) begin
            _EVAL_44 <= 1'h0;
          end else begin
            _EVAL_44 <= _EVAL_46;
          end
        end else begin
          _EVAL_44 <= _EVAL_46;
        end
      end
    end
    if (_EVAL_6) begin
      _EVAL_56 <= 2'h0;
    end else begin
      if (_EVAL_42) begin
        _EVAL_56 <= _EVAL_43;
      end
    end
  end
endmodule
