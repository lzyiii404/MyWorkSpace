//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_79(
  output        _EVAL,
  output [4:0]  _EVAL_0,
  input  [31:0] _EVAL_1,
  output [31:0] _EVAL_2,
  input  [31:0] _EVAL_3,
  input  [7:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  output [2:0]  _EVAL_7,
  output [7:0]  _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input  [7:0]  _EVAL_11,
  input  [7:0]  _EVAL_12,
  output [31:0] _EVAL_13,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  output [7:0]  _EVAL_17,
  output [31:0] _EVAL_18,
  input         _EVAL_19,
  input  [1:0]  _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input  [2:0]  _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input  [2:0]  _EVAL_29,
  input  [7:0]  _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  output [3:0]  _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input  [1:0]  _EVAL_36,
  input  [31:0] _EVAL_37,
  output [3:0]  _EVAL_38,
  input  [4:0]  _EVAL_39,
  output        _EVAL_40,
  output [2:0]  _EVAL_41,
  output [1:0]  _EVAL_42,
  input  [31:0] _EVAL_43,
  input  [3:0]  _EVAL_44,
  output        _EVAL_45,
  output [1:0]  _EVAL_46,
  input  [2:0]  _EVAL_47,
  output        _EVAL_48,
  output        _EVAL_49
);
  wire  axi42tl__EVAL;
  wire  axi42tl__EVAL_0;
  wire [31:0] axi42tl__EVAL_1;
  wire  axi42tl__EVAL_2;
  wire [31:0] axi42tl__EVAL_3;
  wire [31:0] axi42tl__EVAL_4;
  wire [1:0] axi42tl__EVAL_5;
  wire  axi42tl__EVAL_6;
  wire  axi42tl__EVAL_7;
  wire [3:0] axi42tl__EVAL_8;
  wire [4:0] axi42tl__EVAL_9;
  wire  axi42tl__EVAL_10;
  wire [1:0] axi42tl__EVAL_11;
  wire [2:0] axi42tl__EVAL_12;
  wire [4:0] axi42tl__EVAL_13;
  wire [31:0] axi42tl__EVAL_14;
  wire  axi42tl__EVAL_15;
  wire [7:0] axi42tl__EVAL_16;
  wire  axi42tl__EVAL_17;
  wire [2:0] axi42tl__EVAL_18;
  wire  axi42tl__EVAL_19;
  wire [3:0] axi42tl__EVAL_20;
  wire  axi42tl__EVAL_21;
  wire [7:0] axi42tl__EVAL_22;
  wire  axi42tl__EVAL_23;
  wire  axi42tl__EVAL_24;
  wire [31:0] axi42tl__EVAL_25;
  wire  axi42tl__EVAL_26;
  wire [2:0] axi42tl__EVAL_27;
  wire  axi42tl__EVAL_28;
  wire [31:0] axi42tl__EVAL_29;
  wire [2:0] axi42tl__EVAL_30;
  wire  axi42tl__EVAL_31;
  wire  axi42tl__EVAL_32;
  wire [2:0] axi42tl__EVAL_33;
  wire  axi42tl__EVAL_34;
  wire  axi42tl__EVAL_35;
  wire  axi42tl__EVAL_36;
  wire [1:0] axi42tl__EVAL_37;
  wire [3:0] axi42tl__EVAL_38;
  wire [31:0] axi42tl__EVAL_39;
  wire  axi42tl__EVAL_40;
  wire [1:0] axi42tl__EVAL_41;
  wire [3:0] axi42tl__EVAL_42;
  wire [1:0] axi42tl__EVAL_43;
  wire  axi42tl__EVAL_44;
  wire [1:0] axi42tl__EVAL_45;
  wire [31:0] buffer__EVAL;
  wire [4:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire [2:0] buffer__EVAL_4;
  wire [3:0] buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [31:0] buffer__EVAL_10;
  wire [2:0] buffer__EVAL_11;
  wire [2:0] buffer__EVAL_12;
  wire [31:0] buffer__EVAL_13;
  wire [4:0] buffer__EVAL_14;
  wire [4:0] buffer__EVAL_15;
  wire [2:0] buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire [31:0] buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire [4:0] buffer__EVAL_20;
  wire [31:0] buffer__EVAL_21;
  wire [3:0] buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire [31:0] buffer__EVAL_24;
  wire [3:0] buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire [2:0] buffer__EVAL_29;
  wire [1:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [2:0] buffer__EVAL_33;
  wire [3:0] buffer__EVAL_34;
  wire  buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [3:0] buffer__EVAL_37;
  wire [3:0] buffer__EVAL_38;
  wire  buffer__EVAL_39;
  wire [1:0] buffer__EVAL_40;
  wire  axi4yank__EVAL;
  wire  axi4yank__EVAL_0;
  wire [1:0] axi4yank__EVAL_1;
  wire  axi4yank__EVAL_2;
  wire  axi4yank__EVAL_3;
  wire [31:0] axi4yank__EVAL_4;
  wire [2:0] axi4yank__EVAL_5;
  wire  axi4yank__EVAL_6;
  wire [6:0] axi4yank__EVAL_7;
  wire [3:0] axi4yank__EVAL_8;
  wire  axi4yank__EVAL_9;
  wire  axi4yank__EVAL_10;
  wire  axi4yank__EVAL_11;
  wire [7:0] axi4yank__EVAL_12;
  wire  axi4yank__EVAL_13;
  wire  axi4yank__EVAL_14;
  wire  axi4yank__EVAL_15;
  wire [1:0] axi4yank__EVAL_16;
  wire  axi4yank__EVAL_17;
  wire  axi4yank__EVAL_18;
  wire [3:0] axi4yank__EVAL_19;
  wire [31:0] axi4yank__EVAL_20;
  wire  axi4yank__EVAL_21;
  wire  axi4yank__EVAL_22;
  wire  axi4yank__EVAL_23;
  wire [1:0] axi4yank__EVAL_24;
  wire [1:0] axi4yank__EVAL_25;
  wire  axi4yank__EVAL_26;
  wire [1:0] axi4yank__EVAL_27;
  wire [6:0] axi4yank__EVAL_28;
  wire [1:0] axi4yank__EVAL_29;
  wire  axi4yank__EVAL_30;
  wire [31:0] axi4yank__EVAL_31;
  wire [1:0] axi4yank__EVAL_32;
  wire [1:0] axi4yank__EVAL_33;
  wire [6:0] axi4yank__EVAL_34;
  wire [7:0] axi4yank__EVAL_35;
  wire [31:0] axi4yank__EVAL_36;
  wire [31:0] axi4yank__EVAL_37;
  wire [1:0] axi4yank__EVAL_38;
  wire [7:0] axi4yank__EVAL_39;
  wire  axi4yank__EVAL_40;
  wire [2:0] axi4yank__EVAL_41;
  wire  axi4yank__EVAL_42;
  wire  axi4yank__EVAL_43;
  wire [31:0] axi4yank__EVAL_44;
  wire  axi4yank__EVAL_45;
  wire  axi4yank__EVAL_46;
  wire [7:0] axi4yank__EVAL_47;
  wire  axi4yank__EVAL_48;
  wire  axi4yank__EVAL_49;
  wire [2:0] axi4yank__EVAL_50;
  wire [6:0] axi4yank__EVAL_51;
  wire [1:0] axi4yank__EVAL_52;
  wire [1:0] axi4yank__EVAL_53;
  wire  axi4yank__EVAL_54;
  wire [1:0] axi4yank__EVAL_55;
  wire [2:0] axi4yank__EVAL_56;
  wire [31:0] axi4yank__EVAL_57;
  wire [31:0] axi4yank__EVAL_58;
  wire [7:0] axi4buf__EVAL;
  wire  axi4buf__EVAL_0;
  wire [7:0] axi4buf__EVAL_1;
  wire [7:0] axi4buf__EVAL_2;
  wire  axi4buf__EVAL_3;
  wire [1:0] axi4buf__EVAL_4;
  wire  axi4buf__EVAL_5;
  wire  axi4buf__EVAL_6;
  wire [2:0] axi4buf__EVAL_7;
  wire [1:0] axi4buf__EVAL_8;
  wire  axi4buf__EVAL_9;
  wire [31:0] axi4buf__EVAL_10;
  wire [7:0] axi4buf__EVAL_11;
  wire [31:0] axi4buf__EVAL_12;
  wire [1:0] axi4buf__EVAL_13;
  wire [31:0] axi4buf__EVAL_14;
  wire  axi4buf__EVAL_15;
  wire [7:0] axi4buf__EVAL_16;
  wire  axi4buf__EVAL_17;
  wire  axi4buf__EVAL_18;
  wire [31:0] axi4buf__EVAL_19;
  wire [7:0] axi4buf__EVAL_20;
  wire [2:0] axi4buf__EVAL_21;
  wire [3:0] axi4buf__EVAL_22;
  wire [31:0] axi4buf__EVAL_23;
  wire [2:0] axi4buf__EVAL_24;
  wire [7:0] axi4buf__EVAL_25;
  wire [31:0] axi4buf__EVAL_26;
  wire  axi4buf__EVAL_27;
  wire [31:0] axi4buf__EVAL_28;
  wire  axi4buf__EVAL_29;
  wire  axi4buf__EVAL_30;
  wire [7:0] axi4buf__EVAL_31;
  wire  axi4buf__EVAL_32;
  wire  axi4buf__EVAL_33;
  wire [7:0] axi4buf__EVAL_34;
  wire [7:0] axi4buf__EVAL_35;
  wire [2:0] axi4buf__EVAL_36;
  wire  axi4buf__EVAL_37;
  wire  axi4buf__EVAL_38;
  wire [1:0] axi4buf__EVAL_39;
  wire [1:0] axi4buf__EVAL_40;
  wire  axi4buf__EVAL_41;
  wire  axi4buf__EVAL_42;
  wire [31:0] axi4buf__EVAL_43;
  wire  axi4buf__EVAL_44;
  wire  axi4buf__EVAL_45;
  wire [1:0] axi4buf__EVAL_46;
  wire  axi4buf__EVAL_47;
  wire  axi4buf__EVAL_48;
  wire [1:0] axi4buf__EVAL_49;
  wire [1:0] axi4buf__EVAL_50;
  wire  axi4buf__EVAL_51;
  wire  axi4buf__EVAL_52;
  wire [3:0] axi4buf__EVAL_53;
  wire  axi4buf__EVAL_54;
  wire [7:0] axi4buf__EVAL_55;
  wire  axi4buf__EVAL_56;
  wire  axi4buf__EVAL_57;
  wire [7:0] axi4buf__EVAL_58;
  wire  axi4frag__EVAL;
  wire  axi4frag__EVAL_0;
  wire  axi4frag__EVAL_1;
  wire [31:0] axi4frag__EVAL_2;
  wire [6:0] axi4frag__EVAL_3;
  wire [2:0] axi4frag__EVAL_4;
  wire  axi4frag__EVAL_5;
  wire [5:0] axi4frag__EVAL_6;
  wire  axi4frag__EVAL_7;
  wire  axi4frag__EVAL_8;
  wire [1:0] axi4frag__EVAL_9;
  wire [6:0] axi4frag__EVAL_10;
  wire [7:0] axi4frag__EVAL_11;
  wire [7:0] axi4frag__EVAL_12;
  wire [1:0] axi4frag__EVAL_13;
  wire [1:0] axi4frag__EVAL_14;
  wire [1:0] axi4frag__EVAL_15;
  wire [31:0] axi4frag__EVAL_16;
  wire  axi4frag__EVAL_17;
  wire  axi4frag__EVAL_18;
  wire  axi4frag__EVAL_19;
  wire [2:0] axi4frag__EVAL_20;
  wire [31:0] axi4frag__EVAL_21;
  wire [2:0] axi4frag__EVAL_22;
  wire  axi4frag__EVAL_23;
  wire [1:0] axi4frag__EVAL_24;
  wire  axi4frag__EVAL_25;
  wire  axi4frag__EVAL_26;
  wire [5:0] axi4frag__EVAL_27;
  wire  axi4frag__EVAL_28;
  wire  axi4frag__EVAL_29;
  wire [3:0] axi4frag__EVAL_30;
  wire [31:0] axi4frag__EVAL_31;
  wire  axi4frag__EVAL_32;
  wire [1:0] axi4frag__EVAL_33;
  wire [3:0] axi4frag__EVAL_34;
  wire  axi4frag__EVAL_35;
  wire  axi4frag__EVAL_36;
  wire [1:0] axi4frag__EVAL_37;
  wire [1:0] axi4frag__EVAL_38;
  wire [6:0] axi4frag__EVAL_39;
  wire [2:0] axi4frag__EVAL_40;
  wire [5:0] axi4frag__EVAL_41;
  wire [7:0] axi4frag__EVAL_42;
  wire [31:0] axi4frag__EVAL_43;
  wire  axi4frag__EVAL_44;
  wire [31:0] axi4frag__EVAL_45;
  wire [5:0] axi4frag__EVAL_46;
  wire [1:0] axi4frag__EVAL_47;
  wire  axi4frag__EVAL_48;
  wire  axi4frag__EVAL_49;
  wire  axi4frag__EVAL_50;
  wire [1:0] axi4frag__EVAL_51;
  wire [1:0] axi4frag__EVAL_52;
  wire  axi4frag__EVAL_53;
  wire [1:0] axi4frag__EVAL_54;
  wire  axi4frag__EVAL_55;
  wire [31:0] axi4frag__EVAL_56;
  wire  axi4frag__EVAL_57;
  wire [1:0] axi4frag__EVAL_58;
  wire [1:0] axi4frag__EVAL_59;
  wire  axi4frag__EVAL_60;
  wire  axi4frag__EVAL_61;
  wire [31:0] axi4frag__EVAL_62;
  wire [6:0] axi4frag__EVAL_63;
  wire [7:0] axi4frag__EVAL_64;
  wire [31:0] fixer__EVAL;
  wire [2:0] fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire [1:0] fixer__EVAL_2;
  wire  fixer__EVAL_3;
  wire [2:0] fixer__EVAL_4;
  wire [4:0] fixer__EVAL_5;
  wire [31:0] fixer__EVAL_6;
  wire [31:0] fixer__EVAL_7;
  wire [2:0] fixer__EVAL_8;
  wire  fixer__EVAL_9;
  wire [4:0] fixer__EVAL_10;
  wire  fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire [31:0] fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire [3:0] fixer__EVAL_15;
  wire [2:0] fixer__EVAL_16;
  wire [4:0] fixer__EVAL_17;
  wire [1:0] fixer__EVAL_18;
  wire [2:0] fixer__EVAL_19;
  wire [31:0] fixer__EVAL_20;
  wire  fixer__EVAL_21;
  wire [3:0] fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire  fixer__EVAL_24;
  wire  fixer__EVAL_25;
  wire [3:0] fixer__EVAL_26;
  wire [4:0] fixer__EVAL_27;
  wire  fixer__EVAL_28;
  wire  fixer__EVAL_29;
  wire [2:0] fixer__EVAL_30;
  wire  fixer__EVAL_31;
  wire [3:0] fixer__EVAL_32;
  wire [3:0] fixer__EVAL_33;
  wire [3:0] fixer__EVAL_34;
  wire  fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire [31:0] fixer__EVAL_37;
  wire  fixer__EVAL_38;
  wire  fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire [5:0] axi4index__EVAL;
  wire  axi4index__EVAL_0;
  wire [31:0] axi4index__EVAL_1;
  wire [1:0] axi4index__EVAL_2;
  wire [2:0] axi4index__EVAL_3;
  wire [7:0] axi4index__EVAL_4;
  wire [31:0] axi4index__EVAL_5;
  wire  axi4index__EVAL_6;
  wire [1:0] axi4index__EVAL_7;
  wire [2:0] axi4index__EVAL_8;
  wire  axi4index__EVAL_9;
  wire [1:0] axi4index__EVAL_10;
  wire [3:0] axi4index__EVAL_11;
  wire [1:0] axi4index__EVAL_12;
  wire [1:0] axi4index__EVAL_13;
  wire [31:0] axi4index__EVAL_14;
  wire [1:0] axi4index__EVAL_15;
  wire [3:0] axi4index__EVAL_16;
  wire [7:0] axi4index__EVAL_17;
  wire [5:0] axi4index__EVAL_18;
  wire [31:0] axi4index__EVAL_19;
  wire [7:0] axi4index__EVAL_20;
  wire  axi4index__EVAL_21;
  wire [7:0] axi4index__EVAL_22;
  wire  axi4index__EVAL_23;
  wire  axi4index__EVAL_24;
  wire  axi4index__EVAL_25;
  wire  axi4index__EVAL_26;
  wire  axi4index__EVAL_27;
  wire [1:0] axi4index__EVAL_28;
  wire  axi4index__EVAL_29;
  wire [7:0] axi4index__EVAL_30;
  wire [7:0] axi4index__EVAL_31;
  wire [7:0] axi4index__EVAL_32;
  wire [1:0] axi4index__EVAL_33;
  wire [31:0] axi4index__EVAL_34;
  wire [31:0] axi4index__EVAL_35;
  wire  axi4index__EVAL_36;
  wire [2:0] axi4index__EVAL_37;
  wire [5:0] axi4index__EVAL_38;
  wire  axi4index__EVAL_39;
  wire [7:0] axi4index__EVAL_40;
  wire  axi4index__EVAL_41;
  wire  axi4index__EVAL_42;
  wire  axi4index__EVAL_43;
  wire  axi4index__EVAL_44;
  wire [1:0] axi4index__EVAL_45;
  wire [1:0] axi4index__EVAL_46;
  wire [1:0] axi4index__EVAL_47;
  wire  axi4index__EVAL_48;
  wire  axi4index__EVAL_49;
  wire [31:0] axi4index__EVAL_50;
  wire  axi4index__EVAL_51;
  wire  axi4index__EVAL_52;
  wire  axi4index__EVAL_53;
  wire [31:0] axi4index__EVAL_54;
  wire  axi4index__EVAL_55;
  wire [5:0] axi4index__EVAL_56;
  wire  axi4index__EVAL_57;
  wire  axi4index__EVAL_58;
  wire [2:0] axi4index__EVAL_59;
  wire [1:0] axi4index__EVAL_60;
  wire [1:0] widget__EVAL;
  wire [3:0] widget__EVAL_0;
  wire  widget__EVAL_1;
  wire  widget__EVAL_2;
  wire  widget__EVAL_3;
  wire  widget__EVAL_4;
  wire  widget__EVAL_5;
  wire [2:0] widget__EVAL_6;
  wire [31:0] widget__EVAL_7;
  wire [31:0] widget__EVAL_8;
  wire  widget__EVAL_9;
  wire  widget__EVAL_10;
  wire  widget__EVAL_11;
  wire [31:0] widget__EVAL_12;
  wire [3:0] widget__EVAL_13;
  wire [4:0] widget__EVAL_14;
  wire [2:0] widget__EVAL_15;
  wire [3:0] widget__EVAL_16;
  wire [2:0] widget__EVAL_17;
  wire  widget__EVAL_18;
  wire  widget__EVAL_19;
  wire  widget__EVAL_20;
  wire [3:0] widget__EVAL_21;
  wire [4:0] widget__EVAL_22;
  wire  widget__EVAL_23;
  wire  widget__EVAL_24;
  wire [31:0] widget__EVAL_25;
  wire  widget__EVAL_26;
  wire  widget__EVAL_27;
  wire [3:0] widget__EVAL_28;
  wire [31:0] widget__EVAL_29;
  wire [4:0] widget__EVAL_30;
  wire [2:0] widget__EVAL_31;
  wire [2:0] widget__EVAL_32;
  wire  widget__EVAL_33;
  wire [31:0] widget__EVAL_34;
  wire [2:0] widget__EVAL_35;
  wire  widget__EVAL_36;
  wire [3:0] widget__EVAL_37;
  wire [4:0] widget__EVAL_38;
  SiFive__EVAL_69 axi42tl (
    ._EVAL(axi42tl__EVAL),
    ._EVAL_0(axi42tl__EVAL_0),
    ._EVAL_1(axi42tl__EVAL_1),
    ._EVAL_2(axi42tl__EVAL_2),
    ._EVAL_3(axi42tl__EVAL_3),
    ._EVAL_4(axi42tl__EVAL_4),
    ._EVAL_5(axi42tl__EVAL_5),
    ._EVAL_6(axi42tl__EVAL_6),
    ._EVAL_7(axi42tl__EVAL_7),
    ._EVAL_8(axi42tl__EVAL_8),
    ._EVAL_9(axi42tl__EVAL_9),
    ._EVAL_10(axi42tl__EVAL_10),
    ._EVAL_11(axi42tl__EVAL_11),
    ._EVAL_12(axi42tl__EVAL_12),
    ._EVAL_13(axi42tl__EVAL_13),
    ._EVAL_14(axi42tl__EVAL_14),
    ._EVAL_15(axi42tl__EVAL_15),
    ._EVAL_16(axi42tl__EVAL_16),
    ._EVAL_17(axi42tl__EVAL_17),
    ._EVAL_18(axi42tl__EVAL_18),
    ._EVAL_19(axi42tl__EVAL_19),
    ._EVAL_20(axi42tl__EVAL_20),
    ._EVAL_21(axi42tl__EVAL_21),
    ._EVAL_22(axi42tl__EVAL_22),
    ._EVAL_23(axi42tl__EVAL_23),
    ._EVAL_24(axi42tl__EVAL_24),
    ._EVAL_25(axi42tl__EVAL_25),
    ._EVAL_26(axi42tl__EVAL_26),
    ._EVAL_27(axi42tl__EVAL_27),
    ._EVAL_28(axi42tl__EVAL_28),
    ._EVAL_29(axi42tl__EVAL_29),
    ._EVAL_30(axi42tl__EVAL_30),
    ._EVAL_31(axi42tl__EVAL_31),
    ._EVAL_32(axi42tl__EVAL_32),
    ._EVAL_33(axi42tl__EVAL_33),
    ._EVAL_34(axi42tl__EVAL_34),
    ._EVAL_35(axi42tl__EVAL_35),
    ._EVAL_36(axi42tl__EVAL_36),
    ._EVAL_37(axi42tl__EVAL_37),
    ._EVAL_38(axi42tl__EVAL_38),
    ._EVAL_39(axi42tl__EVAL_39),
    ._EVAL_40(axi42tl__EVAL_40),
    ._EVAL_41(axi42tl__EVAL_41),
    ._EVAL_42(axi42tl__EVAL_42),
    ._EVAL_43(axi42tl__EVAL_43),
    ._EVAL_44(axi42tl__EVAL_44),
    ._EVAL_45(axi42tl__EVAL_45)
  );
  SiFive__EVAL_62 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40)
  );
  SiFive__EVAL_71 axi4yank (
    ._EVAL(axi4yank__EVAL),
    ._EVAL_0(axi4yank__EVAL_0),
    ._EVAL_1(axi4yank__EVAL_1),
    ._EVAL_2(axi4yank__EVAL_2),
    ._EVAL_3(axi4yank__EVAL_3),
    ._EVAL_4(axi4yank__EVAL_4),
    ._EVAL_5(axi4yank__EVAL_5),
    ._EVAL_6(axi4yank__EVAL_6),
    ._EVAL_7(axi4yank__EVAL_7),
    ._EVAL_8(axi4yank__EVAL_8),
    ._EVAL_9(axi4yank__EVAL_9),
    ._EVAL_10(axi4yank__EVAL_10),
    ._EVAL_11(axi4yank__EVAL_11),
    ._EVAL_12(axi4yank__EVAL_12),
    ._EVAL_13(axi4yank__EVAL_13),
    ._EVAL_14(axi4yank__EVAL_14),
    ._EVAL_15(axi4yank__EVAL_15),
    ._EVAL_16(axi4yank__EVAL_16),
    ._EVAL_17(axi4yank__EVAL_17),
    ._EVAL_18(axi4yank__EVAL_18),
    ._EVAL_19(axi4yank__EVAL_19),
    ._EVAL_20(axi4yank__EVAL_20),
    ._EVAL_21(axi4yank__EVAL_21),
    ._EVAL_22(axi4yank__EVAL_22),
    ._EVAL_23(axi4yank__EVAL_23),
    ._EVAL_24(axi4yank__EVAL_24),
    ._EVAL_25(axi4yank__EVAL_25),
    ._EVAL_26(axi4yank__EVAL_26),
    ._EVAL_27(axi4yank__EVAL_27),
    ._EVAL_28(axi4yank__EVAL_28),
    ._EVAL_29(axi4yank__EVAL_29),
    ._EVAL_30(axi4yank__EVAL_30),
    ._EVAL_31(axi4yank__EVAL_31),
    ._EVAL_32(axi4yank__EVAL_32),
    ._EVAL_33(axi4yank__EVAL_33),
    ._EVAL_34(axi4yank__EVAL_34),
    ._EVAL_35(axi4yank__EVAL_35),
    ._EVAL_36(axi4yank__EVAL_36),
    ._EVAL_37(axi4yank__EVAL_37),
    ._EVAL_38(axi4yank__EVAL_38),
    ._EVAL_39(axi4yank__EVAL_39),
    ._EVAL_40(axi4yank__EVAL_40),
    ._EVAL_41(axi4yank__EVAL_41),
    ._EVAL_42(axi4yank__EVAL_42),
    ._EVAL_43(axi4yank__EVAL_43),
    ._EVAL_44(axi4yank__EVAL_44),
    ._EVAL_45(axi4yank__EVAL_45),
    ._EVAL_46(axi4yank__EVAL_46),
    ._EVAL_47(axi4yank__EVAL_47),
    ._EVAL_48(axi4yank__EVAL_48),
    ._EVAL_49(axi4yank__EVAL_49),
    ._EVAL_50(axi4yank__EVAL_50),
    ._EVAL_51(axi4yank__EVAL_51),
    ._EVAL_52(axi4yank__EVAL_52),
    ._EVAL_53(axi4yank__EVAL_53),
    ._EVAL_54(axi4yank__EVAL_54),
    ._EVAL_55(axi4yank__EVAL_55),
    ._EVAL_56(axi4yank__EVAL_56),
    ._EVAL_57(axi4yank__EVAL_57),
    ._EVAL_58(axi4yank__EVAL_58)
  );
  SiFive__EVAL_78 axi4buf (
    ._EVAL(axi4buf__EVAL),
    ._EVAL_0(axi4buf__EVAL_0),
    ._EVAL_1(axi4buf__EVAL_1),
    ._EVAL_2(axi4buf__EVAL_2),
    ._EVAL_3(axi4buf__EVAL_3),
    ._EVAL_4(axi4buf__EVAL_4),
    ._EVAL_5(axi4buf__EVAL_5),
    ._EVAL_6(axi4buf__EVAL_6),
    ._EVAL_7(axi4buf__EVAL_7),
    ._EVAL_8(axi4buf__EVAL_8),
    ._EVAL_9(axi4buf__EVAL_9),
    ._EVAL_10(axi4buf__EVAL_10),
    ._EVAL_11(axi4buf__EVAL_11),
    ._EVAL_12(axi4buf__EVAL_12),
    ._EVAL_13(axi4buf__EVAL_13),
    ._EVAL_14(axi4buf__EVAL_14),
    ._EVAL_15(axi4buf__EVAL_15),
    ._EVAL_16(axi4buf__EVAL_16),
    ._EVAL_17(axi4buf__EVAL_17),
    ._EVAL_18(axi4buf__EVAL_18),
    ._EVAL_19(axi4buf__EVAL_19),
    ._EVAL_20(axi4buf__EVAL_20),
    ._EVAL_21(axi4buf__EVAL_21),
    ._EVAL_22(axi4buf__EVAL_22),
    ._EVAL_23(axi4buf__EVAL_23),
    ._EVAL_24(axi4buf__EVAL_24),
    ._EVAL_25(axi4buf__EVAL_25),
    ._EVAL_26(axi4buf__EVAL_26),
    ._EVAL_27(axi4buf__EVAL_27),
    ._EVAL_28(axi4buf__EVAL_28),
    ._EVAL_29(axi4buf__EVAL_29),
    ._EVAL_30(axi4buf__EVAL_30),
    ._EVAL_31(axi4buf__EVAL_31),
    ._EVAL_32(axi4buf__EVAL_32),
    ._EVAL_33(axi4buf__EVAL_33),
    ._EVAL_34(axi4buf__EVAL_34),
    ._EVAL_35(axi4buf__EVAL_35),
    ._EVAL_36(axi4buf__EVAL_36),
    ._EVAL_37(axi4buf__EVAL_37),
    ._EVAL_38(axi4buf__EVAL_38),
    ._EVAL_39(axi4buf__EVAL_39),
    ._EVAL_40(axi4buf__EVAL_40),
    ._EVAL_41(axi4buf__EVAL_41),
    ._EVAL_42(axi4buf__EVAL_42),
    ._EVAL_43(axi4buf__EVAL_43),
    ._EVAL_44(axi4buf__EVAL_44),
    ._EVAL_45(axi4buf__EVAL_45),
    ._EVAL_46(axi4buf__EVAL_46),
    ._EVAL_47(axi4buf__EVAL_47),
    ._EVAL_48(axi4buf__EVAL_48),
    ._EVAL_49(axi4buf__EVAL_49),
    ._EVAL_50(axi4buf__EVAL_50),
    ._EVAL_51(axi4buf__EVAL_51),
    ._EVAL_52(axi4buf__EVAL_52),
    ._EVAL_53(axi4buf__EVAL_53),
    ._EVAL_54(axi4buf__EVAL_54),
    ._EVAL_55(axi4buf__EVAL_55),
    ._EVAL_56(axi4buf__EVAL_56),
    ._EVAL_57(axi4buf__EVAL_57),
    ._EVAL_58(axi4buf__EVAL_58)
  );
  SiFive__EVAL_73 axi4frag (
    ._EVAL(axi4frag__EVAL),
    ._EVAL_0(axi4frag__EVAL_0),
    ._EVAL_1(axi4frag__EVAL_1),
    ._EVAL_2(axi4frag__EVAL_2),
    ._EVAL_3(axi4frag__EVAL_3),
    ._EVAL_4(axi4frag__EVAL_4),
    ._EVAL_5(axi4frag__EVAL_5),
    ._EVAL_6(axi4frag__EVAL_6),
    ._EVAL_7(axi4frag__EVAL_7),
    ._EVAL_8(axi4frag__EVAL_8),
    ._EVAL_9(axi4frag__EVAL_9),
    ._EVAL_10(axi4frag__EVAL_10),
    ._EVAL_11(axi4frag__EVAL_11),
    ._EVAL_12(axi4frag__EVAL_12),
    ._EVAL_13(axi4frag__EVAL_13),
    ._EVAL_14(axi4frag__EVAL_14),
    ._EVAL_15(axi4frag__EVAL_15),
    ._EVAL_16(axi4frag__EVAL_16),
    ._EVAL_17(axi4frag__EVAL_17),
    ._EVAL_18(axi4frag__EVAL_18),
    ._EVAL_19(axi4frag__EVAL_19),
    ._EVAL_20(axi4frag__EVAL_20),
    ._EVAL_21(axi4frag__EVAL_21),
    ._EVAL_22(axi4frag__EVAL_22),
    ._EVAL_23(axi4frag__EVAL_23),
    ._EVAL_24(axi4frag__EVAL_24),
    ._EVAL_25(axi4frag__EVAL_25),
    ._EVAL_26(axi4frag__EVAL_26),
    ._EVAL_27(axi4frag__EVAL_27),
    ._EVAL_28(axi4frag__EVAL_28),
    ._EVAL_29(axi4frag__EVAL_29),
    ._EVAL_30(axi4frag__EVAL_30),
    ._EVAL_31(axi4frag__EVAL_31),
    ._EVAL_32(axi4frag__EVAL_32),
    ._EVAL_33(axi4frag__EVAL_33),
    ._EVAL_34(axi4frag__EVAL_34),
    ._EVAL_35(axi4frag__EVAL_35),
    ._EVAL_36(axi4frag__EVAL_36),
    ._EVAL_37(axi4frag__EVAL_37),
    ._EVAL_38(axi4frag__EVAL_38),
    ._EVAL_39(axi4frag__EVAL_39),
    ._EVAL_40(axi4frag__EVAL_40),
    ._EVAL_41(axi4frag__EVAL_41),
    ._EVAL_42(axi4frag__EVAL_42),
    ._EVAL_43(axi4frag__EVAL_43),
    ._EVAL_44(axi4frag__EVAL_44),
    ._EVAL_45(axi4frag__EVAL_45),
    ._EVAL_46(axi4frag__EVAL_46),
    ._EVAL_47(axi4frag__EVAL_47),
    ._EVAL_48(axi4frag__EVAL_48),
    ._EVAL_49(axi4frag__EVAL_49),
    ._EVAL_50(axi4frag__EVAL_50),
    ._EVAL_51(axi4frag__EVAL_51),
    ._EVAL_52(axi4frag__EVAL_52),
    ._EVAL_53(axi4frag__EVAL_53),
    ._EVAL_54(axi4frag__EVAL_54),
    ._EVAL_55(axi4frag__EVAL_55),
    ._EVAL_56(axi4frag__EVAL_56),
    ._EVAL_57(axi4frag__EVAL_57),
    ._EVAL_58(axi4frag__EVAL_58),
    ._EVAL_59(axi4frag__EVAL_59),
    ._EVAL_60(axi4frag__EVAL_60),
    ._EVAL_61(axi4frag__EVAL_61),
    ._EVAL_62(axi4frag__EVAL_62),
    ._EVAL_63(axi4frag__EVAL_63),
    ._EVAL_64(axi4frag__EVAL_64)
  );
  SiFive__EVAL_64 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40)
  );
  SiFive__EVAL_74 axi4index (
    ._EVAL(axi4index__EVAL),
    ._EVAL_0(axi4index__EVAL_0),
    ._EVAL_1(axi4index__EVAL_1),
    ._EVAL_2(axi4index__EVAL_2),
    ._EVAL_3(axi4index__EVAL_3),
    ._EVAL_4(axi4index__EVAL_4),
    ._EVAL_5(axi4index__EVAL_5),
    ._EVAL_6(axi4index__EVAL_6),
    ._EVAL_7(axi4index__EVAL_7),
    ._EVAL_8(axi4index__EVAL_8),
    ._EVAL_9(axi4index__EVAL_9),
    ._EVAL_10(axi4index__EVAL_10),
    ._EVAL_11(axi4index__EVAL_11),
    ._EVAL_12(axi4index__EVAL_12),
    ._EVAL_13(axi4index__EVAL_13),
    ._EVAL_14(axi4index__EVAL_14),
    ._EVAL_15(axi4index__EVAL_15),
    ._EVAL_16(axi4index__EVAL_16),
    ._EVAL_17(axi4index__EVAL_17),
    ._EVAL_18(axi4index__EVAL_18),
    ._EVAL_19(axi4index__EVAL_19),
    ._EVAL_20(axi4index__EVAL_20),
    ._EVAL_21(axi4index__EVAL_21),
    ._EVAL_22(axi4index__EVAL_22),
    ._EVAL_23(axi4index__EVAL_23),
    ._EVAL_24(axi4index__EVAL_24),
    ._EVAL_25(axi4index__EVAL_25),
    ._EVAL_26(axi4index__EVAL_26),
    ._EVAL_27(axi4index__EVAL_27),
    ._EVAL_28(axi4index__EVAL_28),
    ._EVAL_29(axi4index__EVAL_29),
    ._EVAL_30(axi4index__EVAL_30),
    ._EVAL_31(axi4index__EVAL_31),
    ._EVAL_32(axi4index__EVAL_32),
    ._EVAL_33(axi4index__EVAL_33),
    ._EVAL_34(axi4index__EVAL_34),
    ._EVAL_35(axi4index__EVAL_35),
    ._EVAL_36(axi4index__EVAL_36),
    ._EVAL_37(axi4index__EVAL_37),
    ._EVAL_38(axi4index__EVAL_38),
    ._EVAL_39(axi4index__EVAL_39),
    ._EVAL_40(axi4index__EVAL_40),
    ._EVAL_41(axi4index__EVAL_41),
    ._EVAL_42(axi4index__EVAL_42),
    ._EVAL_43(axi4index__EVAL_43),
    ._EVAL_44(axi4index__EVAL_44),
    ._EVAL_45(axi4index__EVAL_45),
    ._EVAL_46(axi4index__EVAL_46),
    ._EVAL_47(axi4index__EVAL_47),
    ._EVAL_48(axi4index__EVAL_48),
    ._EVAL_49(axi4index__EVAL_49),
    ._EVAL_50(axi4index__EVAL_50),
    ._EVAL_51(axi4index__EVAL_51),
    ._EVAL_52(axi4index__EVAL_52),
    ._EVAL_53(axi4index__EVAL_53),
    ._EVAL_54(axi4index__EVAL_54),
    ._EVAL_55(axi4index__EVAL_55),
    ._EVAL_56(axi4index__EVAL_56),
    ._EVAL_57(axi4index__EVAL_57),
    ._EVAL_58(axi4index__EVAL_58),
    ._EVAL_59(axi4index__EVAL_59),
    ._EVAL_60(axi4index__EVAL_60)
  );
  SiFive__EVAL_66 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36),
    ._EVAL_37(widget__EVAL_37),
    ._EVAL_38(widget__EVAL_38)
  );
  assign axi42tl__EVAL_16 = axi4yank__EVAL_35;
  assign _EVAL = axi4buf__EVAL_56;
  assign axi4buf__EVAL_51 = _EVAL_26;
  assign axi4index__EVAL_38 = axi4frag__EVAL_41;
  assign buffer__EVAL_1 = fixer__EVAL_3;
  assign _EVAL_41 = buffer__EVAL_33;
  assign axi4buf__EVAL_45 = _EVAL_10;
  assign axi4frag__EVAL_7 = axi4index__EVAL_57;
  assign axi4index__EVAL_52 = axi4frag__EVAL_61;
  assign axi4yank__EVAL_16 = axi4frag__EVAL_14;
  assign axi4yank__EVAL_7 = axi4frag__EVAL_10;
  assign widget__EVAL_9 = _EVAL_6;
  assign axi4index__EVAL_18 = axi4frag__EVAL_46;
  assign buffer__EVAL_40 = _EVAL_36;
  assign axi4frag__EVAL_57 = axi4index__EVAL_41;
  assign axi4buf__EVAL_34 = _EVAL_11;
  assign fixer__EVAL_17 = widget__EVAL_30;
  assign fixer__EVAL_15 = widget__EVAL_0;
  assign axi42tl__EVAL_5 = axi4yank__EVAL_32;
  assign axi4index__EVAL_20 = axi4buf__EVAL_35;
  assign axi42tl__EVAL_26 = axi4yank__EVAL_2;
  assign widget__EVAL_10 = fixer__EVAL_24;
  assign axi42tl__EVAL_13 = widget__EVAL_22;
  assign axi4frag__EVAL_53 = axi4index__EVAL_25;
  assign axi4index__EVAL_6 = axi4buf__EVAL_18;
  assign fixer__EVAL_0 = widget__EVAL_6;
  assign axi4buf__EVAL_14 = _EVAL_3;
  assign buffer__EVAL_25 = _EVAL_44;
  assign axi4index__EVAL_27 = axi4frag__EVAL_23;
  assign axi4index__EVAL_17 = axi4buf__EVAL_2;
  assign axi4frag__EVAL_26 = _EVAL_19;
  assign axi4yank__EVAL_6 = _EVAL_19;
  assign _EVAL_49 = axi4buf__EVAL_37;
  assign axi4buf__EVAL_43 = axi4index__EVAL_1;
  assign axi42tl__EVAL_15 = axi4yank__EVAL_15;
  assign axi42tl__EVAL_38 = widget__EVAL_16;
  assign axi4yank__EVAL_46 = axi42tl__EVAL;
  assign axi4buf__EVAL_40 = _EVAL_15;
  assign axi4yank__EVAL_27 = axi42tl__EVAL_41;
  assign fixer__EVAL_12 = widget__EVAL_24;
  assign axi4buf__EVAL_7 = _EVAL_29;
  assign fixer__EVAL_5 = buffer__EVAL_14;
  assign _EVAL_9 = buffer__EVAL_3;
  assign fixer__EVAL_38 = widget__EVAL_19;
  assign axi4index__EVAL_33 = axi4frag__EVAL_52;
  assign axi4frag__EVAL_58 = axi4index__EVAL_45;
  assign axi4buf__EVAL_3 = axi4index__EVAL_9;
  assign axi4index__EVAL_24 = axi4buf__EVAL_52;
  assign axi4yank__EVAL_24 = axi42tl__EVAL_45;
  assign axi4yank__EVAL_23 = axi4frag__EVAL_0;
  assign widget__EVAL_29 = fixer__EVAL;
  assign axi4yank__EVAL_1 = axi4frag__EVAL_37;
  assign axi42tl__EVAL_0 = widget__EVAL_23;
  assign fixer__EVAL_28 = _EVAL_6;
  assign axi4frag__EVAL_51 = axi4yank__EVAL_52;
  assign axi4buf__EVAL_39 = _EVAL_20;
  assign _EVAL_7 = buffer__EVAL_11;
  assign axi4yank__EVAL_31 = axi4frag__EVAL_56;
  assign widget__EVAL_33 = fixer__EVAL_35;
  assign axi4frag__EVAL_59 = axi4index__EVAL_13;
  assign axi4index__EVAL_15 = axi4buf__EVAL_50;
  assign fixer__EVAL_20 = widget__EVAL_25;
  assign axi4frag__EVAL_45 = axi4index__EVAL_5;
  assign axi4index__EVAL_8 = axi4buf__EVAL_24;
  assign _EVAL_18 = buffer__EVAL_18;
  assign axi4frag__EVAL_43 = axi4yank__EVAL_58;
  assign axi42tl__EVAL_28 = _EVAL_19;
  assign axi4index__EVAL_53 = axi4buf__EVAL_41;
  assign axi4yank__EVAL_43 = axi42tl__EVAL_10;
  assign buffer__EVAL_9 = _EVAL_5;
  assign buffer__EVAL_23 = fixer__EVAL_36;
  assign axi4buf__EVAL_49 = axi4index__EVAL_60;
  assign axi4frag__EVAL_25 = axi4index__EVAL_44;
  assign widget__EVAL_34 = axi42tl__EVAL_29;
  assign _EVAL_17 = axi4buf__EVAL_11;
  assign buffer__EVAL_26 = _EVAL_35;
  assign fixer__EVAL_32 = widget__EVAL_37;
  assign axi4buf__EVAL_0 = axi4index__EVAL_48;
  assign axi4frag__EVAL_18 = axi4index__EVAL_39;
  assign axi4index__EVAL_58 = axi4frag__EVAL_29;
  assign buffer__EVAL = fixer__EVAL_37;
  assign buffer__EVAL_32 = fixer__EVAL_14;
  assign axi4yank__EVAL_21 = axi4frag__EVAL_50;
  assign axi4buf__EVAL_54 = _EVAL_23;
  assign _EVAL_46 = axi4buf__EVAL_13;
  assign axi4index__EVAL_26 = axi4frag__EVAL_35;
  assign axi42tl__EVAL_12 = axi4yank__EVAL_50;
  assign axi4buf__EVAL_12 = _EVAL_1;
  assign axi42tl__EVAL_23 = axi4yank__EVAL_22;
  assign fixer__EVAL_40 = buffer__EVAL_17;
  assign axi4frag__EVAL_22 = axi4index__EVAL_59;
  assign fixer__EVAL_7 = buffer__EVAL_21;
  assign widget__EVAL_21 = axi42tl__EVAL_8;
  assign axi4frag__EVAL_28 = axi4yank__EVAL_11;
  assign axi4buf__EVAL_42 = _EVAL_14;
  assign fixer__EVAL_11 = buffer__EVAL_6;
  assign fixer__EVAL_23 = buffer__EVAL_8;
  assign axi4index__EVAL_22 = axi4buf__EVAL_55;
  assign axi4yank__EVAL_5 = axi4frag__EVAL_4;
  assign axi4yank__EVAL_12 = axi4frag__EVAL_42;
  assign fixer__EVAL_21 = _EVAL_19;
  assign axi4index__EVAL_37 = axi4buf__EVAL_21;
  assign axi4yank__EVAL_0 = axi42tl__EVAL_34;
  assign fixer__EVAL_2 = buffer__EVAL_30;
  assign axi4frag__EVAL_54 = axi4yank__EVAL_53;
  assign widget__EVAL_17 = axi42tl__EVAL_27;
  assign _EVAL_45 = buffer__EVAL_39;
  assign axi4index__EVAL_7 = axi4frag__EVAL_13;
  assign fixer__EVAL_31 = buffer__EVAL_36;
  assign axi42tl__EVAL_6 = widget__EVAL_5;
  assign axi42tl__EVAL_33 = axi4yank__EVAL_41;
  assign buffer__EVAL_7 = _EVAL_6;
  assign axi4buf__EVAL_27 = axi4index__EVAL_43;
  assign axi4yank__EVAL_39 = axi4frag__EVAL_12;
  assign axi4index__EVAL_28 = axi4buf__EVAL_4;
  assign _EVAL_31 = buffer__EVAL_31;
  assign axi4index__EVAL_54 = axi4frag__EVAL_16;
  assign buffer__EVAL_4 = fixer__EVAL_4;
  assign axi4frag__EVAL_63 = axi4yank__EVAL_51;
  assign _EVAL_13 = axi4buf__EVAL_19;
  assign axi4buf__EVAL_29 = axi4index__EVAL_21;
  assign axi4buf__EVAL_16 = _EVAL_4;
  assign axi42tl__EVAL_22 = axi4yank__EVAL_47;
  assign axi42tl__EVAL_32 = widget__EVAL_27;
  assign axi4buf__EVAL_25 = axi4index__EVAL_31;
  assign widget__EVAL_35 = axi42tl__EVAL_18;
  assign axi4frag__EVAL_31 = axi4index__EVAL_19;
  assign axi4frag__EVAL_17 = axi4index__EVAL_0;
  assign _EVAL_21 = axi4buf__EVAL_47;
  assign axi4frag__EVAL_27 = axi4index__EVAL;
  assign _EVAL_32 = axi4buf__EVAL_48;
  assign axi4buf__EVAL_36 = _EVAL_24;
  assign axi4yank__EVAL_37 = axi42tl__EVAL_39;
  assign axi4index__EVAL_32 = axi4buf__EVAL_58;
  assign widget__EVAL_4 = fixer__EVAL_29;
  assign axi4yank__EVAL_48 = axi4frag__EVAL_44;
  assign buffer__EVAL_38 = fixer__EVAL_22;
  assign axi42tl__EVAL_36 = widget__EVAL_3;
  assign buffer__EVAL_29 = fixer__EVAL_19;
  assign axi4frag__EVAL_47 = axi4yank__EVAL_33;
  assign axi4yank__EVAL_14 = axi42tl__EVAL_21;
  assign axi4buf__EVAL_32 = _EVAL_19;
  assign widget__EVAL_14 = fixer__EVAL_10;
  assign fixer__EVAL_1 = buffer__EVAL_2;
  assign axi4frag__EVAL_8 = axi4yank__EVAL_30;
  assign axi4buf__EVAL_44 = axi4index__EVAL_55;
  assign axi4index__EVAL_34 = axi4buf__EVAL_28;
  assign axi4frag__EVAL_5 = axi4yank__EVAL_45;
  assign buffer__EVAL_10 = fixer__EVAL_6;
  assign axi42tl__EVAL_35 = axi4yank__EVAL_49;
  assign widget__EVAL_11 = fixer__EVAL_25;
  assign widget__EVAL_38 = axi42tl__EVAL_9;
  assign axi4buf__EVAL_20 = axi4index__EVAL_30;
  assign fixer__EVAL_8 = widget__EVAL_32;
  assign axi4index__EVAL_47 = axi4frag__EVAL_33;
  assign _EVAL_33 = buffer__EVAL_5;
  assign _EVAL_40 = axi4buf__EVAL_57;
  assign fixer__EVAL_39 = widget__EVAL_18;
  assign fixer__EVAL_13 = widget__EVAL_7;
  assign widget__EVAL_2 = _EVAL_19;
  assign axi4index__EVAL_10 = axi4frag__EVAL_15;
  assign axi4frag__EVAL_49 = axi4yank__EVAL_26;
  assign axi4index__EVAL_11 = axi4buf__EVAL_53;
  assign axi42tl__EVAL_1 = widget__EVAL_12;
  assign _EVAL_8 = axi4buf__EVAL;
  assign axi4buf__EVAL_5 = _EVAL_34;
  assign buffer__EVAL_34 = fixer__EVAL_26;
  assign axi4frag__EVAL_38 = axi4yank__EVAL_25;
  assign axi4yank__EVAL_56 = axi4frag__EVAL_40;
  assign axi42tl__EVAL_3 = axi4yank__EVAL_4;
  assign axi4frag__EVAL_9 = axi4index__EVAL_46;
  assign widget__EVAL_15 = fixer__EVAL_16;
  assign axi4buf__EVAL_46 = axi4index__EVAL_12;
  assign axi4yank__EVAL_54 = axi4frag__EVAL_32;
  assign _EVAL_0 = buffer__EVAL_0;
  assign widget__EVAL = fixer__EVAL_18;
  assign axi4index__EVAL_42 = axi4frag__EVAL;
  assign buffer__EVAL_35 = _EVAL_25;
  assign axi4buf__EVAL_1 = _EVAL_30;
  assign axi42tl__EVAL_44 = axi4yank__EVAL_13;
  assign axi4frag__EVAL_36 = axi4yank__EVAL_10;
  assign axi4index__EVAL_23 = axi4buf__EVAL_17;
  assign buffer__EVAL_16 = _EVAL_47;
  assign _EVAL_42 = axi4buf__EVAL_8;
  assign _EVAL_2 = buffer__EVAL_13;
  assign axi42tl__EVAL_30 = widget__EVAL_31;
  assign fixer__EVAL_30 = buffer__EVAL_12;
  assign axi4frag__EVAL_11 = axi4index__EVAL_40;
  assign buffer__EVAL_27 = _EVAL_22;
  assign buffer__EVAL_24 = _EVAL_37;
  assign axi4buf__EVAL_33 = _EVAL_6;
  assign axi4frag__EVAL_6 = axi4index__EVAL_56;
  assign buffer__EVAL_19 = _EVAL_27;
  assign axi4yank__EVAL_44 = axi4frag__EVAL_2;
  assign axi42tl__EVAL_4 = axi4yank__EVAL_36;
  assign axi42tl__EVAL_25 = axi4yank__EVAL_57;
  assign axi4yank__EVAL = axi42tl__EVAL_19;
  assign buffer__EVAL_15 = _EVAL_39;
  assign axi4yank__EVAL_9 = axi42tl__EVAL_17;
  assign axi4frag__EVAL_1 = _EVAL_6;
  assign buffer__EVAL_20 = fixer__EVAL_27;
  assign axi4index__EVAL_29 = axi4buf__EVAL_38;
  assign axi4frag__EVAL_39 = axi4yank__EVAL_34;
  assign axi4index__EVAL_14 = axi4buf__EVAL_23;
  assign axi4yank__EVAL_17 = axi4frag__EVAL_48;
  assign axi4yank__EVAL_28 = axi4frag__EVAL_3;
  assign widget__EVAL_26 = axi42tl__EVAL_40;
  assign axi4frag__EVAL_62 = axi4index__EVAL_50;
  assign axi4index__EVAL_36 = axi4buf__EVAL_30;
  assign axi4index__EVAL_49 = axi4frag__EVAL_55;
  assign axi4buf__EVAL_31 = _EVAL_12;
  assign axi4yank__EVAL_40 = _EVAL_6;
  assign axi4frag__EVAL_60 = axi4yank__EVAL_18;
  assign axi42tl__EVAL_2 = axi4yank__EVAL_42;
  assign axi4index__EVAL_35 = axi4buf__EVAL_26;
  assign axi4buf__EVAL_10 = _EVAL_43;
  assign axi4yank__EVAL_19 = axi4frag__EVAL_34;
  assign axi4buf__EVAL_6 = _EVAL_28;
  assign widget__EVAL_20 = axi42tl__EVAL_31;
  assign axi4frag__EVAL_30 = axi4index__EVAL_16;
  assign widget__EVAL_28 = axi42tl__EVAL_20;
  assign widget__EVAL_36 = axi42tl__EVAL_7;
  assign axi4buf__EVAL_9 = axi4index__EVAL_51;
  assign widget__EVAL_13 = fixer__EVAL_34;
  assign axi4frag__EVAL_24 = axi4index__EVAL_2;
  assign axi4yank__EVAL_20 = axi4frag__EVAL_21;
  assign axi42tl__EVAL_11 = axi4yank__EVAL_29;
  assign axi4yank__EVAL_38 = axi42tl__EVAL_37;
  assign axi4buf__EVAL_22 = _EVAL_16;
  assign axi4frag__EVAL_20 = axi4index__EVAL_3;
  assign axi4yank__EVAL_55 = axi42tl__EVAL_43;
  assign axi42tl__EVAL_24 = _EVAL_6;
  assign axi42tl__EVAL_42 = axi4yank__EVAL_8;
  assign _EVAL_48 = axi4buf__EVAL_15;
  assign widget__EVAL_1 = fixer__EVAL_9;
  assign fixer__EVAL_33 = buffer__EVAL_22;
  assign axi4frag__EVAL_64 = axi4index__EVAL_4;
  assign buffer__EVAL_28 = _EVAL_19;
  assign _EVAL_38 = buffer__EVAL_37;
  assign widget__EVAL_8 = axi42tl__EVAL_14;
  assign axi4yank__EVAL_3 = axi4frag__EVAL_19;
endmodule
