//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_174_assert(
  input         _EVAL,
  input  [29:0] _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [6:0]  _EVAL_12,
  input  [6:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_24;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_46;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_99;
  reg [31:0] _RAND_2;
  reg [6:0] _EVAL_118;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_128;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_155;
  reg [31:0] _RAND_5;
  reg [3:0] _EVAL_163;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_179;
  reg [31:0] _RAND_7;
  reg [29:0] _EVAL_216;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_226;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_237;
  reg [31:0] _RAND_10;
  reg [72:0] _EVAL_239;
  reg [95:0] _RAND_11;
  reg [2:0] _EVAL_253;
  reg [31:0] _RAND_12;
  reg [6:0] _EVAL_270;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_285;
  reg [31:0] _RAND_14;
  wire  _EVAL_166;
  wire  _EVAL_188;
  wire  _EVAL_211;
  wire  _EVAL_194;
  wire  _EVAL_159;
  wire  _EVAL_44;
  wire [127:0] _EVAL_141;
  wire [127:0] _EVAL_100;
  wire [72:0] _EVAL_150;
  wire [72:0] _EVAL_203;
  wire [72:0] _EVAL_41;
  wire  _EVAL_262;
  wire  _EVAL_149;
  wire  _EVAL_39;
  wire  _EVAL_299;
  wire  _EVAL_151;
  wire  _EVAL_233;
  wire [29:0] _EVAL_293;
  wire [30:0] _EVAL_225;
  wire [30:0] _EVAL_196;
  wire  _EVAL_279;
  wire  _EVAL_199;
  wire  _EVAL_80;
  wire [127:0] _EVAL_84;
  wire [127:0] _EVAL_89;
  wire [72:0] _EVAL_114;
  wire  _EVAL_142;
  wire  _EVAL_55;
  wire  _EVAL_22;
  wire  _EVAL_186;
  wire  _EVAL_124;
  wire [3:0] _EVAL_221;
  wire  _EVAL_300;
  wire  _EVAL_204;
  wire [3:0] _EVAL_231;
  wire  _EVAL_206;
  wire  _EVAL_254;
  wire  _EVAL_174;
  wire  _EVAL_284;
  wire [72:0] _EVAL_290;
  wire [72:0] _EVAL_127;
  wire  _EVAL_79;
  wire  _EVAL_20;
  wire  _EVAL_286;
  wire  _EVAL_120;
  wire  _EVAL_227;
  wire [12:0] _EVAL_103;
  wire [5:0] _EVAL_244;
  wire [5:0] _EVAL_201;
  wire [3:0] _EVAL_191;
  wire [3:0] _EVAL_220;
  wire  _EVAL_21;
  wire [2:0] _EVAL_182;
  wire  _EVAL_154;
  wire  _EVAL_148;
  wire  _EVAL_27;
  wire  _EVAL_77;
  wire  _EVAL_278;
  wire  _EVAL_125;
  wire  _EVAL_82;
  wire  _EVAL_205;
  wire  _EVAL_222;
  wire  _EVAL_268;
  wire  _EVAL_298;
  wire  _EVAL_133;
  wire  _EVAL_71;
  wire [3:0] _EVAL_250;
  wire  _EVAL_289;
  wire  _EVAL_60;
  wire [1:0] _EVAL_97;
  wire [1:0] _EVAL_109;
  wire  _EVAL_245;
  wire [3:0] _EVAL_73;
  wire  _EVAL_116;
  wire  _EVAL_247;
  wire  _EVAL_224;
  wire  _EVAL_145;
  wire  _EVAL_292;
  wire  _EVAL_183;
  wire  _EVAL_94;
  wire  _EVAL_192;
  wire  _EVAL_132;
  wire  _EVAL_294;
  wire  _EVAL_126;
  wire  _EVAL_58;
  wire [12:0] _EVAL_144;
  wire  _EVAL_202;
  wire [30:0] _EVAL_110;
  wire  _EVAL_235;
  wire  _EVAL_53;
  wire  _EVAL_184;
  wire  _EVAL_62;
  wire  _EVAL_158;
  wire  _EVAL_261;
  wire  _EVAL_181;
  wire  _EVAL_189;
  wire  _EVAL_123;
  wire [2:0] _EVAL_217;
  wire  _EVAL_91;
  wire  _EVAL_280;
  wire  _EVAL_56;
  wire  _EVAL_63;
  wire  _EVAL_161;
  wire  _EVAL_87;
  wire  _EVAL_302;
  wire  _EVAL_136;
  wire  _EVAL_162;
  wire  _EVAL_295;
  wire  _EVAL_98;
  wire  _EVAL_287;
  wire  _EVAL_83;
  wire  _EVAL_122;
  wire  _EVAL_76;
  wire  _EVAL_42;
  wire  _EVAL_156;
  wire  _EVAL_236;
  wire  _EVAL_119;
  wire  _EVAL_113;
  wire  _EVAL_92;
  wire  _EVAL_112;
  wire  _EVAL_215;
  wire  _EVAL_240;
  wire  _EVAL_93;
  wire  _EVAL_303;
  wire  _EVAL_105;
  wire  _EVAL_212;
  wire  _EVAL_272;
  wire  _EVAL_180;
  wire  _EVAL_219;
  wire  _EVAL_18;
  wire  _EVAL_177;
  wire [3:0] _EVAL_283;
  wire [3:0] _EVAL_130;
  wire [3:0] _EVAL_255;
  wire  _EVAL_96;
  wire  _EVAL_230;
  wire  _EVAL_57;
  wire  _EVAL_241;
  wire  _EVAL_195;
  wire  _EVAL_198;
  wire  _EVAL_274;
  wire  _EVAL_264;
  wire  _EVAL_101;
  wire  _EVAL_117;
  wire  _EVAL_228;
  wire  _EVAL_61;
  wire  _EVAL_175;
  wire [72:0] _EVAL_115;
  wire [72:0] _EVAL_121;
  wire  _EVAL_54;
  wire  _EVAL_267;
  wire [5:0] _EVAL_246;
  wire [5:0] _EVAL_157;
  wire [3:0] _EVAL_281;
  wire  _EVAL_17;
  wire  _EVAL_51;
  wire  _EVAL_95;
  wire  _EVAL_29;
  wire  _EVAL_165;
  wire  _EVAL_47;
  wire  _EVAL_31;
  wire  _EVAL_200;
  wire  _EVAL_23;
  wire  _EVAL_172;
  wire  _EVAL_36;
  wire  _EVAL_288;
  wire  _EVAL_170;
  wire  _EVAL_249;
  wire  _EVAL_131;
  wire  _EVAL_187;
  wire  _EVAL_242;
  wire  _EVAL_258;
  wire  _EVAL_64;
  wire  _EVAL_104;
  wire [29:0] _EVAL_271;
  wire [29:0] _EVAL_213;
  wire  _EVAL_173;
  wire  _EVAL_291;
  wire  _EVAL_190;
  wire  _EVAL_296;
  wire  _EVAL_30;
  wire  _EVAL_108;
  wire  _EVAL_164;
  wire  _EVAL_210;
  wire [31:0] _EVAL_223;
  wire  _EVAL_297;
  wire  _EVAL_214;
  wire  _EVAL_35;
  wire  _EVAL_33;
  wire  _EVAL_111;
  wire  _EVAL_38;
  wire  _EVAL_59;
  wire  _EVAL_171;
  wire  _EVAL_234;
  wire  _EVAL_207;
  wire [3:0] _EVAL_45;
  wire  _EVAL_65;
  wire  _EVAL_160;
  wire  _EVAL_74;
  wire  _EVAL_185;
  wire  _EVAL_140;
  wire  _EVAL_106;
  wire  _EVAL_134;
  wire  _EVAL_107;
  wire  _EVAL_88;
  wire [3:0] _EVAL_229;
  wire  _EVAL_138;
  wire  _EVAL_143;
  wire  _EVAL_256;
  wire  _EVAL_273;
  wire  _EVAL_168;
  wire  _EVAL_49;
  wire  _EVAL_266;
  wire  _EVAL_218;
  wire  _EVAL_251;
  wire  _EVAL_238;
  wire  _EVAL_197;
  wire  _EVAL_129;
  wire  _EVAL_167;
  wire  _EVAL_48;
  wire  _EVAL_260;
  wire  _EVAL_81;
  wire  _EVAL_50;
  wire  _EVAL_169;
  wire  _EVAL_248;
  wire  _EVAL_176;
  wire  _EVAL_243;
  wire  _EVAL_277;
  wire  _EVAL_68;
  wire  _EVAL_252;
  wire  _EVAL_86;
  wire  _EVAL_37;
  wire  _EVAL_139;
  wire  _EVAL_208;
  wire  _EVAL_52;
  wire  _EVAL_28;
  wire  _EVAL_85;
  wire  _EVAL_232;
  wire  _EVAL_102;
  wire  _EVAL_34;
  wire  _EVAL_301;
  wire  _EVAL_25;
  wire  _EVAL_70;
  wire  _EVAL_259;
  wire  _EVAL_69;
  wire  _EVAL_193;
  wire  _EVAL_265;
  wire  _EVAL_282;
  wire  _EVAL_178;
  wire  _EVAL_26;
  wire  _EVAL_66;
  wire  _EVAL_257;
  wire  _EVAL_152;
  wire  _EVAL_209;
  wire  _EVAL_275;
  wire  _EVAL_40;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_166 = _EVAL_16 & _EVAL_11;
  assign _EVAL_188 = _EVAL_128 == 4'h0;
  assign _EVAL_211 = _EVAL_166 & _EVAL_188;
  assign _EVAL_194 = _EVAL_3 == 3'h6;
  assign _EVAL_159 = _EVAL_194 == 1'h0;
  assign _EVAL_44 = _EVAL_211 & _EVAL_159;
  assign _EVAL_141 = 128'h1 << _EVAL_13;
  assign _EVAL_100 = _EVAL_44 ? _EVAL_141 : 128'h0;
  assign _EVAL_150 = _EVAL_100[72:0];
  assign _EVAL_203 = ~ _EVAL_150;
  assign _EVAL_41 = _EVAL_239 >> _EVAL_12;
  assign _EVAL_262 = _EVAL_41[0];
  assign _EVAL_149 = _EVAL_262 == 1'h0;
  assign _EVAL_39 = _EVAL_149 | _EVAL;
  assign _EVAL_299 = _EVAL_39 == 1'h0;
  assign _EVAL_151 = _EVAL_163 == 4'h0;
  assign _EVAL_233 = _EVAL_151 == 1'h0;
  assign _EVAL_293 = _EVAL_0 ^ 30'h20000000;
  assign _EVAL_225 = {1'b0,$signed(_EVAL_293)};
  assign _EVAL_196 = $signed(_EVAL_225) & $signed(-31'sh2000);
  assign _EVAL_279 = _EVAL_14 & _EVAL_8;
  assign _EVAL_199 = _EVAL_99 == 4'h0;
  assign _EVAL_80 = _EVAL_279 & _EVAL_199;
  assign _EVAL_84 = 128'h1 << _EVAL_12;
  assign _EVAL_89 = _EVAL_80 ? _EVAL_84 : 128'h0;
  assign _EVAL_114 = _EVAL_89[72:0];
  assign _EVAL_142 = _EVAL_114 != _EVAL_150;
  assign _EVAL_55 = _EVAL_114 != 73'h0;
  assign _EVAL_22 = _EVAL_55 == 1'h0;
  assign _EVAL_186 = _EVAL_142 | _EVAL_22;
  assign _EVAL_124 = _EVAL_12 == 7'h48;
  assign _EVAL_221 = _EVAL_163 - 4'h1;
  assign _EVAL_300 = _EVAL_15 == 1'h0;
  assign _EVAL_204 = _EVAL_300 | _EVAL_7;
  assign _EVAL_231 = _EVAL_99 - 4'h1;
  assign _EVAL_206 = _EVAL_6 == _EVAL_46;
  assign _EVAL_254 = _EVAL_206 | _EVAL;
  assign _EVAL_174 = _EVAL_254 == 1'h0;
  assign _EVAL_284 = _EVAL_4 <= 3'h3;
  assign _EVAL_290 = _EVAL_114 | _EVAL_239;
  assign _EVAL_127 = _EVAL_290 >> _EVAL_13;
  assign _EVAL_79 = _EVAL_127[0];
  assign _EVAL_20 = _EVAL_79 | _EVAL;
  assign _EVAL_286 = _EVAL_20 == 1'h0;
  assign _EVAL_120 = _EVAL_3 == 3'h1;
  assign _EVAL_227 = _EVAL_3[0];
  assign _EVAL_103 = 13'h3f << _EVAL_5;
  assign _EVAL_244 = _EVAL_103[5:0];
  assign _EVAL_201 = ~ _EVAL_244;
  assign _EVAL_191 = _EVAL_201[5:2];
  assign _EVAL_220 = _EVAL_13[6:3];
  assign _EVAL_21 = _EVAL_220 == 4'h8;
  assign _EVAL_182 = _EVAL_13[2:0];
  assign _EVAL_154 = 3'h1 <= _EVAL_182;
  assign _EVAL_148 = _EVAL_21 & _EVAL_154;
  assign _EVAL_27 = _EVAL_0[1];
  assign _EVAL_77 = _EVAL_239 != 73'h0;
  assign _EVAL_278 = _EVAL_77 == 1'h0;
  assign _EVAL_125 = plusarg_reader_out == 32'h0;
  assign _EVAL_82 = _EVAL_278 | _EVAL_125;
  assign _EVAL_205 = _EVAL_179 < plusarg_reader_out;
  assign _EVAL_222 = _EVAL_82 | _EVAL_205;
  assign _EVAL_268 = _EVAL_222 | _EVAL;
  assign _EVAL_298 = _EVAL_268 == 1'h0;
  assign _EVAL_133 = _EVAL_5 == _EVAL_253;
  assign _EVAL_71 = _EVAL_133 | _EVAL;
  assign _EVAL_250 = _EVAL_12[6:3];
  assign _EVAL_289 = _EVAL_250 == 4'h3;
  assign _EVAL_60 = _EVAL_1[0];
  assign _EVAL_97 = 2'h1 << _EVAL_60;
  assign _EVAL_109 = _EVAL_97 | 2'h1;
  assign _EVAL_245 = _EVAL_109[1];
  assign _EVAL_73 = ~ _EVAL_9;
  assign _EVAL_116 = _EVAL_73 == 4'h0;
  assign _EVAL_247 = _EVAL_116 | _EVAL;
  assign _EVAL_224 = _EVAL_247 == 1'h0;
  assign _EVAL_145 = _EVAL_300 | _EVAL;
  assign _EVAL_292 = _EVAL_145 == 1'h0;
  assign _EVAL_183 = _EVAL_204 | _EVAL;
  assign _EVAL_94 = _EVAL_183 == 1'h0;
  assign _EVAL_192 = _EVAL_12 == _EVAL_118;
  assign _EVAL_132 = _EVAL_109[0];
  assign _EVAL_294 = _EVAL_0[0];
  assign _EVAL_126 = _EVAL_27 & _EVAL_294;
  assign _EVAL_58 = _EVAL_132 & _EVAL_126;
  assign _EVAL_144 = 13'h3f << _EVAL_1;
  assign _EVAL_202 = _EVAL_1 <= 3'h6;
  assign _EVAL_110 = $signed(_EVAL_196);
  assign _EVAL_235 = $signed(_EVAL_110) == $signed(31'sh0);
  assign _EVAL_53 = _EVAL_202 & _EVAL_235;
  assign _EVAL_184 = _EVAL_53 | _EVAL;
  assign _EVAL_62 = _EVAL_184 == 1'h0;
  assign _EVAL_158 = _EVAL_3 == 3'h4;
  assign _EVAL_261 = _EVAL_11 & _EVAL_158;
  assign _EVAL_181 = _EVAL_220 == 4'h0;
  assign _EVAL_189 = _EVAL_12 == 7'h20;
  assign _EVAL_123 = _EVAL_6 == 3'h4;
  assign _EVAL_217 = _EVAL_12[2:0];
  assign _EVAL_91 = 3'h1 <= _EVAL_217;
  assign _EVAL_280 = _EVAL_13 == 7'h48;
  assign _EVAL_56 = _EVAL_13 == 7'h40;
  assign _EVAL_63 = _EVAL_280 | _EVAL_56;
  assign _EVAL_161 = _EVAL_63 | _EVAL_148;
  assign _EVAL_87 = _EVAL_13 == 7'h20;
  assign _EVAL_302 = _EVAL_161 | _EVAL_87;
  assign _EVAL_136 = _EVAL_302 | _EVAL_181;
  assign _EVAL_162 = _EVAL_220 == 4'h1;
  assign _EVAL_295 = _EVAL_136 | _EVAL_162;
  assign _EVAL_98 = _EVAL_220 == 4'h2;
  assign _EVAL_287 = _EVAL_295 | _EVAL_98;
  assign _EVAL_83 = _EVAL_220 == 4'h3;
  assign _EVAL_122 = _EVAL_287 | _EVAL_83;
  assign _EVAL_76 = _EVAL_122 | _EVAL;
  assign _EVAL_42 = _EVAL_76 == 1'h0;
  assign _EVAL_156 = _EVAL_1 >= 3'h2;
  assign _EVAL_236 = _EVAL_245 & _EVAL_27;
  assign _EVAL_119 = _EVAL_156 | _EVAL_236;
  assign _EVAL_113 = _EVAL_119 | _EVAL_58;
  assign _EVAL_92 = _EVAL_294 == 1'h0;
  assign _EVAL_112 = _EVAL_27 & _EVAL_92;
  assign _EVAL_215 = _EVAL_132 & _EVAL_112;
  assign _EVAL_240 = _EVAL_119 | _EVAL_215;
  assign _EVAL_93 = _EVAL_27 == 1'h0;
  assign _EVAL_303 = _EVAL_245 & _EVAL_93;
  assign _EVAL_105 = _EVAL_156 | _EVAL_303;
  assign _EVAL_212 = _EVAL_93 & _EVAL_294;
  assign _EVAL_272 = _EVAL_132 & _EVAL_212;
  assign _EVAL_180 = _EVAL_105 | _EVAL_272;
  assign _EVAL_219 = _EVAL_93 & _EVAL_92;
  assign _EVAL_18 = _EVAL_132 & _EVAL_219;
  assign _EVAL_177 = _EVAL_105 | _EVAL_18;
  assign _EVAL_283 = {_EVAL_113,_EVAL_240,_EVAL_180,_EVAL_177};
  assign _EVAL_130 = ~ _EVAL_283;
  assign _EVAL_255 = _EVAL_9 & _EVAL_130;
  assign _EVAL_96 = _EVAL_255 == 4'h0;
  assign _EVAL_230 = _EVAL_96 | _EVAL;
  assign _EVAL_57 = _EVAL_284 | _EVAL;
  assign _EVAL_241 = _EVAL_4 <= 3'h4;
  assign _EVAL_195 = _EVAL_241 | _EVAL;
  assign _EVAL_198 = _EVAL_4 == _EVAL_285;
  assign _EVAL_274 = _EVAL_198 | _EVAL;
  assign _EVAL_264 = _EVAL_9 == _EVAL_283;
  assign _EVAL_101 = _EVAL_264 | _EVAL;
  assign _EVAL_117 = _EVAL_101 == 1'h0;
  assign _EVAL_228 = _EVAL_250 == 4'h8;
  assign _EVAL_61 = _EVAL_10 == 1'h0;
  assign _EVAL_175 = _EVAL_61 | _EVAL;
  assign _EVAL_115 = _EVAL_239 | _EVAL_114;
  assign _EVAL_121 = _EVAL_115 & _EVAL_203;
  assign _EVAL_54 = _EVAL_6[2];
  assign _EVAL_267 = _EVAL_54 == 1'h0;
  assign _EVAL_246 = _EVAL_144[5:0];
  assign _EVAL_157 = ~ _EVAL_246;
  assign _EVAL_281 = _EVAL_157[5:2];
  assign _EVAL_17 = _EVAL == 1'h0;
  assign _EVAL_51 = _EVAL_0 == _EVAL_216;
  assign _EVAL_95 = _EVAL_12 == 7'h40;
  assign _EVAL_29 = _EVAL_124 | _EVAL_95;
  assign _EVAL_165 = _EVAL_228 & _EVAL_91;
  assign _EVAL_47 = _EVAL_29 | _EVAL_165;
  assign _EVAL_31 = _EVAL_47 | _EVAL_189;
  assign _EVAL_200 = _EVAL_250 == 4'h0;
  assign _EVAL_23 = _EVAL_31 | _EVAL_200;
  assign _EVAL_172 = _EVAL_250 == 4'h1;
  assign _EVAL_36 = _EVAL_23 | _EVAL_172;
  assign _EVAL_288 = _EVAL_250 == 4'h2;
  assign _EVAL_170 = _EVAL_36 | _EVAL_288;
  assign _EVAL_249 = _EVAL_170 | _EVAL_289;
  assign _EVAL_131 = _EVAL_6 == 3'h1;
  assign _EVAL_187 = _EVAL_71 == 1'h0;
  assign _EVAL_242 = _EVAL_279 | _EVAL_166;
  assign _EVAL_258 = _EVAL_4 <= 3'h2;
  assign _EVAL_64 = _EVAL_258 | _EVAL;
  assign _EVAL_104 = _EVAL_64 == 1'h0;
  assign _EVAL_271 = {{24'd0}, _EVAL_157};
  assign _EVAL_213 = _EVAL_0 & _EVAL_271;
  assign _EVAL_173 = _EVAL_213 == 30'h0;
  assign _EVAL_291 = _EVAL_173 | _EVAL;
  assign _EVAL_190 = _EVAL_274 == 1'h0;
  assign _EVAL_296 = _EVAL_3 == 3'h0;
  assign _EVAL_30 = _EVAL_192 | _EVAL;
  assign _EVAL_108 = _EVAL_30 == 1'h0;
  assign _EVAL_164 = _EVAL_3 == _EVAL_226;
  assign _EVAL_210 = _EVAL_164 | _EVAL;
  assign _EVAL_223 = _EVAL_179 + 32'h1;
  assign _EVAL_297 = _EVAL_11 & _EVAL_120;
  assign _EVAL_214 = _EVAL_175 == 1'h0;
  assign _EVAL_35 = _EVAL_3 <= 3'h6;
  assign _EVAL_33 = _EVAL_35 | _EVAL;
  assign _EVAL_111 = _EVAL_33 == 1'h0;
  assign _EVAL_38 = 3'h6 == _EVAL_1;
  assign _EVAL_59 = _EVAL_95 ? _EVAL_38 : 1'h0;
  assign _EVAL_171 = _EVAL_59 | _EVAL;
  assign _EVAL_234 = _EVAL_171 == 1'h0;
  assign _EVAL_207 = _EVAL_155 == 4'h0;
  assign _EVAL_45 = _EVAL_155 - 4'h1;
  assign _EVAL_65 = _EVAL_3 == 3'h2;
  assign _EVAL_160 = _EVAL_11 & _EVAL_65;
  assign _EVAL_74 = _EVAL_15 == _EVAL_24;
  assign _EVAL_185 = _EVAL_74 | _EVAL;
  assign _EVAL_140 = _EVAL_185 == 1'h0;
  assign _EVAL_106 = _EVAL_6 == 3'h6;
  assign _EVAL_134 = _EVAL_13 == _EVAL_270;
  assign _EVAL_107 = _EVAL_134 | _EVAL;
  assign _EVAL_88 = _EVAL_107 == 1'h0;
  assign _EVAL_229 = _EVAL_128 - 4'h1;
  assign _EVAL_138 = _EVAL_7 == 1'h0;
  assign _EVAL_143 = _EVAL_51 | _EVAL;
  assign _EVAL_256 = _EVAL_143 == 1'h0;
  assign _EVAL_273 = _EVAL_5 >= 3'h2;
  assign _EVAL_168 = _EVAL_166 & _EVAL_151;
  assign _EVAL_49 = _EVAL_4 == 3'h0;
  assign _EVAL_266 = _EVAL_156 | _EVAL;
  assign _EVAL_218 = _EVAL_49 | _EVAL;
  assign _EVAL_251 = _EVAL_218 == 1'h0;
  assign _EVAL_238 = _EVAL_273 | _EVAL;
  assign _EVAL_197 = _EVAL_238 == 1'h0;
  assign _EVAL_129 = _EVAL_230 == 1'h0;
  assign _EVAL_167 = _EVAL_3 == 3'h5;
  assign _EVAL_48 = _EVAL_8 & _EVAL_123;
  assign _EVAL_260 = _EVAL_8 & _EVAL_106;
  assign _EVAL_81 = _EVAL_1 == _EVAL_237;
  assign _EVAL_50 = _EVAL_81 | _EVAL;
  assign _EVAL_169 = _EVAL_50 == 1'h0;
  assign _EVAL_248 = _EVAL_279 & _EVAL_207;
  assign _EVAL_176 = _EVAL_4 != 3'h0;
  assign _EVAL_243 = _EVAL_176 | _EVAL;
  assign _EVAL_277 = _EVAL_6 == 3'h7;
  assign _EVAL_68 = _EVAL_8 & _EVAL_277;
  assign _EVAL_252 = _EVAL_291 == 1'h0;
  assign _EVAL_86 = _EVAL_195 == 1'h0;
  assign _EVAL_37 = _EVAL_186 | _EVAL;
  assign _EVAL_139 = _EVAL_138 | _EVAL;
  assign _EVAL_208 = _EVAL_266 == 1'h0;
  assign _EVAL_52 = _EVAL_207 == 1'h0;
  assign _EVAL_28 = _EVAL_6 == 3'h3;
  assign _EVAL_85 = _EVAL_8 & _EVAL_28;
  assign _EVAL_232 = _EVAL_6 == 3'h0;
  assign _EVAL_102 = _EVAL_37 == 1'h0;
  assign _EVAL_34 = _EVAL_6 == 3'h2;
  assign _EVAL_301 = _EVAL_210 == 1'h0;
  assign _EVAL_25 = _EVAL_11 & _EVAL_296;
  assign _EVAL_70 = _EVAL_249 | _EVAL;
  assign _EVAL_259 = _EVAL_70 == 1'h0;
  assign _EVAL_69 = _EVAL_11 & _EVAL_194;
  assign _EVAL_193 = _EVAL_8 & _EVAL_52;
  assign _EVAL_265 = _EVAL_8 & _EVAL_34;
  assign _EVAL_282 = _EVAL_8 & _EVAL_131;
  assign _EVAL_178 = _EVAL_243 == 1'h0;
  assign _EVAL_26 = _EVAL_139 == 1'h0;
  assign _EVAL_66 = _EVAL_6 == 3'h5;
  assign _EVAL_257 = _EVAL_8 & _EVAL_232;
  assign _EVAL_152 = _EVAL_57 == 1'h0;
  assign _EVAL_209 = _EVAL_8 & _EVAL_66;
  assign _EVAL_275 = _EVAL_11 & _EVAL_233;
  assign _EVAL_40 = _EVAL_11 & _EVAL_167;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_46 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_99 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_118 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_128 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_155 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_163 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_179 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_216 = _RAND_8[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_226 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_237 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {3{`RANDOM}};
  _EVAL_239 = _RAND_11[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_253 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_270 = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_285 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_168) begin
      _EVAL_24 <= _EVAL_15;
    end
    if (_EVAL_248) begin
      _EVAL_46 <= _EVAL_6;
    end
    if (_EVAL) begin
      _EVAL_99 <= 4'h0;
    end else begin
      if (_EVAL_279) begin
        if (_EVAL_199) begin
          if (_EVAL_267) begin
            _EVAL_99 <= _EVAL_281;
          end else begin
            _EVAL_99 <= 4'h0;
          end
        end else begin
          _EVAL_99 <= _EVAL_231;
        end
      end
    end
    if (_EVAL_248) begin
      _EVAL_118 <= _EVAL_12;
    end
    if (_EVAL) begin
      _EVAL_128 <= 4'h0;
    end else begin
      if (_EVAL_166) begin
        if (_EVAL_188) begin
          if (_EVAL_227) begin
            _EVAL_128 <= _EVAL_191;
          end else begin
            _EVAL_128 <= 4'h0;
          end
        end else begin
          _EVAL_128 <= _EVAL_229;
        end
      end
    end
    if (_EVAL) begin
      _EVAL_155 <= 4'h0;
    end else begin
      if (_EVAL_279) begin
        if (_EVAL_207) begin
          if (_EVAL_267) begin
            _EVAL_155 <= _EVAL_281;
          end else begin
            _EVAL_155 <= 4'h0;
          end
        end else begin
          _EVAL_155 <= _EVAL_45;
        end
      end
    end
    if (_EVAL) begin
      _EVAL_163 <= 4'h0;
    end else begin
      if (_EVAL_166) begin
        if (_EVAL_151) begin
          if (_EVAL_227) begin
            _EVAL_163 <= _EVAL_191;
          end else begin
            _EVAL_163 <= 4'h0;
          end
        end else begin
          _EVAL_163 <= _EVAL_221;
        end
      end
    end
    if (_EVAL) begin
      _EVAL_179 <= 32'h0;
    end else begin
      if (_EVAL_242) begin
        _EVAL_179 <= 32'h0;
      end else begin
        _EVAL_179 <= _EVAL_223;
      end
    end
    if (_EVAL_248) begin
      _EVAL_216 <= _EVAL_0;
    end
    if (_EVAL_168) begin
      _EVAL_226 <= _EVAL_3;
    end
    if (_EVAL_248) begin
      _EVAL_237 <= _EVAL_1;
    end
    if (_EVAL) begin
      _EVAL_239 <= 73'h0;
    end else begin
      _EVAL_239 <= _EVAL_121;
    end
    if (_EVAL_168) begin
      _EVAL_253 <= _EVAL_5;
    end
    if (_EVAL_168) begin
      _EVAL_270 <= _EVAL_13;
    end
    if (_EVAL_248) begin
      _EVAL_285 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4c01675)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3f5fd3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21363f0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69d145a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(427a432a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da395c87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4254e652)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e896b66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb76387e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67133d4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acde396b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d43d71a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23ffc8fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e7b0483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92090e90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f6deb2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff34e542)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8170401b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea738e92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35d6b96e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(410e2acc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e06f794)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaf70bc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12175d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(331676fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14bc7a9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f56aa3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd4d46e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8534be21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c76f87a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f67b6f1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348ce2eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d6949bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fd8293e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9befbee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ae23bce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611eaded)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47ee6db7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c2667e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ed650a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e508ba18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eeed3a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc30fc5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5882e54b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f85f298)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c62a279e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4afffc43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63ec63ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae751c10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf40994)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5952c9f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29b3020b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90496b5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a6a2d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9081bc73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df546678)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7097df35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f8518c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7fe7db5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e66323ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f76fa691)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d64c5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af003c97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d305e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be600f1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(239b2ed4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd8abca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45cac533)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77091135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee7f18d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33b1301d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1413c8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8948afe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(590cafee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fbd7eea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63a4d8e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7660b70d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6028884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbed6fa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6774dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
