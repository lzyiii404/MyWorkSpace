//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_175(
  input         _EVAL,
  output [31:0] _EVAL_0,
  output        _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [6:0]  _EVAL_4,
  output [2:0]  _EVAL_5,
  input  [6:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  output [6:0]  _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  output [2:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  input         _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  output [3:0]  _EVAL_20,
  input  [29:0] _EVAL_21,
  input  [31:0] _EVAL_22,
  output        _EVAL_23,
  output [2:0]  _EVAL_24,
  output        _EVAL_25,
  input  [3:0]  _EVAL_26,
  input         _EVAL_27,
  output [29:0] _EVAL_28,
  output [6:0]  _EVAL_29,
  input  [2:0]  _EVAL_30,
  input         _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [2:0]  _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  output [31:0] _EVAL_36
);
  assign _EVAL_19 = _EVAL_3;
  assign _EVAL_5 = _EVAL_12;
  assign _EVAL_23 = _EVAL;
  assign _EVAL_7 = _EVAL_8;
  assign _EVAL_20 = _EVAL_26;
  assign _EVAL_24 = _EVAL_33;
  assign _EVAL_29 = _EVAL_4;
  assign _EVAL_36 = _EVAL_14;
  assign _EVAL_11 = _EVAL_32;
  assign _EVAL_0 = _EVAL_22;
  assign _EVAL_16 = _EVAL_2;
  assign _EVAL_34 = _EVAL_35;
  assign _EVAL_13 = _EVAL_30;
  assign _EVAL_1 = _EVAL_17;
  assign _EVAL_18 = _EVAL_10;
  assign _EVAL_28 = _EVAL_21;
  assign _EVAL_25 = _EVAL_31;
  assign _EVAL_9 = _EVAL_6;
endmodule
