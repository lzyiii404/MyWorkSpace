//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module AXI4Shuffler(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire  Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire  Queue_io_deq_bits;
  wire [31:0] plusarg_reader_out;
  wire  MaxPeriodFibonacciLFSR__EVAL;
  wire  MaxPeriodFibonacciLFSR__EVAL_0;
  wire  MaxPeriodFibonacciLFSR__EVAL_1;
  wire  MaxPeriodFibonacciLFSR__EVAL_2;
  wire  MaxPeriodFibonacciLFSR__EVAL_3;
  wire  MaxPeriodFibonacciLFSR__EVAL_4;
  wire  MaxPeriodFibonacciLFSR__EVAL_5;
  wire  MaxPeriodFibonacciLFSR__EVAL_6;
  wire  MaxPeriodFibonacciLFSR__EVAL_7;
  wire  MaxPeriodFibonacciLFSR__EVAL_8;
  wire  MaxPeriodFibonacciLFSR__EVAL_9;
  wire  MaxPeriodFibonacciLFSR__EVAL_10;
  wire  MaxPeriodFibonacciLFSR__EVAL_11;
  wire  MaxPeriodFibonacciLFSR__EVAL_12;
  wire  MaxPeriodFibonacciLFSR__EVAL_13;
  wire  MaxPeriodFibonacciLFSR__EVAL_14;
  wire  MaxPeriodFibonacciLFSR__EVAL_15;
  wire  MaxPeriodFibonacciLFSR__EVAL_16;
  wire  MaxPeriodFibonacciLFSR__EVAL_17;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire  Queue_1_io_enq_bits_data_id;
  wire [29:0] Queue_1_io_enq_bits_data_addr;
  wire [7:0] Queue_1_io_enq_bits_data_len;
  wire [2:0] Queue_1_io_enq_bits_data_size;
  wire [1:0] Queue_1_io_enq_bits_data_burst;
  wire  Queue_1_io_enq_bits_data_lock;
  wire [3:0] Queue_1_io_enq_bits_data_cache;
  wire [2:0] Queue_1_io_enq_bits_data_prot;
  wire [3:0] Queue_1_io_enq_bits_data_qos;
  wire [31:0] Queue_1_io_enq_bits_timestamp;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire  Queue_1_io_deq_bits_data_id;
  wire [29:0] Queue_1_io_deq_bits_data_addr;
  wire [7:0] Queue_1_io_deq_bits_data_len;
  wire [2:0] Queue_1_io_deq_bits_data_size;
  wire [1:0] Queue_1_io_deq_bits_data_burst;
  wire  Queue_1_io_deq_bits_data_lock;
  wire [3:0] Queue_1_io_deq_bits_data_cache;
  wire [2:0] Queue_1_io_deq_bits_data_prot;
  wire [3:0] Queue_1_io_deq_bits_data_qos;
  wire [31:0] Queue_1_io_deq_bits_timestamp;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire  Queue_2_io_enq_bits_data_id;
  wire [29:0] Queue_2_io_enq_bits_data_addr;
  wire [7:0] Queue_2_io_enq_bits_data_len;
  wire [2:0] Queue_2_io_enq_bits_data_size;
  wire [1:0] Queue_2_io_enq_bits_data_burst;
  wire  Queue_2_io_enq_bits_data_lock;
  wire [3:0] Queue_2_io_enq_bits_data_cache;
  wire [2:0] Queue_2_io_enq_bits_data_prot;
  wire [3:0] Queue_2_io_enq_bits_data_qos;
  wire [31:0] Queue_2_io_enq_bits_timestamp;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire  Queue_2_io_deq_bits_data_id;
  wire [29:0] Queue_2_io_deq_bits_data_addr;
  wire [7:0] Queue_2_io_deq_bits_data_len;
  wire [2:0] Queue_2_io_deq_bits_data_size;
  wire [1:0] Queue_2_io_deq_bits_data_burst;
  wire  Queue_2_io_deq_bits_data_lock;
  wire [3:0] Queue_2_io_deq_bits_data_cache;
  wire [2:0] Queue_2_io_deq_bits_data_prot;
  wire [3:0] Queue_2_io_deq_bits_data_qos;
  wire [31:0] Queue_2_io_deq_bits_timestamp;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire  Queue_3_io_enq_bits_id;
  wire [29:0] Queue_3_io_enq_bits_addr;
  wire [7:0] Queue_3_io_enq_bits_len;
  wire [2:0] Queue_3_io_enq_bits_size;
  wire [1:0] Queue_3_io_enq_bits_burst;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire  Queue_3_io_deq_bits_id;
  wire [29:0] Queue_3_io_deq_bits_addr;
  wire [7:0] Queue_3_io_deq_bits_len;
  wire [2:0] Queue_3_io_deq_bits_size;
  wire [1:0] Queue_3_io_deq_bits_burst;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire  Queue_4_io_enq_bits;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire  Queue_4_io_deq_bits;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire  Queue_5_io_enq_bits_id;
  wire [29:0] Queue_5_io_enq_bits_addr;
  wire [7:0] Queue_5_io_enq_bits_len;
  wire [2:0] Queue_5_io_enq_bits_size;
  wire [1:0] Queue_5_io_enq_bits_burst;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire  Queue_5_io_deq_bits_id;
  wire [29:0] Queue_5_io_deq_bits_addr;
  wire [7:0] Queue_5_io_deq_bits_len;
  wire [2:0] Queue_5_io_deq_bits_size;
  wire [1:0] Queue_5_io_deq_bits_burst;
  wire  Queue_6_clock;
  wire  Queue_6_reset;
  wire  Queue_6_io_enq_ready;
  wire  Queue_6_io_enq_valid;
  wire [31:0] Queue_6_io_enq_bits_data;
  wire [3:0] Queue_6_io_enq_bits_strb;
  wire  Queue_6_io_enq_bits_last;
  wire  Queue_6_io_deq_ready;
  wire  Queue_6_io_deq_valid;
  wire [31:0] Queue_6_io_deq_bits_data;
  wire [3:0] Queue_6_io_deq_bits_strb;
  wire  Queue_6_io_deq_bits_last;
  wire  Queue_7_clock;
  wire  Queue_7_reset;
  wire  Queue_7_io_enq_ready;
  wire  Queue_7_io_enq_valid;
  wire [31:0] Queue_7_io_enq_bits_data;
  wire [3:0] Queue_7_io_enq_bits_strb;
  wire  Queue_7_io_enq_bits_last;
  wire  Queue_7_io_deq_ready;
  wire  Queue_7_io_deq_valid;
  wire [31:0] Queue_7_io_deq_bits_data;
  wire [3:0] Queue_7_io_deq_bits_strb;
  wire  Queue_7_io_deq_bits_last;
  wire [31:0] plusarg_reader_1_out;
  wire  MaxPeriodFibonacciLFSR_1__EVAL;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_17;
  wire  Queue_8_clock;
  wire  Queue_8_reset;
  wire  Queue_8_io_enq_ready;
  wire  Queue_8_io_enq_valid;
  wire  Queue_8_io_enq_bits_data_id;
  wire [29:0] Queue_8_io_enq_bits_data_addr;
  wire [7:0] Queue_8_io_enq_bits_data_len;
  wire [2:0] Queue_8_io_enq_bits_data_size;
  wire [1:0] Queue_8_io_enq_bits_data_burst;
  wire  Queue_8_io_enq_bits_data_lock;
  wire [3:0] Queue_8_io_enq_bits_data_cache;
  wire [2:0] Queue_8_io_enq_bits_data_prot;
  wire [3:0] Queue_8_io_enq_bits_data_qos;
  wire [31:0] Queue_8_io_enq_bits_timestamp;
  wire  Queue_8_io_deq_ready;
  wire  Queue_8_io_deq_valid;
  wire  Queue_8_io_deq_bits_data_id;
  wire [29:0] Queue_8_io_deq_bits_data_addr;
  wire [7:0] Queue_8_io_deq_bits_data_len;
  wire [2:0] Queue_8_io_deq_bits_data_size;
  wire [1:0] Queue_8_io_deq_bits_data_burst;
  wire  Queue_8_io_deq_bits_data_lock;
  wire [3:0] Queue_8_io_deq_bits_data_cache;
  wire [2:0] Queue_8_io_deq_bits_data_prot;
  wire [3:0] Queue_8_io_deq_bits_data_qos;
  wire [31:0] Queue_8_io_deq_bits_timestamp;
  wire  Queue_9_clock;
  wire  Queue_9_reset;
  wire  Queue_9_io_enq_ready;
  wire  Queue_9_io_enq_valid;
  wire  Queue_9_io_enq_bits_data_id;
  wire [29:0] Queue_9_io_enq_bits_data_addr;
  wire [7:0] Queue_9_io_enq_bits_data_len;
  wire [2:0] Queue_9_io_enq_bits_data_size;
  wire [1:0] Queue_9_io_enq_bits_data_burst;
  wire  Queue_9_io_enq_bits_data_lock;
  wire [3:0] Queue_9_io_enq_bits_data_cache;
  wire [2:0] Queue_9_io_enq_bits_data_prot;
  wire [3:0] Queue_9_io_enq_bits_data_qos;
  wire [31:0] Queue_9_io_enq_bits_timestamp;
  wire  Queue_9_io_deq_ready;
  wire  Queue_9_io_deq_valid;
  wire  Queue_9_io_deq_bits_data_id;
  wire [29:0] Queue_9_io_deq_bits_data_addr;
  wire [7:0] Queue_9_io_deq_bits_data_len;
  wire [2:0] Queue_9_io_deq_bits_data_size;
  wire [1:0] Queue_9_io_deq_bits_data_burst;
  wire  Queue_9_io_deq_bits_data_lock;
  wire [3:0] Queue_9_io_deq_bits_data_cache;
  wire [2:0] Queue_9_io_deq_bits_data_prot;
  wire [3:0] Queue_9_io_deq_bits_data_qos;
  wire [31:0] Queue_9_io_deq_bits_timestamp;
  wire  Queue_10_clock;
  wire  Queue_10_reset;
  wire  Queue_10_io_enq_ready;
  wire  Queue_10_io_enq_valid;
  wire  Queue_10_io_enq_bits_id;
  wire [29:0] Queue_10_io_enq_bits_addr;
  wire [7:0] Queue_10_io_enq_bits_len;
  wire [2:0] Queue_10_io_enq_bits_size;
  wire [1:0] Queue_10_io_enq_bits_burst;
  wire  Queue_10_io_deq_ready;
  wire  Queue_10_io_deq_valid;
  wire  Queue_10_io_deq_bits_id;
  wire [29:0] Queue_10_io_deq_bits_addr;
  wire [7:0] Queue_10_io_deq_bits_len;
  wire [2:0] Queue_10_io_deq_bits_size;
  wire [1:0] Queue_10_io_deq_bits_burst;
  wire [31:0] plusarg_reader_2_out;
  wire  MaxPeriodFibonacciLFSR_2__EVAL;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_17;
  wire  Queue_11_clock;
  wire  Queue_11_reset;
  wire  Queue_11_io_enq_ready;
  wire  Queue_11_io_enq_valid;
  wire [1:0] Queue_11_io_enq_bits_data_resp;
  wire [31:0] Queue_11_io_enq_bits_timestamp;
  wire  Queue_11_io_deq_ready;
  wire  Queue_11_io_deq_valid;
  wire  Queue_11_io_deq_bits_data_id;
  wire [1:0] Queue_11_io_deq_bits_data_resp;
  wire [31:0] Queue_11_io_deq_bits_timestamp;
  wire  Queue_12_clock;
  wire  Queue_12_reset;
  wire  Queue_12_io_enq_ready;
  wire  Queue_12_io_enq_valid;
  wire [1:0] Queue_12_io_enq_bits_data_resp;
  wire [31:0] Queue_12_io_enq_bits_timestamp;
  wire  Queue_12_io_deq_ready;
  wire  Queue_12_io_deq_valid;
  wire  Queue_12_io_deq_bits_data_id;
  wire [1:0] Queue_12_io_deq_bits_data_resp;
  wire [31:0] Queue_12_io_deq_bits_timestamp;
  wire  Queue_13_clock;
  wire  Queue_13_reset;
  wire  Queue_13_io_enq_ready;
  wire  Queue_13_io_enq_valid;
  wire  Queue_13_io_enq_bits_id;
  wire [1:0] Queue_13_io_enq_bits_resp;
  wire  Queue_13_io_deq_ready;
  wire  Queue_13_io_deq_valid;
  wire  Queue_13_io_deq_bits_id;
  wire [1:0] Queue_13_io_deq_bits_resp;
  wire [31:0] plusarg_reader_3_out;
  wire  MaxPeriodFibonacciLFSR_3__EVAL;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_17;
  wire  Queue_14_clock;
  wire  Queue_14_reset;
  wire  Queue_14_io_enq_ready;
  wire  Queue_14_io_enq_valid;
  wire [31:0] Queue_14_io_enq_bits_data_data;
  wire [1:0] Queue_14_io_enq_bits_data_resp;
  wire  Queue_14_io_enq_bits_data_last;
  wire [31:0] Queue_14_io_enq_bits_timestamp;
  wire  Queue_14_io_deq_ready;
  wire  Queue_14_io_deq_valid;
  wire  Queue_14_io_deq_bits_data_id;
  wire [31:0] Queue_14_io_deq_bits_data_data;
  wire [1:0] Queue_14_io_deq_bits_data_resp;
  wire  Queue_14_io_deq_bits_data_last;
  wire [31:0] Queue_14_io_deq_bits_timestamp;
  wire  Queue_15_clock;
  wire  Queue_15_reset;
  wire  Queue_15_io_enq_ready;
  wire  Queue_15_io_enq_valid;
  wire [31:0] Queue_15_io_enq_bits_data_data;
  wire [1:0] Queue_15_io_enq_bits_data_resp;
  wire  Queue_15_io_enq_bits_data_last;
  wire [31:0] Queue_15_io_enq_bits_timestamp;
  wire  Queue_15_io_deq_ready;
  wire  Queue_15_io_deq_valid;
  wire  Queue_15_io_deq_bits_data_id;
  wire [31:0] Queue_15_io_deq_bits_data_data;
  wire [1:0] Queue_15_io_deq_bits_data_resp;
  wire  Queue_15_io_deq_bits_data_last;
  wire [31:0] Queue_15_io_deq_bits_timestamp;
  wire  Queue_16_clock;
  wire  Queue_16_reset;
  wire  Queue_16_io_enq_ready;
  wire  Queue_16_io_enq_valid;
  wire  Queue_16_io_enq_bits_id;
  wire [31:0] Queue_16_io_enq_bits_data;
  wire [1:0] Queue_16_io_enq_bits_resp;
  wire  Queue_16_io_enq_bits_last;
  wire  Queue_16_io_deq_ready;
  wire  Queue_16_io_deq_valid;
  wire  Queue_16_io_deq_bits_id;
  wire [31:0] Queue_16_io_deq_bits_data;
  wire [1:0] Queue_16_io_deq_bits_resp;
  wire  Queue_16_io_deq_bits_last;
  wire  _T_71_1;
  wire  _T_71_0;
  wire  _GEN_3;
  wire [7:0] _T_19;
  wire [15:0] _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_39;
  wire  _T_40;
  wire  _T_41;
  wire  _T_42;
  wire  _T_43;
  wire [7:0] _T_51;
  wire [15:0] _T_59;
  wire  _T_60;
  wire  _T_9;
  wire  _T_64;
  wire  _T_65;
  wire  _T_6;
  reg [31:0] _T_10;
  reg [31:0] _RAND_0;
  wire [31:0] _T_12;
  wire  _T_63;
  wire [1:0] _T_68;
  wire [31:0] _GEN_32;
  wire [1:0] _T_73;
  wire  _T_75;
  wire  _T_76;
  wire  _T_81;
  wire  _T_82;
  wire  _T_83;
  wire  _T_79_ready;
  reg  _T_92;
  reg [31:0] _RAND_1;
  wire  _T_93;
  wire  _T_87;
  wire  _T_88;
  wire  _T_89;
  wire [1:0] _T_95;
  reg [1:0] _T_102;
  reg [31:0] _RAND_2;
  wire [1:0] _T_103;
  wire [1:0] _T_104;
  wire [3:0] _T_105;
  wire [2:0] _T_106;
  wire [3:0] _GEN_33;
  wire [3:0] _T_107;
  wire [2:0] _T_109;
  wire [3:0] _T_110;
  wire [3:0] _GEN_34;
  wire [3:0] _T_111;
  wire [1:0] _T_112;
  wire [1:0] _T_113;
  wire [1:0] _T_114;
  wire [1:0] _T_115;
  wire  _T_124;
  reg  _T_157_0;
  reg [31:0] _RAND_3;
  wire  _T_159_0;
  wire  _T_160;
  wire  _T_125;
  reg  _T_157_1;
  reg [31:0] _RAND_4;
  wire  _T_159_1;
  wire  _T_161;
  wire  _T_94;
  wire  _T_97;
  wire  _T_99;
  wire  _T_100;
  wire  _T_116;
  wire  _T_117;
  wire [1:0] _T_118;
  wire [2:0] _T_119;
  wire [1:0] _T_120;
  wire [1:0] _T_121;
  wire  _T_127;
  wire  _T_128;
  wire  _T_131;
  wire  _T_133;
  wire  _T_136;
  wire  _T_137;
  wire  _T_140;
  wire  _T_141;
  wire  _T_142;
  wire  _T_143;
  wire  _T_145;
  wire  _T_147;
  wire  _T_148;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _T_167;
  wire  _T_152;
  wire  _T_154;
  wire  _T_158_0;
  wire  _T_158_1;
  wire [2:0] _T_80_bits_prot;
  wire [3:0] _T_80_bits_qos;
  wire  _T_80_bits_lock;
  wire [3:0] _T_80_bits_cache;
  wire [2:0] _T_80_bits_size;
  wire [1:0] _T_80_bits_burst;
  wire  _T_80_bits_id;
  wire [29:0] _T_80_bits_addr;
  wire [7:0] _T_80_bits_len;
  wire [55:0] _T_175;
  wire [55:0] _T_176;
  wire [2:0] _T_86_bits_prot;
  wire [3:0] _T_86_bits_qos;
  wire  _T_86_bits_lock;
  wire [3:0] _T_86_bits_cache;
  wire [2:0] _T_86_bits_size;
  wire [1:0] _T_86_bits_burst;
  wire  _T_86_bits_id;
  wire [29:0] _T_86_bits_addr;
  wire [7:0] _T_86_bits_len;
  wire [55:0] _T_184;
  wire [55:0] _T_185;
  wire [55:0] _T_186;
  wire  _T_199_ready;
  wire  _T_198_valid;
  wire  _T_4_bits;
  wire  _T_204_0;
  wire  _T_204_1;
  wire  _GEN_8;
  wire  _T_205;
  wire  _T_4_valid;
  wire [1:0] _T_209;
  wire  _T_211;
  wire  _T_212;
  wire  _T_213;
  wire  _T_200_bits;
  wire [31:0] _T_219_0_data;
  wire [3:0] _T_219_0_strb;
  wire  _T_219_0_last;
  wire [31:0] _T_219_1_data;
  wire [3:0] _T_219_1_strb;
  wire  _T_219_1_last;
  wire  _GEN_14;
  wire  _T_218_0;
  wire  _T_218_1;
  wire  _GEN_16;
  wire  _T_220;
  wire  _T_200_valid;
  wire [1:0] _T_224;
  wire  _T_226;
  wire  _T_227;
  wire  _T_228;
  wire  _T_233;
  reg [31:0] _T_234;
  reg [31:0] _RAND_5;
  wire [31:0] _T_236;
  wire [7:0] _T_243;
  wire [15:0] _T_251;
  wire  _T_252;
  wire  _T_253;
  wire  _T_254;
  wire  _T_255;
  wire  _T_256;
  wire  _T_257;
  wire  _T_258;
  wire  _T_259;
  wire  _T_260;
  wire  _T_261;
  wire  _T_262;
  wire  _T_263;
  wire  _T_264;
  wire  _T_265;
  wire  _T_266;
  wire  _T_267;
  wire [7:0] _T_275;
  wire [15:0] _T_283;
  wire  _T_284;
  wire  _T_286;
  wire  _T_287;
  wire  _T_295_1;
  wire  _T_295_0;
  wire  _GEN_20;
  wire [1:0] _T_292;
  wire [31:0] _GEN_35;
  wire [1:0] _T_297;
  wire  _T_299;
  wire  _T_300;
  wire  _T_305;
  wire  _T_306;
  wire  _T_307;
  wire  _T_303_ready;
  reg  _T_316;
  reg [31:0] _RAND_6;
  wire  _T_317;
  wire  _T_311;
  wire  _T_312;
  wire  _T_313;
  wire [1:0] _T_319;
  reg [1:0] _T_326;
  reg [31:0] _RAND_7;
  wire [1:0] _T_327;
  wire [1:0] _T_328;
  wire [3:0] _T_329;
  wire [2:0] _T_330;
  wire [3:0] _GEN_36;
  wire [3:0] _T_331;
  wire [2:0] _T_333;
  wire [3:0] _T_334;
  wire [3:0] _GEN_37;
  wire [3:0] _T_335;
  wire [1:0] _T_336;
  wire [1:0] _T_337;
  wire [1:0] _T_338;
  wire [1:0] _T_339;
  wire  _T_348;
  reg  _T_381_0;
  reg [31:0] _RAND_8;
  wire  _T_383_0;
  wire  _T_384;
  wire  _T_349;
  reg  _T_381_1;
  reg [31:0] _RAND_9;
  wire  _T_383_1;
  wire  _T_385;
  wire  _T_318;
  wire  _T_321;
  wire  _T_323;
  wire  _T_324;
  wire  _T_340;
  wire  _T_341;
  wire [1:0] _T_342;
  wire [2:0] _T_343;
  wire [1:0] _T_344;
  wire [1:0] _T_345;
  wire  _T_351;
  wire  _T_352;
  wire  _T_355;
  wire  _T_357;
  wire  _T_360;
  wire  _T_361;
  wire  _T_364;
  wire  _T_365;
  wire  _T_366;
  wire  _T_367;
  wire  _T_369;
  wire  _T_371;
  wire  _T_372;
  wire  _T_387;
  wire  _T_388;
  wire  _T_389;
  wire  _T_391;
  wire  _T_376;
  wire  _T_378;
  wire  _T_382_0;
  wire  _T_382_1;
  wire [2:0] _T_304_bits_prot;
  wire [3:0] _T_304_bits_qos;
  wire  _T_304_bits_lock;
  wire [3:0] _T_304_bits_cache;
  wire [2:0] _T_304_bits_size;
  wire [1:0] _T_304_bits_burst;
  wire  _T_304_bits_id;
  wire [29:0] _T_304_bits_addr;
  wire [7:0] _T_304_bits_len;
  wire [55:0] _T_399;
  wire [55:0] _T_400;
  wire [2:0] _T_310_bits_prot;
  wire [3:0] _T_310_bits_qos;
  wire  _T_310_bits_lock;
  wire [3:0] _T_310_bits_cache;
  wire [2:0] _T_310_bits_size;
  wire [1:0] _T_310_bits_burst;
  wire  _T_310_bits_id;
  wire [29:0] _T_310_bits_addr;
  wire [7:0] _T_310_bits_len;
  wire [55:0] _T_408;
  wire [55:0] _T_409;
  wire [55:0] _T_410;
  wire  _T_424;
  reg [31:0] _T_425;
  reg [31:0] _RAND_10;
  wire [31:0] _T_427;
  wire [7:0] _T_434;
  wire [15:0] _T_442;
  wire  _T_443;
  wire  _T_444;
  wire  _T_445;
  wire  _T_446;
  wire  _T_447;
  wire  _T_448;
  wire  _T_449;
  wire  _T_450;
  wire  _T_451;
  wire  _T_452;
  wire  _T_453;
  wire  _T_454;
  wire  _T_455;
  wire  _T_456;
  wire  _T_457;
  wire  _T_458;
  wire [7:0] _T_466;
  wire [15:0] _T_474;
  wire [1:0] _T_483;
  wire [31:0] _GEN_38;
  wire  _T_496;
  wire  _T_497;
  wire  _T_498;
  wire  _T_494_ready;
  reg  _T_507;
  reg [31:0] _RAND_11;
  wire  _T_508;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire [1:0] _T_510;
  reg [1:0] _T_517;
  reg [31:0] _RAND_12;
  wire [1:0] _T_518;
  wire [1:0] _T_519;
  wire [3:0] _T_520;
  wire [2:0] _T_521;
  wire [3:0] _GEN_39;
  wire [3:0] _T_522;
  wire [2:0] _T_524;
  wire [3:0] _T_525;
  wire [3:0] _GEN_40;
  wire [3:0] _T_526;
  wire [1:0] _T_527;
  wire [1:0] _T_528;
  wire [1:0] _T_529;
  wire [1:0] _T_530;
  wire  _T_539;
  reg  _T_572_0;
  reg [31:0] _RAND_13;
  wire  _T_574_0;
  wire  _T_575;
  wire  _T_540;
  reg  _T_572_1;
  reg [31:0] _RAND_14;
  wire  _T_574_1;
  wire  _T_576;
  wire  _T_509;
  wire  _T_512;
  wire  _T_514;
  wire  _T_515;
  wire  _T_531;
  wire  _T_532;
  wire [1:0] _T_533;
  wire [2:0] _T_534;
  wire [1:0] _T_535;
  wire [1:0] _T_536;
  wire  _T_542;
  wire  _T_543;
  wire  _T_546;
  wire  _T_548;
  wire  _T_551;
  wire  _T_552;
  wire  _T_555;
  wire  _T_556;
  wire  _T_557;
  wire  _T_558;
  wire  _T_560;
  wire  _T_562;
  wire  _T_563;
  wire  _T_578;
  wire  _T_579;
  wire  _T_580;
  wire  _T_582;
  wire  _T_567;
  wire  _T_569;
  wire  _T_573_0;
  wire  _T_573_1;
  wire  _T_495_bits_id;
  wire [1:0] _T_495_bits_resp;
  wire [2:0] _T_583;
  wire [2:0] _T_584;
  wire  _T_501_bits_id;
  wire [1:0] _T_501_bits_resp;
  wire [2:0] _T_585;
  wire [2:0] _T_586;
  wire [2:0] _T_587;
  wire  _T_594;
  reg [31:0] _T_595;
  reg [31:0] _RAND_15;
  wire [31:0] _T_597;
  wire [7:0] _T_604;
  wire [15:0] _T_612;
  wire  _T_613;
  wire  _T_614;
  wire  _T_615;
  wire  _T_616;
  wire  _T_617;
  wire  _T_618;
  wire  _T_619;
  wire  _T_620;
  wire  _T_621;
  wire  _T_622;
  wire  _T_623;
  wire  _T_624;
  wire  _T_625;
  wire  _T_626;
  wire  _T_627;
  wire  _T_628;
  wire [7:0] _T_636;
  wire [15:0] _T_644;
  wire [1:0] _T_653;
  wire [31:0] _GEN_41;
  wire  _T_666;
  wire  _T_667;
  wire  _T_668;
  wire  _T_664_ready;
  reg  _T_677;
  reg [31:0] _RAND_16;
  wire  _T_678;
  wire  _T_672;
  wire  _T_673;
  wire  _T_674;
  wire [1:0] _T_680;
  reg [1:0] _T_687;
  reg [31:0] _RAND_17;
  wire [1:0] _T_688;
  wire [1:0] _T_689;
  wire [3:0] _T_690;
  wire [2:0] _T_691;
  wire [3:0] _GEN_42;
  wire [3:0] _T_692;
  wire [2:0] _T_694;
  wire [3:0] _T_695;
  wire [3:0] _GEN_43;
  wire [3:0] _T_696;
  wire [1:0] _T_697;
  wire [1:0] _T_698;
  wire [1:0] _T_699;
  wire [1:0] _T_700;
  wire  _T_709;
  reg  _T_742_0;
  reg [31:0] _RAND_18;
  wire  _T_744_0;
  wire  _T_745;
  wire  _T_710;
  reg  _T_742_1;
  reg [31:0] _RAND_19;
  wire  _T_744_1;
  wire  _T_746;
  wire  _T_679;
  wire  _T_682;
  wire  _T_684;
  wire  _T_685;
  wire  _T_701;
  wire  _T_702;
  wire [1:0] _T_703;
  wire [2:0] _T_704;
  wire [1:0] _T_705;
  wire [1:0] _T_706;
  wire  _T_712;
  wire  _T_713;
  wire  _T_716;
  wire  _T_718;
  wire  _T_721;
  wire  _T_722;
  wire  _T_725;
  wire  _T_726;
  wire  _T_727;
  wire  _T_728;
  wire  _T_730;
  wire  _T_732;
  wire  _T_733;
  wire  _T_748;
  wire  _T_749;
  wire  _T_750;
  wire  _T_752;
  wire  _T_737;
  wire  _T_739;
  wire  _T_743_0;
  wire  _T_743_1;
  wire [1:0] _T_665_bits_resp;
  wire  _T_665_bits_last;
  wire  _T_665_bits_id;
  wire [31:0] _T_665_bits_data;
  wire [35:0] _T_755;
  wire [35:0] _T_756;
  wire [1:0] _T_671_bits_resp;
  wire  _T_671_bits_last;
  wire  _T_671_bits_id;
  wire [31:0] _T_671_bits_data;
  wire [35:0] _T_759;
  wire [35:0] _T_760;
  wire [35:0] _T_761;
  Queue_85 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR (
    ._EVAL(MaxPeriodFibonacciLFSR__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR__EVAL_17)
  );
  Queue_86 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data_id(Queue_1_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_1_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_1_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_1_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_1_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_1_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_1_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_1_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_1_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_1_io_enq_bits_timestamp),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data_id(Queue_1_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_1_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_1_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_1_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_1_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_1_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_1_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_1_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_1_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_1_io_deq_bits_timestamp)
  );
  Queue_86 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data_id(Queue_2_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_2_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_2_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_2_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_2_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_2_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_2_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_2_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_2_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_2_io_enq_bits_timestamp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data_id(Queue_2_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_2_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_2_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_2_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_2_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_2_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_2_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_2_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_2_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_2_io_deq_bits_timestamp)
  );
  Queue_88 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_len(Queue_3_io_enq_bits_len),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_burst(Queue_3_io_enq_bits_burst),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_len(Queue_3_io_deq_bits_len),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_burst(Queue_3_io_deq_bits_burst)
  );
  Queue_85 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  Queue_88 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_id(Queue_5_io_enq_bits_id),
    .io_enq_bits_addr(Queue_5_io_enq_bits_addr),
    .io_enq_bits_len(Queue_5_io_enq_bits_len),
    .io_enq_bits_size(Queue_5_io_enq_bits_size),
    .io_enq_bits_burst(Queue_5_io_enq_bits_burst),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_id(Queue_5_io_deq_bits_id),
    .io_deq_bits_addr(Queue_5_io_deq_bits_addr),
    .io_deq_bits_len(Queue_5_io_deq_bits_len),
    .io_deq_bits_size(Queue_5_io_deq_bits_size),
    .io_deq_bits_burst(Queue_5_io_deq_bits_burst)
  );
  Queue_91 Queue_6 (
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits_data(Queue_6_io_enq_bits_data),
    .io_enq_bits_strb(Queue_6_io_enq_bits_strb),
    .io_enq_bits_last(Queue_6_io_enq_bits_last),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits_data(Queue_6_io_deq_bits_data),
    .io_deq_bits_strb(Queue_6_io_deq_bits_strb),
    .io_deq_bits_last(Queue_6_io_deq_bits_last)
  );
  Queue_91 Queue_7 (
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits_data(Queue_7_io_enq_bits_data),
    .io_enq_bits_strb(Queue_7_io_enq_bits_strb),
    .io_enq_bits_last(Queue_7_io_enq_bits_last),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits_data(Queue_7_io_deq_bits_data),
    .io_deq_bits_strb(Queue_7_io_deq_bits_strb),
    .io_deq_bits_last(Queue_7_io_deq_bits_last)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 (
    .out(plusarg_reader_1_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_1 (
    ._EVAL(MaxPeriodFibonacciLFSR_1__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_1__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_1__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_1__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_1__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_1__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_1__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_1__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_1__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_1__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_1__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_1__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_1__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_1__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_1__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_1__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_1__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_1__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_1__EVAL_17)
  );
  Queue_86 Queue_8 (
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits_data_id(Queue_8_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_8_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_8_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_8_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_8_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_8_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_8_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_8_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_8_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_8_io_enq_bits_timestamp),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits_data_id(Queue_8_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_8_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_8_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_8_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_8_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_8_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_8_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_8_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_8_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_8_io_deq_bits_timestamp)
  );
  Queue_86 Queue_9 (
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits_data_id(Queue_9_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_9_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_9_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_9_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_9_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_9_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_9_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_9_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_9_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_9_io_enq_bits_timestamp),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits_data_id(Queue_9_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_9_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_9_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_9_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_9_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_9_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_9_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_9_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_9_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_9_io_deq_bits_timestamp)
  );
  Queue_88 Queue_10 (
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits_id(Queue_10_io_enq_bits_id),
    .io_enq_bits_addr(Queue_10_io_enq_bits_addr),
    .io_enq_bits_len(Queue_10_io_enq_bits_len),
    .io_enq_bits_size(Queue_10_io_enq_bits_size),
    .io_enq_bits_burst(Queue_10_io_enq_bits_burst),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits_id(Queue_10_io_deq_bits_id),
    .io_deq_bits_addr(Queue_10_io_deq_bits_addr),
    .io_deq_bits_len(Queue_10_io_deq_bits_len),
    .io_deq_bits_size(Queue_10_io_deq_bits_size),
    .io_deq_bits_burst(Queue_10_io_deq_bits_burst)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_2 (
    .out(plusarg_reader_2_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_2 (
    ._EVAL(MaxPeriodFibonacciLFSR_2__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_2__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_2__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_2__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_2__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_2__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_2__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_2__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_2__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_2__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_2__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_2__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_2__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_2__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_2__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_2__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_2__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_2__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_2__EVAL_17)
  );
  Queue_96 Queue_11 (
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits_data_resp(Queue_11_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_11_io_enq_bits_timestamp),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits_data_id(Queue_11_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_11_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_11_io_deq_bits_timestamp)
  );
  Queue_96 Queue_12 (
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits_data_resp(Queue_12_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_12_io_enq_bits_timestamp),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits_data_id(Queue_12_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_12_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_12_io_deq_bits_timestamp)
  );
  Queue_98 Queue_13 (
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits_id(Queue_13_io_enq_bits_id),
    .io_enq_bits_resp(Queue_13_io_enq_bits_resp),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits_id(Queue_13_io_deq_bits_id),
    .io_deq_bits_resp(Queue_13_io_deq_bits_resp)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_3 (
    .out(plusarg_reader_3_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_3 (
    ._EVAL(MaxPeriodFibonacciLFSR_3__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_3__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_3__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_3__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_3__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_3__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_3__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_3__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_3__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_3__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_3__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_3__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_3__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_3__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_3__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_3__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_3__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_3__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_3__EVAL_17)
  );
  Queue_99 Queue_14 (
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits_data_data(Queue_14_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_14_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_14_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_14_io_enq_bits_timestamp),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits_data_id(Queue_14_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_14_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_14_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_14_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_14_io_deq_bits_timestamp)
  );
  Queue_99 Queue_15 (
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits_data_data(Queue_15_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_15_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_15_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_15_io_enq_bits_timestamp),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits_data_id(Queue_15_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_15_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_15_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_15_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_15_io_deq_bits_timestamp)
  );
  Queue_101 Queue_16 (
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits_id(Queue_16_io_enq_bits_id),
    .io_enq_bits_data(Queue_16_io_enq_bits_data),
    .io_enq_bits_resp(Queue_16_io_enq_bits_resp),
    .io_enq_bits_last(Queue_16_io_enq_bits_last),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits_id(Queue_16_io_deq_bits_id),
    .io_deq_bits_data(Queue_16_io_deq_bits_data),
    .io_deq_bits_resp(Queue_16_io_deq_bits_resp),
    .io_deq_bits_last(Queue_16_io_deq_bits_last)
  );
  assign _T_71_1 = Queue_2_io_enq_ready;
  assign _T_71_0 = Queue_1_io_enq_ready;
  assign _GEN_3 = auto_in_aw_bits_id ? _T_71_1 : _T_71_0;
  assign _T_19 = {MaxPeriodFibonacciLFSR__EVAL_12,MaxPeriodFibonacciLFSR__EVAL_11,MaxPeriodFibonacciLFSR__EVAL_3,MaxPeriodFibonacciLFSR__EVAL_16,MaxPeriodFibonacciLFSR__EVAL_8,MaxPeriodFibonacciLFSR__EVAL_10,MaxPeriodFibonacciLFSR__EVAL_14,MaxPeriodFibonacciLFSR__EVAL_7};
  assign _T_27 = {MaxPeriodFibonacciLFSR__EVAL_0,MaxPeriodFibonacciLFSR__EVAL_17,MaxPeriodFibonacciLFSR__EVAL_1,MaxPeriodFibonacciLFSR__EVAL,MaxPeriodFibonacciLFSR__EVAL_5,MaxPeriodFibonacciLFSR__EVAL_4,MaxPeriodFibonacciLFSR__EVAL_6,MaxPeriodFibonacciLFSR__EVAL_2,_T_19};
  assign _T_28 = _T_27[0];
  assign _T_29 = _T_27[1];
  assign _T_30 = _T_27[2];
  assign _T_31 = _T_27[3];
  assign _T_32 = _T_27[4];
  assign _T_33 = _T_27[5];
  assign _T_34 = _T_27[6];
  assign _T_35 = _T_27[7];
  assign _T_36 = _T_27[8];
  assign _T_37 = _T_27[9];
  assign _T_38 = _T_27[10];
  assign _T_39 = _T_27[11];
  assign _T_40 = _T_27[12];
  assign _T_41 = _T_27[13];
  assign _T_42 = _T_27[14];
  assign _T_43 = _T_27[15];
  assign _T_51 = {_T_36,_T_37,_T_38,_T_39,_T_40,_T_41,_T_42,_T_43};
  assign _T_59 = {_T_28,_T_29,_T_30,_T_31,_T_32,_T_33,_T_34,_T_35,_T_51};
  assign _T_60 = 16'h3fff <= _T_59;
  assign _T_9 = plusarg_reader_out[0];
  assign _T_64 = _T_60 | _T_9;
  assign _T_65 = _GEN_3 & _T_64;
  assign _T_6 = auto_in_aw_valid & Queue_io_enq_ready;
  assign _T_12 = _T_10 + 32'h1;
  assign _T_63 = _T_6 & _T_64;
  assign _T_68 = _T_59[1:0];
  assign _GEN_32 = {{30'd0}, _T_68};
  assign _T_73 = 2'h1 << auto_in_aw_bits_id;
  assign _T_75 = _T_73[0];
  assign _T_76 = _T_73[1];
  assign _T_81 = Queue_1_io_deq_bits_timestamp <= _T_10;
  assign _T_82 = _T_81 | _T_9;
  assign _T_83 = Queue_1_io_deq_valid & _T_82;
  assign _T_79_ready = Queue_3_io_enq_ready;
  assign _T_93 = _T_92 == 1'h0;
  assign _T_87 = Queue_2_io_deq_bits_timestamp <= _T_10;
  assign _T_88 = _T_87 | _T_9;
  assign _T_89 = Queue_2_io_deq_valid & _T_88;
  assign _T_95 = {_T_89,_T_83};
  assign _T_103 = ~ _T_102;
  assign _T_104 = _T_95 & _T_103;
  assign _T_105 = {_T_104,_T_89,_T_83};
  assign _T_106 = _T_105[3:1];
  assign _GEN_33 = {{1'd0}, _T_106};
  assign _T_107 = _T_105 | _GEN_33;
  assign _T_109 = _T_107[3:1];
  assign _T_110 = {_T_102, 2'h0};
  assign _GEN_34 = {{1'd0}, _T_109};
  assign _T_111 = _GEN_34 | _T_110;
  assign _T_112 = _T_111[3:2];
  assign _T_113 = _T_111[1:0];
  assign _T_114 = _T_112 & _T_113;
  assign _T_115 = ~ _T_114;
  assign _T_124 = _T_115[0];
  assign _T_159_0 = _T_93 ? _T_124 : _T_157_0;
  assign _T_160 = _T_79_ready & _T_159_0;
  assign _T_125 = _T_115[1];
  assign _T_159_1 = _T_93 ? _T_125 : _T_157_1;
  assign _T_161 = _T_79_ready & _T_159_1;
  assign _T_94 = _T_93 & _T_79_ready;
  assign _T_97 = _T_95 == _T_95;
  assign _T_99 = _T_97 | reset;
  assign _T_100 = _T_99 == 1'h0;
  assign _T_116 = _T_95 != 2'h0;
  assign _T_117 = _T_94 & _T_116;
  assign _T_118 = _T_115 & _T_95;
  assign _T_119 = {_T_118, 1'h0};
  assign _T_120 = _T_119[1:0];
  assign _T_121 = _T_118 | _T_120;
  assign _T_127 = _T_124 & _T_83;
  assign _T_128 = _T_125 & _T_89;
  assign _T_131 = _T_127 | _T_128;
  assign _T_133 = _T_127 == 1'h0;
  assign _T_136 = _T_128 == 1'h0;
  assign _T_137 = _T_133 | _T_136;
  assign _T_140 = _T_137 | reset;
  assign _T_141 = _T_140 == 1'h0;
  assign _T_142 = _T_83 | _T_89;
  assign _T_143 = _T_142 == 1'h0;
  assign _T_145 = _T_143 | _T_131;
  assign _T_147 = _T_145 | reset;
  assign _T_148 = _T_147 == 1'h0;
  assign _T_163 = _T_157_0 ? _T_83 : 1'h0;
  assign _T_164 = _T_157_1 ? _T_89 : 1'h0;
  assign _T_165 = _T_163 | _T_164;
  assign _T_167 = _T_93 ? _T_142 : _T_165;
  assign _T_152 = _T_79_ready & _T_167;
  assign _T_154 = _T_92 - _T_152;
  assign _T_158_0 = _T_93 ? _T_127 : _T_157_0;
  assign _T_158_1 = _T_93 ? _T_128 : _T_157_1;
  assign _T_80_bits_prot = Queue_1_io_deq_bits_data_prot;
  assign _T_80_bits_qos = Queue_1_io_deq_bits_data_qos;
  assign _T_80_bits_lock = Queue_1_io_deq_bits_data_lock;
  assign _T_80_bits_cache = Queue_1_io_deq_bits_data_cache;
  assign _T_80_bits_size = Queue_1_io_deq_bits_data_size;
  assign _T_80_bits_burst = Queue_1_io_deq_bits_data_burst;
  assign _T_80_bits_id = Queue_1_io_deq_bits_data_id;
  assign _T_80_bits_addr = Queue_1_io_deq_bits_data_addr;
  assign _T_80_bits_len = Queue_1_io_deq_bits_data_len;
  assign _T_175 = {_T_80_bits_id,_T_80_bits_addr,_T_80_bits_len,_T_80_bits_size,_T_80_bits_burst,_T_80_bits_lock,_T_80_bits_cache,_T_80_bits_prot,_T_80_bits_qos};
  assign _T_176 = _T_158_0 ? _T_175 : 56'h0;
  assign _T_86_bits_prot = Queue_2_io_deq_bits_data_prot;
  assign _T_86_bits_qos = Queue_2_io_deq_bits_data_qos;
  assign _T_86_bits_lock = Queue_2_io_deq_bits_data_lock;
  assign _T_86_bits_cache = Queue_2_io_deq_bits_data_cache;
  assign _T_86_bits_size = Queue_2_io_deq_bits_data_size;
  assign _T_86_bits_burst = Queue_2_io_deq_bits_data_burst;
  assign _T_86_bits_id = Queue_2_io_deq_bits_data_id;
  assign _T_86_bits_addr = Queue_2_io_deq_bits_data_addr;
  assign _T_86_bits_len = Queue_2_io_deq_bits_data_len;
  assign _T_184 = {_T_86_bits_id,_T_86_bits_addr,_T_86_bits_len,_T_86_bits_size,_T_86_bits_burst,_T_86_bits_lock,_T_86_bits_cache,_T_86_bits_prot,_T_86_bits_qos};
  assign _T_185 = _T_158_1 ? _T_184 : 56'h0;
  assign _T_186 = _T_176 | _T_185;
  assign _T_199_ready = Queue_5_io_enq_ready;
  assign _T_198_valid = Queue_3_io_deq_valid;
  assign _T_4_bits = Queue_io_deq_bits;
  assign _T_204_0 = Queue_6_io_enq_ready;
  assign _T_204_1 = Queue_7_io_enq_ready;
  assign _GEN_8 = _T_4_bits ? _T_204_1 : _T_204_0;
  assign _T_205 = auto_in_w_bits_last & _GEN_8;
  assign _T_4_valid = Queue_io_deq_valid;
  assign _T_209 = 2'h1 << _T_4_bits;
  assign _T_211 = _T_209[0];
  assign _T_212 = _T_209[1];
  assign _T_213 = _T_4_valid & auto_in_w_valid;
  assign _T_200_bits = Queue_4_io_deq_bits;
  assign _T_219_0_data = Queue_6_io_deq_bits_data;
  assign _T_219_0_strb = Queue_6_io_deq_bits_strb;
  assign _T_219_0_last = Queue_6_io_deq_bits_last;
  assign _T_219_1_data = Queue_7_io_deq_bits_data;
  assign _T_219_1_strb = Queue_7_io_deq_bits_strb;
  assign _T_219_1_last = Queue_7_io_deq_bits_last;
  assign _GEN_14 = _T_200_bits ? _T_219_1_last : _T_219_0_last;
  assign _T_218_0 = Queue_6_io_deq_valid;
  assign _T_218_1 = Queue_7_io_deq_valid;
  assign _GEN_16 = _T_200_bits ? _T_218_1 : _T_218_0;
  assign _T_220 = _GEN_14 & _GEN_16;
  assign _T_200_valid = Queue_4_io_deq_valid;
  assign _T_224 = 2'h1 << _T_200_bits;
  assign _T_226 = _T_224[0];
  assign _T_227 = _T_224[1];
  assign _T_228 = _T_200_valid & auto_out_w_ready;
  assign _T_233 = plusarg_reader_1_out[0];
  assign _T_236 = _T_234 + 32'h1;
  assign _T_243 = {MaxPeriodFibonacciLFSR_1__EVAL_12,MaxPeriodFibonacciLFSR_1__EVAL_11,MaxPeriodFibonacciLFSR_1__EVAL_3,MaxPeriodFibonacciLFSR_1__EVAL_16,MaxPeriodFibonacciLFSR_1__EVAL_8,MaxPeriodFibonacciLFSR_1__EVAL_10,MaxPeriodFibonacciLFSR_1__EVAL_14,MaxPeriodFibonacciLFSR_1__EVAL_7};
  assign _T_251 = {MaxPeriodFibonacciLFSR_1__EVAL_0,MaxPeriodFibonacciLFSR_1__EVAL_17,MaxPeriodFibonacciLFSR_1__EVAL_1,MaxPeriodFibonacciLFSR_1__EVAL,MaxPeriodFibonacciLFSR_1__EVAL_5,MaxPeriodFibonacciLFSR_1__EVAL_4,MaxPeriodFibonacciLFSR_1__EVAL_6,MaxPeriodFibonacciLFSR_1__EVAL_2,_T_243};
  assign _T_252 = _T_251[0];
  assign _T_253 = _T_251[1];
  assign _T_254 = _T_251[2];
  assign _T_255 = _T_251[3];
  assign _T_256 = _T_251[4];
  assign _T_257 = _T_251[5];
  assign _T_258 = _T_251[6];
  assign _T_259 = _T_251[7];
  assign _T_260 = _T_251[8];
  assign _T_261 = _T_251[9];
  assign _T_262 = _T_251[10];
  assign _T_263 = _T_251[11];
  assign _T_264 = _T_251[12];
  assign _T_265 = _T_251[13];
  assign _T_266 = _T_251[14];
  assign _T_267 = _T_251[15];
  assign _T_275 = {_T_260,_T_261,_T_262,_T_263,_T_264,_T_265,_T_266,_T_267};
  assign _T_283 = {_T_252,_T_253,_T_254,_T_255,_T_256,_T_257,_T_258,_T_259,_T_275};
  assign _T_284 = 16'h3fff <= _T_283;
  assign _T_286 = _T_284 | _T_233;
  assign _T_287 = auto_in_ar_valid & _T_286;
  assign _T_295_1 = Queue_9_io_enq_ready;
  assign _T_295_0 = Queue_8_io_enq_ready;
  assign _GEN_20 = auto_in_ar_bits_id ? _T_295_1 : _T_295_0;
  assign _T_292 = _T_283[1:0];
  assign _GEN_35 = {{30'd0}, _T_292};
  assign _T_297 = 2'h1 << auto_in_ar_bits_id;
  assign _T_299 = _T_297[0];
  assign _T_300 = _T_297[1];
  assign _T_305 = Queue_8_io_deq_bits_timestamp <= _T_234;
  assign _T_306 = _T_305 | _T_233;
  assign _T_307 = Queue_8_io_deq_valid & _T_306;
  assign _T_303_ready = Queue_10_io_enq_ready;
  assign _T_317 = _T_316 == 1'h0;
  assign _T_311 = Queue_9_io_deq_bits_timestamp <= _T_234;
  assign _T_312 = _T_311 | _T_233;
  assign _T_313 = Queue_9_io_deq_valid & _T_312;
  assign _T_319 = {_T_313,_T_307};
  assign _T_327 = ~ _T_326;
  assign _T_328 = _T_319 & _T_327;
  assign _T_329 = {_T_328,_T_313,_T_307};
  assign _T_330 = _T_329[3:1];
  assign _GEN_36 = {{1'd0}, _T_330};
  assign _T_331 = _T_329 | _GEN_36;
  assign _T_333 = _T_331[3:1];
  assign _T_334 = {_T_326, 2'h0};
  assign _GEN_37 = {{1'd0}, _T_333};
  assign _T_335 = _GEN_37 | _T_334;
  assign _T_336 = _T_335[3:2];
  assign _T_337 = _T_335[1:0];
  assign _T_338 = _T_336 & _T_337;
  assign _T_339 = ~ _T_338;
  assign _T_348 = _T_339[0];
  assign _T_383_0 = _T_317 ? _T_348 : _T_381_0;
  assign _T_384 = _T_303_ready & _T_383_0;
  assign _T_349 = _T_339[1];
  assign _T_383_1 = _T_317 ? _T_349 : _T_381_1;
  assign _T_385 = _T_303_ready & _T_383_1;
  assign _T_318 = _T_317 & _T_303_ready;
  assign _T_321 = _T_319 == _T_319;
  assign _T_323 = _T_321 | reset;
  assign _T_324 = _T_323 == 1'h0;
  assign _T_340 = _T_319 != 2'h0;
  assign _T_341 = _T_318 & _T_340;
  assign _T_342 = _T_339 & _T_319;
  assign _T_343 = {_T_342, 1'h0};
  assign _T_344 = _T_343[1:0];
  assign _T_345 = _T_342 | _T_344;
  assign _T_351 = _T_348 & _T_307;
  assign _T_352 = _T_349 & _T_313;
  assign _T_355 = _T_351 | _T_352;
  assign _T_357 = _T_351 == 1'h0;
  assign _T_360 = _T_352 == 1'h0;
  assign _T_361 = _T_357 | _T_360;
  assign _T_364 = _T_361 | reset;
  assign _T_365 = _T_364 == 1'h0;
  assign _T_366 = _T_307 | _T_313;
  assign _T_367 = _T_366 == 1'h0;
  assign _T_369 = _T_367 | _T_355;
  assign _T_371 = _T_369 | reset;
  assign _T_372 = _T_371 == 1'h0;
  assign _T_387 = _T_381_0 ? _T_307 : 1'h0;
  assign _T_388 = _T_381_1 ? _T_313 : 1'h0;
  assign _T_389 = _T_387 | _T_388;
  assign _T_391 = _T_317 ? _T_366 : _T_389;
  assign _T_376 = _T_303_ready & _T_391;
  assign _T_378 = _T_316 - _T_376;
  assign _T_382_0 = _T_317 ? _T_351 : _T_381_0;
  assign _T_382_1 = _T_317 ? _T_352 : _T_381_1;
  assign _T_304_bits_prot = Queue_8_io_deq_bits_data_prot;
  assign _T_304_bits_qos = Queue_8_io_deq_bits_data_qos;
  assign _T_304_bits_lock = Queue_8_io_deq_bits_data_lock;
  assign _T_304_bits_cache = Queue_8_io_deq_bits_data_cache;
  assign _T_304_bits_size = Queue_8_io_deq_bits_data_size;
  assign _T_304_bits_burst = Queue_8_io_deq_bits_data_burst;
  assign _T_304_bits_id = Queue_8_io_deq_bits_data_id;
  assign _T_304_bits_addr = Queue_8_io_deq_bits_data_addr;
  assign _T_304_bits_len = Queue_8_io_deq_bits_data_len;
  assign _T_399 = {_T_304_bits_id,_T_304_bits_addr,_T_304_bits_len,_T_304_bits_size,_T_304_bits_burst,_T_304_bits_lock,_T_304_bits_cache,_T_304_bits_prot,_T_304_bits_qos};
  assign _T_400 = _T_382_0 ? _T_399 : 56'h0;
  assign _T_310_bits_prot = Queue_9_io_deq_bits_data_prot;
  assign _T_310_bits_qos = Queue_9_io_deq_bits_data_qos;
  assign _T_310_bits_lock = Queue_9_io_deq_bits_data_lock;
  assign _T_310_bits_cache = Queue_9_io_deq_bits_data_cache;
  assign _T_310_bits_size = Queue_9_io_deq_bits_data_size;
  assign _T_310_bits_burst = Queue_9_io_deq_bits_data_burst;
  assign _T_310_bits_id = Queue_9_io_deq_bits_data_id;
  assign _T_310_bits_addr = Queue_9_io_deq_bits_data_addr;
  assign _T_310_bits_len = Queue_9_io_deq_bits_data_len;
  assign _T_408 = {_T_310_bits_id,_T_310_bits_addr,_T_310_bits_len,_T_310_bits_size,_T_310_bits_burst,_T_310_bits_lock,_T_310_bits_cache,_T_310_bits_prot,_T_310_bits_qos};
  assign _T_409 = _T_382_1 ? _T_408 : 56'h0;
  assign _T_410 = _T_400 | _T_409;
  assign _T_424 = plusarg_reader_2_out[0];
  assign _T_427 = _T_425 + 32'h1;
  assign _T_434 = {MaxPeriodFibonacciLFSR_2__EVAL_12,MaxPeriodFibonacciLFSR_2__EVAL_11,MaxPeriodFibonacciLFSR_2__EVAL_3,MaxPeriodFibonacciLFSR_2__EVAL_16,MaxPeriodFibonacciLFSR_2__EVAL_8,MaxPeriodFibonacciLFSR_2__EVAL_10,MaxPeriodFibonacciLFSR_2__EVAL_14,MaxPeriodFibonacciLFSR_2__EVAL_7};
  assign _T_442 = {MaxPeriodFibonacciLFSR_2__EVAL_0,MaxPeriodFibonacciLFSR_2__EVAL_17,MaxPeriodFibonacciLFSR_2__EVAL_1,MaxPeriodFibonacciLFSR_2__EVAL,MaxPeriodFibonacciLFSR_2__EVAL_5,MaxPeriodFibonacciLFSR_2__EVAL_4,MaxPeriodFibonacciLFSR_2__EVAL_6,MaxPeriodFibonacciLFSR_2__EVAL_2,_T_434};
  assign _T_443 = _T_442[0];
  assign _T_444 = _T_442[1];
  assign _T_445 = _T_442[2];
  assign _T_446 = _T_442[3];
  assign _T_447 = _T_442[4];
  assign _T_448 = _T_442[5];
  assign _T_449 = _T_442[6];
  assign _T_450 = _T_442[7];
  assign _T_451 = _T_442[8];
  assign _T_452 = _T_442[9];
  assign _T_453 = _T_442[10];
  assign _T_454 = _T_442[11];
  assign _T_455 = _T_442[12];
  assign _T_456 = _T_442[13];
  assign _T_457 = _T_442[14];
  assign _T_458 = _T_442[15];
  assign _T_466 = {_T_451,_T_452,_T_453,_T_454,_T_455,_T_456,_T_457,_T_458};
  assign _T_474 = {_T_443,_T_444,_T_445,_T_446,_T_447,_T_448,_T_449,_T_450,_T_466};
  assign _T_483 = _T_474[1:0];
  assign _GEN_38 = {{30'd0}, _T_483};
  assign _T_496 = Queue_11_io_deq_bits_timestamp <= _T_425;
  assign _T_497 = _T_496 | _T_424;
  assign _T_498 = Queue_11_io_deq_valid & _T_497;
  assign _T_494_ready = Queue_13_io_enq_ready;
  assign _T_508 = _T_507 == 1'h0;
  assign _T_502 = Queue_12_io_deq_bits_timestamp <= _T_425;
  assign _T_503 = _T_502 | _T_424;
  assign _T_504 = Queue_12_io_deq_valid & _T_503;
  assign _T_510 = {_T_504,_T_498};
  assign _T_518 = ~ _T_517;
  assign _T_519 = _T_510 & _T_518;
  assign _T_520 = {_T_519,_T_504,_T_498};
  assign _T_521 = _T_520[3:1];
  assign _GEN_39 = {{1'd0}, _T_521};
  assign _T_522 = _T_520 | _GEN_39;
  assign _T_524 = _T_522[3:1];
  assign _T_525 = {_T_517, 2'h0};
  assign _GEN_40 = {{1'd0}, _T_524};
  assign _T_526 = _GEN_40 | _T_525;
  assign _T_527 = _T_526[3:2];
  assign _T_528 = _T_526[1:0];
  assign _T_529 = _T_527 & _T_528;
  assign _T_530 = ~ _T_529;
  assign _T_539 = _T_530[0];
  assign _T_574_0 = _T_508 ? _T_539 : _T_572_0;
  assign _T_575 = _T_494_ready & _T_574_0;
  assign _T_540 = _T_530[1];
  assign _T_574_1 = _T_508 ? _T_540 : _T_572_1;
  assign _T_576 = _T_494_ready & _T_574_1;
  assign _T_509 = _T_508 & _T_494_ready;
  assign _T_512 = _T_510 == _T_510;
  assign _T_514 = _T_512 | reset;
  assign _T_515 = _T_514 == 1'h0;
  assign _T_531 = _T_510 != 2'h0;
  assign _T_532 = _T_509 & _T_531;
  assign _T_533 = _T_530 & _T_510;
  assign _T_534 = {_T_533, 1'h0};
  assign _T_535 = _T_534[1:0];
  assign _T_536 = _T_533 | _T_535;
  assign _T_542 = _T_539 & _T_498;
  assign _T_543 = _T_540 & _T_504;
  assign _T_546 = _T_542 | _T_543;
  assign _T_548 = _T_542 == 1'h0;
  assign _T_551 = _T_543 == 1'h0;
  assign _T_552 = _T_548 | _T_551;
  assign _T_555 = _T_552 | reset;
  assign _T_556 = _T_555 == 1'h0;
  assign _T_557 = _T_498 | _T_504;
  assign _T_558 = _T_557 == 1'h0;
  assign _T_560 = _T_558 | _T_546;
  assign _T_562 = _T_560 | reset;
  assign _T_563 = _T_562 == 1'h0;
  assign _T_578 = _T_572_0 ? _T_498 : 1'h0;
  assign _T_579 = _T_572_1 ? _T_504 : 1'h0;
  assign _T_580 = _T_578 | _T_579;
  assign _T_582 = _T_508 ? _T_557 : _T_580;
  assign _T_567 = _T_494_ready & _T_582;
  assign _T_569 = _T_507 - _T_567;
  assign _T_573_0 = _T_508 ? _T_542 : _T_572_0;
  assign _T_573_1 = _T_508 ? _T_543 : _T_572_1;
  assign _T_495_bits_id = Queue_11_io_deq_bits_data_id;
  assign _T_495_bits_resp = Queue_11_io_deq_bits_data_resp;
  assign _T_583 = {_T_495_bits_id,_T_495_bits_resp};
  assign _T_584 = _T_573_0 ? _T_583 : 3'h0;
  assign _T_501_bits_id = Queue_12_io_deq_bits_data_id;
  assign _T_501_bits_resp = Queue_12_io_deq_bits_data_resp;
  assign _T_585 = {_T_501_bits_id,_T_501_bits_resp};
  assign _T_586 = _T_573_1 ? _T_585 : 3'h0;
  assign _T_587 = _T_584 | _T_586;
  assign _T_594 = plusarg_reader_3_out[0];
  assign _T_597 = _T_595 + 32'h1;
  assign _T_604 = {MaxPeriodFibonacciLFSR_3__EVAL_12,MaxPeriodFibonacciLFSR_3__EVAL_11,MaxPeriodFibonacciLFSR_3__EVAL_3,MaxPeriodFibonacciLFSR_3__EVAL_16,MaxPeriodFibonacciLFSR_3__EVAL_8,MaxPeriodFibonacciLFSR_3__EVAL_10,MaxPeriodFibonacciLFSR_3__EVAL_14,MaxPeriodFibonacciLFSR_3__EVAL_7};
  assign _T_612 = {MaxPeriodFibonacciLFSR_3__EVAL_0,MaxPeriodFibonacciLFSR_3__EVAL_17,MaxPeriodFibonacciLFSR_3__EVAL_1,MaxPeriodFibonacciLFSR_3__EVAL,MaxPeriodFibonacciLFSR_3__EVAL_5,MaxPeriodFibonacciLFSR_3__EVAL_4,MaxPeriodFibonacciLFSR_3__EVAL_6,MaxPeriodFibonacciLFSR_3__EVAL_2,_T_604};
  assign _T_613 = _T_612[0];
  assign _T_614 = _T_612[1];
  assign _T_615 = _T_612[2];
  assign _T_616 = _T_612[3];
  assign _T_617 = _T_612[4];
  assign _T_618 = _T_612[5];
  assign _T_619 = _T_612[6];
  assign _T_620 = _T_612[7];
  assign _T_621 = _T_612[8];
  assign _T_622 = _T_612[9];
  assign _T_623 = _T_612[10];
  assign _T_624 = _T_612[11];
  assign _T_625 = _T_612[12];
  assign _T_626 = _T_612[13];
  assign _T_627 = _T_612[14];
  assign _T_628 = _T_612[15];
  assign _T_636 = {_T_621,_T_622,_T_623,_T_624,_T_625,_T_626,_T_627,_T_628};
  assign _T_644 = {_T_613,_T_614,_T_615,_T_616,_T_617,_T_618,_T_619,_T_620,_T_636};
  assign _T_653 = _T_644[1:0];
  assign _GEN_41 = {{30'd0}, _T_653};
  assign _T_666 = Queue_14_io_deq_bits_timestamp <= _T_595;
  assign _T_667 = _T_666 | _T_594;
  assign _T_668 = Queue_14_io_deq_valid & _T_667;
  assign _T_664_ready = Queue_16_io_enq_ready;
  assign _T_678 = _T_677 == 1'h0;
  assign _T_672 = Queue_15_io_deq_bits_timestamp <= _T_595;
  assign _T_673 = _T_672 | _T_594;
  assign _T_674 = Queue_15_io_deq_valid & _T_673;
  assign _T_680 = {_T_674,_T_668};
  assign _T_688 = ~ _T_687;
  assign _T_689 = _T_680 & _T_688;
  assign _T_690 = {_T_689,_T_674,_T_668};
  assign _T_691 = _T_690[3:1];
  assign _GEN_42 = {{1'd0}, _T_691};
  assign _T_692 = _T_690 | _GEN_42;
  assign _T_694 = _T_692[3:1];
  assign _T_695 = {_T_687, 2'h0};
  assign _GEN_43 = {{1'd0}, _T_694};
  assign _T_696 = _GEN_43 | _T_695;
  assign _T_697 = _T_696[3:2];
  assign _T_698 = _T_696[1:0];
  assign _T_699 = _T_697 & _T_698;
  assign _T_700 = ~ _T_699;
  assign _T_709 = _T_700[0];
  assign _T_744_0 = _T_678 ? _T_709 : _T_742_0;
  assign _T_745 = _T_664_ready & _T_744_0;
  assign _T_710 = _T_700[1];
  assign _T_744_1 = _T_678 ? _T_710 : _T_742_1;
  assign _T_746 = _T_664_ready & _T_744_1;
  assign _T_679 = _T_678 & _T_664_ready;
  assign _T_682 = _T_680 == _T_680;
  assign _T_684 = _T_682 | reset;
  assign _T_685 = _T_684 == 1'h0;
  assign _T_701 = _T_680 != 2'h0;
  assign _T_702 = _T_679 & _T_701;
  assign _T_703 = _T_700 & _T_680;
  assign _T_704 = {_T_703, 1'h0};
  assign _T_705 = _T_704[1:0];
  assign _T_706 = _T_703 | _T_705;
  assign _T_712 = _T_709 & _T_668;
  assign _T_713 = _T_710 & _T_674;
  assign _T_716 = _T_712 | _T_713;
  assign _T_718 = _T_712 == 1'h0;
  assign _T_721 = _T_713 == 1'h0;
  assign _T_722 = _T_718 | _T_721;
  assign _T_725 = _T_722 | reset;
  assign _T_726 = _T_725 == 1'h0;
  assign _T_727 = _T_668 | _T_674;
  assign _T_728 = _T_727 == 1'h0;
  assign _T_730 = _T_728 | _T_716;
  assign _T_732 = _T_730 | reset;
  assign _T_733 = _T_732 == 1'h0;
  assign _T_748 = _T_742_0 ? _T_668 : 1'h0;
  assign _T_749 = _T_742_1 ? _T_674 : 1'h0;
  assign _T_750 = _T_748 | _T_749;
  assign _T_752 = _T_678 ? _T_727 : _T_750;
  assign _T_737 = _T_664_ready & _T_752;
  assign _T_739 = _T_677 - _T_737;
  assign _T_743_0 = _T_678 ? _T_712 : _T_742_0;
  assign _T_743_1 = _T_678 ? _T_713 : _T_742_1;
  assign _T_665_bits_resp = Queue_14_io_deq_bits_data_resp;
  assign _T_665_bits_last = Queue_14_io_deq_bits_data_last;
  assign _T_665_bits_id = Queue_14_io_deq_bits_data_id;
  assign _T_665_bits_data = Queue_14_io_deq_bits_data_data;
  assign _T_755 = {_T_665_bits_id,_T_665_bits_data,_T_665_bits_resp,_T_665_bits_last};
  assign _T_756 = _T_743_0 ? _T_755 : 36'h0;
  assign _T_671_bits_resp = Queue_15_io_deq_bits_data_resp;
  assign _T_671_bits_last = Queue_15_io_deq_bits_data_last;
  assign _T_671_bits_id = Queue_15_io_deq_bits_data_id;
  assign _T_671_bits_data = Queue_15_io_deq_bits_data_data;
  assign _T_759 = {_T_671_bits_id,_T_671_bits_data,_T_671_bits_resp,_T_671_bits_last};
  assign _T_760 = _T_743_1 ? _T_759 : 36'h0;
  assign _T_761 = _T_756 | _T_760;
  assign auto_in_aw_ready = Queue_io_enq_ready & _T_65;
  assign auto_in_w_ready = _GEN_8 & _T_4_valid;
  assign auto_in_b_valid = Queue_13_io_deq_valid;
  assign auto_in_b_bits_id = Queue_13_io_deq_bits_id;
  assign auto_in_b_bits_resp = Queue_13_io_deq_bits_resp;
  assign auto_in_ar_ready = _GEN_20 & _T_286;
  assign auto_in_r_valid = Queue_16_io_deq_valid;
  assign auto_in_r_bits_id = Queue_16_io_deq_bits_id;
  assign auto_in_r_bits_data = Queue_16_io_deq_bits_data;
  assign auto_in_r_bits_resp = Queue_16_io_deq_bits_resp;
  assign auto_in_r_bits_last = Queue_16_io_deq_bits_last;
  assign auto_out_aw_valid = Queue_5_io_deq_valid;
  assign auto_out_aw_bits_id = Queue_5_io_deq_bits_id;
  assign auto_out_aw_bits_addr = Queue_5_io_deq_bits_addr;
  assign auto_out_aw_bits_len = Queue_5_io_deq_bits_len;
  assign auto_out_aw_bits_size = Queue_5_io_deq_bits_size;
  assign auto_out_aw_bits_burst = Queue_5_io_deq_bits_burst;
  assign auto_out_w_valid = _T_200_valid & _GEN_16;
  assign auto_out_w_bits_data = _T_200_bits ? _T_219_1_data : _T_219_0_data;
  assign auto_out_w_bits_strb = _T_200_bits ? _T_219_1_strb : _T_219_0_strb;
  assign auto_out_w_bits_last = _T_200_bits ? _T_219_1_last : _T_219_0_last;
  assign auto_out_b_ready = Queue_11_io_enq_ready;
  assign auto_out_ar_valid = Queue_10_io_deq_valid;
  assign auto_out_ar_bits_id = Queue_10_io_deq_bits_id;
  assign auto_out_ar_bits_addr = Queue_10_io_deq_bits_addr;
  assign auto_out_ar_bits_len = Queue_10_io_deq_bits_len;
  assign auto_out_ar_bits_size = Queue_10_io_deq_bits_size;
  assign auto_out_ar_bits_burst = Queue_10_io_deq_bits_burst;
  assign auto_out_r_ready = Queue_14_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_aw_valid & _T_65;
  assign Queue_io_enq_bits = auto_in_aw_bits_id;
  assign Queue_io_deq_ready = _T_205 & auto_in_w_valid;
  assign MaxPeriodFibonacciLFSR__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR__EVAL_9 = 1'h1;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_63 & _T_75;
  assign Queue_1_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_1_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_1_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_1_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_1_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_1_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_1_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_1_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_1_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_1_io_enq_bits_timestamp = _T_12 + _GEN_32;
  assign Queue_1_io_deq_ready = _T_160 & _T_82;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = _T_63 & _T_76;
  assign Queue_2_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_2_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_2_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_2_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_2_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_2_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_2_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_2_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_2_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_2_io_enq_bits_timestamp = _T_12 + _GEN_32;
  assign Queue_2_io_deq_ready = _T_161 & _T_88;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = _T_93 ? _T_142 : _T_165;
  assign Queue_3_io_enq_bits_id = _T_186[55];
  assign Queue_3_io_enq_bits_addr = _T_186[54:25];
  assign Queue_3_io_enq_bits_len = _T_186[24:17];
  assign Queue_3_io_enq_bits_size = _T_186[16:14];
  assign Queue_3_io_enq_bits_burst = _T_186[13:12];
  assign Queue_3_io_deq_ready = Queue_4_io_enq_ready & _T_199_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = _T_198_valid & _T_199_ready;
  assign Queue_4_io_enq_bits = Queue_3_io_deq_bits_id;
  assign Queue_4_io_deq_ready = _T_220 & auto_out_w_ready;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_5_io_enq_valid = _T_198_valid & Queue_4_io_enq_ready;
  assign Queue_5_io_enq_bits_id = Queue_3_io_deq_bits_id;
  assign Queue_5_io_enq_bits_addr = Queue_3_io_deq_bits_addr;
  assign Queue_5_io_enq_bits_len = Queue_3_io_deq_bits_len;
  assign Queue_5_io_enq_bits_size = Queue_3_io_deq_bits_size;
  assign Queue_5_io_enq_bits_burst = Queue_3_io_deq_bits_burst;
  assign Queue_5_io_deq_ready = auto_out_aw_ready;
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_6_io_enq_valid = _T_213 & _T_211;
  assign Queue_6_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_6_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_6_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_6_io_deq_ready = _T_228 & _T_226;
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_7_io_enq_valid = _T_213 & _T_212;
  assign Queue_7_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_7_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_7_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_7_io_deq_ready = _T_228 & _T_227;
  assign MaxPeriodFibonacciLFSR_1__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR_1__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR_1__EVAL_9 = 1'h1;
  assign Queue_8_clock = clock;
  assign Queue_8_reset = reset;
  assign Queue_8_io_enq_valid = _T_287 & _T_299;
  assign Queue_8_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_8_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_8_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_8_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_8_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_8_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_8_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_8_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_8_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_8_io_enq_bits_timestamp = _T_236 + _GEN_35;
  assign Queue_8_io_deq_ready = _T_384 & _T_306;
  assign Queue_9_clock = clock;
  assign Queue_9_reset = reset;
  assign Queue_9_io_enq_valid = _T_287 & _T_300;
  assign Queue_9_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_9_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_9_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_9_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_9_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_9_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_9_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_9_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_9_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_9_io_enq_bits_timestamp = _T_236 + _GEN_35;
  assign Queue_9_io_deq_ready = _T_385 & _T_312;
  assign Queue_10_clock = clock;
  assign Queue_10_reset = reset;
  assign Queue_10_io_enq_valid = _T_317 ? _T_366 : _T_389;
  assign Queue_10_io_enq_bits_id = _T_410[55];
  assign Queue_10_io_enq_bits_addr = _T_410[54:25];
  assign Queue_10_io_enq_bits_len = _T_410[24:17];
  assign Queue_10_io_enq_bits_size = _T_410[16:14];
  assign Queue_10_io_enq_bits_burst = _T_410[13:12];
  assign Queue_10_io_deq_ready = auto_out_ar_ready;
  assign MaxPeriodFibonacciLFSR_2__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR_2__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR_2__EVAL_9 = 1'h1;
  assign Queue_11_clock = clock;
  assign Queue_11_reset = reset;
  assign Queue_11_io_enq_valid = auto_out_b_valid;
  assign Queue_11_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_11_io_enq_bits_timestamp = _T_427 + _GEN_38;
  assign Queue_11_io_deq_ready = _T_575 & _T_497;
  assign Queue_12_clock = clock;
  assign Queue_12_reset = reset;
  assign Queue_12_io_enq_valid = 1'h0;
  assign Queue_12_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_12_io_enq_bits_timestamp = _T_427 + _GEN_38;
  assign Queue_12_io_deq_ready = _T_576 & _T_503;
  assign Queue_13_clock = clock;
  assign Queue_13_reset = reset;
  assign Queue_13_io_enq_valid = _T_508 ? _T_557 : _T_580;
  assign Queue_13_io_enq_bits_id = _T_587[2];
  assign Queue_13_io_enq_bits_resp = _T_587[1:0];
  assign Queue_13_io_deq_ready = auto_in_b_ready;
  assign MaxPeriodFibonacciLFSR_3__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR_3__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR_3__EVAL_9 = 1'h1;
  assign Queue_14_clock = clock;
  assign Queue_14_reset = reset;
  assign Queue_14_io_enq_valid = auto_out_r_valid;
  assign Queue_14_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_14_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_14_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_14_io_enq_bits_timestamp = _T_597 + _GEN_41;
  assign Queue_14_io_deq_ready = _T_745 & _T_667;
  assign Queue_15_clock = clock;
  assign Queue_15_reset = reset;
  assign Queue_15_io_enq_valid = 1'h0;
  assign Queue_15_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_15_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_15_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_15_io_enq_bits_timestamp = _T_597 + _GEN_41;
  assign Queue_15_io_deq_ready = _T_746 & _T_673;
  assign Queue_16_clock = clock;
  assign Queue_16_reset = reset;
  assign Queue_16_io_enq_valid = _T_678 ? _T_727 : _T_750;
  assign Queue_16_io_enq_bits_id = _T_761[35];
  assign Queue_16_io_enq_bits_data = _T_761[34:3];
  assign Queue_16_io_enq_bits_resp = _T_761[2:1];
  assign Queue_16_io_enq_bits_last = _T_761[0];
  assign Queue_16_io_deq_ready = auto_in_r_ready;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_92 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_102 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_157_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_157_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_234 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_316 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_326 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_381_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_381_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_425 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_507 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_517 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_572_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_572_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_595 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_677 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_687 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_742_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_742_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_10 <= 32'h0;
    end else begin
      _T_10 <= _T_12;
    end
    if (reset) begin
      _T_92 <= 1'h0;
    end else begin
      if (_T_94) begin
        _T_92 <= 1'h0;
      end else begin
        _T_92 <= _T_154;
      end
    end
    if (reset) begin
      _T_102 <= 2'h3;
    end else begin
      if (_T_117) begin
        _T_102 <= _T_121;
      end
    end
    if (reset) begin
      _T_157_0 <= 1'h0;
    end else begin
      if (_T_93) begin
        _T_157_0 <= _T_127;
      end
    end
    if (reset) begin
      _T_157_1 <= 1'h0;
    end else begin
      if (_T_93) begin
        _T_157_1 <= _T_128;
      end
    end
    if (reset) begin
      _T_234 <= 32'h0;
    end else begin
      _T_234 <= _T_236;
    end
    if (reset) begin
      _T_316 <= 1'h0;
    end else begin
      if (_T_318) begin
        _T_316 <= 1'h0;
      end else begin
        _T_316 <= _T_378;
      end
    end
    if (reset) begin
      _T_326 <= 2'h3;
    end else begin
      if (_T_341) begin
        _T_326 <= _T_345;
      end
    end
    if (reset) begin
      _T_381_0 <= 1'h0;
    end else begin
      if (_T_317) begin
        _T_381_0 <= _T_351;
      end
    end
    if (reset) begin
      _T_381_1 <= 1'h0;
    end else begin
      if (_T_317) begin
        _T_381_1 <= _T_352;
      end
    end
    if (reset) begin
      _T_425 <= 32'h0;
    end else begin
      _T_425 <= _T_427;
    end
    if (reset) begin
      _T_507 <= 1'h0;
    end else begin
      if (_T_509) begin
        _T_507 <= 1'h0;
      end else begin
        _T_507 <= _T_569;
      end
    end
    if (reset) begin
      _T_517 <= 2'h3;
    end else begin
      if (_T_532) begin
        _T_517 <= _T_536;
      end
    end
    if (reset) begin
      _T_572_0 <= 1'h0;
    end else begin
      if (_T_508) begin
        _T_572_0 <= _T_542;
      end
    end
    if (reset) begin
      _T_572_1 <= 1'h0;
    end else begin
      if (_T_508) begin
        _T_572_1 <= _T_543;
      end
    end
    if (reset) begin
      _T_595 <= 32'h0;
    end else begin
      _T_595 <= _T_597;
    end
    if (reset) begin
      _T_677 <= 1'h0;
    end else begin
      if (_T_679) begin
        _T_677 <= 1'h0;
      end else begin
        _T_677 <= _T_739;
      end
    end
    if (reset) begin
      _T_687 <= 2'h3;
    end else begin
      if (_T_702) begin
        _T_687 <= _T_706;
      end
    end
    if (reset) begin
      _T_742_0 <= 1'h0;
    end else begin
      if (_T_678) begin
        _T_742_0 <= _T_712;
      end
    end
    if (reset) begin
      _T_742_1 <= 1'h0;
    end else begin
      if (_T_678) begin
        _T_742_1 <= _T_713;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_141) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_148) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_324) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_365) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_372) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_372) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_515) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_515) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_556) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_563) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_563) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_685) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_685) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_726) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_726) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_733) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_733) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
