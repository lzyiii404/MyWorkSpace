//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_322_assert(
  input  [8:0]  _EVAL,
  input  [8:0]  _EVAL_1,
  input  [7:0]  _EVAL_2,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_12,
  input         _EVAL_15,
  input  [2:0]  _EVAL_17,
  input  [2:0]  _EVAL_19,
  input         _EVAL_21,
  input  [2:0]  _EVAL_26,
  input         _EVAL_30,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_36
);
  wire  TLMonitor__EVAL;
  wire [8:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire [2:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [2:0] TLMonitor__EVAL_7;
  wire [8:0] TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire [31:0] TLMonitor__EVAL_12;
  wire [7:0] TLMonitor__EVAL_13;
  wire [2:0] TLMonitor__EVAL_14;
  wire  TLMonitor__EVAL_15;
  wire [2:0] TLMonitor__EVAL_16;
  SiFive__EVAL_321_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16)
  );
  assign TLMonitor__EVAL_12 = _EVAL_8;
  assign TLMonitor__EVAL = _EVAL_6;
  assign TLMonitor__EVAL_4 = _EVAL_12;
  assign TLMonitor__EVAL_3 = _EVAL_33;
  assign TLMonitor__EVAL_5 = _EVAL_30;
  assign TLMonitor__EVAL_11 = _EVAL_5;
  assign TLMonitor__EVAL_16 = _EVAL_17;
  assign TLMonitor__EVAL_15 = _EVAL_15;
  assign TLMonitor__EVAL_2 = _EVAL_9;
  assign TLMonitor__EVAL_0 = _EVAL_1;
  assign TLMonitor__EVAL_6 = _EVAL_36;
  assign TLMonitor__EVAL_13 = _EVAL_2;
  assign TLMonitor__EVAL_8 = _EVAL;
  assign TLMonitor__EVAL_14 = _EVAL_19;
  assign TLMonitor__EVAL_7 = _EVAL_26;
  assign TLMonitor__EVAL_9 = _EVAL_21;
  assign TLMonitor__EVAL_1 = _EVAL_32;
  assign TLMonitor__EVAL_10 = _EVAL_4;

endmodule
