//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_63_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [4:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [31:0] _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  input  [4:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_62;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_68;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_72;
  reg [31:0] _RAND_2;
  reg  _EVAL_89;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_97;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_110;
  reg [31:0] _RAND_5;
  reg [5:0] _EVAL_113;
  reg [31:0] _RAND_6;
  reg  _EVAL_173;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_179;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_208;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_215;
  reg [31:0] _RAND_10;
  reg [4:0] _EVAL_276;
  reg [31:0] _RAND_11;
  reg [5:0] _EVAL_282;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_286;
  reg [31:0] _RAND_13;
  reg [5:0] _EVAL_341;
  reg [31:0] _RAND_14;
  reg [31:0] _EVAL_347;
  reg [31:0] _RAND_15;
  reg [4:0] _EVAL_358;
  reg [31:0] _RAND_16;
  wire [31:0] _EVAL_29;
  wire [32:0] _EVAL_54;
  wire [31:0] _EVAL_65;
  wire  _EVAL_80;
  wire  _EVAL_90;
  wire  _EVAL_354;
  wire  _EVAL_142;
  wire  _EVAL_202;
  wire  _EVAL_337;
  wire [32:0] _EVAL_314;
  wire [32:0] _EVAL_237;
  wire  _EVAL_216;
  wire [31:0] _EVAL_299;
  wire [32:0] _EVAL_166;
  wire [32:0] _EVAL_128;
  wire [32:0] _EVAL_108;
  wire  _EVAL_352;
  wire  _EVAL_125;
  wire [31:0] _EVAL_196;
  wire [32:0] _EVAL_288;
  wire [32:0] _EVAL_243;
  wire [32:0] _EVAL_96;
  wire  _EVAL_228;
  wire  _EVAL_51;
  wire [31:0] _EVAL_278;
  wire [32:0] _EVAL_201;
  wire [32:0] _EVAL_293;
  wire [32:0] _EVAL_88;
  wire  _EVAL_294;
  wire  _EVAL_292;
  wire [32:0] _EVAL_124;
  wire [32:0] _EVAL_265;
  wire [32:0] _EVAL_325;
  wire  _EVAL_279;
  wire  _EVAL_58;
  wire [31:0] _EVAL_167;
  wire [32:0] _EVAL_246;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_123;
  wire  _EVAL_38;
  wire  _EVAL_304;
  wire [31:0] _EVAL_268;
  wire [32:0] _EVAL_187;
  wire [32:0] _EVAL_181;
  wire [32:0] _EVAL_253;
  wire  _EVAL_99;
  wire  _EVAL_162;
  wire [31:0] _EVAL_46;
  wire [32:0] _EVAL_164;
  wire [32:0] _EVAL_194;
  wire [32:0] _EVAL_171;
  wire  _EVAL_36;
  wire  _EVAL_95;
  wire  _EVAL_44;
  wire  _EVAL_356;
  wire [31:0] _EVAL_47;
  wire [32:0] _EVAL_259;
  wire [32:0] _EVAL_195;
  wire [32:0] _EVAL_317;
  wire  _EVAL_226;
  wire  _EVAL_298;
  wire  _EVAL_78;
  wire  _EVAL_207;
  wire  _EVAL_104;
  wire  _EVAL_322;
  wire  _EVAL_45;
  wire [31:0] _EVAL_136;
  wire [31:0] _EVAL_34;
  wire  _EVAL_20;
  wire  _EVAL_241;
  wire  _EVAL_119;
  wire  _EVAL_234;
  wire  _EVAL_301;
  wire  _EVAL_61;
  wire [31:0] _EVAL_262;
  wire [31:0] _EVAL_232;
  wire  _EVAL_204;
  wire  _EVAL_93;
  wire  _EVAL_116;
  wire  _EVAL_217;
  wire  _EVAL_257;
  wire  _EVAL_158;
  wire  _EVAL_145;
  wire  _EVAL_329;
  wire  _EVAL_218;
  wire  _EVAL_26;
  wire [1:0] _EVAL_19;
  wire  _EVAL_60;
  wire  _EVAL_149;
  wire  _EVAL_281;
  wire  _EVAL_252;
  wire  _EVAL_320;
  wire  _EVAL_345;
  wire  _EVAL_236;
  wire  _EVAL_315;
  wire [31:0] _EVAL_319;
  wire [31:0] _EVAL_71;
  wire  _EVAL_40;
  wire  _EVAL_83;
  wire  _EVAL_206;
  wire  _EVAL_247;
  wire  _EVAL_326;
  wire  _EVAL_280;
  wire  _EVAL_22;
  wire  _EVAL_102;
  wire  _EVAL_190;
  wire [31:0] _EVAL_336;
  wire  _EVAL_254;
  wire  _EVAL_24;
  wire  _EVAL_227;
  wire [22:0] _EVAL_316;
  wire [7:0] _EVAL_107;
  wire [7:0] _EVAL_305;
  wire [5:0] _EVAL_342;
  wire [5:0] _EVAL_184;
  wire  _EVAL_94;
  wire  _EVAL_115;
  wire  _EVAL_250;
  wire  _EVAL_175;
  wire  _EVAL_147;
  wire  _EVAL_235;
  wire  _EVAL_77;
  wire  _EVAL_66;
  wire  _EVAL_85;
  wire  _EVAL_308;
  wire  _EVAL_284;
  wire [1:0] _EVAL_300;
  wire [1:0] _EVAL_210;
  wire  _EVAL_258;
  wire [3:0] _EVAL_172;
  wire  _EVAL_238;
  wire  _EVAL_303;
  wire  _EVAL_63;
  wire  _EVAL_30;
  wire  _EVAL_69;
  wire  _EVAL_255;
  wire  _EVAL_333;
  wire  _EVAL_28;
  wire  _EVAL_39;
  wire  _EVAL_127;
  wire  _EVAL_87;
  wire  _EVAL_209;
  wire  _EVAL_214;
  wire  _EVAL_321;
  wire  _EVAL_150;
  wire  _EVAL_200;
  wire  _EVAL_283;
  wire  _EVAL_343;
  wire  _EVAL_248;
  wire  _EVAL_188;
  wire [1:0] _EVAL_106;
  wire  _EVAL_165;
  wire  _EVAL_230;
  wire  _EVAL_355;
  wire  _EVAL_312;
  wire  _EVAL_327;
  wire  _EVAL_178;
  wire  _EVAL_224;
  wire  _EVAL_273;
  wire  _EVAL_122;
  wire  _EVAL_211;
  wire  _EVAL_153;
  wire  _EVAL_244;
  wire  _EVAL_161;
  wire  _EVAL_213;
  wire  _EVAL_48;
  wire  _EVAL_130;
  wire  _EVAL_331;
  wire  _EVAL_290;
  wire  _EVAL_82;
  wire  _EVAL_43;
  wire  _EVAL_21;
  wire  _EVAL_186;
  wire  _EVAL_306;
  wire  _EVAL_353;
  wire  _EVAL_318;
  wire  _EVAL_339;
  wire  _EVAL_260;
  wire [3:0] _EVAL_239;
  wire [3:0] _EVAL_357;
  wire [3:0] _EVAL_267;
  wire  _EVAL_240;
  wire  _EVAL_131;
  wire  _EVAL_140;
  wire  _EVAL_148;
  wire  _EVAL_160;
  wire  _EVAL_197;
  wire  _EVAL_137;
  wire  _EVAL_275;
  wire  _EVAL_157;
  wire  _EVAL_291;
  wire  _EVAL_219;
  wire  _EVAL_330;
  wire  _EVAL_338;
  wire  _EVAL_135;
  wire  _EVAL_121;
  wire [22:0] _EVAL_328;
  wire [7:0] _EVAL_302;
  wire [7:0] _EVAL_350;
  wire  _EVAL_49;
  wire  _EVAL_192;
  wire  _EVAL_134;
  wire  _EVAL_351;
  wire [5:0] _EVAL_203;
  wire  _EVAL_139;
  wire  _EVAL_79;
  wire  _EVAL_155;
  wire  _EVAL_53;
  wire  _EVAL_245;
  wire  _EVAL_27;
  wire  _EVAL_92;
  wire  _EVAL_118;
  wire  _EVAL_289;
  wire  _EVAL_74;
  wire  _EVAL_205;
  wire  _EVAL_231;
  wire  _EVAL_266;
  wire  _EVAL_311;
  wire [31:0] _EVAL_223;
  wire [31:0] _EVAL_109;
  wire  _EVAL_120;
  wire  _EVAL_117;
  wire  _EVAL_222;
  wire  _EVAL_42;
  wire  _EVAL_183;
  wire  _EVAL_277;
  wire  _EVAL_346;
  wire  _EVAL_169;
  wire  _EVAL_274;
  wire  _EVAL_272;
  wire  _EVAL_324;
  wire  _EVAL_31;
  wire  _EVAL_98;
  wire  _EVAL_198;
  wire  _EVAL_310;
  wire  _EVAL_271;
  wire  _EVAL_100;
  wire  _EVAL_86;
  wire  _EVAL_309;
  wire  _EVAL_152;
  wire  _EVAL_159;
  wire  _EVAL_182;
  wire  _EVAL_105;
  wire  _EVAL_91;
  wire  _EVAL_307;
  wire  _EVAL_193;
  wire  _EVAL_249;
  wire  _EVAL_103;
  wire  _EVAL_111;
  wire  _EVAL_269;
  wire  _EVAL_23;
  wire  _EVAL_70;
  wire  _EVAL_56;
  wire [31:0] _EVAL_76;
  wire  _EVAL_334;
  wire  _EVAL_256;
  wire  _EVAL_220;
  wire  _EVAL_344;
  wire  _EVAL_251;
  wire  _EVAL_132;
  wire  _EVAL_189;
  wire  _EVAL_185;
  wire [5:0] _EVAL_112;
  wire  _EVAL_270;
  wire  _EVAL_313;
  wire  _EVAL_323;
  wire  _EVAL_138;
  wire  _EVAL_154;
  wire  _EVAL_126;
  wire  _EVAL_332;
  wire  _EVAL_295;
  wire  _EVAL_146;
  wire  _EVAL_229;
  wire [31:0] _EVAL_64;
  wire [31:0] _EVAL_55;
  wire  _EVAL_129;
  wire  _EVAL_296;
  wire  _EVAL_177;
  wire  _EVAL_168;
  wire  _EVAL_263;
  wire  _EVAL_151;
  wire  _EVAL_174;
  wire  _EVAL_348;
  wire  _EVAL_261;
  wire  _EVAL_143;
  wire  _EVAL_297;
  wire  _EVAL_141;
  wire  _EVAL_73;
  wire [5:0] _EVAL_349;
  wire  _EVAL_340;
  wire  _EVAL_114;
  wire [5:0] _EVAL_144;
  wire  _EVAL_37;
  wire  _EVAL_52;
  wire  _EVAL_84;
  wire  _EVAL_335;
  wire  _EVAL_191;
  wire  _EVAL_212;
  wire  _EVAL_180;
  wire  _EVAL_156;
  wire  _EVAL_57;
  wire  _EVAL_264;
  wire  _EVAL_233;
  wire  _EVAL_285;
  wire  _EVAL_41;
  wire  _EVAL_50;
  wire  _EVAL_133;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_29 = _EVAL_15 ^ 32'h40000000;
  assign _EVAL_54 = {1'b0,$signed(_EVAL_29)};
  assign _EVAL_65 = _EVAL_68 >> _EVAL_12;
  assign _EVAL_80 = _EVAL_65[0];
  assign _EVAL_90 = _EVAL_80 == 1'h0;
  assign _EVAL_354 = _EVAL_90 | _EVAL_17;
  assign _EVAL_142 = _EVAL_354 == 1'h0;
  assign _EVAL_202 = _EVAL_2 <= 2'h2;
  assign _EVAL_337 = _EVAL_16 <= 4'h6;
  assign _EVAL_314 = $signed(_EVAL_54) & $signed(-33'sh2000);
  assign _EVAL_237 = $signed(_EVAL_314);
  assign _EVAL_216 = $signed(_EVAL_237) == $signed(33'sh0);
  assign _EVAL_299 = _EVAL_15 ^ 32'h80000000;
  assign _EVAL_166 = {1'b0,$signed(_EVAL_299)};
  assign _EVAL_128 = $signed(_EVAL_166) & $signed(-33'sh20000);
  assign _EVAL_108 = $signed(_EVAL_128);
  assign _EVAL_352 = $signed(_EVAL_108) == $signed(33'sh0);
  assign _EVAL_125 = _EVAL_216 | _EVAL_352;
  assign _EVAL_196 = _EVAL_15 ^ 32'hc000000;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_196)};
  assign _EVAL_243 = $signed(_EVAL_288) & $signed(-33'sh4000000);
  assign _EVAL_96 = $signed(_EVAL_243);
  assign _EVAL_228 = $signed(_EVAL_96) == $signed(33'sh0);
  assign _EVAL_51 = _EVAL_125 | _EVAL_228;
  assign _EVAL_278 = _EVAL_15 ^ 32'h2000000;
  assign _EVAL_201 = {1'b0,$signed(_EVAL_278)};
  assign _EVAL_293 = $signed(_EVAL_201) & $signed(-33'sh10000);
  assign _EVAL_88 = $signed(_EVAL_293);
  assign _EVAL_294 = $signed(_EVAL_88) == $signed(33'sh0);
  assign _EVAL_292 = _EVAL_51 | _EVAL_294;
  assign _EVAL_124 = {1'b0,$signed(_EVAL_15)};
  assign _EVAL_265 = $signed(_EVAL_124) & $signed(-33'sh5000);
  assign _EVAL_325 = $signed(_EVAL_265);
  assign _EVAL_279 = $signed(_EVAL_325) == $signed(33'sh0);
  assign _EVAL_58 = _EVAL_292 | _EVAL_279;
  assign _EVAL_167 = _EVAL_15 ^ 32'h1800000;
  assign _EVAL_246 = {1'b0,$signed(_EVAL_167)};
  assign _EVAL_163 = $signed(_EVAL_246) & $signed(-33'sh8000);
  assign _EVAL_123 = $signed(_EVAL_163);
  assign _EVAL_38 = $signed(_EVAL_123) == $signed(33'sh0);
  assign _EVAL_304 = _EVAL_58 | _EVAL_38;
  assign _EVAL_268 = _EVAL_15 ^ 32'h1900000;
  assign _EVAL_187 = {1'b0,$signed(_EVAL_268)};
  assign _EVAL_181 = $signed(_EVAL_187) & $signed(-33'sh2000);
  assign _EVAL_253 = $signed(_EVAL_181);
  assign _EVAL_99 = $signed(_EVAL_253) == $signed(33'sh0);
  assign _EVAL_162 = _EVAL_304 | _EVAL_99;
  assign _EVAL_46 = _EVAL_15 ^ 32'h20000000;
  assign _EVAL_164 = {1'b0,$signed(_EVAL_46)};
  assign _EVAL_194 = $signed(_EVAL_164) & $signed(-33'sh2000);
  assign _EVAL_171 = $signed(_EVAL_194);
  assign _EVAL_36 = $signed(_EVAL_171) == $signed(33'sh0);
  assign _EVAL_95 = _EVAL_162 | _EVAL_36;
  assign _EVAL_44 = _EVAL_337 & _EVAL_95;
  assign _EVAL_356 = _EVAL_16 <= 4'h8;
  assign _EVAL_47 = _EVAL_15 ^ 32'h3000;
  assign _EVAL_259 = {1'b0,$signed(_EVAL_47)};
  assign _EVAL_195 = $signed(_EVAL_259) & $signed(-33'sh1000);
  assign _EVAL_317 = $signed(_EVAL_195);
  assign _EVAL_226 = $signed(_EVAL_317) == $signed(33'sh0);
  assign _EVAL_298 = _EVAL_356 & _EVAL_226;
  assign _EVAL_78 = _EVAL_44 | _EVAL_298;
  assign _EVAL_207 = _EVAL_78 | _EVAL_17;
  assign _EVAL_104 = _EVAL_13 & _EVAL_11;
  assign _EVAL_322 = _EVAL_72 == 6'h0;
  assign _EVAL_45 = _EVAL_104 & _EVAL_322;
  assign _EVAL_136 = 32'h1 << _EVAL_12;
  assign _EVAL_34 = _EVAL_45 ? _EVAL_136 : 32'h0;
  assign _EVAL_20 = _EVAL_6 & _EVAL_7;
  assign _EVAL_241 = _EVAL_113 == 6'h0;
  assign _EVAL_119 = _EVAL_20 & _EVAL_241;
  assign _EVAL_234 = _EVAL_5 == 3'h6;
  assign _EVAL_301 = _EVAL_234 == 1'h0;
  assign _EVAL_61 = _EVAL_119 & _EVAL_301;
  assign _EVAL_262 = 32'h1 << _EVAL_18;
  assign _EVAL_232 = _EVAL_61 ? _EVAL_262 : 32'h0;
  assign _EVAL_204 = _EVAL_34 != _EVAL_232;
  assign _EVAL_93 = _EVAL_34 != 32'h0;
  assign _EVAL_116 = _EVAL_93 == 1'h0;
  assign _EVAL_217 = _EVAL_204 | _EVAL_116;
  assign _EVAL_257 = _EVAL_217 | _EVAL_17;
  assign _EVAL_158 = _EVAL_4 == 3'h1;
  assign _EVAL_145 = _EVAL_337 & _EVAL_352;
  assign _EVAL_329 = _EVAL_145 | _EVAL_17;
  assign _EVAL_218 = _EVAL_4 == _EVAL_62;
  assign _EVAL_26 = _EVAL_3 <= 3'h3;
  assign _EVAL_19 = _EVAL_18[4:3];
  assign _EVAL_60 = _EVAL_19 == 2'h0;
  assign _EVAL_149 = _EVAL_19 == 2'h1;
  assign _EVAL_281 = _EVAL_60 | _EVAL_149;
  assign _EVAL_252 = _EVAL_19 == 2'h2;
  assign _EVAL_320 = _EVAL_281 | _EVAL_252;
  assign _EVAL_345 = _EVAL_19 == 2'h3;
  assign _EVAL_236 = _EVAL_320 | _EVAL_345;
  assign _EVAL_315 = _EVAL_236 | _EVAL_17;
  assign _EVAL_319 = _EVAL_34 | _EVAL_68;
  assign _EVAL_71 = _EVAL_319 >> _EVAL_18;
  assign _EVAL_40 = _EVAL_71[0];
  assign _EVAL_83 = _EVAL_5 <= 3'h6;
  assign _EVAL_206 = _EVAL_83 | _EVAL_17;
  assign _EVAL_247 = _EVAL_17 == 1'h0;
  assign _EVAL_326 = _EVAL_11 & _EVAL_158;
  assign _EVAL_280 = _EVAL_16[0];
  assign _EVAL_22 = _EVAL_9 == _EVAL_215;
  assign _EVAL_102 = _EVAL_22 | _EVAL_17;
  assign _EVAL_190 = _EVAL_104 | _EVAL_20;
  assign _EVAL_336 = _EVAL_286 + 32'h1;
  assign _EVAL_254 = _EVAL_282 == 6'h0;
  assign _EVAL_24 = _EVAL_341 == 6'h0;
  assign _EVAL_227 = _EVAL_5[0];
  assign _EVAL_316 = 23'hff << _EVAL_9;
  assign _EVAL_107 = _EVAL_316[7:0];
  assign _EVAL_305 = ~ _EVAL_107;
  assign _EVAL_342 = _EVAL_305[7:2];
  assign _EVAL_184 = _EVAL_341 - 6'h1;
  assign _EVAL_94 = _EVAL_18 == _EVAL_276;
  assign _EVAL_115 = _EVAL_16 <= 4'h2;
  assign _EVAL_250 = _EVAL_226 | _EVAL_228;
  assign _EVAL_175 = _EVAL_250 | _EVAL_294;
  assign _EVAL_147 = _EVAL_175 | _EVAL_279;
  assign _EVAL_235 = _EVAL_147 | _EVAL_38;
  assign _EVAL_77 = _EVAL_235 | _EVAL_99;
  assign _EVAL_66 = _EVAL_77 | _EVAL_36;
  assign _EVAL_85 = _EVAL_115 & _EVAL_66;
  assign _EVAL_308 = _EVAL_85 | _EVAL_17;
  assign _EVAL_284 = _EVAL_308 == 1'h0;
  assign _EVAL_300 = 2'h1 << _EVAL_280;
  assign _EVAL_210 = _EVAL_300 | 2'h1;
  assign _EVAL_258 = _EVAL_210[1];
  assign _EVAL_172 = ~ _EVAL_8;
  assign _EVAL_238 = _EVAL_172 == 4'h0;
  assign _EVAL_303 = _EVAL_238 | _EVAL_17;
  assign _EVAL_63 = _EVAL_303 == 1'h0;
  assign _EVAL_30 = _EVAL_15[1];
  assign _EVAL_69 = _EVAL_15[0];
  assign _EVAL_255 = _EVAL_30 & _EVAL_69;
  assign _EVAL_333 = _EVAL_3 == _EVAL_110;
  assign _EVAL_28 = _EVAL_333 | _EVAL_17;
  assign _EVAL_39 = _EVAL_15 == _EVAL_347;
  assign _EVAL_127 = _EVAL_39 | _EVAL_17;
  assign _EVAL_87 = _EVAL_127 == 1'h0;
  assign _EVAL_209 = _EVAL_4 == 3'h2;
  assign _EVAL_214 = _EVAL_26 | _EVAL_17;
  assign _EVAL_321 = _EVAL_214 == 1'h0;
  assign _EVAL_150 = _EVAL_30 == 1'h0;
  assign _EVAL_200 = _EVAL_3 <= 3'h4;
  assign _EVAL_283 = _EVAL_200 | _EVAL_17;
  assign _EVAL_343 = _EVAL_283 == 1'h0;
  assign _EVAL_248 = _EVAL_4[2];
  assign _EVAL_188 = _EVAL_298 | _EVAL_17;
  assign _EVAL_106 = _EVAL_12[4:3];
  assign _EVAL_165 = _EVAL_106 == 2'h0;
  assign _EVAL_230 = _EVAL_106 == 2'h1;
  assign _EVAL_355 = _EVAL_165 | _EVAL_230;
  assign _EVAL_312 = _EVAL_106 == 2'h2;
  assign _EVAL_327 = _EVAL_355 | _EVAL_312;
  assign _EVAL_178 = _EVAL_106 == 2'h3;
  assign _EVAL_224 = _EVAL_327 | _EVAL_178;
  assign _EVAL_273 = _EVAL_224 | _EVAL_17;
  assign _EVAL_122 = _EVAL_254 == 1'h0;
  assign _EVAL_211 = _EVAL_16 >= 4'h2;
  assign _EVAL_153 = _EVAL_258 & _EVAL_30;
  assign _EVAL_244 = _EVAL_211 | _EVAL_153;
  assign _EVAL_161 = _EVAL_210[0];
  assign _EVAL_213 = _EVAL_161 & _EVAL_255;
  assign _EVAL_48 = _EVAL_244 | _EVAL_213;
  assign _EVAL_130 = _EVAL_69 == 1'h0;
  assign _EVAL_331 = _EVAL_30 & _EVAL_130;
  assign _EVAL_290 = _EVAL_161 & _EVAL_331;
  assign _EVAL_82 = _EVAL_244 | _EVAL_290;
  assign _EVAL_43 = _EVAL_258 & _EVAL_150;
  assign _EVAL_21 = _EVAL_211 | _EVAL_43;
  assign _EVAL_186 = _EVAL_150 & _EVAL_69;
  assign _EVAL_306 = _EVAL_161 & _EVAL_186;
  assign _EVAL_353 = _EVAL_21 | _EVAL_306;
  assign _EVAL_318 = _EVAL_150 & _EVAL_130;
  assign _EVAL_339 = _EVAL_161 & _EVAL_318;
  assign _EVAL_260 = _EVAL_21 | _EVAL_339;
  assign _EVAL_239 = {_EVAL_48,_EVAL_82,_EVAL_353,_EVAL_260};
  assign _EVAL_357 = ~ _EVAL_239;
  assign _EVAL_267 = _EVAL_8 & _EVAL_357;
  assign _EVAL_240 = _EVAL_5 == 3'h0;
  assign _EVAL_131 = _EVAL_40 | _EVAL_17;
  assign _EVAL_140 = _EVAL_131 == 1'h0;
  assign _EVAL_148 = _EVAL_2 != 2'h2;
  assign _EVAL_160 = _EVAL_5 == 3'h5;
  assign _EVAL_197 = _EVAL_7 & _EVAL_160;
  assign _EVAL_137 = _EVAL_16 == _EVAL_208;
  assign _EVAL_275 = _EVAL_4 == 3'h5;
  assign _EVAL_157 = _EVAL_267 == 4'h0;
  assign _EVAL_291 = _EVAL_68 != 32'h0;
  assign _EVAL_219 = _EVAL_291 == 1'h0;
  assign _EVAL_330 = plusarg_reader_out == 32'h0;
  assign _EVAL_338 = _EVAL_219 | _EVAL_330;
  assign _EVAL_135 = _EVAL_286 < plusarg_reader_out;
  assign _EVAL_121 = _EVAL_338 | _EVAL_135;
  assign _EVAL_328 = 23'hff << _EVAL_16;
  assign _EVAL_302 = _EVAL_328[7:0];
  assign _EVAL_350 = ~ _EVAL_302;
  assign _EVAL_49 = _EVAL_5 == _EVAL_97;
  assign _EVAL_192 = _EVAL_49 | _EVAL_17;
  assign _EVAL_134 = _EVAL_192 == 1'h0;
  assign _EVAL_351 = _EVAL_137 | _EVAL_17;
  assign _EVAL_203 = _EVAL_350[7:2];
  assign _EVAL_139 = _EVAL_0 == 1'h0;
  assign _EVAL_79 = _EVAL_10 == 1'h0;
  assign _EVAL_155 = _EVAL_79 | _EVAL_17;
  assign _EVAL_53 = _EVAL_155 == 1'h0;
  assign _EVAL_245 = _EVAL_1 == 1'h0;
  assign _EVAL_27 = _EVAL_245 | _EVAL_17;
  assign _EVAL_92 = _EVAL_27 == 1'h0;
  assign _EVAL_118 = _EVAL_2 == _EVAL_179;
  assign _EVAL_289 = _EVAL_118 | _EVAL_17;
  assign _EVAL_74 = _EVAL_202 | _EVAL_17;
  assign _EVAL_205 = _EVAL_74 == 1'h0;
  assign _EVAL_231 = _EVAL_157 | _EVAL_17;
  assign _EVAL_266 = _EVAL_4 == 3'h3;
  assign _EVAL_311 = _EVAL_11 & _EVAL_266;
  assign _EVAL_223 = {{24'd0}, _EVAL_350};
  assign _EVAL_109 = _EVAL_15 & _EVAL_223;
  assign _EVAL_120 = _EVAL_211 | _EVAL_17;
  assign _EVAL_117 = _EVAL_120 == 1'h0;
  assign _EVAL_222 = _EVAL_248 == 1'h0;
  assign _EVAL_42 = _EVAL_109 == 32'h0;
  assign _EVAL_183 = _EVAL_42 | _EVAL_17;
  assign _EVAL_277 = _EVAL_14 == _EVAL_89;
  assign _EVAL_346 = _EVAL_277 | _EVAL_17;
  assign _EVAL_169 = _EVAL_2 == 2'h0;
  assign _EVAL_274 = _EVAL_169 | _EVAL_17;
  assign _EVAL_272 = _EVAL_121 | _EVAL_17;
  assign _EVAL_324 = _EVAL_4 == 3'h0;
  assign _EVAL_31 = _EVAL_11 & _EVAL_324;
  assign _EVAL_98 = _EVAL_207 == 1'h0;
  assign _EVAL_198 = _EVAL_12 == _EVAL_358;
  assign _EVAL_310 = _EVAL_198 | _EVAL_17;
  assign _EVAL_271 = _EVAL_310 == 1'h0;
  assign _EVAL_100 = _EVAL_9 >= 4'h2;
  assign _EVAL_86 = _EVAL_100 | _EVAL_17;
  assign _EVAL_309 = _EVAL_86 == 1'h0;
  assign _EVAL_152 = _EVAL_8 == _EVAL_239;
  assign _EVAL_159 = _EVAL_152 | _EVAL_17;
  assign _EVAL_182 = _EVAL_159 == 1'h0;
  assign _EVAL_105 = _EVAL_218 | _EVAL_17;
  assign _EVAL_91 = _EVAL_28 == 1'h0;
  assign _EVAL_307 = _EVAL_4 == 3'h6;
  assign _EVAL_193 = _EVAL_11 & _EVAL_307;
  assign _EVAL_249 = _EVAL_4 == 3'h7;
  assign _EVAL_103 = _EVAL_11 & _EVAL_249;
  assign _EVAL_111 = _EVAL_139 | _EVAL_17;
  assign _EVAL_269 = _EVAL_111 == 1'h0;
  assign _EVAL_23 = _EVAL_3 != 3'h0;
  assign _EVAL_70 = _EVAL_329 == 1'h0;
  assign _EVAL_56 = _EVAL_351 == 1'h0;
  assign _EVAL_76 = ~ _EVAL_232;
  assign _EVAL_334 = _EVAL_231 == 1'h0;
  assign _EVAL_256 = _EVAL_104 & _EVAL_254;
  assign _EVAL_220 = _EVAL_3 <= 3'h2;
  assign _EVAL_344 = _EVAL_220 | _EVAL_17;
  assign _EVAL_251 = _EVAL_344 == 1'h0;
  assign _EVAL_132 = _EVAL_139 | _EVAL_10;
  assign _EVAL_189 = _EVAL_132 | _EVAL_17;
  assign _EVAL_185 = _EVAL_189 == 1'h0;
  assign _EVAL_112 = _EVAL_72 - 6'h1;
  assign _EVAL_270 = _EVAL_24 == 1'h0;
  assign _EVAL_313 = _EVAL_7 & _EVAL_270;
  assign _EVAL_323 = _EVAL_346 == 1'h0;
  assign _EVAL_138 = _EVAL_94 | _EVAL_17;
  assign _EVAL_154 = _EVAL_138 == 1'h0;
  assign _EVAL_126 = _EVAL_7 & _EVAL_234;
  assign _EVAL_332 = _EVAL_289 == 1'h0;
  assign _EVAL_295 = _EVAL_188 == 1'h0;
  assign _EVAL_146 = _EVAL_20 & _EVAL_24;
  assign _EVAL_229 = _EVAL_11 & _EVAL_275;
  assign _EVAL_64 = _EVAL_68 | _EVAL_34;
  assign _EVAL_55 = _EVAL_64 & _EVAL_76;
  assign _EVAL_129 = _EVAL_23 | _EVAL_17;
  assign _EVAL_296 = _EVAL_129 == 1'h0;
  assign _EVAL_177 = _EVAL_4 == 3'h4;
  assign _EVAL_168 = _EVAL_0 == _EVAL_173;
  assign _EVAL_263 = _EVAL_168 | _EVAL_17;
  assign _EVAL_151 = _EVAL_263 == 1'h0;
  assign _EVAL_174 = _EVAL_148 | _EVAL_17;
  assign _EVAL_348 = _EVAL_174 == 1'h0;
  assign _EVAL_261 = _EVAL_11 & _EVAL_209;
  assign _EVAL_143 = _EVAL_274 == 1'h0;
  assign _EVAL_297 = _EVAL_102 == 1'h0;
  assign _EVAL_141 = _EVAL_206 == 1'h0;
  assign _EVAL_73 = _EVAL_5 == 3'h2;
  assign _EVAL_349 = _EVAL_282 - 6'h1;
  assign _EVAL_340 = _EVAL_5 == 3'h1;
  assign _EVAL_114 = _EVAL_7 & _EVAL_340;
  assign _EVAL_144 = _EVAL_113 - 6'h1;
  assign _EVAL_37 = _EVAL_272 == 1'h0;
  assign _EVAL_52 = _EVAL_7 & _EVAL_240;
  assign _EVAL_84 = _EVAL_3 == 3'h0;
  assign _EVAL_335 = _EVAL_5 == 3'h4;
  assign _EVAL_191 = _EVAL_7 & _EVAL_335;
  assign _EVAL_212 = _EVAL_84 | _EVAL_17;
  assign _EVAL_180 = _EVAL_212 == 1'h0;
  assign _EVAL_156 = _EVAL_315 == 1'h0;
  assign _EVAL_57 = _EVAL_7 & _EVAL_73;
  assign _EVAL_264 = _EVAL_105 == 1'h0;
  assign _EVAL_233 = _EVAL_273 == 1'h0;
  assign _EVAL_285 = _EVAL_257 == 1'h0;
  assign _EVAL_41 = _EVAL_183 == 1'h0;
  assign _EVAL_50 = _EVAL_11 & _EVAL_177;
  assign _EVAL_133 = _EVAL_11 & _EVAL_122;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_62 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_68 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_72 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_89 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_97 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_110 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_113 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_173 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_179 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_208 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_215 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_276 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_282 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_286 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_341 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_347 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_358 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_256) begin
      _EVAL_62 <= _EVAL_4;
    end
    if (_EVAL_17) begin
      _EVAL_68 <= 32'h0;
    end else begin
      _EVAL_68 <= _EVAL_55;
    end
    if (_EVAL_17) begin
      _EVAL_72 <= 6'h0;
    end else begin
      if (_EVAL_104) begin
        if (_EVAL_322) begin
          if (_EVAL_222) begin
            _EVAL_72 <= _EVAL_203;
          end else begin
            _EVAL_72 <= 6'h0;
          end
        end else begin
          _EVAL_72 <= _EVAL_112;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_89 <= _EVAL_14;
    end
    if (_EVAL_146) begin
      _EVAL_97 <= _EVAL_5;
    end
    if (_EVAL_256) begin
      _EVAL_110 <= _EVAL_3;
    end
    if (_EVAL_17) begin
      _EVAL_113 <= 6'h0;
    end else begin
      if (_EVAL_20) begin
        if (_EVAL_241) begin
          if (_EVAL_227) begin
            _EVAL_113 <= _EVAL_342;
          end else begin
            _EVAL_113 <= 6'h0;
          end
        end else begin
          _EVAL_113 <= _EVAL_144;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_173 <= _EVAL_0;
    end
    if (_EVAL_146) begin
      _EVAL_179 <= _EVAL_2;
    end
    if (_EVAL_256) begin
      _EVAL_208 <= _EVAL_16;
    end
    if (_EVAL_146) begin
      _EVAL_215 <= _EVAL_9;
    end
    if (_EVAL_146) begin
      _EVAL_276 <= _EVAL_18;
    end
    if (_EVAL_17) begin
      _EVAL_282 <= 6'h0;
    end else begin
      if (_EVAL_104) begin
        if (_EVAL_254) begin
          if (_EVAL_222) begin
            _EVAL_282 <= _EVAL_203;
          end else begin
            _EVAL_282 <= 6'h0;
          end
        end else begin
          _EVAL_282 <= _EVAL_349;
        end
      end
    end
    if (_EVAL_17) begin
      _EVAL_286 <= 32'h0;
    end else begin
      if (_EVAL_190) begin
        _EVAL_286 <= 32'h0;
      end else begin
        _EVAL_286 <= _EVAL_336;
      end
    end
    if (_EVAL_17) begin
      _EVAL_341 <= 6'h0;
    end else begin
      if (_EVAL_20) begin
        if (_EVAL_24) begin
          if (_EVAL_227) begin
            _EVAL_341 <= _EVAL_342;
          end else begin
            _EVAL_341 <= 6'h0;
          end
        end else begin
          _EVAL_341 <= _EVAL_184;
        end
      end
    end
    if (_EVAL_256) begin
      _EVAL_347 <= _EVAL_15;
    end
    if (_EVAL_256) begin
      _EVAL_358 <= _EVAL_12;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1dd550e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(660b30be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a23ea2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9042e666)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71458110)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c5212f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de3339e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da218473)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(202a215d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f95bbebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79134b6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cacc5850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef572148)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678b46f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_334) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bedb786)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_332) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d768650f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bac23fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88d37b13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f21c4e2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa14d889)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca10ea70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e952bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4951dd6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2866091f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc1ef5d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6ffaecb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2abe3d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(550155a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de9d9679)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bce4f4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a71d052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4800919a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cf0fd7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30ba5fcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8306b55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(490cd8c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee4e639e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_343) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9d5f800)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f5e6a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b502d2a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f255773e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ec6b862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(789e9b9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fcb015e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fe81767)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd4ca62b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9e0bad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(403cc4f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ed7eb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59b245c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28a140c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb1ec8ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce402863)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(759bde87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38a54e07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bae2349)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65f9ab85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa454c69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(703be1f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca7a317b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a90676b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(691d23fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72736b86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4185a999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(954f6433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(625f2f75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ddbed9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(102af7fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16b65b29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ebe1894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(836e2418)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4315dc09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae982efe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d56af879)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c96992f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(136f27fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7dac0dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fca77980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(498dab41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d4e40ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90ec5dd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93f1638)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_343) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e80abd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73265b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bd65dac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a35bfae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eecdcb93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38a7a3f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
