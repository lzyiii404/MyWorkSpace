//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_276(
  output        _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  output [6:0]  _EVAL_3,
  output        _EVAL_4,
  output [2:0]  _EVAL_5,
  output [31:0] _EVAL_6,
  output [6:0]  _EVAL_7,
  output [1:0]  _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  output [1:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output [31:0] _EVAL_15,
  output        _EVAL_16,
  output [2:0]  _EVAL_17,
  input  [6:0]  _EVAL_18,
  input  [1:0]  _EVAL_19,
  input  [2:0]  _EVAL_20,
  output        _EVAL_21,
  input  [31:0] _EVAL_22,
  output [1:0]  _EVAL_23,
  output        _EVAL_24,
  input  [1:0]  _EVAL_25,
  output        _EVAL_26,
  output [2:0]  _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30
);
  reg [1:0] _EVAL_32;
  reg [31:0] _RAND_0;
  reg  _EVAL_34;
  reg [31:0] _RAND_1;
  reg  _EVAL_39;
  reg [31:0] _RAND_2;
  reg [6:0] _EVAL_40;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_46;
  reg [31:0] _RAND_4;
  reg [31:0] _EVAL_47;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_48;
  reg [31:0] _RAND_6;
  reg  _EVAL_49;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_50;
  reg [31:0] _RAND_8;
  wire  _EVAL_36;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_45;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [1:0] _EVAL_35;
  assign _EVAL_36 = _EVAL_46[1];
  assign _EVAL_51 = _EVAL_36 == 1'h0;
  assign _EVAL_52 = _EVAL_46 == _EVAL_19;
  assign _EVAL_45 = _EVAL_19[0];
  assign _EVAL_41 = _EVAL_36 != _EVAL_45;
  assign _EVAL_42 = _EVAL_26 & _EVAL_28;
  assign _EVAL_43 = _EVAL_46[0];
  assign _EVAL_35 = {_EVAL_43,_EVAL_51};
  assign _EVAL_17 = _EVAL_48;
  assign _EVAL_26 = _EVAL_52 ? _EVAL_13 : _EVAL_41;
  assign _EVAL_12 = _EVAL_46;
  assign _EVAL_4 = _EVAL_29;
  assign _EVAL_3 = _EVAL_18;
  assign _EVAL_7 = _EVAL_40;
  assign _EVAL_30 = _EVAL_20;
  assign _EVAL_27 = _EVAL_2;
  assign _EVAL_16 = _EVAL_0;
  assign _EVAL_9 = _EVAL_39;
  assign _EVAL_23 = _EVAL_32;
  assign _EVAL_8 = _EVAL_25;
  assign _EVAL_21 = _EVAL_49;
  assign _EVAL_5 = _EVAL_50;
  assign _EVAL_10 = _EVAL_14;
  assign _EVAL_24 = _EVAL_28;
  assign _EVAL = _EVAL_34;
  assign _EVAL_15 = _EVAL_47;
  assign _EVAL_6 = _EVAL_22;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_34 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_40 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_46 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_47 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_48 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_49 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_50 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_11) begin
    if (_EVAL_52) begin
      _EVAL_32 <= _EVAL_25;
    end
    if (_EVAL_52) begin
      _EVAL_34 <= _EVAL_29;
    end
    if (_EVAL_52) begin
      _EVAL_39 <= _EVAL_0;
    end
    if (_EVAL_52) begin
      _EVAL_40 <= _EVAL_18;
    end
    if (_EVAL_1) begin
      _EVAL_46 <= 2'h0;
    end else begin
      if (_EVAL_42) begin
        _EVAL_46 <= _EVAL_35;
      end
    end
    if (_EVAL_52) begin
      _EVAL_47 <= _EVAL_22;
    end
    if (_EVAL_52) begin
      _EVAL_48 <= _EVAL_20;
    end
    if (_EVAL_52) begin
      _EVAL_49 <= _EVAL_14;
    end
    if (_EVAL_52) begin
      _EVAL_50 <= _EVAL_2;
    end
  end
endmodule
