//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_284(
  output        _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  output [31:0] _EVAL_2,
  output        _EVAL_3,
  input  [31:0] _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  input  [4:0]  _EVAL_11,
  output [31:0] _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output [31:0] _EVAL_17,
  input         _EVAL_18,
  output [31:0] _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input  [31:0] _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  output [31:0] _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  input  [5:0]  _EVAL_35,
  input  [31:0] _EVAL_36,
  input  [5:0]  _EVAL_37,
  input  [5:0]  _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input  [4:0]  _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  output        _EVAL_50,
  output        _EVAL_51,
  input         _EVAL_52,
  output        _EVAL_53,
  input         _EVAL_54,
  output        _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  output        _EVAL_58,
  output        _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  output [31:0] _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  input  [31:0] _EVAL_65,
  output        _EVAL_66,
  output        _EVAL_67,
  output        _EVAL_68,
  input  [31:0] _EVAL_69,
  input  [31:0] _EVAL_70,
  output [4:0]  _EVAL_71,
  input  [1:0]  _EVAL_72,
  output        _EVAL_73,
  output        _EVAL_74,
  input         _EVAL_75,
  output [5:0]  _EVAL_76,
  input         _EVAL_77,
  output        _EVAL_78,
  output [1:0]  _EVAL_79,
  input         _EVAL_80,
  output [5:0]  _EVAL_81,
  input         _EVAL_82,
  output [5:0]  _EVAL_83,
  output [4:0]  _EVAL_84,
  output [1:0]  _EVAL_85,
  output        _EVAL_86,
  output        _EVAL_87,
  input         _EVAL_88,
  output        _EVAL_89,
  input         _EVAL_90
);
  assign _EVAL_78 = _EVAL_40;
  assign _EVAL_76 = _EVAL_35;
  assign _EVAL_83 = _EVAL_37;
  assign _EVAL_84 = _EVAL_11;
  assign _EVAL_19 = _EVAL_23;
  assign _EVAL_59 = _EVAL_46;
  assign _EVAL_15 = _EVAL_14;
  assign _EVAL_33 = _EVAL_29;
  assign _EVAL_79 = _EVAL_1;
  assign _EVAL_10 = _EVAL_90;
  assign _EVAL_66 = _EVAL_88;
  assign _EVAL = _EVAL_43;
  assign _EVAL_68 = _EVAL_34;
  assign _EVAL_81 = _EVAL_38;
  assign _EVAL_55 = _EVAL_61;
  assign _EVAL_25 = _EVAL_60;
  assign _EVAL_7 = _EVAL_39;
  assign _EVAL_85 = _EVAL_72;
  assign _EVAL_32 = _EVAL_69;
  assign _EVAL_28 = _EVAL_47;
  assign _EVAL_86 = _EVAL_0;
  assign _EVAL_48 = _EVAL_63;
  assign _EVAL_6 = _EVAL_41;
  assign _EVAL_73 = _EVAL_54;
  assign _EVAL_31 = _EVAL_75;
  assign _EVAL_13 = _EVAL_57;
  assign _EVAL_87 = _EVAL_49;
  assign _EVAL_67 = _EVAL_8;
  assign _EVAL_27 = _EVAL_22;
  assign _EVAL_12 = _EVAL_36;
  assign _EVAL_16 = _EVAL_64;
  assign _EVAL_2 = _EVAL_65;
  assign _EVAL_5 = _EVAL_82;
  assign _EVAL_21 = _EVAL_52;
  assign _EVAL_58 = _EVAL_30;
  assign _EVAL_17 = _EVAL_4;
  assign _EVAL_74 = _EVAL_44;
  assign _EVAL_51 = _EVAL_77;
  assign _EVAL_3 = _EVAL_42;
  assign _EVAL_20 = _EVAL_9;
  assign _EVAL_53 = _EVAL_56;
  assign _EVAL_71 = _EVAL_45;
  assign _EVAL_26 = _EVAL_80;
  assign _EVAL_89 = _EVAL_18;
  assign _EVAL_50 = _EVAL_24;
  assign _EVAL_62 = _EVAL_70;
endmodule
