//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_82(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  output        _EVAL_4,
  output [2:0]  _EVAL_5,
  output [5:0]  _EVAL_6,
  output [31:0] _EVAL_7,
  input  [31:0] _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [5:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  output [3:0]  _EVAL_17,
  output [3:0]  _EVAL_18,
  input  [3:0]  _EVAL_19,
  input         _EVAL_20
);
  reg [3:0] _EVAL_25 [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] _EVAL_25__EVAL_26_data;
  wire  _EVAL_25__EVAL_26_addr;
  wire [3:0] _EVAL_25__EVAL_27_data;
  wire  _EVAL_25__EVAL_27_addr;
  wire  _EVAL_25__EVAL_27_mask;
  wire  _EVAL_25__EVAL_27_en;
  reg [31:0] _EVAL_28 [0:1];
  reg [31:0] _RAND_1;
  wire [31:0] _EVAL_28__EVAL_29_data;
  wire  _EVAL_28__EVAL_29_addr;
  wire [31:0] _EVAL_28__EVAL_30_data;
  wire  _EVAL_28__EVAL_30_addr;
  wire  _EVAL_28__EVAL_30_mask;
  wire  _EVAL_28__EVAL_30_en;
  reg [2:0] _EVAL_33 [0:1];
  reg [31:0] _RAND_2;
  wire [2:0] _EVAL_33__EVAL_34_data;
  wire  _EVAL_33__EVAL_34_addr;
  wire [2:0] _EVAL_33__EVAL_35_data;
  wire  _EVAL_33__EVAL_35_addr;
  wire  _EVAL_33__EVAL_35_mask;
  wire  _EVAL_33__EVAL_35_en;
  reg  _EVAL_38 [0:1];
  reg [31:0] _RAND_3;
  wire  _EVAL_38__EVAL_39_data;
  wire  _EVAL_38__EVAL_39_addr;
  wire  _EVAL_38__EVAL_40_data;
  wire  _EVAL_38__EVAL_40_addr;
  wire  _EVAL_38__EVAL_40_mask;
  wire  _EVAL_38__EVAL_40_en;
  reg [2:0] _EVAL_42 [0:1];
  reg [31:0] _RAND_4;
  wire [2:0] _EVAL_42__EVAL_43_data;
  wire  _EVAL_42__EVAL_43_addr;
  wire [2:0] _EVAL_42__EVAL_44_data;
  wire  _EVAL_42__EVAL_44_addr;
  wire  _EVAL_42__EVAL_44_mask;
  wire  _EVAL_42__EVAL_44_en;
  reg [5:0] _EVAL_49 [0:1];
  reg [31:0] _RAND_5;
  wire [5:0] _EVAL_49__EVAL_50_data;
  wire  _EVAL_49__EVAL_50_addr;
  wire [5:0] _EVAL_49__EVAL_51_data;
  wire  _EVAL_49__EVAL_51_addr;
  wire  _EVAL_49__EVAL_51_mask;
  wire  _EVAL_49__EVAL_51_en;
  reg [31:0] _EVAL_53 [0:1];
  reg [31:0] _RAND_6;
  wire [31:0] _EVAL_53__EVAL_54_data;
  wire  _EVAL_53__EVAL_54_addr;
  wire [31:0] _EVAL_53__EVAL_55_data;
  wire  _EVAL_53__EVAL_55_addr;
  wire  _EVAL_53__EVAL_55_mask;
  wire  _EVAL_53__EVAL_55_en;
  reg [3:0] _EVAL_58 [0:1];
  reg [31:0] _RAND_7;
  wire [3:0] _EVAL_58__EVAL_59_data;
  wire  _EVAL_58__EVAL_59_addr;
  wire [3:0] _EVAL_58__EVAL_60_data;
  wire  _EVAL_58__EVAL_60_addr;
  wire  _EVAL_58__EVAL_60_mask;
  wire  _EVAL_58__EVAL_60_en;
  reg  _EVAL_22;
  reg [31:0] _RAND_8;
  reg  _EVAL_37;
  reg [31:0] _RAND_9;
  reg  _EVAL_48;
  reg [31:0] _RAND_10;
  wire  _EVAL_56;
  wire  _EVAL_45;
  wire  _EVAL_23;
  wire  _EVAL_52;
  wire  _EVAL_46;
  wire  _EVAL_57;
  wire  _EVAL_36;
  wire  _EVAL_21;
  wire  _EVAL_47;
  assign _EVAL_25__EVAL_26_addr = _EVAL_22;
  assign _EVAL_25__EVAL_26_data = _EVAL_25[_EVAL_25__EVAL_26_addr];
  assign _EVAL_25__EVAL_27_data = _EVAL_13;
  assign _EVAL_25__EVAL_27_addr = _EVAL_48;
  assign _EVAL_25__EVAL_27_mask = 1'h1;
  assign _EVAL_25__EVAL_27_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_28__EVAL_29_addr = _EVAL_22;
  assign _EVAL_28__EVAL_29_data = _EVAL_28[_EVAL_28__EVAL_29_addr];
  assign _EVAL_28__EVAL_30_data = _EVAL_8;
  assign _EVAL_28__EVAL_30_addr = _EVAL_48;
  assign _EVAL_28__EVAL_30_mask = 1'h1;
  assign _EVAL_28__EVAL_30_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_33__EVAL_34_addr = _EVAL_22;
  assign _EVAL_33__EVAL_34_data = _EVAL_33[_EVAL_33__EVAL_34_addr];
  assign _EVAL_33__EVAL_35_data = _EVAL_15;
  assign _EVAL_33__EVAL_35_addr = _EVAL_48;
  assign _EVAL_33__EVAL_35_mask = 1'h1;
  assign _EVAL_33__EVAL_35_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_38__EVAL_39_addr = _EVAL_22;
  assign _EVAL_38__EVAL_39_data = _EVAL_38[_EVAL_38__EVAL_39_addr];
  assign _EVAL_38__EVAL_40_data = _EVAL_11;
  assign _EVAL_38__EVAL_40_addr = _EVAL_48;
  assign _EVAL_38__EVAL_40_mask = 1'h1;
  assign _EVAL_38__EVAL_40_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_42__EVAL_43_addr = _EVAL_22;
  assign _EVAL_42__EVAL_43_data = _EVAL_42[_EVAL_42__EVAL_43_addr];
  assign _EVAL_42__EVAL_44_data = _EVAL_2;
  assign _EVAL_42__EVAL_44_addr = _EVAL_48;
  assign _EVAL_42__EVAL_44_mask = 1'h1;
  assign _EVAL_42__EVAL_44_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_49__EVAL_50_addr = _EVAL_22;
  assign _EVAL_49__EVAL_50_data = _EVAL_49[_EVAL_49__EVAL_50_addr];
  assign _EVAL_49__EVAL_51_data = _EVAL_12;
  assign _EVAL_49__EVAL_51_addr = _EVAL_48;
  assign _EVAL_49__EVAL_51_mask = 1'h1;
  assign _EVAL_49__EVAL_51_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_53__EVAL_54_addr = _EVAL_22;
  assign _EVAL_53__EVAL_54_data = _EVAL_53[_EVAL_53__EVAL_54_addr];
  assign _EVAL_53__EVAL_55_data = _EVAL_3;
  assign _EVAL_53__EVAL_55_addr = _EVAL_48;
  assign _EVAL_53__EVAL_55_mask = 1'h1;
  assign _EVAL_53__EVAL_55_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_58__EVAL_59_addr = _EVAL_22;
  assign _EVAL_58__EVAL_59_data = _EVAL_58[_EVAL_58__EVAL_59_addr];
  assign _EVAL_58__EVAL_60_data = _EVAL_19;
  assign _EVAL_58__EVAL_60_addr = _EVAL_48;
  assign _EVAL_58__EVAL_60_mask = 1'h1;
  assign _EVAL_58__EVAL_60_en = _EVAL_4 & _EVAL_20;
  assign _EVAL_56 = _EVAL_4 & _EVAL_20;
  assign _EVAL_45 = _EVAL_10 & _EVAL_1;
  assign _EVAL_23 = _EVAL_56 != _EVAL_45;
  assign _EVAL_52 = _EVAL_37 == 1'h0;
  assign _EVAL_46 = _EVAL_48 == _EVAL_22;
  assign _EVAL_57 = _EVAL_46 & _EVAL_37;
  assign _EVAL_36 = _EVAL_48 + 1'h1;
  assign _EVAL_21 = _EVAL_22 + 1'h1;
  assign _EVAL_47 = _EVAL_46 & _EVAL_52;
  assign _EVAL_7 = _EVAL_28__EVAL_29_data;
  assign _EVAL_17 = _EVAL_58__EVAL_59_data;
  assign _EVAL_9 = _EVAL_38__EVAL_39_data;
  assign _EVAL_6 = _EVAL_49__EVAL_50_data;
  assign _EVAL_18 = _EVAL_25__EVAL_26_data;
  assign _EVAL_1 = _EVAL_47 == 1'h0;
  assign _EVAL = _EVAL_42__EVAL_43_data;
  assign _EVAL_16 = _EVAL_53__EVAL_54_data;
  assign _EVAL_4 = _EVAL_57 == 1'h0;
  assign _EVAL_5 = _EVAL_33__EVAL_34_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_25[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_28[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_33[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_38[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_42[initvar] = _RAND_4[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_49[initvar] = _RAND_5[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_53[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_58[initvar] = _RAND_7[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_22 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_37 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_48 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if(_EVAL_25__EVAL_27_en & _EVAL_25__EVAL_27_mask) begin
      _EVAL_25[_EVAL_25__EVAL_27_addr] <= _EVAL_25__EVAL_27_data;
    end
    if(_EVAL_28__EVAL_30_en & _EVAL_28__EVAL_30_mask) begin
      _EVAL_28[_EVAL_28__EVAL_30_addr] <= _EVAL_28__EVAL_30_data;
    end
    if(_EVAL_33__EVAL_35_en & _EVAL_33__EVAL_35_mask) begin
      _EVAL_33[_EVAL_33__EVAL_35_addr] <= _EVAL_33__EVAL_35_data;
    end
    if(_EVAL_38__EVAL_40_en & _EVAL_38__EVAL_40_mask) begin
      _EVAL_38[_EVAL_38__EVAL_40_addr] <= _EVAL_38__EVAL_40_data;
    end
    if(_EVAL_42__EVAL_44_en & _EVAL_42__EVAL_44_mask) begin
      _EVAL_42[_EVAL_42__EVAL_44_addr] <= _EVAL_42__EVAL_44_data;
    end
    if(_EVAL_49__EVAL_51_en & _EVAL_49__EVAL_51_mask) begin
      _EVAL_49[_EVAL_49__EVAL_51_addr] <= _EVAL_49__EVAL_51_data;
    end
    if(_EVAL_53__EVAL_55_en & _EVAL_53__EVAL_55_mask) begin
      _EVAL_53[_EVAL_53__EVAL_55_addr] <= _EVAL_53__EVAL_55_data;
    end
    if(_EVAL_58__EVAL_60_en & _EVAL_58__EVAL_60_mask) begin
      _EVAL_58[_EVAL_58__EVAL_60_addr] <= _EVAL_58__EVAL_60_data;
    end
    if (_EVAL_0) begin
      _EVAL_22 <= 1'h0;
    end else begin
      if (_EVAL_45) begin
        _EVAL_22 <= _EVAL_21;
      end
    end
    if (_EVAL_0) begin
      _EVAL_37 <= 1'h0;
    end else begin
      if (_EVAL_23) begin
        _EVAL_37 <= _EVAL_56;
      end
    end
    if (_EVAL_0) begin
      _EVAL_48 <= 1'h0;
    end else begin
      if (_EVAL_56) begin
        _EVAL_48 <= _EVAL_36;
      end
    end
  end
endmodule
