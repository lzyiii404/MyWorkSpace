//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_263_assert(
  input  [7:0]  _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [1:0]  _EVAL_3,
  input         _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [31:0] _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input  [2:0]  _EVAL_18,
  input  [31:0] _EVAL_19,
  input         _EVAL_20,
  input  [2:0]  _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [2:0]  _EVAL_25,
  input  [2:0]  _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input  [1:0]  _EVAL_29,
  input         _EVAL_30,
  input  [2:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  input         _EVAL_33
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_94;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_117;
  reg [31:0] _RAND_1;
  reg [31:0] _EVAL_194;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_238;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_252;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_266;
  reg [31:0] _RAND_5;
  reg  _EVAL_283;
  reg [31:0] _RAND_6;
  reg [4:0] _EVAL_318;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_327;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_340;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_345;
  reg [31:0] _RAND_10;
  reg [4:0] _EVAL_354;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_359;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_379;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_384;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_391;
  reg [31:0] _RAND_15;
  reg [31:0] _EVAL_398;
  reg [31:0] _RAND_16;
  reg [1:0] _EVAL_401;
  reg [31:0] _RAND_17;
  reg [3:0] _EVAL_408;
  reg [31:0] _RAND_18;
  reg [31:0] _EVAL_443;
  reg [31:0] _RAND_19;
  reg [2:0] _EVAL_464;
  reg [31:0] _RAND_20;
  reg [4:0] _EVAL_485;
  reg [31:0] _RAND_21;
  reg [7:0] _EVAL_490;
  reg [31:0] _RAND_22;
  reg [2:0] _EVAL_506;
  reg [31:0] _RAND_23;
  reg  _EVAL_525;
  reg [31:0] _RAND_24;
  reg [3:0] _EVAL_585;
  reg [31:0] _RAND_25;
  reg [2:0] _EVAL_609;
  reg [31:0] _RAND_26;
  reg [1:0] _EVAL_616;
  reg [31:0] _RAND_27;
  wire [31:0] _EVAL_256;
  wire  _EVAL_557;
  wire [1:0] _EVAL_560;
  wire [3:0] _EVAL_424;
  wire [2:0] _EVAL_556;
  wire [2:0] _EVAL_465;
  wire  _EVAL_328;
  wire  _EVAL_376;
  wire  _EVAL_453;
  wire  _EVAL_292;
  wire  _EVAL_347;
  wire [22:0] _EVAL_280;
  wire [7:0] _EVAL_413;
  wire  _EVAL_166;
  wire  _EVAL_540;
  wire  _EVAL_563;
  wire  _EVAL_299;
  wire  _EVAL_115;
  wire  _EVAL_623;
  wire  _EVAL_314;
  wire  _EVAL_41;
  wire  _EVAL_326;
  wire [7:0] _EVAL_134;
  wire [7:0] _EVAL_472;
  wire [7:0] _EVAL_248;
  wire  _EVAL_554;
  wire  _EVAL_46;
  wire  _EVAL_123;
  wire [22:0] _EVAL_389;
  wire [7:0] _EVAL_49;
  wire [7:0] _EVAL_366;
  wire [4:0] _EVAL_574;
  wire [4:0] _EVAL_532;
  wire  _EVAL_415;
  wire  _EVAL_84;
  wire  _EVAL_497;
  wire  _EVAL_411;
  wire  _EVAL_122;
  wire  _EVAL_162;
  wire [32:0] _EVAL_630;
  wire [32:0] _EVAL_551;
  wire  _EVAL_508;
  wire  _EVAL_476;
  wire  _EVAL_276;
  wire [7:0] _EVAL_615;
  wire [7:0] _EVAL_631;
  wire [7:0] _EVAL_450;
  wire  _EVAL_304;
  wire  _EVAL_349;
  wire  _EVAL_285;
  wire  _EVAL_469;
  wire  _EVAL_267;
  wire  _EVAL_109;
  wire  _EVAL_614;
  wire  _EVAL_462;
  wire  _EVAL_576;
  wire  _EVAL_565;
  wire  _EVAL_483;
  wire [7:0] _EVAL_503;
  wire [31:0] _EVAL_629;
  wire  _EVAL_143;
  wire [31:0] _EVAL_480;
  wire [32:0] _EVAL_518;
  wire [32:0] _EVAL_152;
  wire [32:0] _EVAL_102;
  wire  _EVAL_206;
  wire [31:0] _EVAL_572;
  wire [32:0] _EVAL_195;
  wire [32:0] _EVAL_535;
  wire [32:0] _EVAL_395;
  wire  _EVAL_114;
  wire  _EVAL_311;
  wire [31:0] _EVAL_357;
  wire [32:0] _EVAL_73;
  wire [32:0] _EVAL_627;
  wire [32:0] _EVAL_87;
  wire  _EVAL_394;
  wire  _EVAL_371;
  wire [31:0] _EVAL_148;
  wire [32:0] _EVAL_265;
  wire [32:0] _EVAL_204;
  wire [32:0] _EVAL_452;
  wire  _EVAL_533;
  wire  _EVAL_255;
  wire  _EVAL_83;
  wire [31:0] _EVAL_81;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_55;
  wire  _EVAL_212;
  wire [31:0] _EVAL_239;
  wire [32:0] _EVAL_498;
  wire [32:0] _EVAL_319;
  wire [32:0] _EVAL_325;
  wire  _EVAL_529;
  wire  _EVAL_182;
  wire  _EVAL_85;
  wire  _EVAL_310;
  wire [31:0] _EVAL_489;
  wire [32:0] _EVAL_571;
  wire [32:0] _EVAL_154;
  wire [32:0] _EVAL_343;
  wire  _EVAL_151;
  wire  _EVAL_396;
  wire [31:0] _EVAL_99;
  wire [32:0] _EVAL_54;
  wire [32:0] _EVAL_367;
  wire [32:0] _EVAL_606;
  wire  _EVAL_215;
  wire  _EVAL_323;
  wire [32:0] _EVAL_397;
  wire [32:0] _EVAL_460;
  wire [32:0] _EVAL_513;
  wire  _EVAL_477;
  wire  _EVAL_137;
  wire [31:0] _EVAL_412;
  wire [32:0] _EVAL_605;
  wire [32:0] _EVAL_546;
  wire [32:0] _EVAL_555;
  wire  _EVAL_405;
  wire  _EVAL_38;
  wire [31:0] _EVAL_127;
  wire [32:0] _EVAL_633;
  wire [32:0] _EVAL_298;
  wire [32:0] _EVAL_579;
  wire  _EVAL_254;
  wire  _EVAL_305;
  wire [31:0] _EVAL_226;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_44;
  wire [32:0] _EVAL_61;
  wire  _EVAL_274;
  wire  _EVAL_235;
  wire  _EVAL_101;
  wire  _EVAL_457;
  wire  _EVAL_227;
  wire  _EVAL_106;
  wire  _EVAL_531;
  wire  _EVAL_404;
  wire  _EVAL_324;
  wire  _EVAL_545;
  wire  _EVAL_423;
  wire  _EVAL_534;
  wire  _EVAL_112;
  wire  _EVAL_372;
  wire  _EVAL_370;
  wire  _EVAL_174;
  wire  _EVAL_604;
  wire  _EVAL_168;
  wire  _EVAL_509;
  wire  _EVAL_589;
  wire  _EVAL_420;
  wire  _EVAL_258;
  wire [31:0] _EVAL_42;
  wire [32:0] _EVAL_399;
  wire [32:0] _EVAL_58;
  wire [32:0] _EVAL_582;
  wire  _EVAL_243;
  wire [32:0] _EVAL_308;
  wire [32:0] _EVAL_217;
  wire [32:0] _EVAL_50;
  wire  _EVAL_80;
  wire  _EVAL_63;
  wire [32:0] _EVAL_315;
  wire [32:0] _EVAL_348;
  wire [32:0] _EVAL_516;
  wire  _EVAL_300;
  wire  _EVAL_288;
  wire  _EVAL_253;
  wire  _EVAL_353;
  wire  _EVAL_186;
  wire  _EVAL_157;
  wire  _EVAL_400;
  wire  _EVAL_528;
  wire  _EVAL_597;
  wire [1:0] _EVAL_56;
  wire [1:0] _EVAL_601;
  wire [1:0] _EVAL_144;
  wire  _EVAL_594;
  wire [31:0] _EVAL_279;
  wire [32:0] _EVAL_281;
  wire [32:0] _EVAL_179;
  wire [32:0] _EVAL_451;
  wire  _EVAL_59;
  wire  _EVAL_142;
  wire [31:0] _EVAL_439;
  wire [32:0] _EVAL_409;
  wire [32:0] _EVAL_189;
  wire [32:0] _EVAL_530;
  wire  _EVAL_113;
  wire  _EVAL_547;
  wire [32:0] _EVAL_224;
  wire  _EVAL_146;
  wire  _EVAL_35;
  wire [31:0] _EVAL_523;
  wire [32:0] _EVAL_620;
  wire [32:0] _EVAL_346;
  wire [32:0] _EVAL_313;
  wire  _EVAL_321;
  wire  _EVAL_337;
  wire [31:0] _EVAL_390;
  wire [32:0] _EVAL_548;
  wire [32:0] _EVAL_332;
  wire [32:0] _EVAL_595;
  wire  _EVAL_602;
  wire  _EVAL_493;
  wire [31:0] _EVAL_336;
  wire [32:0] _EVAL_96;
  wire [32:0] _EVAL_558;
  wire [32:0] _EVAL_192;
  wire  _EVAL_632;
  wire  _EVAL_329;
  wire  _EVAL_559;
  wire  _EVAL_297;
  wire  _EVAL_75;
  wire  _EVAL_590;
  wire [31:0] _EVAL_36;
  wire [32:0] _EVAL_147;
  wire [32:0] _EVAL_592;
  wire [31:0] _EVAL_500;
  wire [32:0] _EVAL_139;
  wire [32:0] _EVAL_138;
  wire [32:0] _EVAL_351;
  wire  _EVAL_286;
  wire  _EVAL_584;
  wire  _EVAL_600;
  wire  _EVAL_495;
  wire [31:0] _EVAL_425;
  wire [32:0] _EVAL_382;
  wire [32:0] _EVAL_225;
  wire [32:0] _EVAL_499;
  wire  _EVAL_339;
  wire  _EVAL_427;
  wire [32:0] _EVAL_536;
  wire [32:0] _EVAL_260;
  wire [32:0] _EVAL_407;
  wire  _EVAL_561;
  wire  _EVAL_338;
  wire [31:0] _EVAL_539;
  wire [32:0] _EVAL_156;
  wire [32:0] _EVAL_51;
  wire [32:0] _EVAL_245;
  wire  _EVAL_612;
  wire  _EVAL_251;
  wire [32:0] _EVAL_473;
  wire  _EVAL_198;
  wire  _EVAL_111;
  wire  _EVAL_335;
  wire  _EVAL_149;
  wire  _EVAL_293;
  wire  _EVAL_211;
  wire  _EVAL_591;
  wire  _EVAL_622;
  wire  _EVAL_242;
  wire  _EVAL_377;
  wire [22:0] _EVAL_131;
  wire [7:0] _EVAL_205;
  wire [7:0] _EVAL_241;
  wire [4:0] _EVAL_155;
  wire  _EVAL_419;
  wire  _EVAL_388;
  wire [7:0] _EVAL_53;
  wire [4:0] _EVAL_124;
  wire [4:0] _EVAL_466;
  wire  _EVAL_587;
  wire  _EVAL_352;
  wire  _EVAL_564;
  wire  _EVAL_237;
  wire  _EVAL_76;
  wire  _EVAL_71;
  wire  _EVAL_468;
  wire  _EVAL_190;
  wire  _EVAL_342;
  wire  _EVAL_567;
  wire  _EVAL_543;
  wire  _EVAL_210;
  wire  _EVAL_141;
  wire  _EVAL_228;
  wire  _EVAL_67;
  wire  _EVAL_507;
  wire  _EVAL_626;
  wire  _EVAL_231;
  wire  _EVAL_475;
  wire  _EVAL_511;
  wire  _EVAL_350;
  wire  _EVAL_333;
  wire  _EVAL_107;
  wire [31:0] _EVAL_140;
  wire [31:0] _EVAL_263;
  wire  _EVAL_440;
  wire  _EVAL_262;
  wire  _EVAL_316;
  wire  _EVAL_184;
  wire  _EVAL_541;
  wire  _EVAL_421;
  wire  _EVAL_431;
  wire  _EVAL_428;
  wire  _EVAL_410;
  wire  _EVAL_145;
  wire  _EVAL_132;
  wire  _EVAL_512;
  wire  _EVAL_57;
  wire  _EVAL_170;
  wire  _EVAL_402;
  wire  _EVAL_422;
  wire  _EVAL_178;
  wire  _EVAL_445;
  wire  _EVAL_458;
  wire  _EVAL_290;
  wire  _EVAL_385;
  wire  _EVAL_271;
  wire  _EVAL_309;
  wire  _EVAL_617;
  wire  _EVAL_278;
  wire  _EVAL_247;
  wire  _EVAL_573;
  wire  _EVAL_355;
  wire  _EVAL_442;
  wire  _EVAL_91;
  wire [7:0] _EVAL_159;
  wire  _EVAL_92;
  wire  _EVAL_517;
  wire  _EVAL_188;
  wire  _EVAL_514;
  wire  _EVAL_393;
  wire  _EVAL_296;
  wire  _EVAL_386;
  wire  _EVAL_455;
  wire  _EVAL_448;
  wire  _EVAL_611;
  wire  _EVAL_575;
  wire  _EVAL_624;
  wire [4:0] _EVAL_553;
  wire  _EVAL_446;
  wire  _EVAL_287;
  wire  _EVAL_625;
  wire  _EVAL_257;
  wire  _EVAL_177;
  wire  _EVAL_486;
  wire  _EVAL_220;
  wire  _EVAL_37;
  wire  _EVAL_77;
  wire  _EVAL_368;
  wire [4:0] _EVAL_97;
  wire  _EVAL_364;
  wire  _EVAL_218;
  wire [1:0] _EVAL_209;
  wire [1:0] _EVAL_417;
  wire [1:0] _EVAL_291;
  wire  _EVAL_596;
  wire  _EVAL_363;
  wire  _EVAL_103;
  wire  _EVAL_196;
  wire  _EVAL_502;
  wire  _EVAL_68;
  wire  _EVAL_416;
  wire  _EVAL_108;
  wire  _EVAL_578;
  wire  _EVAL_581;
  wire  _EVAL_330;
  wire  _EVAL_52;
  wire  _EVAL_521;
  wire  _EVAL_89;
  wire  _EVAL_418;
  wire  _EVAL_383;
  wire  _EVAL_136;
  wire  _EVAL_599;
  wire [1:0] _EVAL_187;
  wire  _EVAL_128;
  wire  _EVAL_361;
  wire [7:0] _EVAL_519;
  wire  _EVAL_334;
  wire  _EVAL_482;
  wire  _EVAL_171;
  wire  _EVAL_232;
  wire  _EVAL_487;
  wire  _EVAL_621;
  wire  _EVAL_373;
  wire [31:0] _EVAL_619;
  wire  _EVAL_356;
  wire  _EVAL_264;
  wire  _EVAL_180;
  wire  _EVAL_331;
  wire  _EVAL_470;
  wire  _EVAL_430;
  wire  _EVAL_358;
  wire  _EVAL_86;
  wire  _EVAL_378;
  wire  _EVAL_344;
  wire [4:0] _EVAL_277;
  wire [1:0] _EVAL_172;
  wire  _EVAL_447;
  wire [4:0] _EVAL_261;
  wire  _EVAL_66;
  wire  _EVAL_569;
  wire  _EVAL_116;
  wire  _EVAL_126;
  wire  _EVAL_181;
  wire  _EVAL_488;
  wire [31:0] _EVAL_214;
  wire  _EVAL_586;
  wire  _EVAL_70;
  wire  _EVAL_294;
  wire  _EVAL_362;
  wire  _EVAL_570;
  wire  _EVAL_289;
  wire  _EVAL_120;
  wire  _EVAL_479;
  wire  _EVAL_303;
  wire  _EVAL_580;
  wire [31:0] _EVAL_484;
  wire [31:0] _EVAL_634;
  wire  _EVAL_491;
  wire  _EVAL_403;
  wire  _EVAL_79;
  wire  _EVAL_95;
  wire  _EVAL_222;
  wire  _EVAL_496;
  wire  _EVAL_454;
  wire  _EVAL_520;
  wire  _EVAL_167;
  wire  _EVAL_164;
  wire  _EVAL_438;
  wire  _EVAL_105;
  wire  _EVAL_153;
  wire  _EVAL_246;
  wire  _EVAL_90;
  wire [1:0] _EVAL_542;
  wire  _EVAL_375;
  wire [4:0] _EVAL_436;
  wire  _EVAL_426;
  wire  _EVAL_110;
  wire  _EVAL_628;
  wire  _EVAL_461;
  wire  _EVAL_550;
  wire  _EVAL_93;
  wire  _EVAL_568;
  wire  _EVAL_88;
  wire  _EVAL_474;
  wire  _EVAL_380;
  wire  _EVAL_150;
  wire  _EVAL_233;
  wire  _EVAL_524;
  wire  _EVAL_434;
  wire  _EVAL_118;
  wire  _EVAL_203;
  wire  _EVAL_125;
  wire  _EVAL_527;
  wire  _EVAL_537;
  wire  _EVAL_320;
  wire  _EVAL_437;
  wire  _EVAL_65;
  wire [7:0] _EVAL_387;
  wire [7:0] _EVAL_229;
  wire  _EVAL_341;
  wire  _EVAL_301;
  wire  _EVAL_269;
  wire [7:0] _EVAL_610;
  wire  _EVAL_259;
  wire  _EVAL_272;
  wire  _EVAL_39;
  wire [7:0] _EVAL_273;
  wire [7:0] _EVAL_467;
  wire  _EVAL_284;
  wire  _EVAL_444;
  wire  _EVAL_98;
  wire  _EVAL_236;
  wire  _EVAL_306;
  wire  _EVAL_169;
  wire  _EVAL_270;
  wire  _EVAL_78;
  wire  _EVAL_197;
  wire  _EVAL_133;
  wire  _EVAL_165;
  wire  _EVAL_100;
  wire  _EVAL_158;
  wire  _EVAL_544;
  wire  _EVAL_244;
  wire  _EVAL_240;
  wire  _EVAL_207;
  wire  _EVAL_199;
  wire  _EVAL_381;
  wire  _EVAL_249;
  wire  _EVAL_121;
  wire  _EVAL_216;
  wire  _EVAL_593;
  wire  _EVAL_161;
  wire  _EVAL_223;
  wire  _EVAL_607;
  wire  _EVAL_275;
  wire  _EVAL_494;
  wire  _EVAL_510;
  wire  _EVAL_200;
  wire  _EVAL_515;
  wire  _EVAL_360;
  wire  _EVAL_588;
  wire  _EVAL_501;
  wire  _EVAL_48;
  wire [1:0] _EVAL_504;
  wire  _EVAL_322;
  wire  _EVAL_613;
  wire  _EVAL_185;
  wire  _EVAL_505;
  wire  _EVAL_193;
  wire  _EVAL_119;
  wire  _EVAL_583;
  wire  _EVAL_478;
  wire  _EVAL_62;
  wire  _EVAL_183;
  wire  _EVAL_282;
  wire  _EVAL_374;
  wire  _EVAL_221;
  wire  _EVAL_538;
  wire  _EVAL_295;
  wire  _EVAL_302;
  wire  _EVAL_43;
  wire  _EVAL_566;
  wire  _EVAL_175;
  wire  _EVAL_230;
  wire  _EVAL_74;
  wire  _EVAL_618;
  wire  _EVAL_191;
  wire  _EVAL_481;
  wire  _EVAL_45;
  wire  _EVAL_562;
  wire  _EVAL_173;
  wire  _EVAL_47;
  wire  _EVAL_307;
  wire  _EVAL_492;
  wire  _EVAL_471;
  wire  _EVAL_522;
  wire  _EVAL_441;
  wire  _EVAL_414;
  wire  _EVAL_526;
  wire  _EVAL_463;
  wire  _EVAL_433;
  wire  _EVAL_176;
  wire  _EVAL_406;
  wire  _EVAL_392;
  wire  _EVAL_34;
  wire  _EVAL_234;
  wire  _EVAL_129;
  wire  _EVAL_312;
  wire  _EVAL_459;
  wire  _EVAL_598;
  wire  _EVAL_64;
  wire  _EVAL_40;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_256 = _EVAL_0 ^ 32'h3000;
  assign _EVAL_557 = _EVAL_5 >= 4'h3;
  assign _EVAL_560 = _EVAL_5[1:0];
  assign _EVAL_424 = 4'h1 << _EVAL_560;
  assign _EVAL_556 = _EVAL_424[2:0];
  assign _EVAL_465 = _EVAL_556 | 3'h1;
  assign _EVAL_328 = _EVAL_465[2];
  assign _EVAL_376 = _EVAL_19[2];
  assign _EVAL_453 = _EVAL_376 == 1'h0;
  assign _EVAL_292 = _EVAL_328 & _EVAL_453;
  assign _EVAL_347 = _EVAL_557 | _EVAL_292;
  assign _EVAL_280 = 23'hff << _EVAL_9;
  assign _EVAL_413 = _EVAL_280[7:0];
  assign _EVAL_166 = _EVAL_32 == 3'h5;
  assign _EVAL_540 = _EVAL_8 & _EVAL_166;
  assign _EVAL_563 = _EVAL_17 == _EVAL_585;
  assign _EVAL_299 = _EVAL_12 & _EVAL_28;
  assign _EVAL_115 = _EVAL_485 == 5'h0;
  assign _EVAL_623 = _EVAL_299 & _EVAL_115;
  assign _EVAL_314 = _EVAL_6 == 3'h6;
  assign _EVAL_41 = _EVAL_314 == 1'h0;
  assign _EVAL_326 = _EVAL_623 & _EVAL_41;
  assign _EVAL_134 = 8'h1 << _EVAL_25;
  assign _EVAL_472 = _EVAL_326 ? _EVAL_134 : 8'h0;
  assign _EVAL_248 = ~ _EVAL_472;
  assign _EVAL_554 = _EVAL_22 & _EVAL_8;
  assign _EVAL_46 = _EVAL_354 == 5'h0;
  assign _EVAL_123 = _EVAL_32[0];
  assign _EVAL_389 = 23'hff << _EVAL_17;
  assign _EVAL_49 = _EVAL_389[7:0];
  assign _EVAL_366 = ~ _EVAL_49;
  assign _EVAL_574 = _EVAL_366[7:3];
  assign _EVAL_532 = _EVAL_354 - 5'h1;
  assign _EVAL_415 = _EVAL_3 == _EVAL_616;
  assign _EVAL_84 = _EVAL_415 | _EVAL_23;
  assign _EVAL_497 = _EVAL_84 == 1'h0;
  assign _EVAL_411 = _EVAL_11 == 1'h0;
  assign _EVAL_122 = _EVAL_411 | _EVAL_24;
  assign _EVAL_162 = _EVAL_122 | _EVAL_23;
  assign _EVAL_630 = {1'b0,$signed(_EVAL_0)};
  assign _EVAL_551 = $signed(_EVAL_630) & $signed(-33'sh1000);
  assign _EVAL_508 = _EVAL_1 & _EVAL_33;
  assign _EVAL_476 = _EVAL_318 == 5'h0;
  assign _EVAL_276 = _EVAL_508 & _EVAL_476;
  assign _EVAL_615 = 8'h1 << _EVAL_26;
  assign _EVAL_631 = _EVAL_276 ? _EVAL_615 : 8'h0;
  assign _EVAL_450 = _EVAL_631 | _EVAL_490;
  assign _EVAL_304 = _EVAL_21 == 3'h0;
  assign _EVAL_349 = 4'h6 == _EVAL_17;
  assign _EVAL_285 = _EVAL_304 ? _EVAL_349 : 1'h0;
  assign _EVAL_469 = _EVAL_285 | _EVAL_23;
  assign _EVAL_267 = _EVAL_557 | _EVAL_23;
  assign _EVAL_109 = _EVAL_465[1];
  assign _EVAL_614 = _EVAL_19[1];
  assign _EVAL_462 = _EVAL_614 == 1'h0;
  assign _EVAL_576 = _EVAL_453 & _EVAL_462;
  assign _EVAL_565 = _EVAL_109 & _EVAL_576;
  assign _EVAL_483 = _EVAL_29 == 2'h0;
  assign _EVAL_503 = ~ _EVAL;
  assign _EVAL_629 = _EVAL_0 ^ 32'h80000000;
  assign _EVAL_143 = _EVAL_376 & _EVAL_462;
  assign _EVAL_480 = _EVAL_19 ^ 32'h40000000;
  assign _EVAL_518 = {1'b0,$signed(_EVAL_480)};
  assign _EVAL_152 = $signed(_EVAL_518) & $signed(-33'sh2000);
  assign _EVAL_102 = $signed(_EVAL_152);
  assign _EVAL_206 = $signed(_EVAL_102) == $signed(33'sh0);
  assign _EVAL_572 = _EVAL_19 ^ 32'h80000000;
  assign _EVAL_195 = {1'b0,$signed(_EVAL_572)};
  assign _EVAL_535 = $signed(_EVAL_195) & $signed(-33'sh20000);
  assign _EVAL_395 = $signed(_EVAL_535);
  assign _EVAL_114 = $signed(_EVAL_395) == $signed(33'sh0);
  assign _EVAL_311 = _EVAL_206 | _EVAL_114;
  assign _EVAL_357 = _EVAL_19 ^ 32'hc000000;
  assign _EVAL_73 = {1'b0,$signed(_EVAL_357)};
  assign _EVAL_627 = $signed(_EVAL_73) & $signed(-33'sh4000000);
  assign _EVAL_87 = $signed(_EVAL_627);
  assign _EVAL_394 = $signed(_EVAL_87) == $signed(33'sh0);
  assign _EVAL_371 = _EVAL_311 | _EVAL_394;
  assign _EVAL_148 = _EVAL_15 ^ 32'h3000;
  assign _EVAL_265 = {1'b0,$signed(_EVAL_148)};
  assign _EVAL_204 = $signed(_EVAL_265) & $signed(-33'sh1000);
  assign _EVAL_452 = $signed(_EVAL_204);
  assign _EVAL_533 = _EVAL_267 == 1'h0;
  assign _EVAL_255 = _EVAL_24 == 1'h0;
  assign _EVAL_83 = _EVAL_255 | _EVAL_23;
  assign _EVAL_81 = _EVAL_15 ^ 32'h40000000;
  assign _EVAL_104 = {1'b0,$signed(_EVAL_81)};
  assign _EVAL_130 = $signed(_EVAL_104) & $signed(-33'sh2000);
  assign _EVAL_55 = $signed(_EVAL_130);
  assign _EVAL_212 = $signed(_EVAL_55) == $signed(33'sh0);
  assign _EVAL_239 = _EVAL_15 ^ 32'h80000000;
  assign _EVAL_498 = {1'b0,$signed(_EVAL_239)};
  assign _EVAL_319 = $signed(_EVAL_498) & $signed(-33'sh20000);
  assign _EVAL_325 = $signed(_EVAL_319);
  assign _EVAL_529 = $signed(_EVAL_325) == $signed(33'sh0);
  assign _EVAL_182 = _EVAL_212 | _EVAL_529;
  assign _EVAL_85 = $signed(_EVAL_452) == $signed(33'sh0);
  assign _EVAL_310 = _EVAL_182 | _EVAL_85;
  assign _EVAL_489 = _EVAL_15 ^ 32'hc000000;
  assign _EVAL_571 = {1'b0,$signed(_EVAL_489)};
  assign _EVAL_154 = $signed(_EVAL_571) & $signed(-33'sh4000000);
  assign _EVAL_343 = $signed(_EVAL_154);
  assign _EVAL_151 = $signed(_EVAL_343) == $signed(33'sh0);
  assign _EVAL_396 = _EVAL_310 | _EVAL_151;
  assign _EVAL_99 = _EVAL_15 ^ 32'h2000000;
  assign _EVAL_54 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_367 = $signed(_EVAL_54) & $signed(-33'sh10000);
  assign _EVAL_606 = $signed(_EVAL_367);
  assign _EVAL_215 = $signed(_EVAL_606) == $signed(33'sh0);
  assign _EVAL_323 = _EVAL_396 | _EVAL_215;
  assign _EVAL_397 = {1'b0,$signed(_EVAL_15)};
  assign _EVAL_460 = $signed(_EVAL_397) & $signed(-33'sh1000);
  assign _EVAL_513 = $signed(_EVAL_460);
  assign _EVAL_477 = $signed(_EVAL_513) == $signed(33'sh0);
  assign _EVAL_137 = _EVAL_323 | _EVAL_477;
  assign _EVAL_412 = _EVAL_15 ^ 32'h1800000;
  assign _EVAL_605 = {1'b0,$signed(_EVAL_412)};
  assign _EVAL_546 = $signed(_EVAL_605) & $signed(-33'sh8000);
  assign _EVAL_555 = $signed(_EVAL_546);
  assign _EVAL_405 = $signed(_EVAL_555) == $signed(33'sh0);
  assign _EVAL_38 = _EVAL_137 | _EVAL_405;
  assign _EVAL_127 = _EVAL_15 ^ 32'h4000;
  assign _EVAL_633 = {1'b0,$signed(_EVAL_127)};
  assign _EVAL_298 = $signed(_EVAL_633) & $signed(-33'sh1000);
  assign _EVAL_579 = $signed(_EVAL_298);
  assign _EVAL_254 = $signed(_EVAL_579) == $signed(33'sh0);
  assign _EVAL_305 = _EVAL_38 | _EVAL_254;
  assign _EVAL_226 = _EVAL_15 ^ 32'h20000000;
  assign _EVAL_163 = {1'b0,$signed(_EVAL_226)};
  assign _EVAL_44 = $signed(_EVAL_163) & $signed(-33'sh2000);
  assign _EVAL_61 = $signed(_EVAL_44);
  assign _EVAL_274 = $signed(_EVAL_61) == $signed(33'sh0);
  assign _EVAL_235 = _EVAL_305 | _EVAL_274;
  assign _EVAL_101 = _EVAL_18 == 3'h5;
  assign _EVAL_457 = 3'h1 <= _EVAL_21;
  assign _EVAL_227 = _EVAL_304 | _EVAL_457;
  assign _EVAL_106 = _EVAL_266 == 5'h0;
  assign _EVAL_531 = _EVAL_106 == 1'h0;
  assign _EVAL_404 = _EVAL_28 & _EVAL_531;
  assign _EVAL_324 = _EVAL_453 & _EVAL_614;
  assign _EVAL_545 = _EVAL_109 & _EVAL_324;
  assign _EVAL_423 = _EVAL_347 | _EVAL_545;
  assign _EVAL_534 = _EVAL_465[0];
  assign _EVAL_112 = _EVAL_19[0];
  assign _EVAL_372 = _EVAL_112 == 1'h0;
  assign _EVAL_370 = _EVAL_324 & _EVAL_372;
  assign _EVAL_174 = _EVAL_534 & _EVAL_370;
  assign _EVAL_604 = _EVAL_423 | _EVAL_174;
  assign _EVAL_168 = _EVAL_2 == 3'h0;
  assign _EVAL_509 = _EVAL_168 | _EVAL_23;
  assign _EVAL_589 = _EVAL_32 == _EVAL_506;
  assign _EVAL_420 = _EVAL_589 | _EVAL_23;
  assign _EVAL_258 = _EVAL_420 == 1'h0;
  assign _EVAL_42 = _EVAL_0 ^ 32'h40000000;
  assign _EVAL_399 = {1'b0,$signed(_EVAL_42)};
  assign _EVAL_58 = $signed(_EVAL_399) & $signed(-33'sh2000);
  assign _EVAL_582 = $signed(_EVAL_58);
  assign _EVAL_243 = $signed(_EVAL_582) == $signed(33'sh0);
  assign _EVAL_308 = {1'b0,$signed(_EVAL_629)};
  assign _EVAL_217 = $signed(_EVAL_308) & $signed(-33'sh20000);
  assign _EVAL_50 = $signed(_EVAL_217);
  assign _EVAL_80 = $signed(_EVAL_50) == $signed(33'sh0);
  assign _EVAL_63 = _EVAL_243 | _EVAL_80;
  assign _EVAL_315 = {1'b0,$signed(_EVAL_256)};
  assign _EVAL_348 = $signed(_EVAL_315) & $signed(-33'sh1000);
  assign _EVAL_516 = $signed(_EVAL_348);
  assign _EVAL_300 = $signed(_EVAL_516) == $signed(33'sh0);
  assign _EVAL_288 = _EVAL_63 | _EVAL_300;
  assign _EVAL_253 = _EVAL_379 == 5'h0;
  assign _EVAL_353 = _EVAL_299 & _EVAL_253;
  assign _EVAL_186 = _EVAL_6[2];
  assign _EVAL_157 = _EVAL_6[1];
  assign _EVAL_400 = _EVAL_157 == 1'h0;
  assign _EVAL_528 = _EVAL_186 & _EVAL_400;
  assign _EVAL_597 = _EVAL_353 & _EVAL_528;
  assign _EVAL_56 = 2'h1 << _EVAL_30;
  assign _EVAL_601 = _EVAL_597 ? _EVAL_56 : 2'h0;
  assign _EVAL_144 = _EVAL_601 | _EVAL_401;
  assign _EVAL_594 = _EVAL_9 >= 4'h3;
  assign _EVAL_279 = _EVAL_0 ^ 32'hc000000;
  assign _EVAL_281 = {1'b0,$signed(_EVAL_279)};
  assign _EVAL_179 = $signed(_EVAL_281) & $signed(-33'sh4000000);
  assign _EVAL_451 = $signed(_EVAL_179);
  assign _EVAL_59 = $signed(_EVAL_451) == $signed(33'sh0);
  assign _EVAL_142 = _EVAL_288 | _EVAL_59;
  assign _EVAL_439 = _EVAL_0 ^ 32'h2000000;
  assign _EVAL_409 = {1'b0,$signed(_EVAL_439)};
  assign _EVAL_189 = $signed(_EVAL_409) & $signed(-33'sh10000);
  assign _EVAL_530 = $signed(_EVAL_189);
  assign _EVAL_113 = $signed(_EVAL_530) == $signed(33'sh0);
  assign _EVAL_547 = _EVAL_142 | _EVAL_113;
  assign _EVAL_224 = $signed(_EVAL_551);
  assign _EVAL_146 = $signed(_EVAL_224) == $signed(33'sh0);
  assign _EVAL_35 = _EVAL_547 | _EVAL_146;
  assign _EVAL_523 = _EVAL_0 ^ 32'h1800000;
  assign _EVAL_620 = {1'b0,$signed(_EVAL_523)};
  assign _EVAL_346 = $signed(_EVAL_620) & $signed(-33'sh8000);
  assign _EVAL_313 = $signed(_EVAL_346);
  assign _EVAL_321 = $signed(_EVAL_313) == $signed(33'sh0);
  assign _EVAL_337 = _EVAL_35 | _EVAL_321;
  assign _EVAL_390 = _EVAL_0 ^ 32'h4000;
  assign _EVAL_548 = {1'b0,$signed(_EVAL_390)};
  assign _EVAL_332 = $signed(_EVAL_548) & $signed(-33'sh1000);
  assign _EVAL_595 = $signed(_EVAL_332);
  assign _EVAL_602 = $signed(_EVAL_595) == $signed(33'sh0);
  assign _EVAL_493 = _EVAL_337 | _EVAL_602;
  assign _EVAL_336 = _EVAL_0 ^ 32'h20000000;
  assign _EVAL_96 = {1'b0,$signed(_EVAL_336)};
  assign _EVAL_558 = $signed(_EVAL_96) & $signed(-33'sh2000);
  assign _EVAL_192 = $signed(_EVAL_558);
  assign _EVAL_632 = $signed(_EVAL_192) == $signed(33'sh0);
  assign _EVAL_329 = _EVAL_493 | _EVAL_632;
  assign _EVAL_559 = _EVAL_329 | _EVAL_23;
  assign _EVAL_297 = _EVAL_227 | _EVAL_23;
  assign _EVAL_75 = _EVAL_297 == 1'h0;
  assign _EVAL_590 = _EVAL_10 == 1'h0;
  assign _EVAL_36 = _EVAL_19 ^ 32'h20000000;
  assign _EVAL_147 = {1'b0,$signed(_EVAL_36)};
  assign _EVAL_592 = $signed(_EVAL_147) & $signed(-33'sh2000);
  assign _EVAL_500 = _EVAL_19 ^ 32'h3000;
  assign _EVAL_139 = {1'b0,$signed(_EVAL_500)};
  assign _EVAL_138 = $signed(_EVAL_139) & $signed(-33'sh1000);
  assign _EVAL_351 = $signed(_EVAL_138);
  assign _EVAL_286 = $signed(_EVAL_351) == $signed(33'sh0);
  assign _EVAL_584 = _EVAL_286 | _EVAL_394;
  assign _EVAL_600 = _EVAL_31 <= 3'h4;
  assign _EVAL_495 = _EVAL_5 <= 4'h2;
  assign _EVAL_425 = _EVAL_19 ^ 32'h2000000;
  assign _EVAL_382 = {1'b0,$signed(_EVAL_425)};
  assign _EVAL_225 = $signed(_EVAL_382) & $signed(-33'sh10000);
  assign _EVAL_499 = $signed(_EVAL_225);
  assign _EVAL_339 = $signed(_EVAL_499) == $signed(33'sh0);
  assign _EVAL_427 = _EVAL_584 | _EVAL_339;
  assign _EVAL_536 = {1'b0,$signed(_EVAL_19)};
  assign _EVAL_260 = $signed(_EVAL_536) & $signed(-33'sh5000);
  assign _EVAL_407 = $signed(_EVAL_260);
  assign _EVAL_561 = $signed(_EVAL_407) == $signed(33'sh0);
  assign _EVAL_338 = _EVAL_427 | _EVAL_561;
  assign _EVAL_539 = _EVAL_19 ^ 32'h1800000;
  assign _EVAL_156 = {1'b0,$signed(_EVAL_539)};
  assign _EVAL_51 = $signed(_EVAL_156) & $signed(-33'sh8000);
  assign _EVAL_245 = $signed(_EVAL_51);
  assign _EVAL_612 = $signed(_EVAL_245) == $signed(33'sh0);
  assign _EVAL_251 = _EVAL_338 | _EVAL_612;
  assign _EVAL_473 = $signed(_EVAL_592);
  assign _EVAL_198 = $signed(_EVAL_473) == $signed(33'sh0);
  assign _EVAL_111 = _EVAL_251 | _EVAL_198;
  assign _EVAL_335 = _EVAL_495 & _EVAL_111;
  assign _EVAL_149 = _EVAL_335 | _EVAL_23;
  assign _EVAL_293 = _EVAL_149 == 1'h0;
  assign _EVAL_211 = _EVAL_31 <= 3'h2;
  assign _EVAL_591 = _EVAL_211 | _EVAL_23;
  assign _EVAL_622 = _EVAL_591 == 1'h0;
  assign _EVAL_242 = _EVAL_32 == 3'h0;
  assign _EVAL_377 = _EVAL_8 & _EVAL_242;
  assign _EVAL_131 = 23'hff << _EVAL_5;
  assign _EVAL_205 = _EVAL_131[7:0];
  assign _EVAL_241 = ~ _EVAL_205;
  assign _EVAL_155 = _EVAL_241[7:3];
  assign _EVAL_419 = _EVAL_324 & _EVAL_112;
  assign _EVAL_388 = _EVAL_6[0];
  assign _EVAL_53 = ~ _EVAL_413;
  assign _EVAL_124 = _EVAL_53[7:3];
  assign _EVAL_466 = _EVAL_266 - 5'h1;
  assign _EVAL_587 = _EVAL_29 <= 2'h2;
  assign _EVAL_352 = _EVAL_328 & _EVAL_376;
  assign _EVAL_564 = _EVAL_557 | _EVAL_352;
  assign _EVAL_237 = _EVAL_376 & _EVAL_614;
  assign _EVAL_76 = _EVAL_109 & _EVAL_237;
  assign _EVAL_71 = _EVAL_564 | _EVAL_76;
  assign _EVAL_468 = _EVAL_237 & _EVAL_112;
  assign _EVAL_190 = _EVAL_534 & _EVAL_468;
  assign _EVAL_342 = _EVAL_71 | _EVAL_190;
  assign _EVAL_567 = _EVAL_3 <= 2'h2;
  assign _EVAL_543 = _EVAL_14 & _EVAL_16;
  assign _EVAL_210 = _EVAL_371 | _EVAL_339;
  assign _EVAL_141 = _EVAL_26 == 3'h0;
  assign _EVAL_228 = 4'h6 == _EVAL_5;
  assign _EVAL_67 = _EVAL_141 ? _EVAL_228 : 1'h0;
  assign _EVAL_507 = _EVAL_5 <= 4'h8;
  assign _EVAL_626 = _EVAL_507 & _EVAL_286;
  assign _EVAL_231 = _EVAL_626 | _EVAL_23;
  assign _EVAL_475 = _EVAL_231 == 1'h0;
  assign _EVAL_511 = 3'h1 <= _EVAL_26;
  assign _EVAL_350 = _EVAL_141 | _EVAL_511;
  assign _EVAL_333 = _EVAL_17 >= 4'h3;
  assign _EVAL_107 = _EVAL_333 | _EVAL_23;
  assign _EVAL_140 = {{24'd0}, _EVAL_366};
  assign _EVAL_263 = _EVAL_15 & _EVAL_140;
  assign _EVAL_440 = _EVAL_263 == 32'h0;
  assign _EVAL_262 = _EVAL_440 | _EVAL_23;
  assign _EVAL_316 = _EVAL_2 == _EVAL_359;
  assign _EVAL_184 = _EVAL_316 | _EVAL_23;
  assign _EVAL_541 = _EVAL_184 == 1'h0;
  assign _EVAL_421 = _EVAL_9 == _EVAL_340;
  assign _EVAL_431 = _EVAL_421 | _EVAL_23;
  assign _EVAL_428 = _EVAL_30 == _EVAL_525;
  assign _EVAL_410 = _EVAL_428 | _EVAL_23;
  assign _EVAL_145 = _EVAL_18 == 3'h0;
  assign _EVAL_132 = _EVAL_237 & _EVAL_372;
  assign _EVAL_512 = _EVAL_534 & _EVAL_132;
  assign _EVAL_57 = _EVAL_71 | _EVAL_512;
  assign _EVAL_170 = _EVAL_109 & _EVAL_143;
  assign _EVAL_402 = _EVAL_564 | _EVAL_170;
  assign _EVAL_422 = _EVAL_143 & _EVAL_112;
  assign _EVAL_178 = _EVAL_534 & _EVAL_422;
  assign _EVAL_445 = _EVAL_402 | _EVAL_178;
  assign _EVAL_458 = _EVAL_143 & _EVAL_372;
  assign _EVAL_290 = _EVAL_534 & _EVAL_458;
  assign _EVAL_385 = _EVAL_402 | _EVAL_290;
  assign _EVAL_271 = _EVAL_534 & _EVAL_419;
  assign _EVAL_309 = _EVAL_423 | _EVAL_271;
  assign _EVAL_617 = _EVAL_347 | _EVAL_565;
  assign _EVAL_278 = _EVAL_576 & _EVAL_112;
  assign _EVAL_247 = _EVAL_534 & _EVAL_278;
  assign _EVAL_573 = _EVAL_617 | _EVAL_247;
  assign _EVAL_355 = _EVAL_576 & _EVAL_372;
  assign _EVAL_442 = _EVAL_534 & _EVAL_355;
  assign _EVAL_91 = _EVAL_617 | _EVAL_442;
  assign _EVAL_159 = {_EVAL_342,_EVAL_57,_EVAL_445,_EVAL_385,_EVAL_309,_EVAL_604,_EVAL_573,_EVAL_91};
  assign _EVAL_92 = _EVAL == _EVAL_159;
  assign _EVAL_517 = _EVAL_92 | _EVAL_23;
  assign _EVAL_188 = _EVAL_517 == 1'h0;
  assign _EVAL_514 = _EVAL_587 | _EVAL_23;
  assign _EVAL_393 = _EVAL_514 == 1'h0;
  assign _EVAL_296 = _EVAL_6 == 3'h4;
  assign _EVAL_386 = _EVAL_28 & _EVAL_296;
  assign _EVAL_455 = _EVAL_7 == 1'h0;
  assign _EVAL_448 = _EVAL_455 | _EVAL_23;
  assign _EVAL_611 = _EVAL_252 == 5'h0;
  assign _EVAL_575 = _EVAL_18[2];
  assign _EVAL_624 = _EVAL_575 == 1'h0;
  assign _EVAL_553 = _EVAL_252 - 5'h1;
  assign _EVAL_446 = _EVAL_631 != 8'h0;
  assign _EVAL_287 = _EVAL_446 == 1'h0;
  assign _EVAL_625 = _EVAL_600 | _EVAL_23;
  assign _EVAL_257 = _EVAL_5 <= 4'h6;
  assign _EVAL_177 = _EVAL_257 & _EVAL_114;
  assign _EVAL_486 = _EVAL_177 | _EVAL_23;
  assign _EVAL_220 = _EVAL_29 != 2'h2;
  assign _EVAL_37 = _EVAL_220 | _EVAL_23;
  assign _EVAL_77 = _EVAL_37 == 1'h0;
  assign _EVAL_368 = _EVAL_32 == 3'h1;
  assign _EVAL_97 = _EVAL_485 - 5'h1;
  assign _EVAL_364 = _EVAL_6 == 3'h5;
  assign _EVAL_218 = _EVAL_28 & _EVAL_364;
  assign _EVAL_209 = 2'h1 << _EVAL_20;
  assign _EVAL_417 = _EVAL_543 ? _EVAL_209 : 2'h0;
  assign _EVAL_291 = ~ _EVAL_417;
  assign _EVAL_596 = _EVAL_31 == 3'h0;
  assign _EVAL_363 = _EVAL_18 == 3'h4;
  assign _EVAL_103 = _EVAL_33 & _EVAL_363;
  assign _EVAL_196 = _EVAL_32 == 3'h7;
  assign _EVAL_502 = _EVAL_384 == 5'h0;
  assign _EVAL_68 = _EVAL_502 == 1'h0;
  assign _EVAL_416 = _EVAL_27 & _EVAL_68;
  assign _EVAL_108 = _EVAL_25 == 3'h0;
  assign _EVAL_578 = 3'h1 <= _EVAL_25;
  assign _EVAL_581 = _EVAL_108 | _EVAL_578;
  assign _EVAL_330 = _EVAL_235 | _EVAL_23;
  assign _EVAL_52 = _EVAL_330 == 1'h0;
  assign _EVAL_521 = _EVAL_6 == 3'h1;
  assign _EVAL_89 = _EVAL_28 & _EVAL_521;
  assign _EVAL_418 = _EVAL_31 <= 3'h3;
  assign _EVAL_383 = _EVAL_418 | _EVAL_23;
  assign _EVAL_136 = _EVAL_31 == _EVAL_391;
  assign _EVAL_599 = _EVAL_136 | _EVAL_23;
  assign _EVAL_187 = _EVAL_144 >> _EVAL_20;
  assign _EVAL_128 = _EVAL_2 <= 3'h5;
  assign _EVAL_361 = _EVAL_18 == 3'h1;
  assign _EVAL_519 = _EVAL_490 >> _EVAL_26;
  assign _EVAL_334 = _EVAL_8 & _EVAL_368;
  assign _EVAL_482 = _EVAL_21 == _EVAL_609;
  assign _EVAL_171 = _EVAL_482 | _EVAL_23;
  assign _EVAL_232 = _EVAL_2 <= 3'h2;
  assign _EVAL_487 = _EVAL_567 | _EVAL_23;
  assign _EVAL_621 = _EVAL_487 == 1'h0;
  assign _EVAL_373 = _EVAL_508 | _EVAL_299;
  assign _EVAL_619 = _EVAL_194 + 32'h1;
  assign _EVAL_356 = _EVAL_0 == _EVAL_443;
  assign _EVAL_264 = _EVAL_590 | _EVAL_23;
  assign _EVAL_180 = _EVAL_264 == 1'h0;
  assign _EVAL_331 = _EVAL_18 == 3'h3;
  assign _EVAL_470 = _EVAL_18 == _EVAL_238;
  assign _EVAL_430 = _EVAL_17 <= 4'h6;
  assign _EVAL_358 = _EVAL_430 & _EVAL_529;
  assign _EVAL_86 = _EVAL_358 | _EVAL_23;
  assign _EVAL_378 = _EVAL_86 == 1'h0;
  assign _EVAL_344 = _EVAL_33 & _EVAL_331;
  assign _EVAL_277 = _EVAL_379 - 5'h1;
  assign _EVAL_172 = _EVAL_401 | _EVAL_601;
  assign _EVAL_447 = _EVAL_28 & _EVAL_314;
  assign _EVAL_261 = _EVAL_318 - 5'h1;
  assign _EVAL_66 = _EVAL_299 & _EVAL_106;
  assign _EVAL_569 = _EVAL_29 == _EVAL_327;
  assign _EVAL_116 = _EVAL_569 | _EVAL_23;
  assign _EVAL_126 = _EVAL_116 == 1'h0;
  assign _EVAL_181 = _EVAL_187[0];
  assign _EVAL_488 = _EVAL_383 == 1'h0;
  assign _EVAL_214 = _EVAL_0 & 32'h3f;
  assign _EVAL_586 = _EVAL_214 == 32'h0;
  assign _EVAL_70 = _EVAL_6 == _EVAL_464;
  assign _EVAL_294 = _EVAL_70 | _EVAL_23;
  assign _EVAL_362 = _EVAL_294 == 1'h0;
  assign _EVAL_570 = _EVAL_232 | _EVAL_23;
  assign _EVAL_289 = _EVAL_6 <= 3'h6;
  assign _EVAL_120 = _EVAL_509 == 1'h0;
  assign _EVAL_479 = _EVAL_503 == 8'h0;
  assign _EVAL_303 = _EVAL_479 | _EVAL_23;
  assign _EVAL_580 = _EVAL_303 == 1'h0;
  assign _EVAL_484 = {{24'd0}, _EVAL_241};
  assign _EVAL_634 = _EVAL_19 & _EVAL_484;
  assign _EVAL_491 = _EVAL_490 != 8'h0;
  assign _EVAL_403 = _EVAL_491 == 1'h0;
  assign _EVAL_79 = plusarg_reader_out == 32'h0;
  assign _EVAL_95 = _EVAL_403 | _EVAL_79;
  assign _EVAL_222 = _EVAL_194 < plusarg_reader_out;
  assign _EVAL_496 = _EVAL_95 | _EVAL_222;
  assign _EVAL_454 = _EVAL_19 == _EVAL_94;
  assign _EVAL_520 = _EVAL_454 | _EVAL_23;
  assign _EVAL_167 = _EVAL_520 == 1'h0;
  assign _EVAL_164 = _EVAL_25 == _EVAL_345;
  assign _EVAL_438 = _EVAL_164 | _EVAL_23;
  assign _EVAL_105 = _EVAL_438 == 1'h0;
  assign _EVAL_153 = _EVAL_128 | _EVAL_23;
  assign _EVAL_246 = _EVAL_519[0];
  assign _EVAL_90 = _EVAL_246 == 1'h0;
  assign _EVAL_542 = _EVAL_401 >> _EVAL_30;
  assign _EVAL_375 = _EVAL_162 == 1'h0;
  assign _EVAL_436 = _EVAL_384 - 5'h1;
  assign _EVAL_426 = _EVAL_15 == _EVAL_398;
  assign _EVAL_110 = _EVAL_356 | _EVAL_23;
  assign _EVAL_628 = _EVAL_110 == 1'h0;
  assign _EVAL_461 = _EVAL_33 & _EVAL_145;
  assign _EVAL_550 = _EVAL_542[0];
  assign _EVAL_93 = _EVAL_550 == 1'h0;
  assign _EVAL_568 = _EVAL_611 == 1'h0;
  assign _EVAL_88 = _EVAL_33 & _EVAL_568;
  assign _EVAL_474 = _EVAL_32 == 3'h4;
  assign _EVAL_380 = _EVAL_8 & _EVAL_474;
  assign _EVAL_150 = _EVAL_631 != _EVAL_472;
  assign _EVAL_233 = _EVAL_594 | _EVAL_23;
  assign _EVAL_524 = _EVAL_411 | _EVAL_23;
  assign _EVAL_434 = _EVAL_524 == 1'h0;
  assign _EVAL_118 = _EVAL_596 | _EVAL_23;
  assign _EVAL_203 = _EVAL_4 & _EVAL_27;
  assign _EVAL_125 = _EVAL_210 | _EVAL_561;
  assign _EVAL_527 = _EVAL_233 == 1'h0;
  assign _EVAL_537 = _EVAL_26 == _EVAL_117;
  assign _EVAL_320 = _EVAL_537 | _EVAL_23;
  assign _EVAL_437 = _EVAL_150 | _EVAL_287;
  assign _EVAL_65 = _EVAL_107 == 1'h0;
  assign _EVAL_387 = _EVAL_490 | _EVAL_631;
  assign _EVAL_229 = _EVAL_387 & _EVAL_248;
  assign _EVAL_341 = _EVAL_448 == 1'h0;
  assign _EVAL_301 = _EVAL_11 == _EVAL_283;
  assign _EVAL_269 = _EVAL_18 == 3'h6;
  assign _EVAL_610 = _EVAL_450 >> _EVAL_25;
  assign _EVAL_259 = _EVAL_610[0];
  assign _EVAL_272 = _EVAL_259 | _EVAL_23;
  assign _EVAL_39 = _EVAL_272 == 1'h0;
  assign _EVAL_273 = ~ _EVAL_159;
  assign _EVAL_467 = _EVAL & _EVAL_273;
  assign _EVAL_284 = _EVAL_467 == 8'h0;
  assign _EVAL_444 = _EVAL_284 | _EVAL_23;
  assign _EVAL_98 = _EVAL_634 == 32'h0;
  assign _EVAL_236 = _EVAL_98 | _EVAL_23;
  assign _EVAL_306 = _EVAL_31 != 3'h0;
  assign _EVAL_169 = _EVAL_306 | _EVAL_23;
  assign _EVAL_270 = _EVAL_169 == 1'h0;
  assign _EVAL_78 = _EVAL_350 | _EVAL_23;
  assign _EVAL_197 = _EVAL_78 == 1'h0;
  assign _EVAL_133 = _EVAL_431 == 1'h0;
  assign _EVAL_165 = _EVAL_444 == 1'h0;
  assign _EVAL_100 = _EVAL_486 == 1'h0;
  assign _EVAL_158 = _EVAL_508 & _EVAL_611;
  assign _EVAL_544 = _EVAL_171 == 1'h0;
  assign _EVAL_244 = _EVAL_6 == 3'h2;
  assign _EVAL_240 = _EVAL_28 & _EVAL_244;
  assign _EVAL_207 = _EVAL_554 & _EVAL_46;
  assign _EVAL_199 = _EVAL_125 | _EVAL_612;
  assign _EVAL_381 = _EVAL_199 | _EVAL_198;
  assign _EVAL_249 = _EVAL_257 & _EVAL_381;
  assign _EVAL_121 = _EVAL_249 | _EVAL_626;
  assign _EVAL_216 = _EVAL_121 | _EVAL_23;
  assign _EVAL_593 = _EVAL_216 == 1'h0;
  assign _EVAL_161 = _EVAL_33 & _EVAL_361;
  assign _EVAL_223 = _EVAL_483 | _EVAL_23;
  assign _EVAL_607 = _EVAL_320 == 1'h0;
  assign _EVAL_275 = _EVAL_6 == 3'h0;
  assign _EVAL_494 = _EVAL_28 & _EVAL_275;
  assign _EVAL_510 = _EVAL_262 == 1'h0;
  assign _EVAL_200 = _EVAL_67 | _EVAL_23;
  assign _EVAL_515 = _EVAL_559 == 1'h0;
  assign _EVAL_360 = _EVAL_181 | _EVAL_23;
  assign _EVAL_588 = _EVAL_93 | _EVAL_23;
  assign _EVAL_501 = _EVAL_18 == 3'h7;
  assign _EVAL_48 = _EVAL_33 & _EVAL_501;
  assign _EVAL_504 = _EVAL_172 & _EVAL_291;
  assign _EVAL_322 = _EVAL_5 == _EVAL_408;
  assign _EVAL_613 = _EVAL_496 | _EVAL_23;
  assign _EVAL_185 = _EVAL_613 == 1'h0;
  assign _EVAL_505 = _EVAL_322 | _EVAL_23;
  assign _EVAL_193 = _EVAL_586 | _EVAL_23;
  assign _EVAL_119 = _EVAL_301 | _EVAL_23;
  assign _EVAL_583 = _EVAL_119 == 1'h0;
  assign _EVAL_478 = _EVAL_193 == 1'h0;
  assign _EVAL_62 = _EVAL_236 == 1'h0;
  assign _EVAL_183 = _EVAL_153 == 1'h0;
  assign _EVAL_282 = _EVAL_426 | _EVAL_23;
  assign _EVAL_374 = _EVAL_410 == 1'h0;
  assign _EVAL_221 = _EVAL_470 | _EVAL_23;
  assign _EVAL_538 = _EVAL_33 & _EVAL_101;
  assign _EVAL_295 = _EVAL_599 == 1'h0;
  assign _EVAL_302 = _EVAL_437 | _EVAL_23;
  assign _EVAL_43 = _EVAL_33 & _EVAL_269;
  assign _EVAL_566 = _EVAL_289 | _EVAL_23;
  assign _EVAL_175 = _EVAL_566 == 1'h0;
  assign _EVAL_230 = _EVAL_32 == 3'h6;
  assign _EVAL_74 = _EVAL_8 & _EVAL_230;
  assign _EVAL_618 = _EVAL_221 == 1'h0;
  assign _EVAL_191 = _EVAL_282 == 1'h0;
  assign _EVAL_481 = _EVAL_223 == 1'h0;
  assign _EVAL_45 = _EVAL_302 == 1'h0;
  assign _EVAL_562 = _EVAL_469 == 1'h0;
  assign _EVAL_173 = _EVAL_18 == 3'h2;
  assign _EVAL_47 = _EVAL_505 == 1'h0;
  assign _EVAL_307 = _EVAL_33 & _EVAL_173;
  assign _EVAL_492 = _EVAL_90 | _EVAL_23;
  assign _EVAL_471 = _EVAL_203 & _EVAL_502;
  assign _EVAL_522 = _EVAL_625 == 1'h0;
  assign _EVAL_441 = _EVAL_46 == 1'h0;
  assign _EVAL_414 = _EVAL_8 & _EVAL_441;
  assign _EVAL_526 = _EVAL_118 == 1'h0;
  assign _EVAL_463 = _EVAL_32 == 3'h2;
  assign _EVAL_433 = _EVAL_200 == 1'h0;
  assign _EVAL_176 = _EVAL_8 & _EVAL_196;
  assign _EVAL_406 = _EVAL_581 | _EVAL_23;
  assign _EVAL_392 = _EVAL_406 == 1'h0;
  assign _EVAL_34 = _EVAL_588 == 1'h0;
  assign _EVAL_234 = _EVAL_360 == 1'h0;
  assign _EVAL_129 = _EVAL_570 == 1'h0;
  assign _EVAL_312 = _EVAL_492 == 1'h0;
  assign _EVAL_459 = _EVAL_563 | _EVAL_23;
  assign _EVAL_598 = _EVAL_83 == 1'h0;
  assign _EVAL_64 = _EVAL_459 == 1'h0;
  assign _EVAL_40 = _EVAL_8 & _EVAL_463;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_94 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_117 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_194 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_238 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_252 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_266 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_283 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_318 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_327 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_340 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_345 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_354 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_359 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_379 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_384 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_391 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_398 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_401 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_408 = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_443 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_464 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_485 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_490 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_506 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_525 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_585 = _RAND_25[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_609 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_616 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_13) begin
    if (_EVAL_158) begin
      _EVAL_94 <= _EVAL_19;
    end
    if (_EVAL_158) begin
      _EVAL_117 <= _EVAL_26;
    end
    if (_EVAL_23) begin
      _EVAL_194 <= 32'h0;
    end else begin
      if (_EVAL_373) begin
        _EVAL_194 <= 32'h0;
      end else begin
        _EVAL_194 <= _EVAL_619;
      end
    end
    if (_EVAL_158) begin
      _EVAL_238 <= _EVAL_18;
    end
    if (_EVAL_23) begin
      _EVAL_252 <= 5'h0;
    end else begin
      if (_EVAL_508) begin
        if (_EVAL_611) begin
          if (_EVAL_624) begin
            _EVAL_252 <= _EVAL_155;
          end else begin
            _EVAL_252 <= 5'h0;
          end
        end else begin
          _EVAL_252 <= _EVAL_553;
        end
      end
    end
    if (_EVAL_23) begin
      _EVAL_266 <= 5'h0;
    end else begin
      if (_EVAL_299) begin
        if (_EVAL_106) begin
          if (_EVAL_388) begin
            _EVAL_266 <= _EVAL_124;
          end else begin
            _EVAL_266 <= 5'h0;
          end
        end else begin
          _EVAL_266 <= _EVAL_466;
        end
      end
    end
    if (_EVAL_66) begin
      _EVAL_283 <= _EVAL_11;
    end
    if (_EVAL_23) begin
      _EVAL_318 <= 5'h0;
    end else begin
      if (_EVAL_508) begin
        if (_EVAL_476) begin
          if (_EVAL_624) begin
            _EVAL_318 <= _EVAL_155;
          end else begin
            _EVAL_318 <= 5'h0;
          end
        end else begin
          _EVAL_318 <= _EVAL_261;
        end
      end
    end
    if (_EVAL_66) begin
      _EVAL_327 <= _EVAL_29;
    end
    if (_EVAL_66) begin
      _EVAL_340 <= _EVAL_9;
    end
    if (_EVAL_66) begin
      _EVAL_345 <= _EVAL_25;
    end
    if (_EVAL_23) begin
      _EVAL_354 <= 5'h0;
    end else begin
      if (_EVAL_554) begin
        if (_EVAL_46) begin
          if (_EVAL_123) begin
            _EVAL_354 <= _EVAL_574;
          end else begin
            _EVAL_354 <= 5'h0;
          end
        end else begin
          _EVAL_354 <= _EVAL_532;
        end
      end
    end
    if (_EVAL_207) begin
      _EVAL_359 <= _EVAL_2;
    end
    if (_EVAL_23) begin
      _EVAL_379 <= 5'h0;
    end else begin
      if (_EVAL_299) begin
        if (_EVAL_253) begin
          if (_EVAL_388) begin
            _EVAL_379 <= _EVAL_124;
          end else begin
            _EVAL_379 <= 5'h0;
          end
        end else begin
          _EVAL_379 <= _EVAL_277;
        end
      end
    end
    if (_EVAL_23) begin
      _EVAL_384 <= 5'h0;
    end else begin
      if (_EVAL_203) begin
        if (_EVAL_502) begin
          _EVAL_384 <= 5'h0;
        end else begin
          _EVAL_384 <= _EVAL_436;
        end
      end
    end
    if (_EVAL_158) begin
      _EVAL_391 <= _EVAL_31;
    end
    if (_EVAL_207) begin
      _EVAL_398 <= _EVAL_15;
    end
    if (_EVAL_23) begin
      _EVAL_401 <= 2'h0;
    end else begin
      _EVAL_401 <= _EVAL_504;
    end
    if (_EVAL_158) begin
      _EVAL_408 <= _EVAL_5;
    end
    if (_EVAL_471) begin
      _EVAL_443 <= _EVAL_0;
    end
    if (_EVAL_66) begin
      _EVAL_464 <= _EVAL_6;
    end
    if (_EVAL_23) begin
      _EVAL_485 <= 5'h0;
    end else begin
      if (_EVAL_299) begin
        if (_EVAL_115) begin
          if (_EVAL_388) begin
            _EVAL_485 <= _EVAL_124;
          end else begin
            _EVAL_485 <= 5'h0;
          end
        end else begin
          _EVAL_485 <= _EVAL_97;
        end
      end
    end
    if (_EVAL_23) begin
      _EVAL_490 <= 8'h0;
    end else begin
      _EVAL_490 <= _EVAL_229;
    end
    if (_EVAL_207) begin
      _EVAL_506 <= _EVAL_32;
    end
    if (_EVAL_66) begin
      _EVAL_525 <= _EVAL_30;
    end
    if (_EVAL_207) begin
      _EVAL_585 <= _EVAL_17;
    end
    if (_EVAL_207) begin
      _EVAL_609 <= _EVAL_21;
    end
    if (_EVAL_471) begin
      _EVAL_616 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6252cea1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_541) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c3dcd73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_522) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22770767)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ab584a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(361b8048)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aca78f84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59236efe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c343447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_607) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70f278a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_618) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bd1cca4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25da6bfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_481) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb3ef15d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_622) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f50458e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53a2e087)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_393) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d1ff78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_580) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15e0c15b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_375) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69ee4c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_393) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_618) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df4a88e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_515) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_543 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_527) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(194b9e5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_583) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_527) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e247023)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4639732c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61915890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_533) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcc82905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b4b12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_515) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72f41a6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_416 & _EVAL_497) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_475) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fefa2cef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_375) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611ad937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24038582)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fbbeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_475) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_478) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74024b40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_541) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d34bff6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c26720c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7457a2a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf72239b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e19edad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c93303b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14f7ee8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_533) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_598) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f71221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_375) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_583) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(906e1f8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_593) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc98bc33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14bcd3bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_562) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eef58e55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50a88347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_481) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed9579b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_621) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(603740f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_393) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6f57e2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa6d2bfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b59a877)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d3f2499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b57f125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_362) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_607) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_393) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b66b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_433) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a6d1a02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64bf43cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33acd05c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_481) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64653bee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_593) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2fcc48a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f77c1c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe971dbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49e609cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_543 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2758751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_580) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bac01fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_527) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d05fe6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c0334aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ca1558)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_622) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b9a218f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a82ce00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_522) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(282745f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_598) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8168e84a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_562) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec8aa2a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52befbfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_544) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f087e6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a853ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_478) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70ed4de3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_416 & _EVAL_628) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c126e681)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830c37a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_598) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e322dc87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18692c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e384a09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_562) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_593) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_598) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(260f0425)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a90d8cd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_434) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1f5269)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_533) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5941c87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98414c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6f5f49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_533) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f243b21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_544) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7278f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c478350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_562) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9771a61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f35ab1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_527) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3d5cd40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_374) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(742a6ba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(262762d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_488) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad7a3683)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_374) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_362) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5d2f934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66b7674c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89e2a28f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc2b8200)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89eb2bb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86ef3830)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(180df7be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_433) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_433) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_527) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d52d801)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(400b42ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9374cfa8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c96a586e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_481) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33b29224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_481) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cacf699)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14ddc250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7ab9949)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e364fbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_481) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64414ed3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c87cfc11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb9864cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_527) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52f97f63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_481) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_416 & _EVAL_628) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a0e5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_434) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2834bd8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_416 & _EVAL_497) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e74623c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_481) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ed7e4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab6811ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d60dfe0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_375) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_593) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bd1b448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_593) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_621) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3a45656)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e79dfa82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87fae5d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25d788b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9472627)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_433) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b7d6cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f12bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bcfc082)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(216c3b48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a7a9d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67c97c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_334 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_622) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12b2618f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_488) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_622) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96554803)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13549432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_593) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f06b0c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7c28023)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4f9249d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816ab2a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
