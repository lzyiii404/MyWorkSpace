//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_121_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [29:0] _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [6:0]  _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [6:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_26;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_35;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_48;
  reg [31:0] _RAND_2;
  reg [5:0] _EVAL_62;
  reg [31:0] _RAND_3;
  reg [5:0] _EVAL_102;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_120;
  reg [31:0] _RAND_5;
  reg [29:0] _EVAL_172;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_205;
  reg [31:0] _RAND_7;
  reg [6:0] _EVAL_209;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_235;
  reg [31:0] _RAND_9;
  reg [31:0] _EVAL_247;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_254;
  reg [31:0] _RAND_11;
  reg  _EVAL_267;
  reg [31:0] _RAND_12;
  reg [72:0] _EVAL_270;
  reg [95:0] _RAND_13;
  reg [3:0] _EVAL_271;
  reg [31:0] _RAND_14;
  reg [5:0] _EVAL_303;
  reg [31:0] _RAND_15;
  reg [1:0] _EVAL_351;
  reg [31:0] _RAND_16;
  wire  _EVAL_137;
  wire  _EVAL_107;
  wire  _EVAL_117;
  wire [3:0] _EVAL_241;
  wire  _EVAL_367;
  wire [2:0] _EVAL_160;
  wire  _EVAL_299;
  wire  _EVAL_119;
  wire  _EVAL_325;
  wire  _EVAL_25;
  wire  _EVAL_255;
  wire  _EVAL_245;
  wire  _EVAL_98;
  wire  _EVAL_244;
  wire  _EVAL_292;
  wire  _EVAL_278;
  wire [127:0] _EVAL_144;
  wire [127:0] _EVAL_243;
  wire [72:0] _EVAL_87;
  wire  _EVAL_362;
  wire  _EVAL_310;
  wire  _EVAL_210;
  wire [1:0] _EVAL_288;
  wire [1:0] _EVAL_263;
  wire  _EVAL_142;
  wire  _EVAL_315;
  wire  _EVAL_162;
  wire  _EVAL_156;
  wire  _EVAL_215;
  wire  _EVAL_317;
  wire  _EVAL_258;
  wire  _EVAL_128;
  wire  _EVAL_248;
  wire  _EVAL_207;
  wire  _EVAL_78;
  wire  _EVAL_208;
  wire  _EVAL_342;
  wire  _EVAL_33;
  wire  _EVAL_301;
  wire  _EVAL_273;
  wire  _EVAL_345;
  wire  _EVAL_356;
  wire  _EVAL_24;
  wire  _EVAL_371;
  wire  _EVAL_281;
  wire  _EVAL_114;
  wire [3:0] _EVAL_29;
  wire [3:0] _EVAL_202;
  wire [3:0] _EVAL_77;
  wire  _EVAL_199;
  wire  _EVAL_67;
  wire  _EVAL_219;
  wire [30:0] _EVAL_94;
  wire [30:0] _EVAL_239;
  wire [30:0] _EVAL_108;
  wire  _EVAL_195;
  wire [29:0] _EVAL_196;
  wire [30:0] _EVAL_192;
  wire [72:0] _EVAL_151;
  wire [22:0] _EVAL_55;
  wire [7:0] _EVAL_136;
  wire [7:0] _EVAL_272;
  wire [29:0] _EVAL_358;
  wire  _EVAL_135;
  wire  _EVAL_256;
  wire  _EVAL_354;
  wire [5:0] _EVAL_90;
  wire [5:0] _EVAL_253;
  wire  _EVAL_50;
  wire  _EVAL_121;
  wire  _EVAL_264;
  wire  _EVAL_131;
  wire  _EVAL_282;
  wire  _EVAL_110;
  wire  _EVAL_28;
  wire [29:0] _EVAL_164;
  wire [30:0] _EVAL_75;
  wire [30:0] _EVAL_181;
  wire [30:0] _EVAL_150;
  wire  _EVAL_340;
  wire  _EVAL_296;
  wire  _EVAL_228;
  wire  _EVAL_279;
  wire [29:0] _EVAL_169;
  wire [30:0] _EVAL_49;
  wire [30:0] _EVAL_159;
  wire [30:0] _EVAL_88;
  wire  _EVAL_116;
  wire  _EVAL_237;
  wire  _EVAL_307;
  wire  _EVAL_41;
  wire  _EVAL_225;
  wire  _EVAL_52;
  wire  _EVAL_313;
  wire [127:0] _EVAL_47;
  wire [127:0] _EVAL_141;
  wire [72:0] _EVAL_106;
  wire [72:0] _EVAL_190;
  wire [72:0] _EVAL_262;
  wire  _EVAL_324;
  wire  _EVAL_124;
  wire  _EVAL_73;
  wire [29:0] _EVAL_132;
  wire [30:0] _EVAL_188;
  wire [30:0] _EVAL_34;
  wire [30:0] _EVAL_129;
  wire  _EVAL_21;
  wire [30:0] _EVAL_126;
  wire [30:0] _EVAL_191;
  wire  _EVAL_236;
  wire  _EVAL_189;
  wire  _EVAL_39;
  wire [29:0] _EVAL_234;
  wire [30:0] _EVAL_139;
  wire [30:0] _EVAL_61;
  wire [30:0] _EVAL_53;
  wire  _EVAL_333;
  wire  _EVAL_212;
  wire  _EVAL_80;
  wire [29:0] _EVAL_173;
  wire [30:0] _EVAL_266;
  wire [30:0] _EVAL_68;
  wire [30:0] _EVAL_185;
  wire  _EVAL_252;
  wire  _EVAL_331;
  wire  _EVAL_155;
  wire  _EVAL_64;
  wire  _EVAL_20;
  wire  _EVAL_166;
  wire  _EVAL_229;
  wire [22:0] _EVAL_182;
  wire [7:0] _EVAL_361;
  wire [7:0] _EVAL_277;
  wire [5:0] _EVAL_218;
  wire  _EVAL_360;
  wire  _EVAL_348;
  wire  _EVAL_60;
  wire  _EVAL_224;
  wire  _EVAL_355;
  wire  _EVAL_147;
  wire  _EVAL_314;
  wire  _EVAL_289;
  wire  _EVAL_183;
  wire  _EVAL_284;
  wire  _EVAL_216;
  wire  _EVAL_31;
  wire  _EVAL_127;
  wire  _EVAL_274;
  wire  _EVAL_369;
  wire  _EVAL_95;
  wire  _EVAL_138;
  wire  _EVAL_122;
  wire  _EVAL_319;
  wire  _EVAL_322;
  wire  _EVAL_339;
  wire  _EVAL_359;
  wire [3:0] _EVAL_276;
  wire  _EVAL_320;
  wire [2:0] _EVAL_349;
  wire  _EVAL_338;
  wire  _EVAL_153;
  wire  _EVAL_99;
  wire  _EVAL_163;
  wire [5:0] _EVAL_285;
  wire  _EVAL_194;
  wire  _EVAL_242;
  wire  _EVAL_347;
  wire  _EVAL_201;
  wire  _EVAL_96;
  wire  _EVAL_148;
  wire  _EVAL_174;
  wire  _EVAL_109;
  wire  _EVAL_353;
  wire  _EVAL_69;
  wire  _EVAL_145;
  wire  _EVAL_154;
  wire  _EVAL_193;
  wire  _EVAL_89;
  wire  _EVAL_306;
  wire  _EVAL_335;
  wire  _EVAL_357;
  wire  _EVAL_58;
  wire  _EVAL_286;
  wire  _EVAL_93;
  wire  _EVAL_186;
  wire  _EVAL_36;
  wire  _EVAL_295;
  wire  _EVAL_125;
  wire  _EVAL_346;
  wire  _EVAL_350;
  wire  _EVAL_38;
  wire  _EVAL_45;
  wire [29:0] _EVAL_220;
  wire  _EVAL_246;
  wire  _EVAL_170;
  wire  _EVAL_309;
  wire  _EVAL_293;
  wire  _EVAL_365;
  wire  _EVAL_175;
  wire  _EVAL_76;
  wire  _EVAL_275;
  wire  _EVAL_140;
  wire  _EVAL_261;
  wire  _EVAL_321;
  wire  _EVAL_206;
  wire  _EVAL_251;
  wire  _EVAL_240;
  wire  _EVAL_323;
  wire  _EVAL_81;
  wire  _EVAL_54;
  wire  _EVAL_334;
  wire  _EVAL_23;
  wire [72:0] _EVAL_318;
  wire [72:0] _EVAL_343;
  wire  _EVAL_149;
  wire  _EVAL_84;
  wire  _EVAL_352;
  wire  _EVAL_312;
  wire  _EVAL_19;
  wire  _EVAL_180;
  wire  _EVAL_198;
  wire  _EVAL_221;
  wire  _EVAL_32;
  wire [5:0] _EVAL_30;
  wire  _EVAL_305;
  wire  _EVAL_213;
  wire  _EVAL_233;
  wire  _EVAL_308;
  wire  _EVAL_167;
  wire  _EVAL_197;
  wire  _EVAL_113;
  wire [72:0] _EVAL_341;
  wire  _EVAL_203;
  wire  _EVAL_130;
  wire  _EVAL_71;
  wire  _EVAL_123;
  wire  _EVAL_134;
  wire  _EVAL_304;
  wire  _EVAL_302;
  wire  _EVAL_370;
  wire [31:0] _EVAL_146;
  wire  _EVAL_63;
  wire  _EVAL_368;
  wire  _EVAL_152;
  wire  _EVAL_298;
  wire  _EVAL_311;
  wire  _EVAL_269;
  wire  _EVAL_265;
  wire  _EVAL_364;
  wire  _EVAL_217;
  wire  _EVAL_104;
  wire  _EVAL_344;
  wire  _EVAL_37;
  wire  _EVAL_232;
  wire [5:0] _EVAL_337;
  wire  _EVAL_316;
  wire  _EVAL_59;
  wire  _EVAL_105;
  wire  _EVAL_250;
  wire  _EVAL_171;
  wire  _EVAL_40;
  wire  _EVAL_187;
  wire  _EVAL_200;
  wire  _EVAL_65;
  wire  _EVAL_101;
  wire  _EVAL_178;
  wire  _EVAL_332;
  wire  _EVAL_51;
  wire  _EVAL_283;
  wire  _EVAL_231;
  wire  _EVAL_329;
  wire  _EVAL_85;
  wire  _EVAL_43;
  wire  _EVAL_91;
  wire  _EVAL_249;
  wire  _EVAL_56;
  wire  _EVAL_300;
  wire  _EVAL_92;
  wire  _EVAL_27;
  wire  _EVAL_44;
  wire  _EVAL_363;
  wire [3:0] _EVAL_100;
  wire  _EVAL_42;
  wire  _EVAL_161;
  wire  _EVAL_158;
  wire  _EVAL_46;
  wire  _EVAL_226;
  wire  _EVAL_168;
  wire  _EVAL_214;
  wire  _EVAL_112;
  wire  _EVAL_118;
  wire  _EVAL_70;
  wire  _EVAL_294;
  wire  _EVAL_157;
  wire  _EVAL_179;
  wire  _EVAL_204;
  wire  _EVAL_280;
  wire  _EVAL_260;
  wire  _EVAL_330;
  wire  _EVAL_257;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_238;
  wire  _EVAL_211;
  wire  _EVAL_297;
  wire  _EVAL_97;
  wire  _EVAL_86;
  wire  _EVAL_103;
  wire  _EVAL_83;
  wire  _EVAL_66;
  wire  _EVAL_328;
  wire  _EVAL_57;
  wire  _EVAL_366;
  wire  _EVAL_79;
  wire  _EVAL_327;
  wire  _EVAL_290;
  wire  _EVAL_227;
  wire  _EVAL_165;
  wire  _EVAL_74;
  wire  _EVAL_111;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_137 = _EVAL_13 == 7'h48;
  assign _EVAL_107 = _EVAL_13 == 7'h40;
  assign _EVAL_117 = _EVAL_137 | _EVAL_107;
  assign _EVAL_241 = _EVAL_13[6:3];
  assign _EVAL_367 = _EVAL_241 == 4'h8;
  assign _EVAL_160 = _EVAL_13[2:0];
  assign _EVAL_299 = 3'h1 <= _EVAL_160;
  assign _EVAL_119 = _EVAL_367 & _EVAL_299;
  assign _EVAL_325 = _EVAL_117 | _EVAL_119;
  assign _EVAL_25 = _EVAL_13 == 7'h20;
  assign _EVAL_255 = _EVAL_325 | _EVAL_25;
  assign _EVAL_245 = _EVAL_241 == 4'h0;
  assign _EVAL_98 = _EVAL_255 | _EVAL_245;
  assign _EVAL_244 = _EVAL_6 & _EVAL_12;
  assign _EVAL_292 = _EVAL_235 == 6'h0;
  assign _EVAL_278 = _EVAL_244 & _EVAL_292;
  assign _EVAL_144 = 128'h1 << _EVAL_18;
  assign _EVAL_243 = _EVAL_278 ? _EVAL_144 : 128'h0;
  assign _EVAL_87 = _EVAL_243[72:0];
  assign _EVAL_362 = _EVAL_87 != 73'h0;
  assign _EVAL_310 = _EVAL_16 >= 4'h2;
  assign _EVAL_210 = _EVAL_16[0];
  assign _EVAL_288 = 2'h1 << _EVAL_210;
  assign _EVAL_263 = _EVAL_288 | 2'h1;
  assign _EVAL_142 = _EVAL_263[1];
  assign _EVAL_315 = _EVAL_9[1];
  assign _EVAL_162 = _EVAL_142 & _EVAL_315;
  assign _EVAL_156 = _EVAL_310 | _EVAL_162;
  assign _EVAL_215 = _EVAL_263[0];
  assign _EVAL_317 = _EVAL_9[0];
  assign _EVAL_258 = _EVAL_315 & _EVAL_317;
  assign _EVAL_128 = _EVAL_215 & _EVAL_258;
  assign _EVAL_248 = _EVAL_156 | _EVAL_128;
  assign _EVAL_207 = _EVAL_317 == 1'h0;
  assign _EVAL_78 = _EVAL_315 & _EVAL_207;
  assign _EVAL_208 = _EVAL_215 & _EVAL_78;
  assign _EVAL_342 = _EVAL_156 | _EVAL_208;
  assign _EVAL_33 = _EVAL_315 == 1'h0;
  assign _EVAL_301 = _EVAL_142 & _EVAL_33;
  assign _EVAL_273 = _EVAL_310 | _EVAL_301;
  assign _EVAL_345 = _EVAL_33 & _EVAL_317;
  assign _EVAL_356 = _EVAL_215 & _EVAL_345;
  assign _EVAL_24 = _EVAL_273 | _EVAL_356;
  assign _EVAL_371 = _EVAL_33 & _EVAL_207;
  assign _EVAL_281 = _EVAL_215 & _EVAL_371;
  assign _EVAL_114 = _EVAL_273 | _EVAL_281;
  assign _EVAL_29 = {_EVAL_248,_EVAL_342,_EVAL_24,_EVAL_114};
  assign _EVAL_202 = ~ _EVAL_29;
  assign _EVAL_77 = _EVAL_0 & _EVAL_202;
  assign _EVAL_199 = _EVAL_77 == 4'h0;
  assign _EVAL_67 = _EVAL_199 | _EVAL_2;
  assign _EVAL_219 = _EVAL_102 == 6'h0;
  assign _EVAL_94 = {1'b0,$signed(_EVAL_9)};
  assign _EVAL_239 = $signed(_EVAL_94) & $signed(-31'sh5000);
  assign _EVAL_108 = $signed(_EVAL_239);
  assign _EVAL_195 = $signed(_EVAL_108) == $signed(31'sh0);
  assign _EVAL_196 = _EVAL_9 ^ 30'h2000000;
  assign _EVAL_192 = {1'b0,$signed(_EVAL_196)};
  assign _EVAL_151 = _EVAL_270 | _EVAL_87;
  assign _EVAL_55 = 23'hff << _EVAL_16;
  assign _EVAL_136 = _EVAL_55[7:0];
  assign _EVAL_272 = ~ _EVAL_136;
  assign _EVAL_358 = {{22'd0}, _EVAL_272};
  assign _EVAL_135 = _EVAL_62 == 6'h0;
  assign _EVAL_256 = _EVAL_11[2];
  assign _EVAL_354 = _EVAL_256 == 1'h0;
  assign _EVAL_90 = _EVAL_272[7:2];
  assign _EVAL_253 = _EVAL_62 - 6'h1;
  assign _EVAL_50 = _EVAL_270 != 73'h0;
  assign _EVAL_121 = _EVAL_50 == 1'h0;
  assign _EVAL_264 = plusarg_reader_out == 32'h0;
  assign _EVAL_131 = _EVAL_121 | _EVAL_264;
  assign _EVAL_282 = _EVAL_247 < plusarg_reader_out;
  assign _EVAL_110 = _EVAL_131 | _EVAL_282;
  assign _EVAL_28 = _EVAL_16 <= 4'h8;
  assign _EVAL_164 = _EVAL_9 ^ 30'h3000;
  assign _EVAL_75 = {1'b0,$signed(_EVAL_164)};
  assign _EVAL_181 = $signed(_EVAL_75) & $signed(-31'sh1000);
  assign _EVAL_150 = $signed(_EVAL_181);
  assign _EVAL_340 = $signed(_EVAL_150) == $signed(31'sh0);
  assign _EVAL_296 = _EVAL_28 & _EVAL_340;
  assign _EVAL_228 = _EVAL_296 | _EVAL_2;
  assign _EVAL_279 = _EVAL_4 == 1'h0;
  assign _EVAL_169 = _EVAL_9 ^ 30'h1900000;
  assign _EVAL_49 = {1'b0,$signed(_EVAL_169)};
  assign _EVAL_159 = $signed(_EVAL_49) & $signed(-31'sh2000);
  assign _EVAL_88 = $signed(_EVAL_159);
  assign _EVAL_116 = $signed(_EVAL_88) == $signed(31'sh0);
  assign _EVAL_237 = _EVAL_3 & _EVAL_10;
  assign _EVAL_307 = _EVAL_303 == 6'h0;
  assign _EVAL_41 = _EVAL_237 & _EVAL_307;
  assign _EVAL_225 = _EVAL_17 == 3'h6;
  assign _EVAL_52 = _EVAL_225 == 1'h0;
  assign _EVAL_313 = _EVAL_41 & _EVAL_52;
  assign _EVAL_47 = 128'h1 << _EVAL_13;
  assign _EVAL_141 = _EVAL_313 ? _EVAL_47 : 128'h0;
  assign _EVAL_106 = _EVAL_141[72:0];
  assign _EVAL_190 = ~ _EVAL_106;
  assign _EVAL_262 = _EVAL_151 & _EVAL_190;
  assign _EVAL_324 = _EVAL_11 == 3'h0;
  assign _EVAL_124 = _EVAL_12 & _EVAL_324;
  assign _EVAL_73 = _EVAL_16 <= 4'h6;
  assign _EVAL_132 = _EVAL_9 ^ 30'hc000000;
  assign _EVAL_188 = {1'b0,$signed(_EVAL_132)};
  assign _EVAL_34 = $signed(_EVAL_188) & $signed(-31'sh4000000);
  assign _EVAL_129 = $signed(_EVAL_34);
  assign _EVAL_21 = $signed(_EVAL_129) == $signed(31'sh0);
  assign _EVAL_126 = $signed(_EVAL_192) & $signed(-31'sh10000);
  assign _EVAL_191 = $signed(_EVAL_126);
  assign _EVAL_236 = $signed(_EVAL_191) == $signed(31'sh0);
  assign _EVAL_189 = _EVAL_21 | _EVAL_236;
  assign _EVAL_39 = _EVAL_189 | _EVAL_195;
  assign _EVAL_234 = _EVAL_9 ^ 30'h1800000;
  assign _EVAL_139 = {1'b0,$signed(_EVAL_234)};
  assign _EVAL_61 = $signed(_EVAL_139) & $signed(-31'sh8000);
  assign _EVAL_53 = $signed(_EVAL_61);
  assign _EVAL_333 = $signed(_EVAL_53) == $signed(31'sh0);
  assign _EVAL_212 = _EVAL_39 | _EVAL_333;
  assign _EVAL_80 = _EVAL_212 | _EVAL_116;
  assign _EVAL_173 = _EVAL_9 ^ 30'h20000000;
  assign _EVAL_266 = {1'b0,$signed(_EVAL_173)};
  assign _EVAL_68 = $signed(_EVAL_266) & $signed(-31'sh2000);
  assign _EVAL_185 = $signed(_EVAL_68);
  assign _EVAL_252 = $signed(_EVAL_185) == $signed(31'sh0);
  assign _EVAL_331 = _EVAL_80 | _EVAL_252;
  assign _EVAL_155 = _EVAL_73 & _EVAL_331;
  assign _EVAL_64 = _EVAL_296 | _EVAL_155;
  assign _EVAL_20 = _EVAL_7 <= 3'h3;
  assign _EVAL_166 = _EVAL_20 | _EVAL_2;
  assign _EVAL_229 = _EVAL_166 == 1'h0;
  assign _EVAL_182 = 23'hff << _EVAL_15;
  assign _EVAL_361 = _EVAL_182[7:0];
  assign _EVAL_277 = ~ _EVAL_361;
  assign _EVAL_218 = _EVAL_277[7:2];
  assign _EVAL_360 = _EVAL_14 == _EVAL_267;
  assign _EVAL_348 = _EVAL_14 == 1'h0;
  assign _EVAL_60 = _EVAL_348 | _EVAL_4;
  assign _EVAL_224 = _EVAL_1 == 2'h0;
  assign _EVAL_355 = _EVAL_8 == 1'h0;
  assign _EVAL_147 = _EVAL_355 | _EVAL_2;
  assign _EVAL_314 = _EVAL_147 == 1'h0;
  assign _EVAL_289 = _EVAL_7 <= 3'h2;
  assign _EVAL_183 = _EVAL_289 | _EVAL_2;
  assign _EVAL_284 = _EVAL_183 == 1'h0;
  assign _EVAL_216 = _EVAL_1 != 2'h2;
  assign _EVAL_31 = _EVAL_216 | _EVAL_2;
  assign _EVAL_127 = _EVAL_31 == 1'h0;
  assign _EVAL_274 = _EVAL_241 == 4'h3;
  assign _EVAL_369 = _EVAL_11 == 3'h7;
  assign _EVAL_95 = _EVAL_64 | _EVAL_2;
  assign _EVAL_138 = _EVAL_95 == 1'h0;
  assign _EVAL_122 = _EVAL_241 == 4'h2;
  assign _EVAL_319 = _EVAL_279 | _EVAL_2;
  assign _EVAL_322 = _EVAL_18 == 7'h48;
  assign _EVAL_339 = _EVAL_18 == 7'h40;
  assign _EVAL_359 = _EVAL_322 | _EVAL_339;
  assign _EVAL_276 = _EVAL_18[6:3];
  assign _EVAL_320 = _EVAL_276 == 4'h8;
  assign _EVAL_349 = _EVAL_18[2:0];
  assign _EVAL_338 = 3'h1 <= _EVAL_349;
  assign _EVAL_153 = _EVAL_320 & _EVAL_338;
  assign _EVAL_99 = _EVAL_359 | _EVAL_153;
  assign _EVAL_163 = _EVAL_17[0];
  assign _EVAL_285 = _EVAL_303 - 6'h1;
  assign _EVAL_194 = _EVAL_0 == _EVAL_29;
  assign _EVAL_242 = _EVAL_17 == 3'h0;
  assign _EVAL_347 = _EVAL_10 & _EVAL_242;
  assign _EVAL_201 = _EVAL_11 == _EVAL_205;
  assign _EVAL_96 = _EVAL_201 | _EVAL_2;
  assign _EVAL_148 = _EVAL_96 == 1'h0;
  assign _EVAL_174 = _EVAL_7 == 3'h0;
  assign _EVAL_109 = _EVAL_174 | _EVAL_2;
  assign _EVAL_353 = _EVAL_109 == 1'h0;
  assign _EVAL_69 = _EVAL_17 == 3'h4;
  assign _EVAL_145 = _EVAL_15 == _EVAL_271;
  assign _EVAL_154 = _EVAL_340 | _EVAL_21;
  assign _EVAL_193 = _EVAL_154 | _EVAL_236;
  assign _EVAL_89 = _EVAL_193 | _EVAL_195;
  assign _EVAL_306 = _EVAL_276 == 4'h0;
  assign _EVAL_335 = _EVAL_18 == 7'h20;
  assign _EVAL_357 = _EVAL_99 | _EVAL_335;
  assign _EVAL_58 = _EVAL_357 | _EVAL_306;
  assign _EVAL_286 = _EVAL_276 == 4'h1;
  assign _EVAL_93 = _EVAL_58 | _EVAL_286;
  assign _EVAL_186 = _EVAL_276 == 4'h2;
  assign _EVAL_36 = _EVAL_93 | _EVAL_186;
  assign _EVAL_295 = _EVAL_276 == 4'h3;
  assign _EVAL_125 = _EVAL_36 | _EVAL_295;
  assign _EVAL_346 = _EVAL_125 | _EVAL_2;
  assign _EVAL_350 = _EVAL_241 == 4'h1;
  assign _EVAL_38 = _EVAL_98 | _EVAL_350;
  assign _EVAL_45 = _EVAL_7 <= 3'h4;
  assign _EVAL_220 = _EVAL_9 & _EVAL_358;
  assign _EVAL_246 = _EVAL_220 == 30'h0;
  assign _EVAL_170 = _EVAL_246 | _EVAL_2;
  assign _EVAL_309 = _EVAL_170 == 1'h0;
  assign _EVAL_293 = _EVAL_1 <= 2'h2;
  assign _EVAL_365 = _EVAL_60 | _EVAL_2;
  assign _EVAL_175 = _EVAL_87 != _EVAL_106;
  assign _EVAL_76 = _EVAL_362 == 1'h0;
  assign _EVAL_275 = _EVAL_175 | _EVAL_76;
  assign _EVAL_140 = _EVAL_16 <= 4'h2;
  assign _EVAL_261 = _EVAL_2 == 1'h0;
  assign _EVAL_321 = _EVAL_7 == _EVAL_48;
  assign _EVAL_206 = _EVAL_321 | _EVAL_2;
  assign _EVAL_251 = _EVAL_206 == 1'h0;
  assign _EVAL_240 = _EVAL_11 == 3'h1;
  assign _EVAL_323 = _EVAL_12 & _EVAL_240;
  assign _EVAL_81 = _EVAL_15 >= 4'h2;
  assign _EVAL_54 = _EVAL_89 | _EVAL_333;
  assign _EVAL_334 = _EVAL_54 | _EVAL_116;
  assign _EVAL_23 = _EVAL_334 | _EVAL_252;
  assign _EVAL_318 = _EVAL_87 | _EVAL_270;
  assign _EVAL_343 = _EVAL_318 >> _EVAL_13;
  assign _EVAL_149 = _EVAL_343[0];
  assign _EVAL_84 = _EVAL_149 | _EVAL_2;
  assign _EVAL_352 = _EVAL_84 == 1'h0;
  assign _EVAL_312 = _EVAL_346 == 1'h0;
  assign _EVAL_19 = _EVAL_17 == _EVAL_254;
  assign _EVAL_180 = _EVAL_19 | _EVAL_2;
  assign _EVAL_198 = _EVAL_180 == 1'h0;
  assign _EVAL_221 = _EVAL_13 == _EVAL_209;
  assign _EVAL_32 = _EVAL_221 | _EVAL_2;
  assign _EVAL_30 = _EVAL_102 - 6'h1;
  assign _EVAL_305 = _EVAL_38 | _EVAL_122;
  assign _EVAL_213 = _EVAL_305 | _EVAL_274;
  assign _EVAL_233 = _EVAL_213 | _EVAL_2;
  assign _EVAL_308 = _EVAL_11 == 3'h4;
  assign _EVAL_167 = _EVAL_12 & _EVAL_308;
  assign _EVAL_197 = _EVAL_10 & _EVAL_69;
  assign _EVAL_113 = _EVAL_10 & _EVAL_225;
  assign _EVAL_341 = _EVAL_270 >> _EVAL_18;
  assign _EVAL_203 = _EVAL_341[0];
  assign _EVAL_130 = _EVAL_203 == 1'h0;
  assign _EVAL_71 = _EVAL_130 | _EVAL_2;
  assign _EVAL_123 = _EVAL_71 == 1'h0;
  assign _EVAL_134 = _EVAL_140 & _EVAL_23;
  assign _EVAL_304 = _EVAL_134 | _EVAL_2;
  assign _EVAL_302 = _EVAL_304 == 1'h0;
  assign _EVAL_370 = _EVAL_244 | _EVAL_237;
  assign _EVAL_146 = _EVAL_247 + 32'h1;
  assign _EVAL_63 = _EVAL_18 == _EVAL_35;
  assign _EVAL_368 = _EVAL_219 == 1'h0;
  assign _EVAL_152 = _EVAL_11 == 3'h3;
  assign _EVAL_298 = _EVAL_12 & _EVAL_152;
  assign _EVAL_311 = _EVAL_224 | _EVAL_2;
  assign _EVAL_269 = _EVAL_9 == _EVAL_172;
  assign _EVAL_265 = _EVAL_269 | _EVAL_2;
  assign _EVAL_364 = _EVAL_63 | _EVAL_2;
  assign _EVAL_217 = _EVAL_17 == 3'h5;
  assign _EVAL_104 = _EVAL_32 == 1'h0;
  assign _EVAL_344 = _EVAL_16 == _EVAL_120;
  assign _EVAL_37 = _EVAL_344 | _EVAL_2;
  assign _EVAL_232 = _EVAL_37 == 1'h0;
  assign _EVAL_337 = _EVAL_235 - 6'h1;
  assign _EVAL_316 = _EVAL_310 | _EVAL_2;
  assign _EVAL_59 = _EVAL_81 | _EVAL_2;
  assign _EVAL_105 = _EVAL_59 == 1'h0;
  assign _EVAL_250 = _EVAL_237 & _EVAL_219;
  assign _EVAL_171 = 4'h6 == _EVAL_16;
  assign _EVAL_40 = _EVAL_339 ? _EVAL_171 : 1'h0;
  assign _EVAL_187 = _EVAL_40 | _EVAL_2;
  assign _EVAL_200 = _EVAL_187 == 1'h0;
  assign _EVAL_65 = _EVAL_7 != 3'h0;
  assign _EVAL_101 = _EVAL_65 | _EVAL_2;
  assign _EVAL_178 = _EVAL_244 & _EVAL_135;
  assign _EVAL_332 = _EVAL_17 == 3'h2;
  assign _EVAL_51 = _EVAL_10 & _EVAL_332;
  assign _EVAL_283 = _EVAL_17 <= 3'h6;
  assign _EVAL_231 = _EVAL_283 | _EVAL_2;
  assign _EVAL_329 = _EVAL_231 == 1'h0;
  assign _EVAL_85 = _EVAL == _EVAL_26;
  assign _EVAL_43 = _EVAL_233 == 1'h0;
  assign _EVAL_91 = _EVAL_135 == 1'h0;
  assign _EVAL_249 = _EVAL_275 | _EVAL_2;
  assign _EVAL_56 = _EVAL_348 | _EVAL_2;
  assign _EVAL_300 = _EVAL_194 | _EVAL_2;
  assign _EVAL_92 = _EVAL_300 == 1'h0;
  assign _EVAL_27 = _EVAL_360 | _EVAL_2;
  assign _EVAL_44 = _EVAL_27 == 1'h0;
  assign _EVAL_363 = _EVAL_249 == 1'h0;
  assign _EVAL_100 = ~ _EVAL_0;
  assign _EVAL_42 = _EVAL_11 == 3'h5;
  assign _EVAL_161 = _EVAL_17 == 3'h1;
  assign _EVAL_158 = _EVAL_10 & _EVAL_161;
  assign _EVAL_46 = _EVAL_85 | _EVAL_2;
  assign _EVAL_226 = _EVAL_100 == 4'h0;
  assign _EVAL_168 = _EVAL_226 | _EVAL_2;
  assign _EVAL_214 = _EVAL_168 == 1'h0;
  assign _EVAL_112 = _EVAL_365 == 1'h0;
  assign _EVAL_118 = _EVAL_56 == 1'h0;
  assign _EVAL_70 = _EVAL_145 | _EVAL_2;
  assign _EVAL_294 = _EVAL_70 == 1'h0;
  assign _EVAL_157 = _EVAL_11 == 3'h2;
  assign _EVAL_179 = _EVAL_319 == 1'h0;
  assign _EVAL_204 = _EVAL_265 == 1'h0;
  assign _EVAL_280 = _EVAL_45 | _EVAL_2;
  assign _EVAL_260 = _EVAL_11 == 3'h6;
  assign _EVAL_330 = _EVAL_228 == 1'h0;
  assign _EVAL_257 = _EVAL_293 | _EVAL_2;
  assign _EVAL_176 = _EVAL_316 == 1'h0;
  assign _EVAL_177 = _EVAL_110 | _EVAL_2;
  assign _EVAL_238 = _EVAL_177 == 1'h0;
  assign _EVAL_211 = _EVAL_101 == 1'h0;
  assign _EVAL_297 = _EVAL_12 & _EVAL_42;
  assign _EVAL_97 = _EVAL_67 == 1'h0;
  assign _EVAL_86 = _EVAL_1 == _EVAL_351;
  assign _EVAL_103 = _EVAL_86 | _EVAL_2;
  assign _EVAL_83 = _EVAL_12 & _EVAL_157;
  assign _EVAL_66 = _EVAL_10 & _EVAL_217;
  assign _EVAL_328 = _EVAL_12 & _EVAL_91;
  assign _EVAL_57 = _EVAL_280 == 1'h0;
  assign _EVAL_366 = _EVAL_257 == 1'h0;
  assign _EVAL_79 = _EVAL_103 == 1'h0;
  assign _EVAL_327 = _EVAL_46 == 1'h0;
  assign _EVAL_290 = _EVAL_311 == 1'h0;
  assign _EVAL_227 = _EVAL_12 & _EVAL_260;
  assign _EVAL_165 = _EVAL_10 & _EVAL_368;
  assign _EVAL_74 = _EVAL_12 & _EVAL_369;
  assign _EVAL_111 = _EVAL_364 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_48 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_62 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_102 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_120 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_172 = _RAND_6[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_205 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_209 = _RAND_8[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_235 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_247 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_254 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_267 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {3{`RANDOM}};
  _EVAL_270 = _RAND_13[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_271 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_303 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_351 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_5) begin
    if (_EVAL_250) begin
      _EVAL_26 <= _EVAL;
    end
    if (_EVAL_178) begin
      _EVAL_35 <= _EVAL_18;
    end
    if (_EVAL_178) begin
      _EVAL_48 <= _EVAL_7;
    end
    if (_EVAL_2) begin
      _EVAL_62 <= 6'h0;
    end else begin
      if (_EVAL_244) begin
        if (_EVAL_135) begin
          if (_EVAL_354) begin
            _EVAL_62 <= _EVAL_90;
          end else begin
            _EVAL_62 <= 6'h0;
          end
        end else begin
          _EVAL_62 <= _EVAL_253;
        end
      end
    end
    if (_EVAL_2) begin
      _EVAL_102 <= 6'h0;
    end else begin
      if (_EVAL_237) begin
        if (_EVAL_219) begin
          if (_EVAL_163) begin
            _EVAL_102 <= _EVAL_218;
          end else begin
            _EVAL_102 <= 6'h0;
          end
        end else begin
          _EVAL_102 <= _EVAL_30;
        end
      end
    end
    if (_EVAL_178) begin
      _EVAL_120 <= _EVAL_16;
    end
    if (_EVAL_178) begin
      _EVAL_172 <= _EVAL_9;
    end
    if (_EVAL_178) begin
      _EVAL_205 <= _EVAL_11;
    end
    if (_EVAL_250) begin
      _EVAL_209 <= _EVAL_13;
    end
    if (_EVAL_2) begin
      _EVAL_235 <= 6'h0;
    end else begin
      if (_EVAL_244) begin
        if (_EVAL_292) begin
          if (_EVAL_354) begin
            _EVAL_235 <= _EVAL_90;
          end else begin
            _EVAL_235 <= 6'h0;
          end
        end else begin
          _EVAL_235 <= _EVAL_337;
        end
      end
    end
    if (_EVAL_2) begin
      _EVAL_247 <= 32'h0;
    end else begin
      if (_EVAL_370) begin
        _EVAL_247 <= 32'h0;
      end else begin
        _EVAL_247 <= _EVAL_146;
      end
    end
    if (_EVAL_250) begin
      _EVAL_254 <= _EVAL_17;
    end
    if (_EVAL_250) begin
      _EVAL_267 <= _EVAL_14;
    end
    if (_EVAL_2) begin
      _EVAL_270 <= 73'h0;
    end else begin
      _EVAL_270 <= _EVAL_262;
    end
    if (_EVAL_250) begin
      _EVAL_271 <= _EVAL_15;
    end
    if (_EVAL_2) begin
      _EVAL_303 <= 6'h0;
    end else begin
      if (_EVAL_237) begin
        if (_EVAL_307) begin
          if (_EVAL_163) begin
            _EVAL_303 <= _EVAL_218;
          end else begin
            _EVAL_303 <= 6'h0;
          end
        end else begin
          _EVAL_303 <= _EVAL_285;
        end
      end
    end
    if (_EVAL_250) begin
      _EVAL_351 <= _EVAL_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb54076)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3976e961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(834b78f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fac5c366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a936f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48671a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fa45eb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef10e62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d61cbfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a67546b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b76301b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4cf5055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c31ee64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588dbf31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472c9bff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20657607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c36915bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b34505b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb46fff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1488a66b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3c947f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4601cae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bda8bb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41bb422c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ede3b35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef2b85d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1705b6f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e39d222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b097bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(770f51eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4337fd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c6d055d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(522e3f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de65256c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61691de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13e497ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d979533)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc7a8141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de98c78a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_329) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcb46a47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f32acee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eba0fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7623faea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(921d29b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1014c15f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7958a3f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b71bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fad31d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f13222c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12017301)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5afd06ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a01f7a17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75e00e62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77ce0d47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69f220b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c73cc2b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c94b8ded)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(482c0d2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbfd156f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e823663b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86958323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9277fbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(753c1f62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74145526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0321c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee7f6063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9384970)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5ac6119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1306952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(549ee43e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a989c54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928fcba7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1feb6378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffcbbb45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eafd1aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82def109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96cc6616)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e34ca659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d1b43a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df624b50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36cfea1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(869d34cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eed0b641)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30d7db54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bb218fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8144a5eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_329) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57b9a694)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c12727a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(252fad29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75965c4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
