//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_228(
  input         _EVAL,
  input         _EVAL_0,
  input  [29:0] _EVAL_1,
  input         _EVAL_2,
  input  [1:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input  [29:0] _EVAL_18,
  input  [1:0]  _EVAL_19,
  input  [31:0] _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [1:0]  _EVAL_25,
  output        _EVAL_26,
  input  [31:0] _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input  [1:0]  _EVAL_35,
  input         _EVAL_36,
  input  [31:0] _EVAL_37,
  input  [1:0]  _EVAL_38,
  input  [31:0] _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input  [29:0] _EVAL_42,
  input  [29:0] _EVAL_43,
  input         _EVAL_44,
  input  [29:0] _EVAL_45,
  input         _EVAL_46,
  input  [29:0] _EVAL_47,
  input         _EVAL_48,
  input  [31:0] _EVAL_49,
  input         _EVAL_50,
  input  [1:0]  _EVAL_51,
  input         _EVAL_52,
  input  [29:0] _EVAL_53,
  input  [31:0] _EVAL_54,
  input         _EVAL_55,
  input  [1:0]  _EVAL_56,
  input  [29:0] _EVAL_57,
  input         _EVAL_58,
  input  [31:0] _EVAL_59
);
  wire [31:0] _EVAL_335;
  wire [31:0] _EVAL_83;
  wire [31:0] _EVAL_331;
  wire [31:0] _EVAL_360;
  wire [31:0] _EVAL_153;
  wire [31:0] _EVAL_357;
  wire [31:0] _EVAL_320;
  wire [31:0] _EVAL_263;
  wire [31:0] _EVAL_110;
  wire [31:0] _EVAL_220;
  wire  _EVAL_203;
  wire  _EVAL_288;
  wire  _EVAL_226;
  wire  _EVAL_142;
  wire  _EVAL_64;
  wire [31:0] _EVAL_240;
  wire  _EVAL_332;
  wire  _EVAL_116;
  wire  _EVAL_202;
  wire [31:0] _EVAL_123;
  wire [31:0] _EVAL_219;
  wire [31:0] _EVAL_307;
  wire [31:0] _EVAL_277;
  wire [31:0] _EVAL_70;
  wire [31:0] _EVAL_271;
  wire [31:0] _EVAL_124;
  wire  _EVAL_218;
  wire  _EVAL_156;
  wire [31:0] _EVAL_155;
  wire [31:0] _EVAL_102;
  wire [31:0] _EVAL_114;
  wire [31:0] _EVAL_160;
  wire  _EVAL_195;
  wire  _EVAL_77;
  wire  _EVAL_338;
  wire  _EVAL_213;
  wire  _EVAL_169;
  wire  _EVAL_79;
  wire  _EVAL_62;
  wire  _EVAL_306;
  wire  _EVAL_217;
  wire  _EVAL_249;
  wire [31:0] _EVAL_111;
  wire [31:0] _EVAL_252;
  wire [31:0] _EVAL_309;
  wire [31:0] _EVAL_211;
  wire [31:0] _EVAL_230;
  wire [31:0] _EVAL_129;
  wire [31:0] _EVAL_192;
  wire  _EVAL_112;
  wire  _EVAL_236;
  wire  _EVAL_88;
  wire  _EVAL_343;
  wire  _EVAL_280;
  wire  _EVAL_93;
  wire  _EVAL_237;
  wire  _EVAL_367;
  wire  _EVAL_242;
  wire  _EVAL_173;
  wire  _EVAL_245;
  wire [31:0] _EVAL_65;
  wire [31:0] _EVAL_336;
  wire [31:0] _EVAL_254;
  wire [31:0] _EVAL_316;
  wire [31:0] _EVAL_89;
  wire [31:0] _EVAL_63;
  wire [31:0] _EVAL_95;
  wire  _EVAL_136;
  wire  _EVAL_138;
  wire  _EVAL_72;
  wire  _EVAL_341;
  wire  _EVAL_91;
  wire  _EVAL_266;
  wire  _EVAL_180;
  wire  _EVAL_297;
  wire  _EVAL_175;
  wire [31:0] _EVAL_246;
  wire [31:0] _EVAL_229;
  wire [31:0] _EVAL_313;
  wire [31:0] _EVAL_283;
  wire [31:0] _EVAL_96;
  wire [31:0] _EVAL_141;
  wire [31:0] _EVAL_233;
  wire  _EVAL_128;
  wire  _EVAL_232;
  wire  _EVAL_120;
  wire  _EVAL_185;
  wire  _EVAL_162;
  wire  _EVAL_348;
  wire  _EVAL_311;
  wire  _EVAL_328;
  wire  _EVAL_74;
  wire  _EVAL_272;
  wire  _EVAL_140;
  wire  _EVAL_349;
  wire  _EVAL_339;
  wire  _EVAL_295;
  wire  _EVAL_256;
  wire  _EVAL_146;
  wire [31:0] _EVAL_204;
  wire [31:0] _EVAL_262;
  wire [31:0] _EVAL_290;
  wire  _EVAL_115;
  wire  _EVAL_355;
  wire [31:0] _EVAL_122;
  wire [31:0] _EVAL_81;
  wire [31:0] _EVAL_168;
  wire [31:0] _EVAL_84;
  wire  _EVAL_118;
  wire  _EVAL_131;
  wire  _EVAL_308;
  wire  _EVAL_67;
  wire  _EVAL_201;
  wire  _EVAL_69;
  wire [31:0] _EVAL_157;
  wire [31:0] _EVAL_261;
  wire  _EVAL_278;
  wire  _EVAL_76;
  wire  _EVAL_119;
  wire  _EVAL_353;
  wire  _EVAL_302;
  wire  _EVAL_98;
  wire [31:0] _EVAL_209;
  wire  _EVAL_148;
  wire  _EVAL_176;
  wire  _EVAL_193;
  wire  _EVAL_294;
  wire  _EVAL_337;
  wire  _EVAL_284;
  wire  _EVAL_258;
  wire  _EVAL_304;
  wire  _EVAL_370;
  wire  _EVAL_158;
  wire  _EVAL_315;
  wire  _EVAL_351;
  wire  _EVAL_342;
  wire  _EVAL_105;
  wire [31:0] _EVAL_224;
  wire [31:0] _EVAL_346;
  wire [31:0] _EVAL_137;
  wire  _EVAL_274;
  wire  _EVAL_188;
  wire  _EVAL_99;
  wire  _EVAL_178;
  wire  _EVAL_235;
  wire  _EVAL_340;
  wire  _EVAL_300;
  wire  _EVAL_196;
  wire  _EVAL_87;
  wire  _EVAL_212;
  assign _EVAL_335 = {_EVAL_45, 2'h0};
  assign _EVAL_83 = ~ _EVAL_335;
  assign _EVAL_331 = _EVAL_83 | 32'h3f;
  assign _EVAL_360 = ~ _EVAL_331;
  assign _EVAL_153 = _EVAL_10 ^ _EVAL_360;
  assign _EVAL_357 = {_EVAL_43, 2'h0};
  assign _EVAL_320 = ~ _EVAL_357;
  assign _EVAL_263 = _EVAL_320 | 32'h3f;
  assign _EVAL_110 = ~ _EVAL_263;
  assign _EVAL_220 = _EVAL_10 ^ _EVAL_110;
  assign _EVAL_203 = _EVAL_38 > 2'h1;
  assign _EVAL_288 = _EVAL_32 == 1'h0;
  assign _EVAL_226 = _EVAL_203 & _EVAL_288;
  assign _EVAL_142 = _EVAL_44 | _EVAL_226;
  assign _EVAL_64 = _EVAL_36 == 1'h0;
  assign _EVAL_240 = ~ _EVAL_20;
  assign _EVAL_332 = _EVAL_24 == 1'h0;
  assign _EVAL_116 = _EVAL_203 & _EVAL_332;
  assign _EVAL_202 = _EVAL_3[1];
  assign _EVAL_123 = {_EVAL_57, 2'h0};
  assign _EVAL_219 = ~ _EVAL_123;
  assign _EVAL_307 = _EVAL_219 | 32'h3f;
  assign _EVAL_277 = ~ _EVAL_307;
  assign _EVAL_70 = _EVAL_10 ^ _EVAL_277;
  assign _EVAL_271 = ~ _EVAL_7;
  assign _EVAL_124 = _EVAL_70 & _EVAL_271;
  assign _EVAL_218 = _EVAL_124 == 32'h0;
  assign _EVAL_156 = _EVAL_3[0];
  assign _EVAL_155 = {_EVAL_1, 2'h0};
  assign _EVAL_102 = ~ _EVAL_155;
  assign _EVAL_114 = _EVAL_102 | 32'h3f;
  assign _EVAL_160 = ~ _EVAL_114;
  assign _EVAL_195 = _EVAL_10 < _EVAL_160;
  assign _EVAL_77 = _EVAL_195 == 1'h0;
  assign _EVAL_338 = _EVAL_10 < _EVAL_277;
  assign _EVAL_213 = _EVAL_77 & _EVAL_338;
  assign _EVAL_169 = _EVAL_156 & _EVAL_213;
  assign _EVAL_79 = _EVAL_202 ? _EVAL_218 : _EVAL_169;
  assign _EVAL_62 = _EVAL_5 == 1'h0;
  assign _EVAL_306 = _EVAL_203 & _EVAL_62;
  assign _EVAL_217 = _EVAL_6 | _EVAL_306;
  assign _EVAL_249 = _EVAL_25[1];
  assign _EVAL_111 = {_EVAL_18, 2'h0};
  assign _EVAL_252 = ~ _EVAL_111;
  assign _EVAL_309 = _EVAL_252 | 32'h3f;
  assign _EVAL_211 = ~ _EVAL_309;
  assign _EVAL_230 = _EVAL_10 ^ _EVAL_211;
  assign _EVAL_129 = ~ _EVAL_27;
  assign _EVAL_192 = _EVAL_230 & _EVAL_129;
  assign _EVAL_112 = _EVAL_192 == 32'h0;
  assign _EVAL_236 = _EVAL_25[0];
  assign _EVAL_88 = _EVAL_338 == 1'h0;
  assign _EVAL_343 = _EVAL_10 < _EVAL_211;
  assign _EVAL_280 = _EVAL_88 & _EVAL_343;
  assign _EVAL_93 = _EVAL_236 & _EVAL_280;
  assign _EVAL_237 = _EVAL_249 ? _EVAL_112 : _EVAL_93;
  assign _EVAL_367 = _EVAL_48 == 1'h0;
  assign _EVAL_242 = _EVAL_203 & _EVAL_367;
  assign _EVAL_173 = _EVAL_14 | _EVAL_242;
  assign _EVAL_245 = _EVAL_19[1];
  assign _EVAL_65 = {_EVAL_53, 2'h0};
  assign _EVAL_336 = ~ _EVAL_65;
  assign _EVAL_254 = _EVAL_336 | 32'h3f;
  assign _EVAL_316 = ~ _EVAL_254;
  assign _EVAL_89 = _EVAL_10 ^ _EVAL_316;
  assign _EVAL_63 = ~ _EVAL_39;
  assign _EVAL_95 = _EVAL_89 & _EVAL_63;
  assign _EVAL_136 = _EVAL_95 == 32'h0;
  assign _EVAL_138 = _EVAL_19[0];
  assign _EVAL_72 = _EVAL_343 == 1'h0;
  assign _EVAL_341 = _EVAL_10 < _EVAL_316;
  assign _EVAL_91 = _EVAL_72 & _EVAL_341;
  assign _EVAL_266 = _EVAL_138 & _EVAL_91;
  assign _EVAL_180 = _EVAL_245 ? _EVAL_136 : _EVAL_266;
  assign _EVAL_297 = _EVAL | _EVAL_116;
  assign _EVAL_175 = _EVAL_8[1];
  assign _EVAL_246 = {_EVAL_42, 2'h0};
  assign _EVAL_229 = ~ _EVAL_246;
  assign _EVAL_313 = _EVAL_229 | 32'h3f;
  assign _EVAL_283 = ~ _EVAL_313;
  assign _EVAL_96 = _EVAL_10 ^ _EVAL_283;
  assign _EVAL_141 = ~ _EVAL_59;
  assign _EVAL_233 = _EVAL_96 & _EVAL_141;
  assign _EVAL_128 = _EVAL_233 == 32'h0;
  assign _EVAL_232 = _EVAL_8[0];
  assign _EVAL_120 = _EVAL_341 == 1'h0;
  assign _EVAL_185 = _EVAL_10 < _EVAL_283;
  assign _EVAL_162 = _EVAL_120 & _EVAL_185;
  assign _EVAL_348 = _EVAL_232 & _EVAL_162;
  assign _EVAL_311 = _EVAL_175 ? _EVAL_128 : _EVAL_348;
  assign _EVAL_328 = _EVAL_29 == 1'h0;
  assign _EVAL_74 = _EVAL_203 & _EVAL_328;
  assign _EVAL_272 = _EVAL_52 | _EVAL_74;
  assign _EVAL_140 = _EVAL_311 ? _EVAL_272 : _EVAL_203;
  assign _EVAL_349 = _EVAL_180 ? _EVAL_297 : _EVAL_140;
  assign _EVAL_339 = _EVAL_237 ? _EVAL_173 : _EVAL_349;
  assign _EVAL_295 = _EVAL_79 ? _EVAL_217 : _EVAL_339;
  assign _EVAL_256 = _EVAL_34 == 1'h0;
  assign _EVAL_146 = _EVAL_51[1];
  assign _EVAL_204 = _EVAL_10 ^ _EVAL_160;
  assign _EVAL_262 = ~ _EVAL_54;
  assign _EVAL_290 = _EVAL_204 & _EVAL_262;
  assign _EVAL_115 = _EVAL_290 == 32'h0;
  assign _EVAL_355 = _EVAL_51[0];
  assign _EVAL_122 = {_EVAL_47, 2'h0};
  assign _EVAL_81 = ~ _EVAL_122;
  assign _EVAL_168 = _EVAL_81 | 32'h3f;
  assign _EVAL_84 = ~ _EVAL_168;
  assign _EVAL_118 = _EVAL_10 < _EVAL_84;
  assign _EVAL_131 = _EVAL_118 == 1'h0;
  assign _EVAL_308 = _EVAL_131 & _EVAL_195;
  assign _EVAL_67 = _EVAL_355 & _EVAL_308;
  assign _EVAL_201 = _EVAL_146 ? _EVAL_115 : _EVAL_67;
  assign _EVAL_69 = _EVAL_17[1];
  assign _EVAL_157 = ~ _EVAL_37;
  assign _EVAL_261 = _EVAL_220 & _EVAL_157;
  assign _EVAL_278 = _EVAL_261 == 32'h0;
  assign _EVAL_76 = _EVAL_17[0];
  assign _EVAL_119 = _EVAL_10 < _EVAL_110;
  assign _EVAL_353 = _EVAL_76 & _EVAL_119;
  assign _EVAL_302 = _EVAL_69 ? _EVAL_278 : _EVAL_353;
  assign _EVAL_98 = _EVAL_35[1];
  assign _EVAL_209 = _EVAL_153 & _EVAL_240;
  assign _EVAL_148 = _EVAL_209 == 32'h0;
  assign _EVAL_176 = _EVAL_35[0];
  assign _EVAL_193 = _EVAL_119 == 1'h0;
  assign _EVAL_294 = _EVAL_10 < _EVAL_360;
  assign _EVAL_337 = _EVAL_193 & _EVAL_294;
  assign _EVAL_284 = _EVAL_176 & _EVAL_337;
  assign _EVAL_258 = _EVAL_98 ? _EVAL_148 : _EVAL_284;
  assign _EVAL_304 = _EVAL_203 & _EVAL_64;
  assign _EVAL_370 = _EVAL_294 == 1'h0;
  assign _EVAL_158 = _EVAL_370 & _EVAL_118;
  assign _EVAL_315 = _EVAL_203 & _EVAL_256;
  assign _EVAL_351 = _EVAL_13 | _EVAL_315;
  assign _EVAL_342 = _EVAL_31 == 1'h0;
  assign _EVAL_105 = _EVAL_56[1];
  assign _EVAL_224 = _EVAL_10 ^ _EVAL_84;
  assign _EVAL_346 = ~ _EVAL_49;
  assign _EVAL_137 = _EVAL_224 & _EVAL_346;
  assign _EVAL_274 = _EVAL_137 == 32'h0;
  assign _EVAL_188 = _EVAL_56[0];
  assign _EVAL_99 = _EVAL_188 & _EVAL_158;
  assign _EVAL_178 = _EVAL_105 ? _EVAL_274 : _EVAL_99;
  assign _EVAL_235 = _EVAL_203 & _EVAL_342;
  assign _EVAL_340 = _EVAL_30 | _EVAL_235;
  assign _EVAL_300 = _EVAL_201 ? _EVAL_351 : _EVAL_295;
  assign _EVAL_196 = _EVAL_178 ? _EVAL_340 : _EVAL_300;
  assign _EVAL_87 = _EVAL_258 ? _EVAL_142 : _EVAL_196;
  assign _EVAL_212 = _EVAL_2 | _EVAL_304;
  assign _EVAL_26 = _EVAL_302 ? _EVAL_212 : _EVAL_87;
endmodule
