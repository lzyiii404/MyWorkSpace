//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_260_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [7:0]  _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [24:0] _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_33;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_37;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_58;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_69;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_71;
  reg [31:0] _RAND_4;
  reg [24:0] _EVAL_106;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_109;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_116;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_156;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_163;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_165;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_181;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_213;
  reg [31:0] _RAND_12;
  reg [7:0] _EVAL_247;
  reg [31:0] _RAND_13;
  wire [1:0] _EVAL_199;
  wire [3:0] _EVAL_138;
  wire [2:0] _EVAL_151;
  wire [2:0] _EVAL_130;
  wire  _EVAL_178;
  wire  _EVAL_230;
  wire  _EVAL_205;
  wire  _EVAL_26;
  wire  _EVAL_41;
  wire  _EVAL_224;
  wire  _EVAL_206;
  wire  _EVAL_44;
  wire  _EVAL_15;
  wire  _EVAL_52;
  wire  _EVAL_134;
  wire  _EVAL_120;
  wire  _EVAL_280;
  wire [7:0] _EVAL_257;
  wire  _EVAL_282;
  wire  _EVAL_168;
  wire  _EVAL_85;
  wire  _EVAL_20;
  wire  _EVAL_131;
  wire  _EVAL_43;
  wire  _EVAL_140;
  wire  _EVAL_234;
  wire [7:0] _EVAL_83;
  wire  _EVAL_215;
  wire  _EVAL_251;
  wire  _EVAL_261;
  wire  _EVAL_28;
  wire  _EVAL_160;
  wire  _EVAL_207;
  wire  _EVAL_158;
  wire  _EVAL_135;
  wire  _EVAL_185;
  wire  _EVAL_72;
  wire  _EVAL_269;
  wire  _EVAL_243;
  wire  _EVAL_278;
  wire  _EVAL_124;
  wire  _EVAL_203;
  wire  _EVAL_148;
  wire [24:0] _EVAL_49;
  wire [25:0] _EVAL_180;
  wire [25:0] _EVAL_173;
  wire [2:0] _EVAL_164;
  wire  _EVAL_240;
  wire  _EVAL_286;
  wire  _EVAL_192;
  wire  _EVAL_136;
  wire  _EVAL_94;
  wire  _EVAL_70;
  wire [7:0] _EVAL_96;
  wire [7:0] _EVAL_118;
  wire  _EVAL_190;
  wire  _EVAL_157;
  wire  _EVAL_54;
  wire [7:0] _EVAL_144;
  wire [7:0] _EVAL_127;
  wire  _EVAL_108;
  wire  _EVAL_183;
  wire  _EVAL_122;
  wire  _EVAL_60;
  wire  _EVAL_211;
  wire  _EVAL_279;
  wire  _EVAL_283;
  wire  _EVAL_210;
  wire  _EVAL_61;
  wire  _EVAL_81;
  wire  _EVAL_162;
  wire [25:0] _EVAL_209;
  wire  _EVAL_80;
  wire  _EVAL_27;
  wire  _EVAL_246;
  wire [7:0] _EVAL_272;
  wire [12:0] _EVAL_21;
  wire  _EVAL_253;
  wire  _EVAL_197;
  wire  _EVAL_114;
  wire [31:0] _EVAL_51;
  wire  _EVAL_182;
  wire  _EVAL_175;
  wire  _EVAL_59;
  wire  _EVAL_267;
  wire [12:0] _EVAL_95;
  wire [5:0] _EVAL_77;
  wire [5:0] _EVAL_98;
  wire [2:0] _EVAL_84;
  wire [2:0] _EVAL_125;
  wire [7:0] _EVAL_256;
  wire  _EVAL_285;
  wire  _EVAL_64;
  wire  _EVAL_75;
  wire  _EVAL_275;
  wire  _EVAL_237;
  wire  _EVAL_172;
  wire  _EVAL_62;
  wire [7:0] _EVAL_260;
  wire  _EVAL_179;
  wire  _EVAL_232;
  wire [24:0] _EVAL_126;
  wire  _EVAL_55;
  wire  _EVAL_145;
  wire  _EVAL_219;
  wire  _EVAL_19;
  wire  _EVAL_34;
  wire  _EVAL_107;
  wire  _EVAL_113;
  wire  _EVAL_88;
  wire  _EVAL_29;
  wire  _EVAL_119;
  wire  _EVAL_233;
  wire  _EVAL_265;
  wire  _EVAL_63;
  wire  _EVAL_66;
  wire  _EVAL_212;
  wire  _EVAL_57;
  wire  _EVAL_137;
  wire  _EVAL_155;
  wire  _EVAL_23;
  wire  _EVAL_274;
  wire  _EVAL_228;
  wire  _EVAL_167;
  wire  _EVAL_218;
  wire  _EVAL_214;
  wire  _EVAL_147;
  wire  _EVAL_186;
  wire  _EVAL_276;
  wire  _EVAL_39;
  wire  _EVAL_146;
  wire  _EVAL_188;
  wire  _EVAL_266;
  wire  _EVAL_252;
  wire  _EVAL_201;
  wire  _EVAL_45;
  wire  _EVAL_254;
  wire  _EVAL_242;
  wire  _EVAL_101;
  wire  _EVAL_184;
  wire  _EVAL_195;
  wire  _EVAL_198;
  wire  _EVAL_226;
  wire  _EVAL_100;
  wire  _EVAL_222;
  wire  _EVAL_91;
  wire  _EVAL_17;
  wire  _EVAL_139;
  wire  _EVAL_112;
  wire  _EVAL_46;
  wire  _EVAL_86;
  wire  _EVAL_30;
  wire  _EVAL_259;
  wire  _EVAL_166;
  wire  _EVAL_110;
  wire  _EVAL_191;
  wire  _EVAL_132;
  wire  _EVAL_225;
  wire  _EVAL_273;
  wire  _EVAL_74;
  wire  _EVAL_90;
  wire  _EVAL_18;
  wire [7:0] _EVAL_238;
  wire [7:0] _EVAL_78;
  wire  _EVAL_149;
  wire  _EVAL_117;
  wire  _EVAL_16;
  wire  _EVAL_53;
  wire  _EVAL_142;
  wire  _EVAL_152;
  wire  _EVAL_171;
  wire  _EVAL_38;
  wire  _EVAL_236;
  wire  _EVAL_35;
  wire  _EVAL_99;
  wire  _EVAL_111;
  wire  _EVAL_202;
  wire  _EVAL_32;
  wire  _EVAL_229;
  wire  _EVAL_277;
  wire  _EVAL_200;
  wire  _EVAL_262;
  wire  _EVAL_40;
  wire [5:0] _EVAL_103;
  wire [5:0] _EVAL_93;
  wire [2:0] _EVAL_216;
  wire [2:0] _EVAL_241;
  wire  _EVAL_161;
  wire [2:0] _EVAL_102;
  wire [7:0] _EVAL_56;
  wire  _EVAL_174;
  wire  _EVAL_133;
  wire  _EVAL_47;
  wire  _EVAL_141;
  wire [24:0] _EVAL_221;
  wire  _EVAL_50;
  wire  _EVAL_87;
  wire  _EVAL_177;
  wire  _EVAL_268;
  wire  _EVAL_235;
  wire  _EVAL_244;
  wire  _EVAL_248;
  wire  _EVAL_270;
  wire  _EVAL_153;
  wire  _EVAL_223;
  wire  _EVAL_193;
  wire  _EVAL_25;
  wire  _EVAL_67;
  wire  _EVAL_284;
  wire  _EVAL_258;
  wire  _EVAL_264;
  wire  _EVAL_22;
  wire  _EVAL_24;
  wire  _EVAL_105;
  wire  _EVAL_143;
  wire  _EVAL_245;
  wire  _EVAL_208;
  wire [7:0] _EVAL_79;
  wire [7:0] _EVAL_169;
  wire  _EVAL_121;
  wire  _EVAL_176;
  wire  _EVAL_271;
  wire  _EVAL_68;
  wire  _EVAL_263;
  wire  _EVAL_42;
  wire  _EVAL_97;
  wire  _EVAL_250;
  wire  _EVAL_154;
  wire  _EVAL_159;
  wire  _EVAL_255;
  wire  _EVAL_115;
  wire  _EVAL_65;
  wire  _EVAL_281;
  wire  _EVAL_150;
  wire  _EVAL_31;
  wire  _EVAL_76;
  wire  _EVAL_239;
  wire  _EVAL_189;
  wire  _EVAL_48;
  wire  _EVAL_36;
  wire  _EVAL_220;
  wire  _EVAL_204;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_199 = _EVAL_4[1:0];
  assign _EVAL_138 = 4'h1 << _EVAL_199;
  assign _EVAL_151 = _EVAL_138[2:0];
  assign _EVAL_130 = _EVAL_151 | 3'h1;
  assign _EVAL_178 = _EVAL_130[0];
  assign _EVAL_230 = _EVAL_9[2];
  assign _EVAL_205 = _EVAL_9[1];
  assign _EVAL_26 = _EVAL_205 == 1'h0;
  assign _EVAL_41 = _EVAL_230 & _EVAL_26;
  assign _EVAL_224 = _EVAL_9[0];
  assign _EVAL_206 = _EVAL_224 == 1'h0;
  assign _EVAL_44 = _EVAL_41 & _EVAL_206;
  assign _EVAL_15 = _EVAL_178 & _EVAL_44;
  assign _EVAL_52 = _EVAL_11 <= 3'h2;
  assign _EVAL_134 = _EVAL_52 | _EVAL_1;
  assign _EVAL_120 = _EVAL_8 == 3'h1;
  assign _EVAL_280 = _EVAL_12 == _EVAL_116;
  assign _EVAL_257 = ~ _EVAL_6;
  assign _EVAL_282 = _EVAL_247 != 8'h0;
  assign _EVAL_168 = _EVAL_282 == 1'h0;
  assign _EVAL_85 = plusarg_reader_out == 32'h0;
  assign _EVAL_20 = _EVAL_168 | _EVAL_85;
  assign _EVAL_131 = _EVAL_5 & _EVAL_2;
  assign _EVAL_43 = _EVAL_33 == 3'h0;
  assign _EVAL_140 = _EVAL_131 & _EVAL_43;
  assign _EVAL_234 = _EVAL_181 < plusarg_reader_out;
  assign _EVAL_83 = _EVAL_247 >> _EVAL_12;
  assign _EVAL_215 = _EVAL_4 >= 3'h3;
  assign _EVAL_251 = _EVAL_130[2];
  assign _EVAL_261 = _EVAL_251 & _EVAL_230;
  assign _EVAL_28 = _EVAL_215 | _EVAL_261;
  assign _EVAL_160 = _EVAL_130[1];
  assign _EVAL_207 = _EVAL_230 & _EVAL_205;
  assign _EVAL_158 = _EVAL_160 & _EVAL_207;
  assign _EVAL_135 = _EVAL_28 | _EVAL_158;
  assign _EVAL_185 = 3'h1 <= _EVAL_0;
  assign _EVAL_72 = _EVAL_8 == 3'h5;
  assign _EVAL_269 = _EVAL_14 & _EVAL_72;
  assign _EVAL_243 = _EVAL_10 == 3'h5;
  assign _EVAL_278 = _EVAL_83[0];
  assign _EVAL_124 = _EVAL_278 == 1'h0;
  assign _EVAL_203 = _EVAL_124 | _EVAL_1;
  assign _EVAL_148 = _EVAL_203 == 1'h0;
  assign _EVAL_49 = _EVAL_9 ^ 25'h1900000;
  assign _EVAL_180 = {1'b0,$signed(_EVAL_49)};
  assign _EVAL_173 = $signed(_EVAL_180) & $signed(-26'sh2000);
  assign _EVAL_164 = _EVAL_58 - 3'h1;
  assign _EVAL_240 = _EVAL_207 & _EVAL_206;
  assign _EVAL_286 = _EVAL_178 & _EVAL_240;
  assign _EVAL_192 = _EVAL_135 | _EVAL_286;
  assign _EVAL_136 = _EVAL_3 & _EVAL_14;
  assign _EVAL_94 = _EVAL_71 == 3'h0;
  assign _EVAL_70 = _EVAL_136 & _EVAL_94;
  assign _EVAL_96 = 8'h1 << _EVAL_12;
  assign _EVAL_118 = _EVAL_70 ? _EVAL_96 : 8'h0;
  assign _EVAL_190 = _EVAL_10 == 3'h6;
  assign _EVAL_157 = _EVAL_190 == 1'h0;
  assign _EVAL_54 = _EVAL_140 & _EVAL_157;
  assign _EVAL_144 = 8'h1 << _EVAL_0;
  assign _EVAL_127 = _EVAL_54 ? _EVAL_144 : 8'h0;
  assign _EVAL_108 = _EVAL_118 != _EVAL_127;
  assign _EVAL_183 = _EVAL_9 == _EVAL_106;
  assign _EVAL_122 = _EVAL_183 | _EVAL_1;
  assign _EVAL_60 = _EVAL_230 == 1'h0;
  assign _EVAL_211 = _EVAL_60 & _EVAL_26;
  assign _EVAL_279 = _EVAL_211 & _EVAL_206;
  assign _EVAL_283 = _EVAL_178 & _EVAL_279;
  assign _EVAL_210 = _EVAL_7 == 1'h0;
  assign _EVAL_61 = _EVAL_210 | _EVAL_1;
  assign _EVAL_81 = _EVAL_61 == 1'h0;
  assign _EVAL_162 = _EVAL_4 <= 3'h6;
  assign _EVAL_209 = $signed(_EVAL_173);
  assign _EVAL_80 = _EVAL_12 == 3'h0;
  assign _EVAL_27 = 3'h6 == _EVAL_4;
  assign _EVAL_246 = _EVAL_80 ? _EVAL_27 : 1'h0;
  assign _EVAL_272 = _EVAL_118 | _EVAL_247;
  assign _EVAL_21 = 13'h3f << _EVAL_13;
  assign _EVAL_253 = _EVAL_10 == _EVAL_165;
  assign _EVAL_197 = _EVAL_253 | _EVAL_1;
  assign _EVAL_114 = _EVAL_136 | _EVAL_131;
  assign _EVAL_51 = _EVAL_181 + 32'h1;
  assign _EVAL_182 = _EVAL_20 | _EVAL_234;
  assign _EVAL_175 = _EVAL_182 | _EVAL_1;
  assign _EVAL_59 = _EVAL_8[2];
  assign _EVAL_267 = _EVAL_59 == 1'h0;
  assign _EVAL_95 = 13'h3f << _EVAL_4;
  assign _EVAL_77 = _EVAL_95[5:0];
  assign _EVAL_98 = ~ _EVAL_77;
  assign _EVAL_84 = _EVAL_98[5:3];
  assign _EVAL_125 = _EVAL_71 - 3'h1;
  assign _EVAL_256 = _EVAL_272 >> _EVAL_0;
  assign _EVAL_285 = _EVAL_118 != 8'h0;
  assign _EVAL_64 = _EVAL_285 == 1'h0;
  assign _EVAL_75 = _EVAL_108 | _EVAL_64;
  assign _EVAL_275 = _EVAL_41 & _EVAL_224;
  assign _EVAL_237 = _EVAL_178 & _EVAL_275;
  assign _EVAL_172 = _EVAL_251 & _EVAL_60;
  assign _EVAL_62 = _EVAL_215 | _EVAL_172;
  assign _EVAL_260 = ~ _EVAL_127;
  assign _EVAL_179 = _EVAL_160 & _EVAL_41;
  assign _EVAL_232 = _EVAL_280 | _EVAL_1;
  assign _EVAL_126 = {{19'd0}, _EVAL_98};
  assign _EVAL_55 = _EVAL_0 == 3'h0;
  assign _EVAL_145 = _EVAL_13 == _EVAL_163;
  assign _EVAL_219 = _EVAL_145 | _EVAL_1;
  assign _EVAL_19 = _EVAL_219 == 1'h0;
  assign _EVAL_34 = _EVAL_60 & _EVAL_205;
  assign _EVAL_107 = _EVAL_160 & _EVAL_34;
  assign _EVAL_113 = _EVAL_8 == 3'h4;
  assign _EVAL_88 = _EVAL_11 != 3'h0;
  assign _EVAL_29 = _EVAL_88 | _EVAL_1;
  assign _EVAL_119 = _EVAL_4 <= 3'h2;
  assign _EVAL_233 = $signed(_EVAL_209) == $signed(26'sh0);
  assign _EVAL_265 = _EVAL_119 & _EVAL_233;
  assign _EVAL_63 = _EVAL_11 == _EVAL_109;
  assign _EVAL_66 = _EVAL_63 | _EVAL_1;
  assign _EVAL_212 = _EVAL_1 == 1'h0;
  assign _EVAL_57 = _EVAL_34 & _EVAL_206;
  assign _EVAL_137 = _EVAL_69 == 3'h0;
  assign _EVAL_155 = _EVAL_137 == 1'h0;
  assign _EVAL_23 = _EVAL_4 == _EVAL_156;
  assign _EVAL_274 = _EVAL_23 | _EVAL_1;
  assign _EVAL_228 = _EVAL_274 == 1'h0;
  assign _EVAL_167 = _EVAL_14 & _EVAL_113;
  assign _EVAL_218 = _EVAL_11 <= 3'h4;
  assign _EVAL_214 = _EVAL_58 == 3'h0;
  assign _EVAL_147 = _EVAL_256[0];
  assign _EVAL_186 = _EVAL_147 | _EVAL_1;
  assign _EVAL_276 = _EVAL_186 == 1'h0;
  assign _EVAL_39 = _EVAL_134 == 1'h0;
  assign _EVAL_146 = _EVAL_28 | _EVAL_179;
  assign _EVAL_188 = _EVAL_8 == 3'h2;
  assign _EVAL_266 = _EVAL_14 & _EVAL_188;
  assign _EVAL_252 = _EVAL_75 | _EVAL_1;
  assign _EVAL_201 = _EVAL_252 == 1'h0;
  assign _EVAL_45 = _EVAL_29 == 1'h0;
  assign _EVAL_254 = _EVAL_131 & _EVAL_137;
  assign _EVAL_242 = _EVAL_207 & _EVAL_224;
  assign _EVAL_101 = _EVAL_178 & _EVAL_242;
  assign _EVAL_184 = _EVAL_246 | _EVAL_1;
  assign _EVAL_195 = _EVAL_184 == 1'h0;
  assign _EVAL_198 = _EVAL_175 == 1'h0;
  assign _EVAL_226 = _EVAL_13 >= 3'h3;
  assign _EVAL_100 = _EVAL_226 | _EVAL_1;
  assign _EVAL_222 = _EVAL_160 & _EVAL_211;
  assign _EVAL_91 = _EVAL_62 | _EVAL_222;
  assign _EVAL_17 = _EVAL_91 | _EVAL_283;
  assign _EVAL_139 = _EVAL_10 <= 3'h6;
  assign _EVAL_112 = _EVAL_139 | _EVAL_1;
  assign _EVAL_46 = _EVAL_112 == 1'h0;
  assign _EVAL_86 = _EVAL_135 | _EVAL_101;
  assign _EVAL_30 = _EVAL_146 | _EVAL_237;
  assign _EVAL_259 = _EVAL_146 | _EVAL_15;
  assign _EVAL_166 = _EVAL_62 | _EVAL_107;
  assign _EVAL_110 = _EVAL_34 & _EVAL_224;
  assign _EVAL_191 = _EVAL_178 & _EVAL_110;
  assign _EVAL_132 = _EVAL_166 | _EVAL_191;
  assign _EVAL_225 = _EVAL_178 & _EVAL_57;
  assign _EVAL_273 = _EVAL_166 | _EVAL_225;
  assign _EVAL_74 = _EVAL_211 & _EVAL_224;
  assign _EVAL_90 = _EVAL_178 & _EVAL_74;
  assign _EVAL_18 = _EVAL_91 | _EVAL_90;
  assign _EVAL_238 = {_EVAL_86,_EVAL_192,_EVAL_30,_EVAL_259,_EVAL_132,_EVAL_273,_EVAL_18,_EVAL_17};
  assign _EVAL_78 = ~ _EVAL_238;
  assign _EVAL_149 = _EVAL_6 == _EVAL_238;
  assign _EVAL_117 = _EVAL_149 | _EVAL_1;
  assign _EVAL_16 = 3'h1 <= _EVAL_12;
  assign _EVAL_53 = _EVAL_80 | _EVAL_16;
  assign _EVAL_142 = _EVAL_8 == 3'h7;
  assign _EVAL_152 = _EVAL_14 & _EVAL_142;
  assign _EVAL_171 = _EVAL_2 & _EVAL_190;
  assign _EVAL_38 = _EVAL_257 == 8'h0;
  assign _EVAL_236 = _EVAL_38 | _EVAL_1;
  assign _EVAL_35 = _EVAL_236 == 1'h0;
  assign _EVAL_99 = _EVAL_53 | _EVAL_1;
  assign _EVAL_111 = _EVAL_99 == 1'h0;
  assign _EVAL_202 = _EVAL_10 == 3'h2;
  assign _EVAL_32 = _EVAL_2 & _EVAL_202;
  assign _EVAL_229 = _EVAL_10 == 3'h4;
  assign _EVAL_277 = _EVAL_55 | _EVAL_185;
  assign _EVAL_200 = _EVAL_277 | _EVAL_1;
  assign _EVAL_262 = _EVAL_200 == 1'h0;
  assign _EVAL_40 = _EVAL_10[0];
  assign _EVAL_103 = _EVAL_21[5:0];
  assign _EVAL_93 = ~ _EVAL_103;
  assign _EVAL_216 = _EVAL_93[5:3];
  assign _EVAL_241 = _EVAL_69 - 3'h1;
  assign _EVAL_161 = _EVAL_232 == 1'h0;
  assign _EVAL_102 = _EVAL_33 - 3'h1;
  assign _EVAL_56 = _EVAL_6 & _EVAL_78;
  assign _EVAL_174 = _EVAL_56 == 8'h0;
  assign _EVAL_133 = _EVAL_2 & _EVAL_243;
  assign _EVAL_47 = _EVAL_0 == _EVAL_213;
  assign _EVAL_141 = _EVAL_2 & _EVAL_155;
  assign _EVAL_221 = _EVAL_9 & _EVAL_126;
  assign _EVAL_50 = _EVAL_221 == 25'h0;
  assign _EVAL_87 = _EVAL_50 | _EVAL_1;
  assign _EVAL_177 = _EVAL_87 == 1'h0;
  assign _EVAL_268 = _EVAL_10 == 3'h1;
  assign _EVAL_235 = _EVAL_2 & _EVAL_268;
  assign _EVAL_244 = _EVAL_11 == 3'h0;
  assign _EVAL_248 = _EVAL_244 | _EVAL_1;
  assign _EVAL_270 = _EVAL_66 == 1'h0;
  assign _EVAL_153 = _EVAL_100 == 1'h0;
  assign _EVAL_223 = _EVAL_2 & _EVAL_229;
  assign _EVAL_193 = _EVAL_214 == 1'h0;
  assign _EVAL_25 = _EVAL_162 & _EVAL_233;
  assign _EVAL_67 = _EVAL_25 | _EVAL_1;
  assign _EVAL_284 = _EVAL_67 == 1'h0;
  assign _EVAL_258 = _EVAL_8 == 3'h0;
  assign _EVAL_264 = _EVAL_14 & _EVAL_120;
  assign _EVAL_22 = _EVAL_136 & _EVAL_214;
  assign _EVAL_24 = _EVAL_8 == 3'h3;
  assign _EVAL_105 = _EVAL_248 == 1'h0;
  assign _EVAL_143 = _EVAL_47 | _EVAL_1;
  assign _EVAL_245 = _EVAL_143 == 1'h0;
  assign _EVAL_208 = _EVAL_218 | _EVAL_1;
  assign _EVAL_79 = _EVAL_247 | _EVAL_118;
  assign _EVAL_169 = _EVAL_79 & _EVAL_260;
  assign _EVAL_121 = _EVAL_208 == 1'h0;
  assign _EVAL_176 = _EVAL_14 & _EVAL_193;
  assign _EVAL_271 = _EVAL_11 <= 3'h3;
  assign _EVAL_68 = _EVAL_117 == 1'h0;
  assign _EVAL_263 = _EVAL_265 | _EVAL_1;
  assign _EVAL_42 = _EVAL_263 == 1'h0;
  assign _EVAL_97 = _EVAL_10 == 3'h0;
  assign _EVAL_250 = _EVAL_2 & _EVAL_97;
  assign _EVAL_154 = _EVAL_8 == _EVAL_37;
  assign _EVAL_159 = _EVAL_215 | _EVAL_1;
  assign _EVAL_255 = _EVAL_159 == 1'h0;
  assign _EVAL_115 = _EVAL_197 == 1'h0;
  assign _EVAL_65 = _EVAL_8 == 3'h6;
  assign _EVAL_281 = _EVAL_271 | _EVAL_1;
  assign _EVAL_150 = _EVAL_154 | _EVAL_1;
  assign _EVAL_31 = _EVAL_281 == 1'h0;
  assign _EVAL_76 = _EVAL_174 | _EVAL_1;
  assign _EVAL_239 = _EVAL_76 == 1'h0;
  assign _EVAL_189 = _EVAL_122 == 1'h0;
  assign _EVAL_48 = _EVAL_14 & _EVAL_65;
  assign _EVAL_36 = _EVAL_14 & _EVAL_24;
  assign _EVAL_220 = _EVAL_14 & _EVAL_258;
  assign _EVAL_204 = _EVAL_150 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_33 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_37 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_58 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_69 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_71 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_106 = _RAND_5[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_109 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_116 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_156 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_163 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_165 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_181 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_213 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_247 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_1) begin
      _EVAL_33 <= 3'h0;
    end else begin
      if (_EVAL_131) begin
        if (_EVAL_43) begin
          if (_EVAL_40) begin
            _EVAL_33 <= _EVAL_216;
          end else begin
            _EVAL_33 <= 3'h0;
          end
        end else begin
          _EVAL_33 <= _EVAL_102;
        end
      end
    end
    if (_EVAL_22) begin
      _EVAL_37 <= _EVAL_8;
    end
    if (_EVAL_1) begin
      _EVAL_58 <= 3'h0;
    end else begin
      if (_EVAL_136) begin
        if (_EVAL_214) begin
          if (_EVAL_267) begin
            _EVAL_58 <= _EVAL_84;
          end else begin
            _EVAL_58 <= 3'h0;
          end
        end else begin
          _EVAL_58 <= _EVAL_164;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_69 <= 3'h0;
    end else begin
      if (_EVAL_131) begin
        if (_EVAL_137) begin
          if (_EVAL_40) begin
            _EVAL_69 <= _EVAL_216;
          end else begin
            _EVAL_69 <= 3'h0;
          end
        end else begin
          _EVAL_69 <= _EVAL_241;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_71 <= 3'h0;
    end else begin
      if (_EVAL_136) begin
        if (_EVAL_94) begin
          if (_EVAL_267) begin
            _EVAL_71 <= _EVAL_84;
          end else begin
            _EVAL_71 <= 3'h0;
          end
        end else begin
          _EVAL_71 <= _EVAL_125;
        end
      end
    end
    if (_EVAL_22) begin
      _EVAL_106 <= _EVAL_9;
    end
    if (_EVAL_22) begin
      _EVAL_109 <= _EVAL_11;
    end
    if (_EVAL_22) begin
      _EVAL_116 <= _EVAL_12;
    end
    if (_EVAL_22) begin
      _EVAL_156 <= _EVAL_4;
    end
    if (_EVAL_254) begin
      _EVAL_163 <= _EVAL_13;
    end
    if (_EVAL_254) begin
      _EVAL_165 <= _EVAL_10;
    end
    if (_EVAL_1) begin
      _EVAL_181 <= 32'h0;
    end else begin
      if (_EVAL_114) begin
        _EVAL_181 <= 32'h0;
      end else begin
        _EVAL_181 <= _EVAL_51;
      end
    end
    if (_EVAL_254) begin
      _EVAL_213 <= _EVAL_0;
    end
    if (_EVAL_1) begin
      _EVAL_247 <= 8'h0;
    end else begin
      _EVAL_247 <= _EVAL_169;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbd294d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab7bc0dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e2728d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc168bfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(598a3ab7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d7cbd51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf4fdc2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b00d5a60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2d08900)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d2a87df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e5bff93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78ec812)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64b3f45b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fca89d97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43007d1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b1287a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34ae7a08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56c925d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fe4f54c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78a9153d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c05cf9fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(379d9dc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bf6114a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1edd4df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa4c4b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43be48d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d65cea8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e791ed27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c1f0c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff24ecff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6410998e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb05745)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf292a26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(915d703b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d96eb9c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e38b2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b026dee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4207bbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b89550f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99944328)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61025bfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4548748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9799aa06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beca18d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1d62cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eba2a820)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b49a6dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(654a451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(268e8c50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac028f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d722dd34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(494c6db7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1e3d808)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d6f28b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac8f64b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a8fbd16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(300a4472)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(119411ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc7a3e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f083e0ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20ed685)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff7bc866)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e914dcff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cd5e7f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3062bbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5b78b2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(773a9e64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf668a83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a1baee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30c9f912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ba39490)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38017101)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
