//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_24(
  output [31:0] _EVAL,
  output [3:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  output [1:0]  _EVAL_3,
  output        _EVAL_4,
  input  [3:0]  _EVAL_5,
  output [30:0] _EVAL_6,
  output [1:0]  _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [30:0] _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input  [7:0]  _EVAL_19,
  output [3:0]  _EVAL_20,
  output [3:0]  _EVAL_21,
  input         _EVAL_22,
  output [31:0] _EVAL_23,
  output [3:0]  _EVAL_24,
  output [3:0]  _EVAL_25,
  output [1:0]  _EVAL_26,
  output [2:0]  _EVAL_27,
  input  [31:0] _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  input  [7:0]  _EVAL_32,
  input  [3:0]  _EVAL_33,
  output [3:0]  _EVAL_34,
  output [3:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  output [7:0]  _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  output [2:0]  _EVAL_40,
  output        _EVAL_41,
  output [3:0]  _EVAL_42,
  input         _EVAL_43,
  input  [2:0]  _EVAL_44,
  output        _EVAL_45,
  output        _EVAL_46,
  input  [3:0]  _EVAL_47,
  input         _EVAL_48,
  output [3:0]  _EVAL_49,
  output [2:0]  _EVAL_50,
  input  [1:0]  _EVAL_51,
  output [7:0]  _EVAL_52,
  input  [30:0] _EVAL_53,
  input  [2:0]  _EVAL_54,
  input         _EVAL_55,
  output        _EVAL_56,
  input         _EVAL_57,
  output        _EVAL_58,
  input         _EVAL_59,
  input  [1:0]  _EVAL_60,
  input         _EVAL_61,
  input  [31:0] _EVAL_62,
  input         _EVAL_63,
  output        _EVAL_64,
  input  [3:0]  _EVAL_65,
  output        _EVAL_66,
  input  [1:0]  _EVAL_67,
  output        _EVAL_68,
  output [30:0] _EVAL_69,
  input  [2:0]  _EVAL_70,
  output        _EVAL_71,
  output [1:0]  _EVAL_72,
  input  [3:0]  _EVAL_73,
  input  [2:0]  _EVAL_74
);
  wire  Queue_2__EVAL;
  wire  Queue_2__EVAL_0;
  wire  Queue_2__EVAL_1;
  wire [3:0] Queue_2__EVAL_2;
  wire [1:0] Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire  Queue_2__EVAL_5;
  wire [1:0] Queue_2__EVAL_6;
  wire [3:0] Queue_2__EVAL_7;
  wire  Queue_2__EVAL_8;
  wire  Queue__EVAL;
  wire [1:0] Queue__EVAL_0;
  wire [2:0] Queue__EVAL_1;
  wire [3:0] Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire [7:0] Queue__EVAL_5;
  wire [3:0] Queue__EVAL_6;
  wire [3:0] Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire [30:0] Queue__EVAL_9;
  wire [2:0] Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire  Queue__EVAL_12;
  wire [2:0] Queue__EVAL_13;
  wire [3:0] Queue__EVAL_14;
  wire [2:0] Queue__EVAL_15;
  wire  Queue__EVAL_16;
  wire [3:0] Queue__EVAL_17;
  wire [7:0] Queue__EVAL_18;
  wire [30:0] Queue__EVAL_19;
  wire  Queue__EVAL_20;
  wire [1:0] Queue__EVAL_21;
  wire [3:0] Queue__EVAL_22;
  wire  Queue_3__EVAL;
  wire [1:0] Queue_3__EVAL_0;
  wire [2:0] Queue_3__EVAL_1;
  wire [3:0] Queue_3__EVAL_2;
  wire  Queue_3__EVAL_3;
  wire  Queue_3__EVAL_4;
  wire [7:0] Queue_3__EVAL_5;
  wire [3:0] Queue_3__EVAL_6;
  wire [3:0] Queue_3__EVAL_7;
  wire  Queue_3__EVAL_8;
  wire [30:0] Queue_3__EVAL_9;
  wire [2:0] Queue_3__EVAL_10;
  wire  Queue_3__EVAL_11;
  wire  Queue_3__EVAL_12;
  wire [2:0] Queue_3__EVAL_13;
  wire [3:0] Queue_3__EVAL_14;
  wire [2:0] Queue_3__EVAL_15;
  wire  Queue_3__EVAL_16;
  wire [3:0] Queue_3__EVAL_17;
  wire [7:0] Queue_3__EVAL_18;
  wire [30:0] Queue_3__EVAL_19;
  wire  Queue_3__EVAL_20;
  wire [1:0] Queue_3__EVAL_21;
  wire [3:0] Queue_3__EVAL_22;
  wire [31:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire [31:0] Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire [3:0] Queue_1__EVAL_8;
  wire  Queue_1__EVAL_9;
  wire [3:0] Queue_1__EVAL_10;
  SiFive__EVAL_23 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6),
    ._EVAL_7(Queue_2__EVAL_7),
    ._EVAL_8(Queue_2__EVAL_8)
  );
  SiFive__EVAL_21 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18),
    ._EVAL_19(Queue__EVAL_19),
    ._EVAL_20(Queue__EVAL_20),
    ._EVAL_21(Queue__EVAL_21),
    ._EVAL_22(Queue__EVAL_22)
  );
  SiFive__EVAL_21 Queue_3 (
    ._EVAL(Queue_3__EVAL),
    ._EVAL_0(Queue_3__EVAL_0),
    ._EVAL_1(Queue_3__EVAL_1),
    ._EVAL_2(Queue_3__EVAL_2),
    ._EVAL_3(Queue_3__EVAL_3),
    ._EVAL_4(Queue_3__EVAL_4),
    ._EVAL_5(Queue_3__EVAL_5),
    ._EVAL_6(Queue_3__EVAL_6),
    ._EVAL_7(Queue_3__EVAL_7),
    ._EVAL_8(Queue_3__EVAL_8),
    ._EVAL_9(Queue_3__EVAL_9),
    ._EVAL_10(Queue_3__EVAL_10),
    ._EVAL_11(Queue_3__EVAL_11),
    ._EVAL_12(Queue_3__EVAL_12),
    ._EVAL_13(Queue_3__EVAL_13),
    ._EVAL_14(Queue_3__EVAL_14),
    ._EVAL_15(Queue_3__EVAL_15),
    ._EVAL_16(Queue_3__EVAL_16),
    ._EVAL_17(Queue_3__EVAL_17),
    ._EVAL_18(Queue_3__EVAL_18),
    ._EVAL_19(Queue_3__EVAL_19),
    ._EVAL_20(Queue_3__EVAL_20),
    ._EVAL_21(Queue_3__EVAL_21),
    ._EVAL_22(Queue_3__EVAL_22)
  );
  SiFive__EVAL_22 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10)
  );
  assign _EVAL_52 = Queue_3__EVAL_5;
  assign _EVAL_72 = Queue_3__EVAL_0;
  assign Queue__EVAL_4 = _EVAL_14;
  assign _EVAL_26 = Queue__EVAL_0;
  assign Queue_3__EVAL_12 = _EVAL_55;
  assign Queue_1__EVAL_9 = _EVAL_8;
  assign _EVAL_27 = Queue_3__EVAL_10;
  assign Queue_2__EVAL_5 = _EVAL_43;
  assign Queue__EVAL_21 = _EVAL_2;
  assign Queue__EVAL_12 = _EVAL_13;
  assign Queue_2__EVAL = _EVAL_38;
  assign Queue_3__EVAL_8 = _EVAL_12;
  assign _EVAL_24 = Queue_1__EVAL_10;
  assign _EVAL_68 = _EVAL_63;
  assign _EVAL_36 = Queue__EVAL_10;
  assign _EVAL_4 = Queue__EVAL_11;
  assign _EVAL_11 = Queue__EVAL_16;
  assign _EVAL_21 = Queue__EVAL_22;
  assign Queue_1__EVAL_0 = _EVAL_48;
  assign Queue__EVAL_17 = _EVAL_33;
  assign Queue__EVAL_19 = _EVAL_53;
  assign _EVAL_56 = Queue_2__EVAL_0;
  assign _EVAL_46 = Queue_3__EVAL_11;
  assign _EVAL_42 = Queue_3__EVAL_7;
  assign Queue_1__EVAL_2 = _EVAL_12;
  assign Queue_3__EVAL_1 = _EVAL_74;
  assign Queue_3__EVAL_2 = _EVAL_10;
  assign _EVAL_7 = _EVAL_67;
  assign _EVAL_0 = Queue__EVAL_7;
  assign _EVAL_50 = Queue__EVAL_15;
  assign _EVAL_30 = Queue_3__EVAL_16;
  assign _EVAL_6 = Queue_3__EVAL_9;
  assign _EVAL_25 = Queue_3__EVAL_14;
  assign Queue_3__EVAL_19 = _EVAL_15;
  assign _EVAL_49 = Queue_2__EVAL_2;
  assign Queue_3__EVAL_13 = _EVAL_70;
  assign Queue__EVAL_18 = _EVAL_19;
  assign Queue_2__EVAL_7 = _EVAL_1;
  assign _EVAL_45 = Queue_1__EVAL_6;
  assign _EVAL_58 = _EVAL_18;
  assign _EVAL_40 = Queue_3__EVAL_15;
  assign _EVAL_41 = Queue_1__EVAL_5;
  assign _EVAL_66 = Queue_1__EVAL_7;
  assign _EVAL_35 = Queue_3__EVAL_22;
  assign Queue_1__EVAL = _EVAL_28;
  assign _EVAL_69 = Queue__EVAL_9;
  assign Queue__EVAL = _EVAL_59;
  assign Queue__EVAL_3 = _EVAL_22;
  assign Queue_3__EVAL_3 = _EVAL_17;
  assign _EVAL_20 = Queue__EVAL_14;
  assign _EVAL_31 = Queue_3__EVAL_20;
  assign Queue__EVAL_6 = _EVAL_47;
  assign _EVAL = Queue_1__EVAL_3;
  assign Queue_3__EVAL_6 = _EVAL_73;
  assign Queue_3__EVAL_17 = _EVAL_65;
  assign Queue_1__EVAL_8 = _EVAL_9;
  assign Queue_3__EVAL_18 = _EVAL_32;
  assign Queue_1__EVAL_4 = _EVAL_14;
  assign _EVAL_37 = Queue__EVAL_5;
  assign _EVAL_23 = _EVAL_62;
  assign Queue_2__EVAL_4 = _EVAL_14;
  assign Queue_2__EVAL_3 = _EVAL_51;
  assign _EVAL_3 = Queue_2__EVAL_6;
  assign _EVAL_71 = Queue__EVAL_20;
  assign Queue__EVAL_2 = _EVAL_5;
  assign Queue_3__EVAL_21 = _EVAL_60;
  assign Queue_3__EVAL_4 = _EVAL_14;
  assign _EVAL_29 = Queue_2__EVAL_1;
  assign _EVAL_64 = _EVAL_61;
  assign _EVAL_34 = _EVAL_16;
  assign Queue_3__EVAL = _EVAL_57;
  assign Queue_2__EVAL_8 = _EVAL_12;
  assign Queue__EVAL_1 = _EVAL_54;
  assign Queue_1__EVAL_1 = _EVAL_39;
  assign Queue__EVAL_13 = _EVAL_44;
  assign Queue__EVAL_8 = _EVAL_12;
endmodule
