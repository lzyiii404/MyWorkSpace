//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_78(
  output [7:0]  _EVAL,
  input         _EVAL_0,
  input  [7:0]  _EVAL_1,
  output [7:0]  _EVAL_2,
  input         _EVAL_3,
  output [1:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  output [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  output [7:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  output [1:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  output        _EVAL_15,
  input  [7:0]  _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  output [31:0] _EVAL_19,
  input  [7:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  input  [3:0]  _EVAL_22,
  output [31:0] _EVAL_23,
  output [2:0]  _EVAL_24,
  input  [7:0]  _EVAL_25,
  output [31:0] _EVAL_26,
  input         _EVAL_27,
  output [31:0] _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  input  [7:0]  _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input  [7:0]  _EVAL_34,
  output [7:0]  _EVAL_35,
  input  [2:0]  _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  input  [1:0]  _EVAL_39,
  input  [1:0]  _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  input  [31:0] _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  input  [1:0]  _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  input  [1:0]  _EVAL_49,
  output [1:0]  _EVAL_50,
  input         _EVAL_51,
  output        _EVAL_52,
  output [3:0]  _EVAL_53,
  input         _EVAL_54,
  output [7:0]  _EVAL_55,
  output        _EVAL_56,
  output        _EVAL_57,
  output [7:0]  _EVAL_58
);
  wire [31:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire [31:0] Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire [3:0] Queue_1__EVAL_8;
  wire  Queue_1__EVAL_9;
  wire [3:0] Queue_1__EVAL_10;
  wire  Queue_3__EVAL;
  wire [7:0] Queue_3__EVAL_0;
  wire  Queue_3__EVAL_1;
  wire [1:0] Queue_3__EVAL_2;
  wire [1:0] Queue_3__EVAL_3;
  wire [31:0] Queue_3__EVAL_4;
  wire [2:0] Queue_3__EVAL_5;
  wire [2:0] Queue_3__EVAL_6;
  wire  Queue_3__EVAL_7;
  wire [31:0] Queue_3__EVAL_8;
  wire [7:0] Queue_3__EVAL_9;
  wire  Queue_3__EVAL_10;
  wire [7:0] Queue_3__EVAL_11;
  wire [7:0] Queue_3__EVAL_12;
  wire  Queue_3__EVAL_13;
  wire  Queue_3__EVAL_14;
  wire [7:0] Queue_4__EVAL;
  wire [1:0] Queue_4__EVAL_0;
  wire  Queue_4__EVAL_1;
  wire [31:0] Queue_4__EVAL_2;
  wire  Queue_4__EVAL_3;
  wire  Queue_4__EVAL_4;
  wire  Queue_4__EVAL_5;
  wire  Queue_4__EVAL_6;
  wire  Queue_4__EVAL_7;
  wire [1:0] Queue_4__EVAL_8;
  wire [31:0] Queue_4__EVAL_9;
  wire  Queue_4__EVAL_10;
  wire [7:0] Queue_4__EVAL_11;
  wire  Queue_4__EVAL_12;
  wire  Queue_2__EVAL;
  wire [7:0] Queue_2__EVAL_0;
  wire  Queue_2__EVAL_1;
  wire  Queue_2__EVAL_2;
  wire [7:0] Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire [1:0] Queue_2__EVAL_5;
  wire [1:0] Queue_2__EVAL_6;
  wire  Queue_2__EVAL_7;
  wire  Queue_2__EVAL_8;
  wire  Queue__EVAL;
  wire [7:0] Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire [1:0] Queue__EVAL_2;
  wire [1:0] Queue__EVAL_3;
  wire [31:0] Queue__EVAL_4;
  wire [2:0] Queue__EVAL_5;
  wire [2:0] Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire [31:0] Queue__EVAL_8;
  wire [7:0] Queue__EVAL_9;
  wire  Queue__EVAL_10;
  wire [7:0] Queue__EVAL_11;
  wire [7:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire  Queue__EVAL_14;
  SiFive__EVAL_22 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10)
  );
  SiFive__EVAL_75 Queue_3 (
    ._EVAL(Queue_3__EVAL),
    ._EVAL_0(Queue_3__EVAL_0),
    ._EVAL_1(Queue_3__EVAL_1),
    ._EVAL_2(Queue_3__EVAL_2),
    ._EVAL_3(Queue_3__EVAL_3),
    ._EVAL_4(Queue_3__EVAL_4),
    ._EVAL_5(Queue_3__EVAL_5),
    ._EVAL_6(Queue_3__EVAL_6),
    ._EVAL_7(Queue_3__EVAL_7),
    ._EVAL_8(Queue_3__EVAL_8),
    ._EVAL_9(Queue_3__EVAL_9),
    ._EVAL_10(Queue_3__EVAL_10),
    ._EVAL_11(Queue_3__EVAL_11),
    ._EVAL_12(Queue_3__EVAL_12),
    ._EVAL_13(Queue_3__EVAL_13),
    ._EVAL_14(Queue_3__EVAL_14)
  );
  SiFive__EVAL_77 Queue_4 (
    ._EVAL(Queue_4__EVAL),
    ._EVAL_0(Queue_4__EVAL_0),
    ._EVAL_1(Queue_4__EVAL_1),
    ._EVAL_2(Queue_4__EVAL_2),
    ._EVAL_3(Queue_4__EVAL_3),
    ._EVAL_4(Queue_4__EVAL_4),
    ._EVAL_5(Queue_4__EVAL_5),
    ._EVAL_6(Queue_4__EVAL_6),
    ._EVAL_7(Queue_4__EVAL_7),
    ._EVAL_8(Queue_4__EVAL_8),
    ._EVAL_9(Queue_4__EVAL_9),
    ._EVAL_10(Queue_4__EVAL_10),
    ._EVAL_11(Queue_4__EVAL_11),
    ._EVAL_12(Queue_4__EVAL_12)
  );
  SiFive__EVAL_76 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6),
    ._EVAL_7(Queue_2__EVAL_7),
    ._EVAL_8(Queue_2__EVAL_8)
  );
  SiFive__EVAL_75 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14)
  );
  assign _EVAL_15 = Queue_1__EVAL_5;
  assign Queue_2__EVAL_0 = _EVAL_25;
  assign Queue_2__EVAL_6 = _EVAL_46;
  assign Queue__EVAL_13 = _EVAL_33;
  assign _EVAL_21 = Queue__EVAL_5;
  assign _EVAL_55 = Queue_3__EVAL_9;
  assign Queue_4__EVAL = _EVAL_20;
  assign _EVAL_19 = Queue_4__EVAL_2;
  assign Queue_2__EVAL_2 = _EVAL_32;
  assign Queue__EVAL_8 = _EVAL_12;
  assign _EVAL_56 = Queue_3__EVAL_14;
  assign _EVAL_26 = Queue_3__EVAL_4;
  assign _EVAL_53 = Queue_1__EVAL_10;
  assign _EVAL_8 = Queue_4__EVAL_8;
  assign _EVAL_35 = Queue__EVAL_9;
  assign _EVAL_23 = Queue_1__EVAL_3;
  assign Queue_3__EVAL_0 = _EVAL_16;
  assign Queue_2__EVAL_8 = _EVAL_5;
  assign Queue_3__EVAL_6 = _EVAL_36;
  assign Queue_4__EVAL_4 = _EVAL_29;
  assign Queue_4__EVAL_5 = _EVAL_54;
  assign _EVAL_48 = Queue_2__EVAL;
  assign Queue_1__EVAL_2 = _EVAL_33;
  assign _EVAL_37 = Queue__EVAL_14;
  assign _EVAL_57 = Queue_4__EVAL_12;
  assign Queue_2__EVAL_7 = _EVAL_33;
  assign Queue_1__EVAL_1 = _EVAL_45;
  assign Queue__EVAL = _EVAL_32;
  assign Queue_3__EVAL_2 = _EVAL_39;
  assign _EVAL = Queue_4__EVAL_11;
  assign Queue_4__EVAL_3 = _EVAL_32;
  assign _EVAL_47 = Queue_4__EVAL_1;
  assign Queue_3__EVAL_1 = _EVAL_3;
  assign Queue_2__EVAL_4 = _EVAL_9;
  assign _EVAL_38 = Queue__EVAL_7;
  assign _EVAL_24 = Queue_3__EVAL_5;
  assign _EVAL_28 = Queue__EVAL_4;
  assign _EVAL_30 = Queue_1__EVAL_7;
  assign Queue_3__EVAL_10 = _EVAL_51;
  assign Queue_1__EVAL_4 = _EVAL_32;
  assign Queue__EVAL_12 = _EVAL_31;
  assign Queue__EVAL_6 = _EVAL_7;
  assign Queue__EVAL_1 = _EVAL_27;
  assign Queue_1__EVAL_8 = _EVAL_22;
  assign _EVAL_50 = Queue__EVAL_3;
  assign _EVAL_58 = Queue_3__EVAL_11;
  assign _EVAL_41 = Queue_4__EVAL_6;
  assign Queue_3__EVAL_8 = _EVAL_14;
  assign Queue__EVAL_2 = _EVAL_40;
  assign Queue__EVAL_0 = _EVAL_1;
  assign _EVAL_4 = Queue_3__EVAL_3;
  assign _EVAL_2 = Queue__EVAL_11;
  assign Queue_1__EVAL_9 = _EVAL_6;
  assign Queue__EVAL_10 = _EVAL_42;
  assign _EVAL_13 = Queue_2__EVAL_5;
  assign Queue_3__EVAL_12 = _EVAL_34;
  assign Queue_4__EVAL_7 = _EVAL_33;
  assign _EVAL_52 = Queue_2__EVAL_1;
  assign _EVAL_11 = Queue_2__EVAL_3;
  assign _EVAL_17 = Queue_1__EVAL_6;
  assign _EVAL_18 = Queue_3__EVAL_7;
  assign Queue_1__EVAL = _EVAL_10;
  assign Queue_4__EVAL_10 = _EVAL_44;
  assign Queue_4__EVAL_9 = _EVAL_43;
  assign Queue_3__EVAL_13 = _EVAL_33;
  assign Queue_3__EVAL = _EVAL_32;
  assign Queue_4__EVAL_0 = _EVAL_49;
  assign Queue_1__EVAL_0 = _EVAL_0;
endmodule
