//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_62(
  input  [31:0] _EVAL,
  output [4:0]  _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  input  [2:0]  _EVAL_4,
  output [3:0]  _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  output [2:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  output [31:0] _EVAL_13,
  output [4:0]  _EVAL_14,
  input  [4:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  output        _EVAL_17,
  output [31:0] _EVAL_18,
  input         _EVAL_19,
  input  [4:0]  _EVAL_20,
  output [31:0] _EVAL_21,
  output [3:0]  _EVAL_22,
  input         _EVAL_23,
  input  [31:0] _EVAL_24,
  input  [3:0]  _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input  [2:0]  _EVAL_29,
  output [1:0]  _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  output [2:0]  _EVAL_33,
  input  [3:0]  _EVAL_34,
  input         _EVAL_35,
  output        _EVAL_36,
  output [3:0]  _EVAL_37,
  input  [3:0]  _EVAL_38,
  output        _EVAL_39,
  input  [1:0]  _EVAL_40
);
  assign _EVAL_30 = _EVAL_40;
  assign _EVAL_0 = _EVAL_20;
  assign _EVAL_5 = _EVAL_34;
  assign _EVAL_11 = _EVAL_29;
  assign _EVAL_13 = _EVAL_10;
  assign _EVAL_17 = _EVAL_35;
  assign _EVAL_6 = _EVAL_26;
  assign _EVAL_39 = _EVAL_1;
  assign _EVAL_14 = _EVAL_15;
  assign _EVAL_3 = _EVAL_23;
  assign _EVAL_21 = _EVAL_24;
  assign _EVAL_22 = _EVAL_25;
  assign _EVAL_12 = _EVAL_16;
  assign _EVAL_37 = _EVAL_38;
  assign _EVAL_2 = _EVAL_9;
  assign _EVAL_36 = _EVAL_27;
  assign _EVAL_18 = _EVAL;
  assign _EVAL_8 = _EVAL_19;
  assign _EVAL_31 = _EVAL_32;
  assign _EVAL_33 = _EVAL_4;
endmodule
