//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_155(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output [14:0] _EVAL_3,
  output [2:0]  _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input  [11:0] _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input  [31:0] _EVAL_10,
  output [2:0]  _EVAL_11,
  output [11:0] _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [2:0]  _EVAL_18,
  output [1:0]  _EVAL_19,
  input  [6:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  output        _EVAL_23,
  input  [2:0]  _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [31:0] _EVAL_26,
  output [3:0]  _EVAL_27,
  input  [14:0] _EVAL_28,
  output [2:0]  _EVAL_29,
  output [6:0]  _EVAL_30,
  input         _EVAL_31,
  input  [3:0]  _EVAL_32
);
  wire [14:0] Repeater__EVAL;
  wire [3:0] Repeater__EVAL_0;
  wire  Repeater__EVAL_1;
  wire  Repeater__EVAL_2;
  wire [6:0] Repeater__EVAL_3;
  wire [3:0] Repeater__EVAL_4;
  wire  Repeater__EVAL_5;
  wire [2:0] Repeater__EVAL_6;
  wire  Repeater__EVAL_7;
  wire  Repeater__EVAL_8;
  wire [2:0] Repeater__EVAL_9;
  wire  Repeater__EVAL_10;
  wire [2:0] Repeater__EVAL_11;
  wire  Repeater__EVAL_12;
  wire  Repeater__EVAL_13;
  wire  Repeater__EVAL_14;
  wire [6:0] Repeater__EVAL_15;
  wire [14:0] Repeater__EVAL_16;
  wire [2:0] Repeater__EVAL_17;
  wire [2:0] Repeater__EVAL_18;
  wire [2:0] Repeater__EVAL_19;
  wire  Repeater__EVAL_20;
  reg  _EVAL_46;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_75;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_115;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_116;
  reg [31:0] _RAND_3;
  reg  _EVAL_120;
  reg [31:0] _RAND_4;
  wire [4:0] _EVAL_123;
  wire [1:0] _EVAL_90;
  wire  _EVAL_57;
  wire  _EVAL_107;
  wire  _EVAL_100;
  wire [3:0] _EVAL_65;
  wire [5:0] _EVAL_34;
  wire [1:0] _EVAL_53;
  wire [5:0] _EVAL_63;
  wire [5:0] _EVAL_89;
  wire [6:0] _EVAL_50;
  wire [6:0] _EVAL_108;
  wire [6:0] _EVAL_96;
  wire [6:0] _EVAL_49;
  wire [6:0] _EVAL_35;
  wire [3:0] _EVAL_55;
  wire  _EVAL_106;
  wire  _EVAL_121;
  wire  _EVAL_41;
  wire  _EVAL_83;
  wire [12:0] _EVAL_82;
  wire [5:0] _EVAL_51;
  wire [5:0] _EVAL_45;
  wire [3:0] _EVAL_40;
  wire [3:0] _EVAL_36;
  wire [3:0] _EVAL_105;
  wire [5:0] _EVAL_56;
  wire [5:0] _EVAL_77;
  wire [5:0] _EVAL_43;
  wire  _EVAL_70;
  wire [2:0] _EVAL_68;
  wire [8:0] _EVAL_37;
  wire [1:0] _EVAL_73;
  wire [1:0] _EVAL_111;
  wire [5:0] _EVAL_60;
  wire [5:0] _EVAL_92;
  wire  _EVAL_86;
  wire  _EVAL_94;
  wire  _EVAL_72;
  wire  _EVAL_84;
  wire  _EVAL_33;
  wire  _EVAL_88;
  wire  _EVAL_76;
  wire  _EVAL_117;
  wire  _EVAL_102;
  wire [2:0] _EVAL_98;
  wire [3:0] _EVAL_71;
  wire [3:0] _EVAL_48;
  wire [1:0] _EVAL_62;
  wire [3:0] _EVAL_110;
  wire [2:0] _EVAL_113;
  wire  _EVAL_67;
  wire  _EVAL_38;
  wire [3:0] _EVAL_66;
  wire [3:0] _EVAL_61;
  wire  _EVAL_47;
  wire  _EVAL_69;
  wire  _EVAL_52;
  wire [1:0] _EVAL_104;
  wire  _EVAL_103;
  wire [1:0] _EVAL_39;
  wire  _EVAL_78;
  wire [2:0] _EVAL_114;
  wire [3:0] _EVAL_119;
  wire [3:0] _EVAL_42;
  wire [5:0] _EVAL_118;
  wire [5:0] _EVAL_109;
  wire  _EVAL_91;
  wire [14:0] _EVAL_99;
  wire [7:0] _EVAL_80;
  SiFive__EVAL_154 Repeater (
    ._EVAL(Repeater__EVAL),
    ._EVAL_0(Repeater__EVAL_0),
    ._EVAL_1(Repeater__EVAL_1),
    ._EVAL_2(Repeater__EVAL_2),
    ._EVAL_3(Repeater__EVAL_3),
    ._EVAL_4(Repeater__EVAL_4),
    ._EVAL_5(Repeater__EVAL_5),
    ._EVAL_6(Repeater__EVAL_6),
    ._EVAL_7(Repeater__EVAL_7),
    ._EVAL_8(Repeater__EVAL_8),
    ._EVAL_9(Repeater__EVAL_9),
    ._EVAL_10(Repeater__EVAL_10),
    ._EVAL_11(Repeater__EVAL_11),
    ._EVAL_12(Repeater__EVAL_12),
    ._EVAL_13(Repeater__EVAL_13),
    ._EVAL_14(Repeater__EVAL_14),
    ._EVAL_15(Repeater__EVAL_15),
    ._EVAL_16(Repeater__EVAL_16),
    ._EVAL_17(Repeater__EVAL_17),
    ._EVAL_18(Repeater__EVAL_18),
    ._EVAL_19(Repeater__EVAL_19),
    ._EVAL_20(Repeater__EVAL_20)
  );
  assign _EVAL_123 = 5'h3 << _EVAL_15;
  assign _EVAL_90 = _EVAL_123[1:0];
  assign _EVAL_57 = _EVAL_25[0];
  assign _EVAL_107 = Repeater__EVAL_1;
  assign _EVAL_100 = _EVAL_0 & _EVAL_107;
  assign _EVAL_65 = _EVAL_7[3:0];
  assign _EVAL_34 = {_EVAL_65, 2'h0};
  assign _EVAL_53 = ~ _EVAL_90;
  assign _EVAL_63 = {{4'd0}, _EVAL_53};
  assign _EVAL_89 = _EVAL_34 | _EVAL_63;
  assign _EVAL_50 = {_EVAL_89, 1'h0};
  assign _EVAL_108 = _EVAL_50 | 7'h1;
  assign _EVAL_96 = {1'h0,_EVAL_89};
  assign _EVAL_49 = ~ _EVAL_96;
  assign _EVAL_35 = _EVAL_108 & _EVAL_49;
  assign _EVAL_55 = _EVAL_35[3:0];
  assign _EVAL_106 = _EVAL_115 == 4'h0;
  assign _EVAL_121 = Repeater__EVAL_11[2];
  assign _EVAL_41 = _EVAL_121 == 1'h0;
  assign _EVAL_83 = _EVAL_41 == 1'h0;
  assign _EVAL_82 = 13'h3f << Repeater__EVAL_6;
  assign _EVAL_51 = _EVAL_82[5:0];
  assign _EVAL_45 = ~ _EVAL_51;
  assign _EVAL_40 = _EVAL_45[5:2];
  assign _EVAL_36 = _EVAL_115 - 4'h1;
  assign _EVAL_105 = _EVAL_106 ? _EVAL_40 : _EVAL_36;
  assign _EVAL_56 = {_EVAL_105, 2'h0};
  assign _EVAL_77 = ~ _EVAL_45;
  assign _EVAL_43 = _EVAL_56 | _EVAL_77;
  assign _EVAL_70 = Repeater__EVAL_6 > 3'h2;
  assign _EVAL_68 = _EVAL_70 ? 3'h2 : Repeater__EVAL_6;
  assign _EVAL_37 = 9'h3 << _EVAL_68;
  assign _EVAL_73 = _EVAL_37[1:0];
  assign _EVAL_111 = ~ _EVAL_73;
  assign _EVAL_60 = {{4'd0}, _EVAL_111};
  assign _EVAL_92 = _EVAL_43 | _EVAL_60;
  assign _EVAL_86 = _EVAL_106 ? _EVAL_46 : _EVAL_120;
  assign _EVAL_94 = _EVAL_86 == 1'h0;
  assign _EVAL_72 = _EVAL_57 == 1'h0;
  assign _EVAL_84 = _EVAL_65 == 4'h0;
  assign _EVAL_33 = _EVAL_84 == 1'h0;
  assign _EVAL_88 = _EVAL_72 & _EVAL_33;
  assign _EVAL_76 = _EVAL_31 | _EVAL_88;
  assign _EVAL_117 = _EVAL_76 & _EVAL_6;
  assign _EVAL_102 = _EVAL_88 == 1'h0;
  assign _EVAL_98 = _EVAL_35[6:4];
  assign _EVAL_71 = {{1'd0}, _EVAL_98};
  assign _EVAL_48 = _EVAL_71 | _EVAL_55;
  assign _EVAL_62 = _EVAL_48[1:0];
  assign _EVAL_110 = 4'h1 << _EVAL_15;
  assign _EVAL_113 = _EVAL_110[2:0];
  assign _EVAL_67 = _EVAL_113[2:2];
  assign _EVAL_38 = _EVAL_57 ? 1'h1 : _EVAL_67;
  assign _EVAL_66 = {{3'd0}, _EVAL_38};
  assign _EVAL_61 = _EVAL_75 - _EVAL_66;
  assign _EVAL_47 = _EVAL_75 == 4'h0;
  assign _EVAL_69 = _EVAL_7[4];
  assign _EVAL_52 = _EVAL_98 != 3'h0;
  assign _EVAL_104 = _EVAL_48[3:2];
  assign _EVAL_103 = _EVAL_104 != 2'h0;
  assign _EVAL_39 = _EVAL_104 | _EVAL_62;
  assign _EVAL_78 = _EVAL_39[1];
  assign _EVAL_114 = {_EVAL_52,_EVAL_103,_EVAL_78};
  assign _EVAL_119 = ~ _EVAL_105;
  assign _EVAL_42 = ~ _EVAL_119;
  assign _EVAL_118 = _EVAL_92 | 6'h3;
  assign _EVAL_109 = ~ _EVAL_118;
  assign _EVAL_91 = _EVAL_42 != 4'h0;
  assign _EVAL_99 = {{9'd0}, _EVAL_109};
  assign _EVAL_80 = {Repeater__EVAL_15,_EVAL_94};
  assign _EVAL_29 = _EVAL_25;
  assign _EVAL_5 = _EVAL_31 | _EVAL_88;
  assign _EVAL_26 = _EVAL_17;
  assign Repeater__EVAL_14 = _EVAL_14;
  assign Repeater__EVAL_2 = _EVAL_2;
  assign _EVAL_19 = _EVAL_68[1:0];
  assign _EVAL_27 = Repeater__EVAL_20 ? 4'hf : _EVAL_32;
  assign _EVAL_12 = {_EVAL_80,_EVAL_42};
  assign _EVAL_9 = _EVAL_6 & _EVAL_102;
  assign _EVAL_13 = Repeater__EVAL_10;
  assign Repeater__EVAL_7 = _EVAL;
  assign Repeater__EVAL = _EVAL_28;
  assign _EVAL_11 = Repeater__EVAL_18;
  assign _EVAL_4 = _EVAL_47 ? _EVAL_114 : _EVAL_116;
  assign Repeater__EVAL_17 = _EVAL_24;
  assign Repeater__EVAL_8 = _EVAL_1;
  assign _EVAL_3 = Repeater__EVAL_16 | _EVAL_99;
  assign _EVAL_16 = _EVAL_10;
  assign Repeater__EVAL_5 = _EVAL_83 & _EVAL_91;
  assign Repeater__EVAL_9 = _EVAL_21;
  assign _EVAL_22 = Repeater__EVAL_11;
  assign _EVAL_23 = Repeater__EVAL_13;
  assign _EVAL_30 = _EVAL_7[11:5];
  assign Repeater__EVAL_3 = _EVAL_20;
  assign Repeater__EVAL_19 = _EVAL_18;
  assign _EVAL_8 = Repeater__EVAL_1;
  assign Repeater__EVAL_0 = _EVAL_32;
  assign Repeater__EVAL_12 = _EVAL_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_46 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_75 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_115 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_116 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_120 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL_1) begin
      _EVAL_46 <= 1'h0;
    end else begin
      if (_EVAL_117) begin
        if (_EVAL_47) begin
          _EVAL_46 <= _EVAL_69;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_75 <= 4'h0;
    end else begin
      if (_EVAL_117) begin
        if (_EVAL_47) begin
          _EVAL_75 <= _EVAL_65;
        end else begin
          _EVAL_75 <= _EVAL_61;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_115 <= 4'h0;
    end else begin
      if (_EVAL_100) begin
        _EVAL_115 <= _EVAL_42;
      end
    end
    if (_EVAL_117) begin
      if (_EVAL_47) begin
        _EVAL_116 <= _EVAL_114;
      end
    end
    if (_EVAL_106) begin
      _EVAL_120 <= _EVAL_46;
    end
  end
endmodule
