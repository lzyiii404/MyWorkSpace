//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_5_assert(
  input  [2:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [31:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input  [7:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input  [3:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  input         _EVAL_20,
  input  [3:0]  _EVAL_21,
  input         _EVAL_22,
  input  [31:0] _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input  [1:0]  _EVAL_27,
  input  [3:0]  _EVAL_28,
  input         _EVAL_29,
  input  [2:0]  _EVAL_30,
  input  [31:0] _EVAL_31,
  input         _EVAL_32
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_43;
  reg [31:0] _RAND_0;
  reg [4:0] _EVAL_58;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_64;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_70;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_95;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_99;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_109;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_169;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_173;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_187;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_211;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_237;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_257;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_323;
  reg [31:0] _RAND_13;
  reg [31:0] _EVAL_343;
  reg [31:0] _RAND_14;
  reg [4:0] _EVAL_387;
  reg [31:0] _RAND_15;
  reg [4:0] _EVAL_450;
  reg [31:0] _RAND_16;
  reg [1:0] _EVAL_488;
  reg [31:0] _RAND_17;
  reg [1:0] _EVAL_491;
  reg [31:0] _RAND_18;
  reg [31:0] _EVAL_509;
  reg [31:0] _RAND_19;
  reg [4:0] _EVAL_561;
  reg [31:0] _RAND_20;
  reg  _EVAL_568;
  reg [31:0] _RAND_21;
  reg [4:0] _EVAL_619;
  reg [31:0] _RAND_22;
  reg [3:0] _EVAL_622;
  reg [31:0] _RAND_23;
  reg [4:0] _EVAL_634;
  reg [31:0] _RAND_24;
  reg [8:0] _EVAL_636;
  reg [31:0] _RAND_25;
  reg  _EVAL_646;
  reg [31:0] _RAND_26;
  reg [3:0] _EVAL_668;
  reg [31:0] _RAND_27;
  wire  _EVAL_367;
  wire  _EVAL_174;
  wire  _EVAL_276;
  wire [15:0] _EVAL_448;
  wire [15:0] _EVAL_555;
  wire [8:0] _EVAL_462;
  wire  _EVAL_290;
  wire  _EVAL_658;
  wire [7:0] _EVAL_152;
  wire  _EVAL_416;
  wire  _EVAL_147;
  wire  _EVAL_136;
  wire  _EVAL_617;
  wire  _EVAL_325;
  wire  _EVAL_566;
  wire [31:0] _EVAL_469;
  wire [32:0] _EVAL_111;
  wire [32:0] _EVAL_85;
  wire [32:0] _EVAL_621;
  wire  _EVAL_119;
  wire [31:0] _EVAL_527;
  wire [32:0] _EVAL_626;
  wire [32:0] _EVAL_504;
  wire [32:0] _EVAL_389;
  wire  _EVAL_269;
  wire  _EVAL_239;
  wire [31:0] _EVAL_368;
  wire [32:0] _EVAL_406;
  wire [32:0] _EVAL_224;
  wire [32:0] _EVAL_374;
  wire  _EVAL_103;
  wire  _EVAL_333;
  wire [31:0] _EVAL_630;
  wire [32:0] _EVAL_34;
  wire [32:0] _EVAL_664;
  wire [32:0] _EVAL_296;
  wire  _EVAL_649;
  wire  _EVAL_559;
  wire [32:0] _EVAL_602;
  wire [32:0] _EVAL_487;
  wire [32:0] _EVAL_362;
  wire  _EVAL_606;
  wire  _EVAL_357;
  wire [31:0] _EVAL_377;
  wire [32:0] _EVAL_394;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_317;
  wire  _EVAL_471;
  wire  _EVAL_507;
  wire [31:0] _EVAL_180;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_393;
  wire [32:0] _EVAL_370;
  wire  _EVAL_304;
  wire  _EVAL_590;
  wire [31:0] _EVAL_141;
  wire [32:0] _EVAL_282;
  wire [32:0] _EVAL_86;
  wire [32:0] _EVAL_196;
  wire  _EVAL_643;
  wire  _EVAL_660;
  wire [31:0] _EVAL_135;
  wire [32:0] _EVAL_403;
  wire [32:0] _EVAL_577;
  wire  _EVAL_353;
  wire  _EVAL_115;
  wire [4:0] _EVAL_298;
  wire  _EVAL_369;
  wire [1:0] _EVAL_68;
  wire [3:0] _EVAL_101;
  wire [2:0] _EVAL_506;
  wire [2:0] _EVAL_199;
  wire  _EVAL_235;
  wire  _EVAL_334;
  wire  _EVAL_49;
  wire  _EVAL_388;
  wire  _EVAL_274;
  wire  _EVAL_319;
  wire  _EVAL_656;
  wire  _EVAL_508;
  wire  _EVAL_314;
  wire  _EVAL_404;
  wire  _EVAL_261;
  wire  _EVAL_539;
  wire  _EVAL_110;
  wire  _EVAL_505;
  wire  _EVAL_277;
  wire  _EVAL_595;
  wire  _EVAL_558;
  wire  _EVAL_591;
  wire  _EVAL_234;
  wire  _EVAL_548;
  wire  _EVAL_513;
  wire  _EVAL_220;
  wire  _EVAL_184;
  wire  _EVAL_456;
  wire  _EVAL_405;
  wire  _EVAL_165;
  wire  _EVAL_364;
  wire  _EVAL_311;
  wire  _EVAL_241;
  wire  _EVAL_162;
  wire  _EVAL_142;
  wire  _EVAL_356;
  wire  _EVAL_243;
  wire  _EVAL_151;
  wire  _EVAL_285;
  wire  _EVAL_73;
  wire  _EVAL_209;
  wire  _EVAL_549;
  wire  _EVAL_320;
  wire  _EVAL_308;
  wire  _EVAL_185;
  wire  _EVAL_263;
  wire  _EVAL_252;
  wire  _EVAL_418;
  wire  _EVAL_248;
  wire  _EVAL_671;
  wire  _EVAL_365;
  wire  _EVAL_391;
  wire  _EVAL_256;
  wire [7:0] _EVAL_193;
  wire [7:0] _EVAL_438;
  wire [7:0] _EVAL_570;
  wire  _EVAL_412;
  wire  _EVAL_597;
  wire  _EVAL_358;
  wire  _EVAL_516;
  wire  _EVAL_593;
  wire  _EVAL_512;
  wire  _EVAL_330;
  wire  _EVAL_114;
  wire  _EVAL_81;
  wire  _EVAL_168;
  wire  _EVAL_378;
  wire  _EVAL_231;
  wire [31:0] _EVAL_611;
  wire  _EVAL_189;
  wire  _EVAL_286;
  wire [2:0] _EVAL_425;
  wire  _EVAL_108;
  wire  _EVAL_586;
  wire  _EVAL_289;
  wire  _EVAL_349;
  wire  _EVAL_473;
  wire  _EVAL_603;
  wire  _EVAL_496;
  wire [15:0] _EVAL_642;
  wire [15:0] _EVAL_219;
  wire [8:0] _EVAL_88;
  wire  _EVAL_588;
  wire  _EVAL_287;
  wire  _EVAL_655;
  wire  _EVAL_259;
  wire  _EVAL_641;
  wire [31:0] _EVAL_175;
  wire [32:0] _EVAL_569;
  wire [32:0] _EVAL_486;
  wire [32:0] _EVAL_443;
  wire  _EVAL_584;
  wire  _EVAL_464;
  wire  _EVAL_544;
  wire  _EVAL_659;
  wire  _EVAL_572;
  wire  _EVAL_321;
  wire  _EVAL_275;
  wire  _EVAL_309;
  wire  _EVAL_492;
  wire [22:0] _EVAL_262;
  wire [7:0] _EVAL_266;
  wire [7:0] _EVAL_562;
  wire [4:0] _EVAL_436;
  wire  _EVAL_520;
  wire [8:0] _EVAL_93;
  wire [8:0] _EVAL_251;
  wire  _EVAL_490;
  wire  _EVAL_116;
  wire  _EVAL_402;
  wire  _EVAL_46;
  wire  _EVAL_650;
  wire  _EVAL_42;
  wire [8:0] _EVAL_542;
  wire [1:0] _EVAL_340;
  wire  _EVAL_587;
  wire  _EVAL_466;
  wire  _EVAL_297;
  wire  _EVAL_533;
  wire [31:0] _EVAL_379;
  wire [32:0] _EVAL_376;
  wire [32:0] _EVAL_255;
  wire [32:0] _EVAL_172;
  wire  _EVAL_214;
  wire  _EVAL_52;
  wire [31:0] _EVAL_47;
  wire [32:0] _EVAL_383;
  wire [1:0] _EVAL_208;
  wire [31:0] _EVAL_153;
  wire  _EVAL_122;
  wire  _EVAL_460;
  wire  _EVAL_327;
  wire  _EVAL_413;
  wire [22:0] _EVAL_439;
  wire [7:0] _EVAL_574;
  wire  _EVAL_40;
  wire  _EVAL_575;
  wire  _EVAL_41;
  wire  _EVAL_518;
  wire  _EVAL_154;
  wire  _EVAL_373;
  wire  _EVAL_74;
  wire  _EVAL_186;
  wire  _EVAL_534;
  wire  _EVAL_210;
  wire  _EVAL_183;
  wire  _EVAL_361;
  wire  _EVAL_546;
  wire [31:0] _EVAL_638;
  wire [7:0] _EVAL_283;
  wire [4:0] _EVAL_381;
  wire [4:0] _EVAL_607;
  wire [31:0] _EVAL_594;
  wire [32:0] _EVAL_76;
  wire [32:0] _EVAL_233;
  wire [32:0] _EVAL_503;
  wire  _EVAL_557;
  wire [31:0] _EVAL_176;
  wire [32:0] _EVAL_435;
  wire [32:0] _EVAL_300;
  wire [32:0] _EVAL_605;
  wire  _EVAL_395;
  wire  _EVAL_665;
  wire [31:0] _EVAL_72;
  wire [32:0] _EVAL_221;
  wire [32:0] _EVAL_223;
  wire [32:0] _EVAL_667;
  wire  _EVAL_167;
  wire  _EVAL_635;
  wire [31:0] _EVAL_480;
  wire [32:0] _EVAL_576;
  wire [32:0] _EVAL_647;
  wire [32:0] _EVAL_158;
  wire  _EVAL_51;
  wire  _EVAL_98;
  wire [31:0] _EVAL_400;
  wire [32:0] _EVAL_206;
  wire [32:0] _EVAL_83;
  wire [32:0] _EVAL_53;
  wire  _EVAL_482;
  wire  _EVAL_84;
  wire [32:0] _EVAL_627;
  wire [32:0] _EVAL_331;
  wire [32:0] _EVAL_215;
  wire  _EVAL_472;
  wire  _EVAL_273;
  wire  _EVAL_560;
  wire  _EVAL_424;
  wire [32:0] _EVAL_91;
  wire [32:0] _EVAL_112;
  wire  _EVAL_531;
  wire  _EVAL_226;
  wire  _EVAL_552;
  wire  _EVAL_337;
  wire  _EVAL_80;
  wire  _EVAL_629;
  wire  _EVAL_344;
  wire  _EVAL_543;
  wire  _EVAL_316;
  wire  _EVAL_582;
  wire  _EVAL_360;
  wire  _EVAL_526;
  wire  _EVAL_547;
  wire  _EVAL_144;
  wire  _EVAL_538;
  wire  _EVAL_522;
  wire  _EVAL_198;
  wire  _EVAL_87;
  wire  _EVAL_493;
  wire  _EVAL_341;
  wire  _EVAL_652;
  wire  _EVAL_218;
  wire  _EVAL_295;
  wire  _EVAL_382;
  wire  _EVAL_645;
  wire  _EVAL_288;
  wire  _EVAL_307;
  wire  _EVAL_213;
  wire [22:0] _EVAL_258;
  wire [7:0] _EVAL_56;
  wire [7:0] _EVAL_514;
  wire [4:0] _EVAL_238;
  wire [4:0] _EVAL_294;
  wire  _EVAL_397;
  wire  _EVAL_69;
  wire  _EVAL_657;
  wire  _EVAL_35;
  wire  _EVAL_511;
  wire  _EVAL_432;
  wire [31:0] _EVAL_225;
  wire [32:0] _EVAL_179;
  wire [32:0] _EVAL_342;
  wire [8:0] _EVAL_417;
  wire  _EVAL_481;
  wire  _EVAL_474;
  wire  _EVAL_236;
  wire [31:0] _EVAL_386;
  wire [32:0] _EVAL_270;
  wire  _EVAL_240;
  wire  _EVAL_65;
  wire  _EVAL_585;
  wire [32:0] _EVAL_579;
  wire  _EVAL_339;
  wire  _EVAL_384;
  wire  _EVAL_354;
  wire  _EVAL_609;
  wire  _EVAL_281;
  wire  _EVAL_434;
  wire  _EVAL_501;
  wire  _EVAL_163;
  wire  _EVAL_500;
  wire  _EVAL_583;
  wire  _EVAL_305;
  wire  _EVAL_431;
  wire  _EVAL_38;
  wire  _EVAL_502;
  wire  _EVAL_573;
  wire  _EVAL_477;
  wire [32:0] _EVAL_127;
  wire [32:0] _EVAL_485;
  wire  _EVAL_524;
  wire  _EVAL_188;
  wire  _EVAL_399;
  wire  _EVAL_444;
  wire [31:0] _EVAL_553;
  wire [32:0] _EVAL_366;
  wire [32:0] _EVAL_616;
  wire [32:0] _EVAL_625;
  wire  _EVAL_128;
  wire [31:0] _EVAL_267;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_254;
  wire [32:0] _EVAL_195;
  wire  _EVAL_249;
  wire  _EVAL_437;
  wire [31:0] _EVAL_312;
  wire [32:0] _EVAL_554;
  wire [32:0] _EVAL_78;
  wire [32:0] _EVAL_644;
  wire  _EVAL_429;
  wire  _EVAL_345;
  wire [32:0] _EVAL_39;
  wire  _EVAL_350;
  wire  _EVAL_517;
  wire [31:0] _EVAL_145;
  wire [32:0] _EVAL_246;
  wire [32:0] _EVAL_57;
  wire [32:0] _EVAL_385;
  wire  _EVAL_371;
  wire  _EVAL_229;
  wire  _EVAL_467;
  wire  _EVAL_293;
  wire  _EVAL_600;
  wire  _EVAL_632;
  wire  _EVAL_355;
  wire  _EVAL_648;
  wire  _EVAL_410;
  wire  _EVAL_244;
  wire  _EVAL_36;
  wire  _EVAL_75;
  wire  _EVAL_279;
  wire  _EVAL_421;
  wire  _EVAL_138;
  wire  _EVAL_63;
  wire  _EVAL_89;
  wire  _EVAL_60;
  wire  _EVAL_161;
  wire  _EVAL_280;
  wire  _EVAL_589;
  wire  _EVAL_302;
  wire  _EVAL_441;
  wire  _EVAL_216;
  wire  _EVAL_537;
  wire [32:0] _EVAL_470;
  wire [32:0] _EVAL_156;
  wire  _EVAL_301;
  wire  _EVAL_401;
  wire [31:0] _EVAL_133;
  wire [31:0] _EVAL_408;
  wire  _EVAL_515;
  wire  _EVAL_310;
  wire  _EVAL_134;
  wire  _EVAL_166;
  wire  _EVAL_227;
  wire  _EVAL_468;
  wire  _EVAL_228;
  wire  _EVAL_409;
  wire  _EVAL_155;
  wire  _EVAL_662;
  wire [1:0] _EVAL_322;
  wire [1:0] _EVAL_499;
  wire [1:0] _EVAL_232;
  wire [1:0] _EVAL_565;
  wire [32:0] _EVAL_61;
  wire  _EVAL_623;
  wire  _EVAL_96;
  wire [31:0] _EVAL_640;
  wire [32:0] _EVAL_663;
  wire [32:0] _EVAL_118;
  wire [32:0] _EVAL_182;
  wire  _EVAL_205;
  wire  _EVAL_171;
  wire [32:0] _EVAL_426;
  wire [32:0] _EVAL_59;
  wire [32:0] _EVAL_45;
  wire  _EVAL_494;
  wire  _EVAL_428;
  wire  _EVAL_615;
  wire  _EVAL_318;
  wire  _EVAL_50;
  wire  _EVAL_102;
  wire  _EVAL_670;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_126;
  wire  _EVAL_71;
  wire [4:0] _EVAL_442;
  wire  _EVAL_124;
  wire [4:0] _EVAL_247;
  wire  _EVAL_217;
  wire [31:0] _EVAL_550;
  wire [32:0] _EVAL_100;
  wire [32:0] _EVAL_146;
  wire [32:0] _EVAL_529;
  wire  _EVAL_48;
  wire  _EVAL_375;
  wire  _EVAL_614;
  wire  _EVAL_571;
  wire  _EVAL_201;
  wire [31:0] _EVAL_303;
  wire [32:0] _EVAL_123;
  wire [32:0] _EVAL_398;
  wire [32:0] _EVAL_82;
  wire  _EVAL_264;
  wire  _EVAL_564;
  wire  _EVAL_620;
  wire  _EVAL_446;
  wire  _EVAL_639;
  wire [2:0] _EVAL_618;
  wire  _EVAL_427;
  wire  _EVAL_592;
  wire  _EVAL_580;
  wire  _EVAL_465;
  wire  _EVAL_521;
  wire  _EVAL_336;
  wire  _EVAL_284;
  wire  _EVAL_242;
  wire [2:0] _EVAL_148;
  wire  _EVAL_272;
  wire  _EVAL_420;
  wire  _EVAL_265;
  wire  _EVAL_351;
  wire  _EVAL_495;
  wire  _EVAL_433;
  wire  _EVAL_445;
  wire  _EVAL_540;
  wire  _EVAL_414;
  wire  _EVAL_440;
  wire  _EVAL_352;
  wire  _EVAL_77;
  wire  _EVAL_207;
  wire  _EVAL_411;
  wire  _EVAL_396;
  wire  _EVAL_497;
  wire [4:0] _EVAL_245;
  wire  _EVAL_528;
  wire  _EVAL_479;
  wire  _EVAL_651;
  wire  _EVAL_140;
  wire  _EVAL_661;
  wire  _EVAL_181;
  wire  _EVAL_536;
  wire  _EVAL_105;
  wire  _EVAL_291;
  wire  _EVAL_332;
  wire  _EVAL_447;
  wire  _EVAL_278;
  wire  _EVAL_463;
  wire  _EVAL_461;
  wire  _EVAL_338;
  wire  _EVAL_525;
  wire  _EVAL_407;
  wire  _EVAL_192;
  wire  _EVAL_458;
  wire  _EVAL_160;
  wire  _EVAL_551;
  wire  _EVAL_599;
  wire  _EVAL_415;
  wire  _EVAL_324;
  wire  _EVAL_131;
  wire [8:0] _EVAL_335;
  wire  _EVAL_556;
  wire  _EVAL_347;
  wire  _EVAL_419;
  wire  _EVAL_392;
  wire  _EVAL_567;
  wire  _EVAL_106;
  wire  _EVAL_510;
  wire  _EVAL_654;
  wire  _EVAL_372;
  wire  _EVAL_107;
  wire [31:0] _EVAL_422;
  wire [31:0] _EVAL_633;
  wire  _EVAL_535;
  wire  _EVAL_612;
  wire  _EVAL_129;
  wire  _EVAL_170;
  wire  _EVAL_523;
  wire  _EVAL_578;
  wire  _EVAL_610;
  wire  _EVAL_653;
  wire  _EVAL_326;
  wire  _EVAL_250;
  wire  _EVAL_608;
  wire  _EVAL_628;
  wire  _EVAL_423;
  wire [4:0] _EVAL_313;
  wire [1:0] _EVAL_203;
  wire [1:0] _EVAL_449;
  wire  _EVAL_624;
  wire  _EVAL_430;
  wire  _EVAL_489;
  wire  _EVAL_476;
  wire  _EVAL_117;
  wire  _EVAL_455;
  wire  _EVAL_222;
  wire  _EVAL_143;
  wire  _EVAL_268;
  wire  _EVAL_178;
  wire  _EVAL_94;
  wire  _EVAL_601;
  wire  _EVAL_260;
  wire  _EVAL_545;
  wire  _EVAL_581;
  wire  _EVAL_197;
  wire  _EVAL_457;
  wire  _EVAL_62;
  wire  _EVAL_79;
  wire  _EVAL_666;
  wire  _EVAL_90;
  wire  _EVAL_125;
  wire  _EVAL_204;
  wire  _EVAL_194;
  wire [8:0] _EVAL_328;
  wire  _EVAL_306;
  wire  _EVAL_315;
  wire  _EVAL_598;
  wire [1:0] _EVAL_359;
  wire  _EVAL_613;
  wire  _EVAL_97;
  wire  _EVAL_348;
  wire  _EVAL_669;
  wire  _EVAL_230;
  wire  _EVAL_498;
  wire  _EVAL_92;
  wire  _EVAL_519;
  wire  _EVAL_459;
  wire  _EVAL_159;
  wire  _EVAL_113;
  wire  _EVAL_363;
  wire  _EVAL_346;
  wire  _EVAL_253;
  wire  _EVAL_120;
  wire [1:0] _EVAL_604;
  wire  _EVAL_202;
  wire  _EVAL_475;
  wire  _EVAL_177;
  wire  _EVAL_452;
  wire  _EVAL_200;
  wire  _EVAL_149;
  wire  _EVAL_191;
  wire  _EVAL_563;
  wire  _EVAL_164;
  wire  _EVAL_67;
  wire  _EVAL_530;
  wire  _EVAL_292;
  wire  _EVAL_478;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_367 = _EVAL_5 & _EVAL_8;
  assign _EVAL_174 = _EVAL_450 == 5'h0;
  assign _EVAL_276 = _EVAL_367 & _EVAL_174;
  assign _EVAL_448 = 16'h1 << _EVAL_28;
  assign _EVAL_555 = _EVAL_276 ? _EVAL_448 : 16'h0;
  assign _EVAL_462 = _EVAL_555[8:0];
  assign _EVAL_290 = _EVAL_462 != 9'h0;
  assign _EVAL_658 = _EVAL_290 == 1'h0;
  assign _EVAL_152 = ~ _EVAL_9;
  assign _EVAL_416 = _EVAL_19 == 3'h0;
  assign _EVAL_147 = _EVAL_30 == 3'h0;
  assign _EVAL_136 = _EVAL_147 | _EVAL_1;
  assign _EVAL_617 = _EVAL_11 == 4'h8;
  assign _EVAL_325 = _EVAL_387 == 5'h0;
  assign _EVAL_566 = _EVAL_325 == 1'h0;
  assign _EVAL_469 = _EVAL_4 ^ 32'h40000000;
  assign _EVAL_111 = {1'b0,$signed(_EVAL_469)};
  assign _EVAL_85 = $signed(_EVAL_111) & $signed(-33'sh2000);
  assign _EVAL_621 = $signed(_EVAL_85);
  assign _EVAL_119 = $signed(_EVAL_621) == $signed(33'sh0);
  assign _EVAL_527 = _EVAL_4 ^ 32'h80000000;
  assign _EVAL_626 = {1'b0,$signed(_EVAL_527)};
  assign _EVAL_504 = $signed(_EVAL_626) & $signed(-33'sh20000);
  assign _EVAL_389 = $signed(_EVAL_504);
  assign _EVAL_269 = $signed(_EVAL_389) == $signed(33'sh0);
  assign _EVAL_239 = _EVAL_119 | _EVAL_269;
  assign _EVAL_368 = _EVAL_4 ^ 32'hc000000;
  assign _EVAL_406 = {1'b0,$signed(_EVAL_368)};
  assign _EVAL_224 = $signed(_EVAL_406) & $signed(-33'sh4000000);
  assign _EVAL_374 = $signed(_EVAL_224);
  assign _EVAL_103 = $signed(_EVAL_374) == $signed(33'sh0);
  assign _EVAL_333 = _EVAL_239 | _EVAL_103;
  assign _EVAL_630 = _EVAL_4 ^ 32'h2000000;
  assign _EVAL_34 = {1'b0,$signed(_EVAL_630)};
  assign _EVAL_664 = $signed(_EVAL_34) & $signed(-33'sh10000);
  assign _EVAL_296 = $signed(_EVAL_664);
  assign _EVAL_649 = $signed(_EVAL_296) == $signed(33'sh0);
  assign _EVAL_559 = _EVAL_333 | _EVAL_649;
  assign _EVAL_602 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_487 = $signed(_EVAL_602) & $signed(-33'sh5000);
  assign _EVAL_362 = $signed(_EVAL_487);
  assign _EVAL_606 = $signed(_EVAL_362) == $signed(33'sh0);
  assign _EVAL_357 = _EVAL_559 | _EVAL_606;
  assign _EVAL_377 = _EVAL_4 ^ 32'h1800000;
  assign _EVAL_394 = {1'b0,$signed(_EVAL_377)};
  assign _EVAL_104 = $signed(_EVAL_394) & $signed(-33'sh8000);
  assign _EVAL_317 = $signed(_EVAL_104);
  assign _EVAL_471 = $signed(_EVAL_317) == $signed(33'sh0);
  assign _EVAL_507 = _EVAL_357 | _EVAL_471;
  assign _EVAL_180 = _EVAL_4 ^ 32'h1900000;
  assign _EVAL_150 = {1'b0,$signed(_EVAL_180)};
  assign _EVAL_393 = $signed(_EVAL_150) & $signed(-33'sh2000);
  assign _EVAL_370 = $signed(_EVAL_393);
  assign _EVAL_304 = $signed(_EVAL_370) == $signed(33'sh0);
  assign _EVAL_590 = _EVAL_507 | _EVAL_304;
  assign _EVAL_141 = _EVAL_4 ^ 32'h20000000;
  assign _EVAL_282 = {1'b0,$signed(_EVAL_141)};
  assign _EVAL_86 = $signed(_EVAL_282) & $signed(-33'sh2000);
  assign _EVAL_196 = $signed(_EVAL_86);
  assign _EVAL_643 = $signed(_EVAL_196) == $signed(33'sh0);
  assign _EVAL_660 = _EVAL_590 | _EVAL_643;
  assign _EVAL_135 = _EVAL_31 ^ 32'hc000000;
  assign _EVAL_403 = {1'b0,$signed(_EVAL_135)};
  assign _EVAL_577 = $signed(_EVAL_403) & $signed(-33'sh4000000);
  assign _EVAL_353 = _EVAL_634 == 5'h0;
  assign _EVAL_115 = _EVAL_32 & _EVAL_20;
  assign _EVAL_298 = _EVAL_634 - 5'h1;
  assign _EVAL_369 = _EVAL_0 >= 4'h3;
  assign _EVAL_68 = _EVAL_0[1:0];
  assign _EVAL_101 = 4'h1 << _EVAL_68;
  assign _EVAL_506 = _EVAL_101[2:0];
  assign _EVAL_199 = _EVAL_506 | 3'h1;
  assign _EVAL_235 = _EVAL_199[2];
  assign _EVAL_334 = _EVAL_4[2];
  assign _EVAL_49 = _EVAL_235 & _EVAL_334;
  assign _EVAL_388 = _EVAL_369 | _EVAL_49;
  assign _EVAL_274 = _EVAL_199[1];
  assign _EVAL_319 = _EVAL_4[1];
  assign _EVAL_656 = _EVAL_334 & _EVAL_319;
  assign _EVAL_508 = _EVAL_274 & _EVAL_656;
  assign _EVAL_314 = _EVAL_388 | _EVAL_508;
  assign _EVAL_404 = _EVAL_199[0];
  assign _EVAL_261 = _EVAL_4[0];
  assign _EVAL_539 = _EVAL_656 & _EVAL_261;
  assign _EVAL_110 = _EVAL_404 & _EVAL_539;
  assign _EVAL_505 = _EVAL_314 | _EVAL_110;
  assign _EVAL_277 = _EVAL_261 == 1'h0;
  assign _EVAL_595 = _EVAL_656 & _EVAL_277;
  assign _EVAL_558 = _EVAL_404 & _EVAL_595;
  assign _EVAL_591 = _EVAL_314 | _EVAL_558;
  assign _EVAL_234 = _EVAL_319 == 1'h0;
  assign _EVAL_548 = _EVAL_334 & _EVAL_234;
  assign _EVAL_513 = _EVAL_274 & _EVAL_548;
  assign _EVAL_220 = _EVAL_388 | _EVAL_513;
  assign _EVAL_184 = _EVAL_548 & _EVAL_261;
  assign _EVAL_456 = _EVAL_404 & _EVAL_184;
  assign _EVAL_405 = _EVAL_220 | _EVAL_456;
  assign _EVAL_165 = _EVAL_548 & _EVAL_277;
  assign _EVAL_364 = _EVAL_404 & _EVAL_165;
  assign _EVAL_311 = _EVAL_220 | _EVAL_364;
  assign _EVAL_241 = _EVAL_334 == 1'h0;
  assign _EVAL_162 = _EVAL_235 & _EVAL_241;
  assign _EVAL_142 = _EVAL_369 | _EVAL_162;
  assign _EVAL_356 = _EVAL_241 & _EVAL_319;
  assign _EVAL_243 = _EVAL_274 & _EVAL_356;
  assign _EVAL_151 = _EVAL_142 | _EVAL_243;
  assign _EVAL_285 = _EVAL_356 & _EVAL_261;
  assign _EVAL_73 = _EVAL_404 & _EVAL_285;
  assign _EVAL_209 = _EVAL_151 | _EVAL_73;
  assign _EVAL_549 = _EVAL_356 & _EVAL_277;
  assign _EVAL_320 = _EVAL_404 & _EVAL_549;
  assign _EVAL_308 = _EVAL_151 | _EVAL_320;
  assign _EVAL_185 = _EVAL_241 & _EVAL_234;
  assign _EVAL_263 = _EVAL_274 & _EVAL_185;
  assign _EVAL_252 = _EVAL_142 | _EVAL_263;
  assign _EVAL_418 = _EVAL_185 & _EVAL_261;
  assign _EVAL_248 = _EVAL_404 & _EVAL_418;
  assign _EVAL_671 = _EVAL_252 | _EVAL_248;
  assign _EVAL_365 = _EVAL_185 & _EVAL_277;
  assign _EVAL_391 = _EVAL_404 & _EVAL_365;
  assign _EVAL_256 = _EVAL_252 | _EVAL_391;
  assign _EVAL_193 = {_EVAL_505,_EVAL_591,_EVAL_405,_EVAL_311,_EVAL_209,_EVAL_308,_EVAL_671,_EVAL_256};
  assign _EVAL_438 = ~ _EVAL_193;
  assign _EVAL_570 = _EVAL_9 & _EVAL_438;
  assign _EVAL_412 = _EVAL_7[3:3];
  assign _EVAL_597 = _EVAL_31 == _EVAL_323;
  assign _EVAL_358 = _EVAL_597 | _EVAL_1;
  assign _EVAL_516 = _EVAL_358 == 1'h0;
  assign _EVAL_593 = _EVAL_353 == 1'h0;
  assign _EVAL_512 = _EVAL_20 & _EVAL_593;
  assign _EVAL_330 = _EVAL_6 & _EVAL_566;
  assign _EVAL_114 = _EVAL_152 == 8'h0;
  assign _EVAL_81 = _EVAL_114 | _EVAL_1;
  assign _EVAL_168 = _EVAL_30 != 3'h0;
  assign _EVAL_378 = _EVAL_2 & _EVAL_6;
  assign _EVAL_231 = _EVAL_367 | _EVAL_378;
  assign _EVAL_611 = _EVAL_509 + 32'h1;
  assign _EVAL_189 = _EVAL_28[3:3];
  assign _EVAL_286 = _EVAL_189 == 1'h0;
  assign _EVAL_425 = _EVAL_28[2:0];
  assign _EVAL_108 = 3'h1 <= _EVAL_425;
  assign _EVAL_586 = _EVAL_286 & _EVAL_108;
  assign _EVAL_289 = _EVAL_561 == 5'h0;
  assign _EVAL_349 = _EVAL_378 & _EVAL_289;
  assign _EVAL_473 = _EVAL_14 == 3'h6;
  assign _EVAL_603 = _EVAL_473 == 1'h0;
  assign _EVAL_496 = _EVAL_349 & _EVAL_603;
  assign _EVAL_642 = 16'h1 << _EVAL_11;
  assign _EVAL_219 = _EVAL_496 ? _EVAL_642 : 16'h0;
  assign _EVAL_88 = _EVAL_219[8:0];
  assign _EVAL_588 = _EVAL_462 != _EVAL_88;
  assign _EVAL_287 = _EVAL_588 | _EVAL_658;
  assign _EVAL_655 = _EVAL_28 == _EVAL_237;
  assign _EVAL_259 = _EVAL_655 | _EVAL_1;
  assign _EVAL_641 = _EVAL_259 == 1'h0;
  assign _EVAL_175 = _EVAL_4 ^ 32'h3000;
  assign _EVAL_569 = {1'b0,$signed(_EVAL_175)};
  assign _EVAL_486 = $signed(_EVAL_569) & $signed(-33'sh1000);
  assign _EVAL_443 = $signed(_EVAL_486);
  assign _EVAL_584 = $signed(_EVAL_443) == $signed(33'sh0);
  assign _EVAL_464 = _EVAL_584 | _EVAL_103;
  assign _EVAL_544 = _EVAL_464 | _EVAL_649;
  assign _EVAL_659 = _EVAL_211 == 5'h0;
  assign _EVAL_572 = _EVAL_659 == 1'h0;
  assign _EVAL_321 = _EVAL_8 & _EVAL_572;
  assign _EVAL_275 = _EVAL_7 == _EVAL_43;
  assign _EVAL_309 = _EVAL_19[2];
  assign _EVAL_492 = _EVAL_309 == 1'h0;
  assign _EVAL_262 = 23'hff << _EVAL_0;
  assign _EVAL_266 = _EVAL_262[7:0];
  assign _EVAL_562 = ~ _EVAL_266;
  assign _EVAL_436 = _EVAL_562[7:3];
  assign _EVAL_520 = _EVAL_10 == 3'h6;
  assign _EVAL_93 = _EVAL_462 | _EVAL_636;
  assign _EVAL_251 = _EVAL_93 >> _EVAL_11;
  assign _EVAL_490 = _EVAL == 3'h0;
  assign _EVAL_116 = _EVAL_490 | _EVAL_1;
  assign _EVAL_402 = _EVAL_18 >= 4'h3;
  assign _EVAL_46 = _EVAL_3 == 1'h0;
  assign _EVAL_650 = _EVAL_46 | _EVAL_1;
  assign _EVAL_42 = _EVAL_650 == 1'h0;
  assign _EVAL_542 = _EVAL_636 | _EVAL_462;
  assign _EVAL_340 = 2'h1 << _EVAL_26;
  assign _EVAL_587 = _EVAL_17 == _EVAL_488;
  assign _EVAL_466 = _EVAL_587 | _EVAL_1;
  assign _EVAL_297 = _EVAL_466 == 1'h0;
  assign _EVAL_533 = _EVAL_12 & _EVAL_24;
  assign _EVAL_379 = _EVAL_31 ^ 32'h20000000;
  assign _EVAL_376 = {1'b0,$signed(_EVAL_379)};
  assign _EVAL_255 = $signed(_EVAL_376) & $signed(-33'sh2000);
  assign _EVAL_172 = $signed(_EVAL_255);
  assign _EVAL_214 = $signed(_EVAL_172) == $signed(33'sh0);
  assign _EVAL_52 = _EVAL_0 <= 4'h8;
  assign _EVAL_47 = _EVAL_31 ^ 32'h4000;
  assign _EVAL_383 = {1'b0,$signed(_EVAL_47)};
  assign _EVAL_208 = _EVAL_95 >> _EVAL_13;
  assign _EVAL_153 = _EVAL_23 & 32'h3f;
  assign _EVAL_122 = _EVAL_153 == 32'h0;
  assign _EVAL_460 = _EVAL_122 | _EVAL_1;
  assign _EVAL_327 = _EVAL_460 == 1'h0;
  assign _EVAL_413 = _EVAL_18 == _EVAL_70;
  assign _EVAL_439 = 23'hff << _EVAL_21;
  assign _EVAL_574 = _EVAL_439[7:0];
  assign _EVAL_40 = _EVAL_619 == 5'h0;
  assign _EVAL_575 = _EVAL_378 & _EVAL_40;
  assign _EVAL_41 = _EVAL_14[2];
  assign _EVAL_518 = _EVAL_14[1];
  assign _EVAL_154 = _EVAL_518 == 1'h0;
  assign _EVAL_373 = _EVAL_41 & _EVAL_154;
  assign _EVAL_74 = _EVAL_575 & _EVAL_373;
  assign _EVAL_186 = _EVAL_19 == 3'h6;
  assign _EVAL_534 = _EVAL_0 <= 4'h6;
  assign _EVAL_210 = _EVAL_534 & _EVAL_660;
  assign _EVAL_183 = _EVAL_168 | _EVAL_1;
  assign _EVAL_361 = _EVAL_27 == _EVAL_491;
  assign _EVAL_546 = _EVAL_361 | _EVAL_1;
  assign _EVAL_638 = _EVAL_31 ^ 32'h1900000;
  assign _EVAL_283 = ~ _EVAL_574;
  assign _EVAL_381 = _EVAL_283[7:3];
  assign _EVAL_607 = _EVAL_619 - 5'h1;
  assign _EVAL_594 = _EVAL_23 ^ 32'h40000000;
  assign _EVAL_76 = {1'b0,$signed(_EVAL_594)};
  assign _EVAL_233 = $signed(_EVAL_76) & $signed(-33'sh2000);
  assign _EVAL_503 = $signed(_EVAL_233);
  assign _EVAL_557 = $signed(_EVAL_503) == $signed(33'sh0);
  assign _EVAL_176 = _EVAL_23 ^ 32'h80000000;
  assign _EVAL_435 = {1'b0,$signed(_EVAL_176)};
  assign _EVAL_300 = $signed(_EVAL_435) & $signed(-33'sh20000);
  assign _EVAL_605 = $signed(_EVAL_300);
  assign _EVAL_395 = $signed(_EVAL_605) == $signed(33'sh0);
  assign _EVAL_665 = _EVAL_557 | _EVAL_395;
  assign _EVAL_72 = _EVAL_23 ^ 32'h3000;
  assign _EVAL_221 = {1'b0,$signed(_EVAL_72)};
  assign _EVAL_223 = $signed(_EVAL_221) & $signed(-33'sh1000);
  assign _EVAL_667 = $signed(_EVAL_223);
  assign _EVAL_167 = $signed(_EVAL_667) == $signed(33'sh0);
  assign _EVAL_635 = _EVAL_665 | _EVAL_167;
  assign _EVAL_480 = _EVAL_23 ^ 32'hc000000;
  assign _EVAL_576 = {1'b0,$signed(_EVAL_480)};
  assign _EVAL_647 = $signed(_EVAL_576) & $signed(-33'sh4000000);
  assign _EVAL_158 = $signed(_EVAL_647);
  assign _EVAL_51 = $signed(_EVAL_158) == $signed(33'sh0);
  assign _EVAL_98 = _EVAL_635 | _EVAL_51;
  assign _EVAL_400 = _EVAL_23 ^ 32'h2000000;
  assign _EVAL_206 = {1'b0,$signed(_EVAL_400)};
  assign _EVAL_83 = $signed(_EVAL_206) & $signed(-33'sh10000);
  assign _EVAL_53 = $signed(_EVAL_83);
  assign _EVAL_482 = $signed(_EVAL_53) == $signed(33'sh0);
  assign _EVAL_84 = _EVAL_98 | _EVAL_482;
  assign _EVAL_627 = {1'b0,$signed(_EVAL_23)};
  assign _EVAL_331 = $signed(_EVAL_627) & $signed(-33'sh1000);
  assign _EVAL_215 = $signed(_EVAL_331);
  assign _EVAL_472 = $signed(_EVAL_215) == $signed(33'sh0);
  assign _EVAL_273 = _EVAL_84 | _EVAL_472;
  assign _EVAL_560 = _EVAL_30 <= 3'h2;
  assign _EVAL_424 = _EVAL_560 | _EVAL_1;
  assign _EVAL_91 = $signed(_EVAL_383) & $signed(-33'sh1000);
  assign _EVAL_112 = $signed(_EVAL_91);
  assign _EVAL_531 = $signed(_EVAL_112) == $signed(33'sh0);
  assign _EVAL_226 = _EVAL_22 == 1'h0;
  assign _EVAL_552 = _EVAL_19 == _EVAL_173;
  assign _EVAL_337 = _EVAL_552 | _EVAL_1;
  assign _EVAL_80 = _EVAL_337 == 1'h0;
  assign _EVAL_629 = _EVAL == _EVAL_187;
  assign _EVAL_344 = _EVAL_629 | _EVAL_1;
  assign _EVAL_543 = _EVAL_344 == 1'h0;
  assign _EVAL_316 = _EVAL_424 == 1'h0;
  assign _EVAL_582 = plusarg_reader_out == 32'h0;
  assign _EVAL_360 = _EVAL_19 == 3'h1;
  assign _EVAL_526 = _EVAL_8 & _EVAL_360;
  assign _EVAL_547 = _EVAL_52 & _EVAL_584;
  assign _EVAL_144 = _EVAL_210 | _EVAL_547;
  assign _EVAL_538 = _EVAL_144 | _EVAL_1;
  assign _EVAL_522 = _EVAL_538 == 1'h0;
  assign _EVAL_198 = _EVAL <= 3'h2;
  assign _EVAL_87 = _EVAL_198 | _EVAL_1;
  assign _EVAL_493 = _EVAL_570 == 8'h0;
  assign _EVAL_341 = _EVAL_493 | _EVAL_1;
  assign _EVAL_652 = _EVAL_341 == 1'h0;
  assign _EVAL_218 = _EVAL_0 == _EVAL_169;
  assign _EVAL_295 = _EVAL_218 | _EVAL_1;
  assign _EVAL_382 = _EVAL_295 == 1'h0;
  assign _EVAL_645 = _EVAL_534 & _EVAL_269;
  assign _EVAL_288 = _EVAL_645 | _EVAL_1;
  assign _EVAL_307 = _EVAL_288 == 1'h0;
  assign _EVAL_213 = _EVAL_14[0];
  assign _EVAL_258 = 23'hff << _EVAL_18;
  assign _EVAL_56 = _EVAL_258[7:0];
  assign _EVAL_514 = ~ _EVAL_56;
  assign _EVAL_238 = _EVAL_514[7:3];
  assign _EVAL_294 = _EVAL_561 - 5'h1;
  assign _EVAL_397 = _EVAL_369 | _EVAL_1;
  assign _EVAL_69 = _EVAL_397 == 1'h0;
  assign _EVAL_657 = _EVAL_14 == 3'h0;
  assign _EVAL_35 = _EVAL_27 <= 2'h2;
  assign _EVAL_511 = _EVAL_35 | _EVAL_1;
  assign _EVAL_432 = _EVAL_511 == 1'h0;
  assign _EVAL_225 = _EVAL_23 ^ 32'h20000000;
  assign _EVAL_179 = {1'b0,$signed(_EVAL_225)};
  assign _EVAL_342 = $signed(_EVAL_179) & $signed(-33'sh2000);
  assign _EVAL_417 = _EVAL_636 >> _EVAL_28;
  assign _EVAL_481 = _EVAL_417[0];
  assign _EVAL_474 = _EVAL_481 == 1'h0;
  assign _EVAL_236 = _EVAL_474 | _EVAL_1;
  assign _EVAL_386 = _EVAL_23 ^ 32'h1800000;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_386)};
  assign _EVAL_240 = _EVAL_636 != 9'h0;
  assign _EVAL_65 = _EVAL_240 == 1'h0;
  assign _EVAL_585 = _EVAL_65 | _EVAL_582;
  assign _EVAL_579 = $signed(_EVAL_342);
  assign _EVAL_339 = $signed(_EVAL_579) == $signed(33'sh0);
  assign _EVAL_384 = _EVAL_21 >= 4'h3;
  assign _EVAL_354 = _EVAL_384 | _EVAL_1;
  assign _EVAL_609 = _EVAL_354 == 1'h0;
  assign _EVAL_281 = _EVAL_7 == 4'h8;
  assign _EVAL_434 = _EVAL <= 3'h5;
  assign _EVAL_501 = _EVAL_434 | _EVAL_1;
  assign _EVAL_163 = _EVAL_23 == _EVAL_343;
  assign _EVAL_500 = _EVAL_163 | _EVAL_1;
  assign _EVAL_583 = _EVAL_208[0];
  assign _EVAL_305 = _EVAL_583 == 1'h0;
  assign _EVAL_431 = _EVAL_305 | _EVAL_1;
  assign _EVAL_38 = _EVAL_431 == 1'h0;
  assign _EVAL_502 = _EVAL_16 == 1'h0;
  assign _EVAL_573 = _EVAL_502 | _EVAL_1;
  assign _EVAL_477 = _EVAL_573 == 1'h0;
  assign _EVAL_127 = $signed(_EVAL_270) & $signed(-33'sh8000);
  assign _EVAL_485 = $signed(_EVAL_127);
  assign _EVAL_524 = $signed(_EVAL_485) == $signed(33'sh0);
  assign _EVAL_188 = _EVAL_30 <= 3'h3;
  assign _EVAL_399 = _EVAL_188 | _EVAL_1;
  assign _EVAL_444 = _EVAL_399 == 1'h0;
  assign _EVAL_553 = _EVAL_31 ^ 32'h40000000;
  assign _EVAL_366 = {1'b0,$signed(_EVAL_553)};
  assign _EVAL_616 = $signed(_EVAL_366) & $signed(-33'sh2000);
  assign _EVAL_625 = $signed(_EVAL_616);
  assign _EVAL_128 = $signed(_EVAL_625) == $signed(33'sh0);
  assign _EVAL_267 = _EVAL_31 ^ 32'h80000000;
  assign _EVAL_130 = {1'b0,$signed(_EVAL_267)};
  assign _EVAL_254 = $signed(_EVAL_130) & $signed(-33'sh20000);
  assign _EVAL_195 = $signed(_EVAL_254);
  assign _EVAL_249 = $signed(_EVAL_195) == $signed(33'sh0);
  assign _EVAL_437 = _EVAL_128 | _EVAL_249;
  assign _EVAL_312 = _EVAL_31 ^ 32'h3000;
  assign _EVAL_554 = {1'b0,$signed(_EVAL_312)};
  assign _EVAL_78 = $signed(_EVAL_554) & $signed(-33'sh1000);
  assign _EVAL_644 = $signed(_EVAL_78);
  assign _EVAL_429 = $signed(_EVAL_644) == $signed(33'sh0);
  assign _EVAL_345 = _EVAL_437 | _EVAL_429;
  assign _EVAL_39 = $signed(_EVAL_577);
  assign _EVAL_350 = $signed(_EVAL_39) == $signed(33'sh0);
  assign _EVAL_517 = _EVAL_345 | _EVAL_350;
  assign _EVAL_145 = _EVAL_31 ^ 32'h2000000;
  assign _EVAL_246 = {1'b0,$signed(_EVAL_145)};
  assign _EVAL_57 = $signed(_EVAL_246) & $signed(-33'sh10000);
  assign _EVAL_385 = $signed(_EVAL_57);
  assign _EVAL_371 = $signed(_EVAL_385) == $signed(33'sh0);
  assign _EVAL_229 = _EVAL_517 | _EVAL_371;
  assign _EVAL_467 = _EVAL_21 <= 4'h6;
  assign _EVAL_293 = _EVAL_467 & _EVAL_249;
  assign _EVAL_600 = _EVAL_293 | _EVAL_1;
  assign _EVAL_632 = _EVAL_600 == 1'h0;
  assign _EVAL_355 = _EVAL_9 == _EVAL_193;
  assign _EVAL_648 = _EVAL_355 | _EVAL_1;
  assign _EVAL_410 = _EVAL_27 == 2'h0;
  assign _EVAL_244 = _EVAL_410 | _EVAL_1;
  assign _EVAL_36 = _EVAL_244 == 1'h0;
  assign _EVAL_75 = _EVAL_502 | _EVAL_3;
  assign _EVAL_279 = _EVAL_75 | _EVAL_1;
  assign _EVAL_421 = _EVAL_0 <= 4'h2;
  assign _EVAL_138 = _EVAL_544 | _EVAL_606;
  assign _EVAL_63 = _EVAL_138 | _EVAL_471;
  assign _EVAL_89 = _EVAL_63 | _EVAL_304;
  assign _EVAL_60 = _EVAL_89 | _EVAL_643;
  assign _EVAL_161 = _EVAL_421 & _EVAL_60;
  assign _EVAL_280 = _EVAL_19 == 3'h5;
  assign _EVAL_589 = _EVAL_8 & _EVAL_280;
  assign _EVAL_302 = _EVAL_116 == 1'h0;
  assign _EVAL_441 = _EVAL_501 == 1'h0;
  assign _EVAL_216 = _EVAL_8 & _EVAL_416;
  assign _EVAL_537 = _EVAL_11 == _EVAL_622;
  assign _EVAL_470 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_156 = $signed(_EVAL_470) & $signed(-33'sh1000);
  assign _EVAL_301 = _EVAL_10 == 3'h0;
  assign _EVAL_401 = _EVAL_24 & _EVAL_301;
  assign _EVAL_133 = {{24'd0}, _EVAL_283};
  assign _EVAL_408 = _EVAL_31 & _EVAL_133;
  assign _EVAL_515 = _EVAL_408 == 32'h0;
  assign _EVAL_310 = _EVAL_515 | _EVAL_1;
  assign _EVAL_134 = _EVAL_310 == 1'h0;
  assign _EVAL_166 = _EVAL_14 == _EVAL_99;
  assign _EVAL_227 = _EVAL_166 | _EVAL_1;
  assign _EVAL_468 = _EVAL_227 == 1'h0;
  assign _EVAL_228 = 4'h6 == _EVAL_21;
  assign _EVAL_409 = _EVAL_28 == 4'h8;
  assign _EVAL_155 = _EVAL_28 == 4'h0;
  assign _EVAL_662 = _EVAL_409 | _EVAL_155;
  assign _EVAL_322 = 2'h1 << _EVAL_13;
  assign _EVAL_499 = _EVAL_74 ? _EVAL_322 : 2'h0;
  assign _EVAL_232 = _EVAL_499 | _EVAL_95;
  assign _EVAL_565 = _EVAL_232 >> _EVAL_26;
  assign _EVAL_61 = $signed(_EVAL_156);
  assign _EVAL_623 = $signed(_EVAL_61) == $signed(33'sh0);
  assign _EVAL_96 = _EVAL_229 | _EVAL_623;
  assign _EVAL_640 = _EVAL_31 ^ 32'h1800000;
  assign _EVAL_663 = {1'b0,$signed(_EVAL_640)};
  assign _EVAL_118 = $signed(_EVAL_663) & $signed(-33'sh8000);
  assign _EVAL_182 = $signed(_EVAL_118);
  assign _EVAL_205 = $signed(_EVAL_182) == $signed(33'sh0);
  assign _EVAL_171 = _EVAL_96 | _EVAL_205;
  assign _EVAL_426 = {1'b0,$signed(_EVAL_638)};
  assign _EVAL_59 = $signed(_EVAL_426) & $signed(-33'sh2000);
  assign _EVAL_45 = $signed(_EVAL_59);
  assign _EVAL_494 = $signed(_EVAL_45) == $signed(33'sh0);
  assign _EVAL_428 = _EVAL_171 | _EVAL_494;
  assign _EVAL_615 = _EVAL_428 | _EVAL_531;
  assign _EVAL_318 = _EVAL_615 | _EVAL_214;
  assign _EVAL_50 = _EVAL_318 | _EVAL_1;
  assign _EVAL_102 = _EVAL_50 == 1'h0;
  assign _EVAL_670 = _EVAL_10 == 3'h5;
  assign _EVAL_483 = _EVAL_21 == _EVAL_668;
  assign _EVAL_484 = _EVAL_251[0];
  assign _EVAL_126 = _EVAL_484 | _EVAL_1;
  assign _EVAL_71 = _EVAL_8 & _EVAL_186;
  assign _EVAL_442 = _EVAL_450 - 5'h1;
  assign _EVAL_124 = _EVAL_648 == 1'h0;
  assign _EVAL_247 = _EVAL_211 - 5'h1;
  assign _EVAL_217 = _EVAL_273 | _EVAL_524;
  assign _EVAL_550 = _EVAL_23 ^ 32'h1900000;
  assign _EVAL_100 = {1'b0,$signed(_EVAL_550)};
  assign _EVAL_146 = $signed(_EVAL_100) & $signed(-33'sh2000);
  assign _EVAL_529 = $signed(_EVAL_146);
  assign _EVAL_48 = $signed(_EVAL_529) == $signed(33'sh0);
  assign _EVAL_375 = _EVAL_217 | _EVAL_48;
  assign _EVAL_614 = _EVAL_30 == _EVAL_109;
  assign _EVAL_571 = _EVAL_614 | _EVAL_1;
  assign _EVAL_201 = _EVAL_14 == 3'h5;
  assign _EVAL_303 = _EVAL_23 ^ 32'h4000;
  assign _EVAL_123 = {1'b0,$signed(_EVAL_303)};
  assign _EVAL_398 = $signed(_EVAL_123) & $signed(-33'sh1000);
  assign _EVAL_82 = $signed(_EVAL_398);
  assign _EVAL_264 = $signed(_EVAL_82) == $signed(33'sh0);
  assign _EVAL_564 = _EVAL_375 | _EVAL_264;
  assign _EVAL_620 = _EVAL_564 | _EVAL_339;
  assign _EVAL_446 = _EVAL_11[3:3];
  assign _EVAL_639 = _EVAL_446 == 1'h0;
  assign _EVAL_618 = _EVAL_11[2:0];
  assign _EVAL_427 = 3'h1 <= _EVAL_618;
  assign _EVAL_592 = _EVAL_639 & _EVAL_427;
  assign _EVAL_580 = _EVAL_14 == 3'h1;
  assign _EVAL_465 = _EVAL_6 & _EVAL_580;
  assign _EVAL_521 = _EVAL_27 != 2'h2;
  assign _EVAL_336 = _EVAL_521 | _EVAL_1;
  assign _EVAL_284 = _EVAL_336 == 1'h0;
  assign _EVAL_242 = _EVAL_6 & _EVAL_473;
  assign _EVAL_148 = _EVAL_7[2:0];
  assign _EVAL_272 = 3'h1 <= _EVAL_148;
  assign _EVAL_420 = _EVAL_29 == 1'h0;
  assign _EVAL_265 = _EVAL_420 | _EVAL_1;
  assign _EVAL_351 = _EVAL_11 == 4'h0;
  assign _EVAL_495 = _EVAL_617 | _EVAL_351;
  assign _EVAL_433 = _EVAL_495 | _EVAL_592;
  assign _EVAL_445 = _EVAL_433 | _EVAL_1;
  assign _EVAL_540 = _EVAL_445 == 1'h0;
  assign _EVAL_414 = _EVAL_17 <= 2'h2;
  assign _EVAL_440 = _EVAL_14 == 3'h4;
  assign _EVAL_352 = _EVAL_6 & _EVAL_440;
  assign _EVAL_77 = _EVAL_24 & _EVAL_520;
  assign _EVAL_207 = _EVAL_24 & _EVAL_670;
  assign _EVAL_411 = _EVAL_236 == 1'h0;
  assign _EVAL_396 = _EVAL_58 == 5'h0;
  assign _EVAL_497 = _EVAL_10[0];
  assign _EVAL_245 = _EVAL_58 - 5'h1;
  assign _EVAL_528 = _EVAL_10 == _EVAL_64;
  assign _EVAL_479 = _EVAL_528 | _EVAL_1;
  assign _EVAL_651 = _EVAL_16 == _EVAL_646;
  assign _EVAL_140 = _EVAL_651 | _EVAL_1;
  assign _EVAL_661 = _EVAL_19 == 3'h3;
  assign _EVAL_181 = _EVAL_19 == 3'h4;
  assign _EVAL_536 = _EVAL_279 == 1'h0;
  assign _EVAL_105 = _EVAL_413 | _EVAL_1;
  assign _EVAL_291 = _EVAL_105 == 1'h0;
  assign _EVAL_332 = _EVAL_14 <= 3'h6;
  assign _EVAL_447 = _EVAL_14 == 3'h2;
  assign _EVAL_278 = _EVAL_6 & _EVAL_447;
  assign _EVAL_463 = _EVAL_19 == 3'h7;
  assign _EVAL_461 = _EVAL_8 & _EVAL_463;
  assign _EVAL_338 = _EVAL_565[0];
  assign _EVAL_525 = _EVAL_338 | _EVAL_1;
  assign _EVAL_407 = _EVAL_4 == _EVAL_257;
  assign _EVAL_192 = _EVAL_407 | _EVAL_1;
  assign _EVAL_458 = _EVAL_547 | _EVAL_1;
  assign _EVAL_160 = _EVAL_126 == 1'h0;
  assign _EVAL_551 = _EVAL_30 <= 3'h4;
  assign _EVAL_599 = _EVAL_551 | _EVAL_1;
  assign _EVAL_415 = _EVAL_599 == 1'h0;
  assign _EVAL_324 = _EVAL_458 == 1'h0;
  assign _EVAL_131 = _EVAL_10 == 3'h7;
  assign _EVAL_335 = ~ _EVAL_88;
  assign _EVAL_556 = _EVAL_479 == 1'h0;
  assign _EVAL_347 = _EVAL_10 == 3'h2;
  assign _EVAL_419 = _EVAL_509 < plusarg_reader_out;
  assign _EVAL_392 = _EVAL_585 | _EVAL_419;
  assign _EVAL_567 = _EVAL_392 | _EVAL_1;
  assign _EVAL_106 = _EVAL_567 == 1'h0;
  assign _EVAL_510 = _EVAL_10 == 3'h1;
  assign _EVAL_654 = _EVAL_414 | _EVAL_1;
  assign _EVAL_372 = _EVAL_654 == 1'h0;
  assign _EVAL_107 = _EVAL_367 & _EVAL_659;
  assign _EVAL_422 = {{24'd0}, _EVAL_562};
  assign _EVAL_633 = _EVAL_4 & _EVAL_422;
  assign _EVAL_535 = _EVAL_633 == 32'h0;
  assign _EVAL_612 = _EVAL_287 | _EVAL_1;
  assign _EVAL_129 = _EVAL_161 | _EVAL_1;
  assign _EVAL_170 = _EVAL_129 == 1'h0;
  assign _EVAL_523 = _EVAL_13 == _EVAL_568;
  assign _EVAL_578 = _EVAL_24 & _EVAL_131;
  assign _EVAL_610 = _EVAL_523 | _EVAL_1;
  assign _EVAL_653 = _EVAL_610 == 1'h0;
  assign _EVAL_326 = _EVAL_10 == 3'h4;
  assign _EVAL_250 = _EVAL_24 & _EVAL_326;
  assign _EVAL_608 = _EVAL_612 == 1'h0;
  assign _EVAL_628 = _EVAL_8 & _EVAL_661;
  assign _EVAL_423 = _EVAL_6 & _EVAL_657;
  assign _EVAL_313 = _EVAL_387 - 5'h1;
  assign _EVAL_203 = _EVAL_15 ? _EVAL_340 : 2'h0;
  assign _EVAL_449 = ~ _EVAL_203;
  assign _EVAL_624 = _EVAL_7 == 4'h0;
  assign _EVAL_430 = _EVAL_624 ? _EVAL_228 : 1'h0;
  assign _EVAL_489 = _EVAL_546 == 1'h0;
  assign _EVAL_476 = _EVAL_226 | _EVAL_1;
  assign _EVAL_117 = _EVAL_476 == 1'h0;
  assign _EVAL_455 = _EVAL_537 | _EVAL_1;
  assign _EVAL_222 = _EVAL_483 | _EVAL_1;
  assign _EVAL_143 = _EVAL_281 | _EVAL_624;
  assign _EVAL_268 = _EVAL_412 == 1'h0;
  assign _EVAL_178 = _EVAL_268 & _EVAL_272;
  assign _EVAL_94 = _EVAL_143 | _EVAL_178;
  assign _EVAL_601 = _EVAL_94 | _EVAL_1;
  assign _EVAL_260 = _EVAL_601 == 1'h0;
  assign _EVAL_545 = 4'h6 == _EVAL_0;
  assign _EVAL_581 = _EVAL_155 ? _EVAL_545 : 1'h0;
  assign _EVAL_197 = _EVAL_581 | _EVAL_1;
  assign _EVAL_457 = _EVAL_396 == 1'h0;
  assign _EVAL_62 = _EVAL_24 & _EVAL_457;
  assign _EVAL_79 = _EVAL_6 & _EVAL_201;
  assign _EVAL_666 = _EVAL_275 | _EVAL_1;
  assign _EVAL_90 = _EVAL_19 == 3'h2;
  assign _EVAL_125 = _EVAL_8 & _EVAL_90;
  assign _EVAL_204 = _EVAL_332 | _EVAL_1;
  assign _EVAL_194 = _EVAL_81 == 1'h0;
  assign _EVAL_328 = _EVAL_542 & _EVAL_335;
  assign _EVAL_306 = _EVAL_662 | _EVAL_586;
  assign _EVAL_315 = _EVAL_455 == 1'h0;
  assign _EVAL_598 = _EVAL_183 == 1'h0;
  assign _EVAL_359 = _EVAL_95 | _EVAL_499;
  assign _EVAL_613 = _EVAL_402 | _EVAL_1;
  assign _EVAL_97 = _EVAL_535 | _EVAL_1;
  assign _EVAL_348 = _EVAL_97 == 1'h0;
  assign _EVAL_669 = _EVAL_666 == 1'h0;
  assign _EVAL_230 = _EVAL_8 & _EVAL_181;
  assign _EVAL_498 = _EVAL_140 == 1'h0;
  assign _EVAL_92 = _EVAL_197 == 1'h0;
  assign _EVAL_519 = _EVAL_525 == 1'h0;
  assign _EVAL_459 = _EVAL_306 | _EVAL_1;
  assign _EVAL_159 = _EVAL_459 == 1'h0;
  assign _EVAL_113 = _EVAL_378 & _EVAL_325;
  assign _EVAL_363 = _EVAL_265 == 1'h0;
  assign _EVAL_346 = _EVAL_87 == 1'h0;
  assign _EVAL_253 = _EVAL_430 | _EVAL_1;
  assign _EVAL_120 = _EVAL_24 & _EVAL_347;
  assign _EVAL_604 = _EVAL_359 & _EVAL_449;
  assign _EVAL_202 = _EVAL_620 | _EVAL_1;
  assign _EVAL_475 = _EVAL_204 == 1'h0;
  assign _EVAL_177 = _EVAL_24 & _EVAL_510;
  assign _EVAL_452 = _EVAL_571 == 1'h0;
  assign _EVAL_200 = _EVAL_202 == 1'h0;
  assign _EVAL_149 = _EVAL_115 & _EVAL_353;
  assign _EVAL_191 = _EVAL_136 == 1'h0;
  assign _EVAL_563 = _EVAL_222 == 1'h0;
  assign _EVAL_164 = _EVAL_533 & _EVAL_396;
  assign _EVAL_67 = _EVAL_253 == 1'h0;
  assign _EVAL_530 = _EVAL_192 == 1'h0;
  assign _EVAL_292 = _EVAL_613 == 1'h0;
  assign _EVAL_478 = _EVAL_500 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_43 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_58 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_70 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_95 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_99 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_109 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_169 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_173 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_187 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_211 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_237 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_257 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_323 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_343 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_387 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_450 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_488 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_491 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_509 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_561 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_568 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_619 = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_622 = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_634 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_636 = _RAND_25[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_646 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_668 = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_25) begin
    if (_EVAL_164) begin
      _EVAL_43 <= _EVAL_7;
    end
    if (_EVAL_1) begin
      _EVAL_58 <= 5'h0;
    end else begin
      if (_EVAL_533) begin
        if (_EVAL_396) begin
          if (_EVAL_497) begin
            _EVAL_58 <= _EVAL_381;
          end else begin
            _EVAL_58 <= 5'h0;
          end
        end else begin
          _EVAL_58 <= _EVAL_245;
        end
      end
    end
    if (_EVAL_164) begin
      _EVAL_64 <= _EVAL_10;
    end
    if (_EVAL_113) begin
      _EVAL_70 <= _EVAL_18;
    end
    if (_EVAL_1) begin
      _EVAL_95 <= 2'h0;
    end else begin
      _EVAL_95 <= _EVAL_604;
    end
    if (_EVAL_113) begin
      _EVAL_99 <= _EVAL_14;
    end
    if (_EVAL_107) begin
      _EVAL_109 <= _EVAL_30;
    end
    if (_EVAL_107) begin
      _EVAL_169 <= _EVAL_0;
    end
    if (_EVAL_107) begin
      _EVAL_173 <= _EVAL_19;
    end
    if (_EVAL_164) begin
      _EVAL_187 <= _EVAL;
    end
    if (_EVAL_1) begin
      _EVAL_211 <= 5'h0;
    end else begin
      if (_EVAL_367) begin
        if (_EVAL_659) begin
          if (_EVAL_492) begin
            _EVAL_211 <= _EVAL_436;
          end else begin
            _EVAL_211 <= 5'h0;
          end
        end else begin
          _EVAL_211 <= _EVAL_247;
        end
      end
    end
    if (_EVAL_107) begin
      _EVAL_237 <= _EVAL_28;
    end
    if (_EVAL_107) begin
      _EVAL_257 <= _EVAL_4;
    end
    if (_EVAL_164) begin
      _EVAL_323 <= _EVAL_31;
    end
    if (_EVAL_149) begin
      _EVAL_343 <= _EVAL_23;
    end
    if (_EVAL_1) begin
      _EVAL_387 <= 5'h0;
    end else begin
      if (_EVAL_378) begin
        if (_EVAL_325) begin
          if (_EVAL_213) begin
            _EVAL_387 <= _EVAL_238;
          end else begin
            _EVAL_387 <= 5'h0;
          end
        end else begin
          _EVAL_387 <= _EVAL_313;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_450 <= 5'h0;
    end else begin
      if (_EVAL_367) begin
        if (_EVAL_174) begin
          if (_EVAL_492) begin
            _EVAL_450 <= _EVAL_436;
          end else begin
            _EVAL_450 <= 5'h0;
          end
        end else begin
          _EVAL_450 <= _EVAL_442;
        end
      end
    end
    if (_EVAL_149) begin
      _EVAL_488 <= _EVAL_17;
    end
    if (_EVAL_113) begin
      _EVAL_491 <= _EVAL_27;
    end
    if (_EVAL_1) begin
      _EVAL_509 <= 32'h0;
    end else begin
      if (_EVAL_231) begin
        _EVAL_509 <= 32'h0;
      end else begin
        _EVAL_509 <= _EVAL_611;
      end
    end
    if (_EVAL_1) begin
      _EVAL_561 <= 5'h0;
    end else begin
      if (_EVAL_378) begin
        if (_EVAL_289) begin
          if (_EVAL_213) begin
            _EVAL_561 <= _EVAL_238;
          end else begin
            _EVAL_561 <= 5'h0;
          end
        end else begin
          _EVAL_561 <= _EVAL_294;
        end
      end
    end
    if (_EVAL_113) begin
      _EVAL_568 <= _EVAL_13;
    end
    if (_EVAL_1) begin
      _EVAL_619 <= 5'h0;
    end else begin
      if (_EVAL_378) begin
        if (_EVAL_40) begin
          if (_EVAL_213) begin
            _EVAL_619 <= _EVAL_238;
          end else begin
            _EVAL_619 <= 5'h0;
          end
        end else begin
          _EVAL_619 <= _EVAL_607;
        end
      end
    end
    if (_EVAL_113) begin
      _EVAL_622 <= _EVAL_11;
    end
    if (_EVAL_1) begin
      _EVAL_634 <= 5'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_353) begin
          _EVAL_634 <= 5'h0;
        end else begin
          _EVAL_634 <= _EVAL_298;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_636 <= 9'h0;
    end else begin
      _EVAL_636 <= _EVAL_328;
    end
    if (_EVAL_113) begin
      _EVAL_646 <= _EVAL_16;
    end
    if (_EVAL_164) begin
      _EVAL_668 <= _EVAL_21;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b823022d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd292967)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_441) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_496 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cf5e85c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35f49693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_540) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50631b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_530) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_536) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_432) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d45a31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e397ea91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_609) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc32cfdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc5ab02f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_441) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39664d0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_522) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adc8fa6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d6ec6d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_519) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af3f9d96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(213faa3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c93409d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_609) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd6897f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46659908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_669) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42240a67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_609) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc99deaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_415) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9d71385)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_536) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9f82b01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41358d3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_556) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab228bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_382) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_498) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e54472)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a82adad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_641) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(865470a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_498) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7bfa46c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a26431f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_536) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e01a8c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39529ffe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_641) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1dfb936)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d7268ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_522) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb26aa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_478) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1560d20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_543) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1c2bb2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_346) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_609) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_598) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b92351)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92c4199d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_346) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88d0145a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a344ed9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_540) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ad9da13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_346) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53d1376e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_540) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b73a62b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_411) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bacb818f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_372) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(814e0328)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1303c48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_540) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2c7719a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1601a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_522) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade3ba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa71e3fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8cacb27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c8b58b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_653) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55294ce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3c4a52c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_653) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e99ed56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68679031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_475) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ffb3f9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f70bcc86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a83c49c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a25c66f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3489e8b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efe45fc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e81073f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dc25373)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92098ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e970b1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6906831c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f340da2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_609) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c4c3768)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_652) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e946274)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_441) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_468) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b15d092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_563) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_477) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64f82939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_522) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2768d659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42f3897f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb1f12ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_432) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55533e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7e963f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a80fe296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bbc41d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c55b7188)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(154a9deb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_540) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a59ac25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_609) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ecb4baf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_475) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a879d53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_522) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(695747f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0914e4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5096735)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_441) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9966346a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6f4aff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_432) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_543) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c0ccb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_608) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cf31ca9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f210d78e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c5eb78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_496 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72ead85c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_382) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90c9da73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(671218e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b977f508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_489) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc7d8f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_669) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c470a22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee5204f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_563) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(253748b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13c4e6c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_468) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df87eb86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_346) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49e234a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_489) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff499e78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9277159)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f67a541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_516) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(953ac23c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4edb33e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bab742ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_415) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9462eb86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_519) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f41a463)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d091301)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_536) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2af4a89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38266bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0c12a06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_372) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9840af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_432) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf449980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d65af737)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_608) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf10615c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cec5fc89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_540) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f30d5df9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_530) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dce1cecc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_609) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1345af5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(708e6a62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dd80080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e4dc12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7f89c17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_411) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e455f60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(774787f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dddeb6c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8b3af4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdeb363e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721d3d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_609) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_477) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_522) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8464716)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d209ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9047aa79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_516) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee4b06b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_478) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e59e437f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
