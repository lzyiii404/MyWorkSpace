//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_185_assert(
  input  [11:0]   _EVAL_20,
  input  [27:0]   _EVAL_51,
  input           _EVAL_58,
  input           _EVAL_59,
  input  [3:0]    _EVAL_69,
  input  [1:0]    _EVAL_79,
  input  [2:0]    _EVAL_86,
  input           _EVAL_105,
  input           _EVAL_131,
  input           _EVAL_142,
  input  [2:0]    _EVAL_143,
  input  [2:0]    _EVAL_663,
  input  [6:0]    _EVAL_3235,
  input  [25:0]   _EVAL_910,
  input           _EVAL_3673,
  input  [1023:0] _EVAL_2999,
  input           _EVAL_2866,
  input           _EVAL_2267,
  input  [31:0]   _EVAL_2124,
  input  [2:0]    _EVAL_3165,
  input           _EVAL_532,
  input           _EVAL_886,
  input           _EVAL_2234,
  input           _EVAL_3059,
  input           _EVAL_2184,
  input           _EVAL_429,
  input           _EVAL_1847,
  input           _EVAL_1531,
  input           _EVAL_1886,
  input           _EVAL_3215,
  input           _EVAL_2610,
  input           _EVAL_3593,
  input           _EVAL_1820,
  input           _EVAL_3152,
  input           _EVAL_2252,
  input           _EVAL_318,
  input           _EVAL_2130,
  input           _EVAL_822,
  input           _EVAL_1515,
  input           _EVAL_2543,
  input           _EVAL_2057,
  input           _EVAL_3820,
  input           _EVAL_2122,
  input           _EVAL_1907,
  input           _EVAL_1328,
  input  [6:0]    _EVAL_1332,
  input           _EVAL_1236,
  input           _EVAL_2001,
  input           _EVAL_829,
  input           _EVAL_1634,
  input           _EVAL_4001,
  input           _EVAL_2940,
  input           _EVAL_3094,
  input           _EVAL_873,
  input           _EVAL_2571,
  input           _EVAL_1201,
  input  [7:0]    _EVAL_638,
  input           _EVAL_938,
  input           _EVAL_2869,
  input           _EVAL_824,
  input           _EVAL_1475,
  input           _EVAL_2835,
  input           _EVAL_2856,
  input           _EVAL_2660,
  input           _EVAL_2713,
  input           _EVAL_2054,
  input           _EVAL_660,
  input           _EVAL_2052,
  input           _EVAL_1355,
  input  [7:0]    _EVAL_3372,
  input           _EVAL_2528,
  input           _EVAL_3594,
  input  [7:0]    _EVAL_695,
  input           _EVAL_2865,
  input           _EVAL_979,
  input           _EVAL_3932,
  input  [7:0]    _EVAL_3055,
  input           _EVAL_3454,
  input           _EVAL_4054,
  input           _EVAL_1944,
  input           _EVAL_3325,
  input           _EVAL_3816,
  input           _EVAL_1533,
  input           _EVAL_3520,
  input           _EVAL_3908,
  input           _EVAL_1107,
  input           _EVAL_985,
  input           _EVAL_3018,
  input           _EVAL_1232,
  input           _EVAL_828,
  input           _EVAL_226,
  input           _EVAL_2048,
  input           _EVAL_845,
  input           _EVAL_3884,
  input           _EVAL_3318,
  input           _EVAL_3508,
  input           _EVAL_3423,
  input  [13:0]   _EVAL_291,
  input           _EVAL_236,
  input           _EVAL_1326,
  input           _EVAL_1337,
  input           _EVAL_1309,
  input           _EVAL_1706,
  input           _EVAL_1548,
  input           _EVAL_2515,
  input           _EVAL_3642,
  input           _EVAL_3679,
  input           _EVAL_3234,
  input           _EVAL_455,
  input           _EVAL_466,
  input           _EVAL_353,
  input           _EVAL_2947,
  input           _EVAL_3628,
  input           _EVAL_2845,
  input           _EVAL_1613,
  input           _EVAL_2825,
  input           _EVAL_851,
  input           _EVAL_3489,
  input           _EVAL_3726,
  input           _EVAL_1880,
  input           _EVAL_3069,
  input           _EVAL_3919,
  input           _EVAL_926,
  input           _EVAL_3043,
  input           _EVAL_415,
  input           _EVAL_265,
  input           _EVAL_1648,
  input           _EVAL_2742,
  input           _EVAL_1230,
  input           _EVAL_2303,
  input           _EVAL_1215,
  input           _EVAL_3088,
  input           _EVAL_2696,
  input  [6:0]    _EVAL_666,
  input           _EVAL_1990,
  input           _EVAL_515,
  input           _EVAL_3117,
  input           _EVAL_1707,
  input           _EVAL_939,
  input           _EVAL_2959,
  input           _EVAL_3744,
  input           _EVAL_3409,
  input           _EVAL_1432,
  input           _EVAL_4041,
  input           _EVAL_4040,
  input           _EVAL_2731,
  input           _EVAL_1064,
  input           _EVAL_1502,
  input           _EVAL_3981,
  input           _EVAL_3873,
  input           _EVAL_1922,
  input           _EVAL_3882,
  input           _EVAL_4062,
  input           _EVAL_3847,
  input           _EVAL_2697,
  input           _EVAL_3707,
  input           _EVAL_2233,
  input           _EVAL_2770,
  input           _EVAL_847,
  input           _EVAL_2567,
  input           _EVAL_2189,
  input           _EVAL_2823,
  input           _EVAL_927,
  input  [126:0]  _EVAL_3572,
  input           _EVAL_1439,
  input           _EVAL_308,
  input           _EVAL_1948,
  input           _EVAL_1235,
  input           _EVAL_1650,
  input           _EVAL_260,
  input           _EVAL_2743,
  input           _EVAL_3682,
  input           _EVAL_2644,
  input           _EVAL_3844,
  input           _EVAL_1957,
  input           _EVAL_3287,
  input           _EVAL_954,
  input           _EVAL_1213,
  input           _EVAL_1216,
  input           _EVAL_612,
  input           _EVAL_3101,
  input           _EVAL_412,
  input           _EVAL_1325,
  input           _EVAL_3350,
  input           _EVAL_3185,
  input           _EVAL_315,
  input           _EVAL_1833,
  input           _EVAL_2097,
  input           _EVAL_2690,
  input           _EVAL_2520,
  input           _EVAL_1013,
  input           _EVAL_1182,
  input           _EVAL_3024,
  input           _EVAL_4009,
  input           _EVAL_691,
  input           _EVAL_2426,
  input           _EVAL_3460,
  input           _EVAL_2302,
  input           _EVAL_1841,
  input           _EVAL_3832,
  input           _EVAL_1400,
  input           _EVAL_3579,
  input           _EVAL_2143,
  input           _EVAL_1240,
  input           _EVAL_3618,
  input           _EVAL_3337,
  input           _EVAL_925,
  input           _EVAL_3213,
  input           _EVAL_667,
  input           _EVAL_1067,
  input           _EVAL_1682,
  input           _EVAL_3539,
  input           _EVAL_3940,
  input           _EVAL_316,
  input           _EVAL_2533,
  input           _EVAL_313,
  input           _EVAL_1225,
  input           _EVAL_295,
  input           _EVAL_1027,
  input           _EVAL_1558,
  input           _EVAL_3064,
  input           _EVAL_1161,
  input           _EVAL_1120,
  input           _EVAL_2608,
  input           _EVAL_1784,
  input           _EVAL_1113,
  input           _EVAL_190,
  input           _EVAL_571,
  input           _EVAL_1655,
  input           _EVAL_815,
  input           _EVAL_1386,
  input           _EVAL_268,
  input           _EVAL_866,
  input           _EVAL_2058,
  input  [126:0]  _EVAL_2527,
  input           _EVAL_3198,
  input           _EVAL_807,
  input           _EVAL_1773,
  input           _EVAL_796,
  input           _EVAL_1205,
  input           _EVAL_3353,
  input           _EVAL_2511,
  input           _EVAL_2903,
  input           _EVAL_3683,
  input           _EVAL_3681,
  input           _EVAL_1015,
  input           _EVAL_1966,
  input           _EVAL_479,
  input           _EVAL_2639,
  input           _EVAL_1472,
  input           _EVAL_3997,
  input           _EVAL_2408,
  input           _EVAL_1178,
  input           _EVAL_2109,
  input           _EVAL_391,
  input           _EVAL_3774,
  input           _EVAL_1311,
  input           _EVAL_2654,
  input           _EVAL_3456,
  input           _EVAL_3842,
  input           _EVAL_1728,
  input           _EVAL_2411,
  input           _EVAL_2015,
  input           _EVAL_2563,
  input           _EVAL_1042,
  input           _EVAL_3650,
  input           _EVAL_3284,
  input           _EVAL_1378,
  input           _EVAL_3214,
  input           _EVAL_3998,
  input           _EVAL_2218,
  input           _EVAL_706,
  input           _EVAL_2099,
  input           _EVAL_541,
  input           _EVAL_1139,
  input           _EVAL_1157,
  input           _EVAL_4061,
  input           _EVAL_3191,
  input           _EVAL_3005,
  input           _EVAL_1461,
  input           _EVAL_1998,
  input           _EVAL_2785,
  input           _EVAL_3669,
  input           _EVAL_1082,
  input           _EVAL_3738,
  input           _EVAL_2603,
  input           _EVAL_1403,
  input           _EVAL_1591,
  input           _EVAL_1510,
  input           _EVAL_3583,
  input           _EVAL_298,
  input           _EVAL_2160,
  input           _EVAL_1187,
  input           _EVAL_3103,
  input           _EVAL_359,
  input           _EVAL_182,
  input           _EVAL_651,
  input           _EVAL_3939,
  input           _EVAL_1663,
  input           _EVAL_3764,
  input           _EVAL_2776,
  input           _EVAL_1446,
  input           _EVAL_1025,
  input           _EVAL_2729,
  input           _EVAL_975,
  input           _EVAL_2439,
  input           _EVAL_2663,
  input           _EVAL_576,
  input           _EVAL_1271,
  input           _EVAL_1842,
  input           _EVAL_2744,
  input           Queue__EVAL_5,
  input           Queue__EVAL_12
);
  wire [2:0] TLMonitor__EVAL;
  wire [2:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire [27:0] TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire [2:0] TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire [1:0] TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire [1:0] TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire [3:0] TLMonitor__EVAL_12;
  wire [11:0] TLMonitor__EVAL_13;
  wire [11:0] TLMonitor__EVAL_14;
  reg  _EVAL_1327;
  reg [31:0] _RAND_0;
  reg [126:0] _EVAL_3531;
  reg [127:0] _RAND_1;
  reg  _EVAL_3861;
  reg [31:0] _RAND_2;
  wire  _EVAL_2645;
  wire  _EVAL_929;
  wire  _EVAL_534;
  wire  _EVAL_3781;
  wire [23:0] _EVAL_2747;
  wire  _EVAL_1249;
  wire  _EVAL_2976;
  wire  _EVAL_1925;
  wire  _EVAL_2558;
  wire  _EVAL_1749;
  wire  _EVAL_843;
  wire  _EVAL_3057;
  wire  _EVAL_367;
  wire  _EVAL_1519;
  wire  _EVAL_974;
  wire [9:0] _EVAL_2638;
  wire [1023:0] _EVAL_1942;
  wire  _EVAL_2990;
  wire  _EVAL_758;
  wire  _EVAL_1381;
  wire  _EVAL_599;
  wire [23:0] _EVAL_3143;
  wire  _EVAL_246;
  wire  _EVAL_1588;
  wire  _EVAL_1647;
  wire  _EVAL_3402;
  wire  _EVAL_3188;
  wire  _EVAL_1300;
  wire  _EVAL_2191;
  wire  _EVAL_3225;
  wire [7:0] _EVAL_1726;
  wire  _EVAL_2817;
  wire [7:0] _EVAL_3261;
  wire  _EVAL_1754;
  wire [7:0] _EVAL_3977;
  wire  _EVAL_779;
  wire [7:0] _EVAL_1379;
  wire [31:0] _EVAL_1377;
  wire [2:0] _EVAL_347;
  wire  _EVAL_1996;
  wire  _EVAL_458;
  wire  _EVAL_3286;
  wire  _EVAL_402;
  wire  _EVAL_2995;
  wire  _EVAL_1545;
  wire  _EVAL_3954;
  wire  _EVAL_948;
  wire  _EVAL_3110;
  wire  _EVAL_911;
  wire  _EVAL_1778;
  wire  _EVAL_3790;
  wire  _EVAL_2551;
  wire  _EVAL_1129;
  wire  _EVAL_889;
  wire  _EVAL_1831;
  wire  _EVAL_1324;
  wire  _EVAL_859;
  wire  _EVAL_1278;
  wire  _EVAL_3154;
  wire  _EVAL_3075;
  wire  _EVAL_3471;
  wire  _EVAL_1252;
  wire  _EVAL_2812;
  wire  _EVAL_3446;
  wire  _EVAL_958;
  wire  _EVAL_3596;
  wire  _EVAL_1806;
  wire  _EVAL_2497;
  wire  _EVAL_905;
  wire  _EVAL_747;
  wire  _EVAL_1307;
  wire  _EVAL_2101;
  wire  _EVAL_1279;
  wire  _EVAL_3194;
  wire  _EVAL_1507;
  wire  _EVAL_3906;
  wire  _EVAL_399;
  wire  _EVAL_1543;
  wire  _EVAL_2961;
  wire  _EVAL_4059;
  wire  _EVAL_3022;
  wire  _EVAL_1605;
  wire  _EVAL_2112;
  wire  _EVAL_806;
  wire  _EVAL_454;
  wire  _EVAL_204;
  wire  _EVAL_1024;
  wire  _EVAL_1275;
  wire  _EVAL_1857;
  wire  _EVAL_3470;
  wire  _EVAL_2674;
  wire  _EVAL_3568;
  wire  _EVAL_3330;
  wire  _EVAL_1470;
  wire  _EVAL_2020;
  wire  _EVAL_2180;
  wire  _EVAL_3652;
  wire  _EVAL_3987;
  wire  _EVAL_2585;
  wire  _EVAL_3901;
  wire  _EVAL_2594;
  wire  _EVAL_2591;
  wire  _EVAL_2219;
  wire  _EVAL_2986;
  wire  _EVAL_1889;
  wire  _EVAL_680;
  wire  _EVAL_4031;
  wire  _EVAL_3812;
  wire  _EVAL_1209;
  wire  _EVAL_998;
  wire  _EVAL_258;
  wire  _EVAL_3238;
  wire  _EVAL_2380;
  wire  _EVAL_827;
  wire  _EVAL_309;
  wire  _EVAL_3558;
  wire  _EVAL_2676;
  wire  _EVAL_1566;
  wire  _EVAL_3207;
  wire  _EVAL_3206;
  wire  _EVAL_1174;
  wire  _EVAL_1643;
  wire  _EVAL_1057;
  wire  _EVAL_1742;
  wire  _EVAL_1417;
  wire  _EVAL_1505;
  wire  _EVAL_1010;
  wire  _EVAL_3048;
  wire  _EVAL_379;
  wire  _EVAL_3377;
  wire  _EVAL_496;
  wire  _EVAL_3889;
  wire  _EVAL_3485;
  wire  _EVAL_2671;
  wire  _EVAL_2650;
  wire  _EVAL_3148;
  wire  _EVAL_3461;
  wire  _EVAL_1497;
  wire  _EVAL_1910;
  wire  _EVAL_508;
  wire  _EVAL_3280;
  wire  _EVAL_2211;
  wire  _EVAL_1681;
  wire  _EVAL_694;
  wire  _EVAL_1180;
  wire  _EVAL_3029;
  wire  _EVAL_183;
  wire  _EVAL_2041;
  wire  _EVAL_1221;
  wire  _EVAL_609;
  wire  _EVAL_2062;
  wire  _EVAL_3621;
  wire  _EVAL_2733;
  wire  _EVAL_1145;
  wire  _EVAL_2583;
  wire  _EVAL_2941;
  wire  _EVAL_2991;
  wire  _EVAL_933;
  wire  _EVAL_692;
  wire  _EVAL_3295;
  wire  _EVAL_2525;
  wire  _EVAL_1638;
  wire  _EVAL_3228;
  wire  _EVAL_3736;
  wire  _EVAL_2319;
  wire  _EVAL_2199;
  wire  _EVAL_743;
  wire  _EVAL_2166;
  wire  _EVAL_1951;
  wire  _EVAL_2685;
  wire  _EVAL_1960;
  wire  _EVAL_3063;
  wire  _EVAL_250;
  wire  _EVAL_1398;
  wire  _EVAL_2699;
  wire  _EVAL_469;
  wire  _EVAL_3562;
  wire  _EVAL_3450;
  wire  _EVAL_431;
  wire  _EVAL_4006;
  wire  _EVAL_804;
  wire  _EVAL_2984;
  wire  _EVAL_2800;
  wire  _EVAL_2091;
  wire  _EVAL_1702;
  wire  _EVAL_2004;
  wire  _EVAL_3272;
  wire  _EVAL_1092;
  wire  _EVAL_3966;
  wire  _EVAL_717;
  wire  _EVAL_3381;
  wire  _EVAL_3856;
  wire  _EVAL_520;
  wire  _EVAL_2794;
  wire  _EVAL_2042;
  wire  _EVAL_1053;
  wire  _EVAL_1383;
  wire  _EVAL_3973;
  wire  _EVAL_1818;
  wire  _EVAL_2501;
  wire  _EVAL_2609;
  wire  _EVAL_3701;
  wire  _EVAL_3196;
  wire  _EVAL_2340;
  wire  _EVAL_3413;
  wire  _EVAL_2978;
  wire  _EVAL_1821;
  wire  _EVAL_2397;
  wire  _EVAL_3897;
  wire  _EVAL_1868;
  wire  _EVAL_649;
  wire  _EVAL_3180;
  wire  _EVAL_3865;
  wire  _EVAL_834;
  wire  _EVAL_3445;
  wire  _EVAL_3458;
  wire  _EVAL_3397;
  wire  _EVAL_2732;
  wire  _EVAL_1744;
  wire  _EVAL_1172;
  wire  _EVAL_3363;
  wire  _EVAL_2263;
  wire  _EVAL_629;
  wire  _EVAL_311;
  wire  _EVAL_266;
  wire  _EVAL_215;
  wire  _EVAL_1695;
  wire  _EVAL_3810;
  wire  _EVAL_4048;
  wire  _EVAL_1724;
  wire  _EVAL_2375;
  wire  _EVAL_3264;
  wire  _EVAL_2339;
  wire  _EVAL_3976;
  wire  _EVAL_1911;
  wire  _EVAL_1335;
  wire  _EVAL_894;
  wire  _EVAL_1862;
  wire  _EVAL_543;
  wire  _EVAL_2266;
  wire  _EVAL_3035;
  wire  _EVAL_1553;
  wire  _EVAL_3779;
  wire  _EVAL_2668;
  wire  _EVAL_3869;
  wire  _EVAL_1894;
  wire  _EVAL_1504;
  wire  _EVAL_2053;
  wire  _EVAL_1476;
  wire  _EVAL_1689;
  wire  _EVAL_356;
  wire  _EVAL_699;
  wire  _EVAL_2445;
  wire  _EVAL_2798;
  wire  _EVAL_1245;
  wire  _EVAL_1775;
  wire  _EVAL_2105;
  wire  _EVAL_3664;
  wire  _EVAL_1666;
  wire [7:0] _EVAL_1045;
  wire  _EVAL_2544;
  wire  _EVAL_1047;
  wire  _EVAL_1040;
  wire  _EVAL_1567;
  wire  _EVAL_2712;
  wire  _EVAL_2560;
  wire  _EVAL_2649;
  wire  _EVAL_2423;
  wire  _EVAL_3104;
  wire  _EVAL_3557;
  wire  _EVAL_2173;
  wire [7:0] _EVAL_1371;
  wire  _EVAL_2283;
  wire  _EVAL_1459;
  wire  _EVAL_1179;
  wire  _EVAL_321;
  wire  _EVAL_3298;
  wire  _EVAL_818;
  wire  _EVAL_637;
  wire  _EVAL_2151;
  wire  _EVAL_1207;
  wire  _EVAL_3376;
  wire  _EVAL_1228;
  wire  _EVAL_4049;
  wire  _EVAL_3093;
  wire  _EVAL_2824;
  wire  _EVAL_721;
  wire  _EVAL_1903;
  wire  _EVAL_2815;
  wire  _EVAL_897;
  wire  _EVAL_611;
  wire  _EVAL_2027;
  wire  _EVAL_1354;
  wire  _EVAL_327;
  wire  _EVAL_3516;
  wire  _EVAL_2179;
  wire  _EVAL_1034;
  wire  _EVAL_1224;
  wire  _EVAL_471;
  wire  _EVAL_2621;
  wire  _EVAL_1522;
  wire  _EVAL_2691;
  wire  _EVAL_1012;
  wire  _EVAL_914;
  wire  _EVAL_3270;
  wire  _EVAL_3000;
  wire  _EVAL_2617;
  wire  _EVAL_966;
  wire  _EVAL_1901;
  wire  _EVAL_477;
  wire  _EVAL_1005;
  wire  _EVAL_3503;
  wire  _EVAL_1078;
  wire  _EVAL_3693;
  wire  _EVAL_980;
  wire  _EVAL_3347;
  wire  _EVAL_919;
  wire  _EVAL_756;
  wire  _EVAL_4019;
  wire  _EVAL_403;
  wire  _EVAL_530;
  wire  _EVAL_2775;
  wire  _EVAL_3795;
  wire  _EVAL_825;
  wire  _EVAL_1079;
  wire  _EVAL_4016;
  wire  _EVAL_1041;
  wire  _EVAL_152;
  wire  _EVAL_3391;
  wire  _EVAL_1735;
  wire  _EVAL_1295;
  wire  _EVAL_4069;
  wire  _EVAL_1701;
  wire  _EVAL_790;
  wire  _EVAL_957;
  wire  _EVAL_2804;
  wire  _EVAL_2072;
  wire  _EVAL_3322;
  wire  _EVAL_1989;
  wire  _EVAL_669;
  wire  _EVAL_3248;
  wire  _EVAL_868;
  wire  _EVAL_3218;
  wire  _EVAL_2369;
  wire  _EVAL_1372;
  wire  _EVAL_1834;
  wire  _EVAL_3140;
  wire  _EVAL_2756;
  wire  _EVAL_3561;
  wire  _EVAL_2083;
  wire  _EVAL_535;
  wire  _EVAL_1048;
  wire  _EVAL_1044;
  wire  _EVAL_3246;
  wire  _EVAL_2996;
  wire  _EVAL_518;
  wire  _EVAL_3163;
  wire  _EVAL_3472;
  wire  _EVAL_3285;
  wire  _EVAL_3455;
  wire  _EVAL_662;
  wire  _EVAL_3914;
  wire  _EVAL_884;
  wire  _EVAL_2241;
  wire  _EVAL_2556;
  wire  _EVAL_392;
  wire  _EVAL_1621;
  wire  _EVAL_1396;
  wire  _EVAL_3468;
  wire  _EVAL_2683;
  wire  _EVAL_2043;
  wire  _EVAL_3988;
  wire  _EVAL_3278;
  wire  _EVAL_551;
  wire  _EVAL_2736;
  wire  _EVAL_858;
  wire  _EVAL_1277;
  wire  _EVAL_755;
  wire  _EVAL_2962;
  wire  _EVAL_2305;
  wire  _EVAL_3927;
  wire  _EVAL_916;
  wire  _EVAL_1645;
  wire  _EVAL_4033;
  wire  _EVAL_2614;
  wire  _EVAL_3770;
  wire  _EVAL_3229;
  wire  _EVAL_3241;
  wire  _EVAL_3537;
  wire  _EVAL_3051;
  wire  _EVAL_3575;
  wire  _EVAL_1629;
  wire  _EVAL_1166;
  wire  _EVAL_3062;
  wire  _EVAL_2273;
  wire  _EVAL_2450;
  wire  _EVAL_302;
  wire  _EVAL_2914;
  wire  _EVAL_1542;
  wire  _EVAL_2980;
  wire  _EVAL_3767;
  wire  _EVAL_3821;
  wire  _EVAL_3352;
  wire  _EVAL_655;
  wire  _EVAL_3937;
  wire  _EVAL_400;
  wire  _EVAL_1490;
  wire  _EVAL_764;
  wire  _EVAL_2195;
  wire  _EVAL_801;
  wire  _EVAL_1143;
  wire  _EVAL_2012;
  wire  _EVAL_2108;
  wire  _EVAL_2808;
  wire  _EVAL_2442;
  wire  _EVAL_3405;
  wire  _EVAL_2943;
  wire  _EVAL_411;
  wire  _EVAL_3394;
  wire  _EVAL_3678;
  wire  _EVAL_2665;
  wire  _EVAL_3974;
  wire  _EVAL_3969;
  wire  _EVAL_2078;
  wire  _EVAL_941;
  wire  _EVAL_2874;
  wire  _EVAL_3249;
  wire  _EVAL_2613;
  wire  _EVAL_264;
  wire  _EVAL_1940;
  wire  _EVAL_1947;
  wire  _EVAL_3145;
  wire  _EVAL_1670;
  wire  _EVAL_1823;
  wire  _EVAL_2249;
  wire  _EVAL_1524;
  wire  _EVAL_2285;
  wire  _EVAL_424;
  wire  _EVAL_646;
  wire  _EVAL_2830;
  wire  _EVAL_984;
  wire  _EVAL_3746;
  wire  _EVAL_2960;
  wire  _EVAL_1054;
  wire  _EVAL_4012;
  wire  _EVAL_3369;
  wire  _EVAL_1885;
  wire [28:0] _EVAL_639;
  wire  _EVAL_2470;
  wire  _EVAL_1631;
  wire  _EVAL_1423;
  wire  _EVAL_856;
  wire  _EVAL_819;
  wire  _EVAL_289;
  wire  _EVAL_2605;
  wire  _EVAL_405;
  wire  _EVAL_1860;
  wire  _EVAL_2489;
  wire  _EVAL_2702;
  wire  _EVAL_3835;
  wire  _EVAL_1969;
  wire  _EVAL_1982;
  wire  _EVAL_1102;
  wire  _EVAL_2465;
  wire  _EVAL_909;
  wire  _EVAL_1686;
  wire  _EVAL_1854;
  wire  _EVAL_478;
  wire  _EVAL_1258;
  wire  _EVAL_546;
  wire  _EVAL_1017;
  wire  _EVAL_3171;
  wire  _EVAL_3054;
  wire  _EVAL_633;
  wire  _EVAL_3818;
  wire  _EVAL_234;
  wire  _EVAL_202;
  wire  _EVAL_2398;
  wire  _EVAL_3001;
  wire  _EVAL_876;
  wire  _EVAL_2873;
  wire  _EVAL_2383;
  wire  _EVAL_2276;
  wire  _EVAL_2030;
  wire [6:0] _EVAL_1119;
  wire  _EVAL_3953;
  wire  _EVAL_3716;
  wire  _EVAL_1404;
  wire  _EVAL_2433;
  wire  _EVAL_3230;
  wire  _EVAL_3782;
  wire  _EVAL_2009;
  wire  _EVAL_3619;
  wire  _EVAL_1481;
  wire  _EVAL_522;
  wire  _EVAL_1642;
  wire  _EVAL_1595;
  wire  _EVAL_1809;
  wire  _EVAL_969;
  wire  _EVAL_661;
  wire  _EVAL_1026;
  wire  _EVAL_848;
  wire  _EVAL_2724;
  wire  _EVAL_2541;
  wire  _EVAL_523;
  wire  _EVAL_2622;
  wire  _EVAL_2693;
  wire  _EVAL_2993;
  wire  _EVAL_169;
  wire  _EVAL_2201;
  wire  _EVAL_554;
  wire  _EVAL_3616;
  wire  _EVAL_3528;
  wire  _EVAL_465;
  wire  _EVAL_2401;
  wire  _EVAL_978;
  wire  _EVAL_3190;
  wire  _EVAL_3653;
  wire  _EVAL_3119;
  wire  _EVAL_1781;
  wire  _EVAL_598;
  wire  _EVAL_3699;
  wire  _EVAL_2954;
  wire  _EVAL_2611;
  wire  _EVAL_3807;
  wire  _EVAL_3052;
  wire  _EVAL_1203;
  wire  _EVAL_1761;
  wire  _EVAL_1620;
  wire  _EVAL_1103;
  wire  _EVAL_3648;
  wire  _EVAL_2658;
  wire  _EVAL_1004;
  wire  _EVAL_3328;
  wire  _EVAL_2194;
  wire  _EVAL_536;
  wire  _EVAL_3462;
  wire  _EVAL_241;
  wire  _EVAL_724;
  wire  _EVAL_3481;
  wire  _EVAL_3574;
  wire  _EVAL_418;
  wire  _EVAL_2985;
  wire  _EVAL_3071;
  wire  _EVAL_2741;
  wire  _EVAL_3320;
  wire  _EVAL_1534;
  wire  _EVAL_2420;
  wire  _EVAL_1923;
  wire  _EVAL_1128;
  wire  _EVAL_3411;
  wire  _EVAL_1950;
  wire  _EVAL_1106;
  wire  _EVAL_1431;
  wire  _EVAL_168;
  wire  _EVAL_3613;
  wire  _EVAL_3827;
  wire  _EVAL_336;
  wire  _EVAL_3933;
  wire  _EVAL_2805;
  wire  _EVAL_1405;
  wire  _EVAL_1099;
  wire  _EVAL_2176;
  wire  _EVAL_2979;
  wire  _EVAL_3960;
  wire  _EVAL_2181;
  wire  _EVAL_181;
  wire  _EVAL_1884;
  wire  _EVAL_2647;
  wire  _EVAL_2386;
  wire  _EVAL_2951;
  wire  _EVAL_872;
  wire  _EVAL_3345;
  wire  _EVAL_1369;
  wire  _EVAL_772;
  wire  _EVAL_1920;
  wire  _EVAL_778;
  wire  _EVAL_1872;
  wire  _EVAL_3789;
  wire  _EVAL_3151;
  wire [3:0] _EVAL_3406;
  wire  _EVAL_813;
  wire  _EVAL_1791;
  wire  _EVAL_357;
  wire  _EVAL_365;
  wire  _EVAL_814;
  wire  _EVAL_935;
  wire  _EVAL_2182;
  wire  _EVAL_2016;
  wire  _EVAL_3438;
  wire  _EVAL_2373;
  wire  _EVAL_2284;
  wire  _EVAL_145;
  wire  _EVAL_992;
  wire  _EVAL_977;
  wire  _EVAL_255;
  wire  _EVAL_2778;
  wire  _EVAL_2259;
  wire  _EVAL_3848;
  wire  _EVAL_297;
  wire  _EVAL_2205;
  wire  _EVAL_2342;
  wire  _EVAL_475;
  wire  _EVAL_1581;
  wire  _EVAL_2587;
  wire  _EVAL_404;
  wire  _EVAL_3210;
  wire  _EVAL_3087;
  wire  _EVAL_3656;
  wire  _EVAL_3565;
  wire  _EVAL_1140;
  wire  _EVAL_2253;
  wire  _EVAL_1110;
  wire  _EVAL_3511;
  wire  _EVAL_949;
  wire  _EVAL_2923;
  wire  _EVAL_2376;
  wire  _EVAL_2506;
  wire  _EVAL_3514;
  wire  _EVAL_567;
  wire  _EVAL_2831;
  wire  _EVAL_3829;
  wire  _EVAL_3120;
  wire  _EVAL_697;
  wire  _EVAL_1976;
  wire  _EVAL_1544;
  wire  _EVAL_4023;
  wire  _EVAL_384;
  wire  _EVAL_1192;
  wire  _EVAL_210;
  wire  _EVAL_3016;
  wire  _EVAL_863;
  wire  _EVAL_300;
  wire  _EVAL_1921;
  wire  _EVAL_3067;
  wire  _EVAL_3173;
  wire  _EVAL_3717;
  wire  _EVAL_3542;
  wire  _EVAL_2780;
  wire  _EVAL_568;
  wire  _EVAL_3332;
  wire  _EVAL_2755;
  wire  _EVAL_2294;
  wire  _EVAL_1420;
  wire  _EVAL_3036;
  wire  _EVAL_2332;
  wire  _EVAL_2922;
  wire  _EVAL_2322;
  wire  _EVAL_953;
  wire  _EVAL_2413;
  wire  _EVAL_2657;
  wire  _EVAL_1867;
  wire  _EVAL_3894;
  wire  _EVAL_1514;
  wire  _EVAL_3611;
  wire  _EVAL_3387;
  wire  _EVAL_2620;
  wire  _EVAL_1963;
  wire  _EVAL_2829;
  wire  _EVAL_1897;
  wire  _EVAL_3079;
  wire  _EVAL_2395;
  wire  _EVAL_2337;
  wire  _EVAL_3530;
  wire  _EVAL_3306;
  wire  _EVAL_3451;
  wire  _EVAL_2258;
  wire  _EVAL_2162;
  wire  _EVAL_2402;
  wire  _EVAL_3949;
  wire  _EVAL_3378;
  wire  _EVAL_3725;
  wire  _EVAL_1191;
  wire  _EVAL_2694;
  wire  _EVAL_2498;
  wire  _EVAL_3339;
  wire  _EVAL_330;
  wire  _EVAL_2906;
  wire  _EVAL_3038;
  wire  _EVAL_2632;
  wire  _EVAL_1683;
  wire  _EVAL_3599;
  wire  _EVAL_3934;
  wire  _EVAL_2293;
  wire  _EVAL_728;
  wire  _EVAL_2580;
  wire  _EVAL_767;
  wire  _EVAL_1575;
  wire  _EVAL_1312;
  wire  _EVAL_504;
  wire  _EVAL_883;
  wire  _EVAL_2530;
  wire  _EVAL_1745;
  wire  _EVAL_1836;
  wire  _EVAL_3208;
  wire  _EVAL_960;
  wire  _EVAL_243;
  wire  _EVAL_358;
  wire  _EVAL_3141;
  wire  _EVAL_2444;
  wire  _EVAL_2792;
  wire  _EVAL_2061;
  wire  _EVAL_2516;
  wire  _EVAL_3095;
  wire  _EVAL_474;
  wire  _EVAL_2711;
  wire  _EVAL_1609;
  wire  _EVAL_2576;
  wire  _EVAL_547;
  wire  _EVAL_1937;
  wire  _EVAL_3806;
  wire  _EVAL_470;
  wire  _EVAL_685;
  wire  _EVAL_3836;
  wire  _EVAL_566;
  wire  _EVAL_784;
  wire  _EVAL_3319;
  wire  _EVAL_1491;
  wire  _EVAL_279;
  wire  _EVAL_656;
  wire  _EVAL_4065;
  wire  _EVAL_2667;
  wire  _EVAL_2636;
  wire  _EVAL_3735;
  wire  _EVAL_696;
  wire  _EVAL_1484;
  wire  _EVAL_2331;
  wire  _EVAL_2196;
  wire  _EVAL_3737;
  wire  _EVAL_1322;
  wire  _EVAL_3440;
  wire  _EVAL_657;
  wire  _EVAL_1618;
  wire  _EVAL_1800;
  wire  _EVAL_2040;
  wire  _EVAL_3441;
  wire  _EVAL_1016;
  wire  _EVAL_686;
  wire  _EVAL_1895;
  wire  _EVAL_3408;
  wire  _EVAL_1766;
  wire  _EVAL_887;
  wire  _EVAL_2087;
  wire  _EVAL_849;
  wire  _EVAL_2726;
  wire  _EVAL_3968;
  wire  _EVAL_498;
  wire  _EVAL_3982;
  wire  _EVAL_1415;
  wire  _EVAL_1817;
  wire  _EVAL_3480;
  wire  _EVAL_3771;
  wire  _EVAL_2044;
  wire  _EVAL_3845;
  wire  _EVAL_2326;
  wire  _EVAL_1426;
  wire  _EVAL_1310;
  wire  _EVAL_1949;
  wire  _EVAL_2757;
  wire  _EVAL_1636;
  wire  _EVAL_763;
  wire  _EVAL_999;
  wire  _EVAL_3326;
  wire  _EVAL_869;
  wire  _EVAL_3162;
  wire  _EVAL_1263;
  wire  _EVAL_3366;
  wire  _EVAL_2348;
  wire  _EVAL_2379;
  wire  _EVAL_332;
  wire  _EVAL_499;
  wire  _EVAL_1538;
  wire  _EVAL_3257;
  wire  _EVAL_3209;
  wire  _EVAL_2740;
  wire  _EVAL_1705;
  wire  _EVAL_2396;
  wire  _EVAL_494;
  wire  _EVAL_3805;
  wire  _EVAL_1829;
  wire  _EVAL_3730;
  wire  _EVAL_2706;
  wire  _EVAL_501;
  wire  _EVAL_2820;
  wire  _EVAL_3582;
  wire  _EVAL_1748;
  wire  _EVAL_550;
  wire  _EVAL_432;
  wire  _EVAL_179;
  wire  _EVAL_198;
  wire  _EVAL_1577;
  wire  _EVAL_3876;
  wire  _EVAL_398;
  wire  _EVAL_3368;
  wire  _EVAL_324;
  wire  _EVAL_3791;
  wire  _EVAL_4035;
  wire  _EVAL_284;
  wire  _EVAL_2928;
  wire  _EVAL_2221;
  wire  _EVAL_1883;
  wire  _EVAL_904;
  wire  _EVAL_340;
  wire  _EVAL_2145;
  wire  _EVAL_3631;
  wire  _EVAL_3697;
  wire  _EVAL_440;
  wire  _EVAL_687;
  wire  _EVAL_635;
  wire  _EVAL_2236;
  wire  _EVAL_2508;
  wire  _EVAL_2363;
  wire  _EVAL_3189;
  wire  _EVAL_3633;
  wire  _EVAL_931;
  wire  _EVAL_442;
  wire  _EVAL_1455;
  wire  _EVAL_319;
  wire  _EVAL_538;
  wire  _EVAL_2540;
  wire  _EVAL_1792;
  wire  _EVAL_3294;
  wire  _EVAL_2407;
  wire  _EVAL_1983;
  wire  _EVAL_719;
  wire  _EVAL_564;
  wire  _EVAL_1155;
  wire  _EVAL_1248;
  wire  _EVAL_2403;
  wire  _EVAL_1935;
  wire  _EVAL_232;
  wire  _EVAL_3872;
  wire  _EVAL_2203;
  wire  _EVAL_2086;
  wire  _EVAL_2534;
  wire  _EVAL_2836;
  wire  _EVAL_2679;
  wire  _EVAL_920;
  wire  _EVAL_2412;
  wire  _EVAL_1715;
  wire  _EVAL_3742;
  wire  _EVAL_1089;
  wire  _EVAL_752;
  wire  _EVAL_3217;
  wire  _EVAL_2428;
  wire  _EVAL_2522;
  wire  _EVAL_3702;
  wire  _EVAL_2859;
  wire  _EVAL_1814;
  wire  _EVAL_2783;
  wire  _EVAL_2547;
  wire  _EVAL_328;
  wire  _EVAL_3819;
  wire  _EVAL_1437;
  wire  _EVAL_3089;
  wire  _EVAL_500;
  wire  _EVAL_1926;
  wire  _EVAL_211;
  wire  _EVAL_2721;
  wire  _EVAL_823;
  wire  _EVAL_1274;
  wire  _EVAL_1813;
  wire  _EVAL_3290;
  wire  _EVAL_388;
  wire  _EVAL_2577;
  wire  _EVAL_3467;
  wire  _EVAL_1188;
  wire  _EVAL_2029;
  wire  _EVAL_1314;
  wire  _EVAL_892;
  wire  _EVAL_2021;
  wire  _EVAL_446;
  wire  _EVAL_2323;
  wire  _EVAL_3935;
  wire  _EVAL_1612;
  wire  _EVAL_413;
  wire  _EVAL_2919;
  wire  _EVAL_2793;
  wire  _EVAL_2884;
  wire  _EVAL_2795;
  wire  _EVAL_1561;
  wire  _EVAL_2643;
  wire  _EVAL_3863;
  wire  _EVAL_3962;
  wire  _EVAL_3643;
  wire  _EVAL_3501;
  wire  _EVAL_3684;
  wire  _EVAL_575;
  wire  _EVAL_1464;
  wire  _EVAL_3797;
  wire  _EVAL_1409;
  wire  _EVAL_2419;
  wire  _EVAL_3634;
  wire  _EVAL_333;
  wire  _EVAL_2080;
  wire  _EVAL_1743;
  wire  _EVAL_3809;
  wire  _EVAL_1729;
  wire  _EVAL_2393;
  wire  _EVAL_1480;
  wire  _EVAL_1616;
  wire  _EVAL_3512;
  wire  _EVAL_1029;
  wire  _EVAL_451;
  wire  _EVAL_2846;
  wire  _EVAL_1554;
  wire  _EVAL_705;
  wire  _EVAL_2357;
  wire  _EVAL_1169;
  wire  _EVAL_882;
  wire  _EVAL_2260;
  wire  _EVAL_1560;
  wire  _EVAL_1646;
  wire  _EVAL_3696;
  wire  _EVAL_3833;
  wire  _EVAL_2344;
  wire  _EVAL_1563;
  wire  _EVAL_2933;
  wire  _EVAL_1869;
  wire  _EVAL_1340;
  wire  _EVAL_1395;
  wire  _EVAL_597;
  wire  _EVAL_934;
  wire  _EVAL_3449;
  wire  _EVAL_3427;
  wire  _EVAL_1846;
  wire  _EVAL_2469;
  wire  _EVAL_776;
  wire  _EVAL_1782;
  wire  _EVAL_3761;
  wire  _EVAL_2452;
  wire  _EVAL_2949;
  wire  _EVAL_1523;
  wire  _EVAL_468;
  wire  _EVAL_1331;
  wire  _EVAL_2901;
  wire  _EVAL_1183;
  wire  _EVAL_997;
  wire  _EVAL_3849;
  wire  _EVAL_3333;
  wire  _EVAL_3685;
  wire  _EVAL_435;
  wire  _EVAL_1688;
  wire  _EVAL_3032;
  wire  _EVAL_740;
  wire  _EVAL_2871;
  wire  _EVAL_1812;
  wire  _EVAL_1787;
  wire  _EVAL_3980;
  wire  _EVAL_2689;
  wire  _EVAL_1152;
  wire  _EVAL_1871;
  wire  _EVAL_2247;
  wire  _EVAL_3128;
  wire  _EVAL_2641;
  wire  _EVAL_1589;
  wire  _EVAL_1691;
  wire [7:0] _EVAL_2900;
  wire  _EVAL_2456;
  wire  _EVAL_1296;
  wire  _EVAL_1158;
  wire  _EVAL_2240;
  wire  _EVAL_2891;
  wire  _EVAL_1457;
  wire  _EVAL_1153;
  wire  _EVAL_526;
  wire  _EVAL_2457;
  wire  _EVAL_2606;
  wire  _EVAL_1084;
  wire  _EVAL_3691;
  wire  _EVAL_3920;
  wire  _EVAL_4000;
  wire  _EVAL_1603;
  wire  _EVAL_3153;
  wire  _EVAL_1630;
  wire  _EVAL_3963;
  wire  _EVAL_1330;
  wire  _EVAL_1281;
  wire  _EVAL_393;
  wire  _EVAL_3417;
  wire  _EVAL_1576;
  wire  _EVAL_4060;
  wire  _EVAL_3524;
  wire  _EVAL_3395;
  wire  _EVAL_3635;
  wire  _EVAL_678;
  wire  _EVAL_166;
  wire  _EVAL_184;
  wire  _EVAL_803;
  wire  _EVAL_2618;
  wire  _EVAL_965;
  wire  _EVAL_175;
  wire  _EVAL_3986;
  wire  _EVAL_1091;
  wire  _EVAL_1694;
  wire  _EVAL_2945;
  wire  _EVAL_3600;
  wire  _EVAL_1445;
  wire  _EVAL_2483;
  wire  _EVAL_1624;
  wire  _EVAL_3654;
  wire  _EVAL_2280;
  wire  _EVAL_2161;
  wire  _EVAL_810;
  wire  _EVAL_2765;
  wire  _EVAL_3116;
  wire  _EVAL_2862;
  wire  _EVAL_1086;
  wire  _EVAL_3068;
  wire  _EVAL_3342;
  wire  _EVAL_2983;
  wire  _EVAL_952;
  wire  _EVAL_3310;
  wire  _EVAL_3754;
  wire  _EVAL_3304;
  wire  _EVAL_205;
  wire  _EVAL_3924;
  wire  _EVAL_3532;
  wire  _EVAL_385;
  wire  _EVAL_502;
  wire  _EVAL_4024;
  wire  _EVAL_1967;
  wire  _EVAL_2904;
  wire  _EVAL_3027;
  wire  _EVAL_1661;
  wire  _EVAL_670;
  wire  _EVAL_2372;
  wire  _EVAL_223;
  wire  _EVAL_256;
  wire  _EVAL_2272;
  wire  _EVAL_2127;
  wire  _EVAL_216;
  wire  _EVAL_3958;
  wire  _EVAL_3164;
  wire  _EVAL_3985;
  wire  _EVAL_3877;
  wire  _EVAL_2566;
  wire  _EVAL_2599;
  wire  _EVAL_1692;
  wire  _EVAL_4046;
  wire  _EVAL_744;
  wire  _EVAL_2974;
  wire  _EVAL_441;
  wire  _EVAL_1840;
  wire  _EVAL_1382;
  wire  _EVAL_1083;
  wire  _EVAL_3763;
  wire  _EVAL_1125;
  wire  _EVAL_3597;
  wire  _EVAL_3121;
  wire  _EVAL_2879;
  wire  _EVAL_3555;
  wire  _EVAL_3487;
  wire  _EVAL_2692;
  wire  _EVAL_290;
  wire  _EVAL_344;
  wire  _EVAL_2505;
  wire  _EVAL_1664;
  wire  _EVAL_2034;
  wire  _EVAL_967;
  wire  _EVAL_2637;
  wire  _EVAL_1530;
  wire  _EVAL_1043;
  wire  _EVAL_2230;
  wire  _EVAL_3479;
  wire  _EVAL_3989;
  wire  _EVAL_2493;
  wire  _EVAL_665;
  wire  _EVAL_3601;
  wire  _EVAL_1499;
  wire  _EVAL_874;
  wire  _EVAL_857;
  wire  _EVAL_877;
  wire  _EVAL_1060;
  wire  _EVAL_3838;
  wire  _EVAL_483;
  wire  _EVAL_936;
  wire  _EVAL_1316;
  wire  _EVAL_4071;
  wire  _EVAL_4004;
  wire  _EVAL_777;
  wire  _EVAL_3676;
  wire  _EVAL_2725;
  wire  _EVAL_1447;
  wire  _EVAL_1000;
  wire  _EVAL_2837;
  wire  _EVAL_982;
  wire  _EVAL_2834;
  wire  _EVAL_1532;
  wire  _EVAL_3639;
  wire  _EVAL_3176;
  wire  _EVAL_1375;
  wire  _EVAL_3144;
  wire  _EVAL_3891;
  wire  _EVAL_1822;
  wire  _EVAL_4022;
  wire  _EVAL_2138;
  wire  _EVAL_3694;
  wire  _EVAL_2014;
  wire  _EVAL_668;
  wire  _EVAL_3871;
  wire  _EVAL_3917;
  wire  _EVAL_164;
  wire  _EVAL_3367;
  wire  _EVAL_766;
  wire  _EVAL_2596;
  wire  _EVAL_2359;
  wire  _EVAL_1364;
  wire  _EVAL_3482;
  wire  _EVAL_1401;
  wire  _EVAL_2681;
  wire  _EVAL_3092;
  wire  _EVAL_702;
  wire  _EVAL_2400;
  wire  _EVAL_196;
  wire  _EVAL_3692;
  wire  _EVAL_1358;
  wire  _EVAL_275;
  wire  _EVAL_1022;
  wire  _EVAL_4037;
  wire  _EVAL_1116;
  wire  _EVAL_1319;
  wire  _EVAL_2312;
  wire  _EVAL_3517;
  wire  _EVAL_1049;
  wire  _EVAL_1031;
  wire  _EVAL_153;
  wire  _EVAL_2264;
  wire  _EVAL_3610;
  wire  _EVAL_2769;
  wire  _EVAL_337;
  wire  _EVAL_2569;
  wire  _EVAL_2759;
  wire  _EVAL_484;
  wire  _EVAL_3885;
  wire  _EVAL_1653;
  wire  _EVAL_3834;
  wire  _EVAL_1755;
  wire  _EVAL_558;
  wire  _EVAL_1912;
  wire  _EVAL_2250;
  wire  _EVAL_1384;
  wire  _EVAL_1065;
  wire  _EVAL_1997;
  wire  _EVAL_544;
  wire  _EVAL_2275;
  wire  _EVAL_991;
  wire  _EVAL_903;
  wire  _EVAL_3496;
  wire  _EVAL_1098;
  wire  _EVAL_3313;
  wire  _EVAL_1961;
  wire  _EVAL_3327;
  wire  _EVAL_1652;
  wire  _EVAL_1659;
  wire  _EVAL_3375;
  wire  _EVAL_3777;
  wire  _EVAL_2855;
  wire  _EVAL_1001;
  wire  _EVAL_2678;
  wire  _EVAL_2630;
  wire  _EVAL_2488;
  wire  _EVAL_1941;
  wire  _EVAL_2753;
  wire  _EVAL_3931;
  wire  _EVAL_456;
  wire  _EVAL_654;
  wire  _EVAL_785;
  wire  _EVAL_2154;
  wire  _EVAL_2992;
  wire  _EVAL_1759;
  wire  _EVAL_3580;
  wire  _EVAL_3392;
  wire  _EVAL_2212;
  wire  _EVAL_789;
  wire  _EVAL_3085;
  wire  _EVAL_783;
  wire  _EVAL_2546;
  wire  _EVAL_3197;
  wire  _EVAL_2039;
  wire  _EVAL_2387;
  wire  _EVAL_2816;
  wire  _EVAL_2069;
  wire  _EVAL_3598;
  wire  _EVAL_2570;
  wire  _EVAL_3212;
  wire  _EVAL_3253;
  wire  _EVAL_2352;
  wire  _EVAL_1428;
  wire  _EVAL_3124;
  wire  _EVAL_3672;
  wire  _EVAL_1964;
  wire  _EVAL_1747;
  wire  _EVAL_1039;
  wire  _EVAL_642;
  wire  _EVAL_2672;
  wire  _EVAL_3567;
  wire  _EVAL_630;
  wire  _EVAL_895;
  wire  _EVAL_3983;
  wire  _EVAL_2406;
  wire  _EVAL_453;
  wire  _EVAL_1105;
  wire  _EVAL_1828;
  wire  _EVAL_1233;
  wire  _EVAL_853;
  wire  _EVAL_2292;
  wire  _EVAL_2695;
  wire  _EVAL_3255;
  wire  _EVAL_2822;
  wire  _EVAL_170;
  wire  _EVAL_3031;
  wire  _EVAL_2512;
  wire  _EVAL_2887;
  wire  _EVAL_2200;
  wire  _EVAL_2222;
  wire  _EVAL_2924;
  wire  _EVAL_1975;
  wire  _EVAL_3170;
  wire  _EVAL_3967;
  wire  _EVAL_738;
  wire  _EVAL_3498;
  wire  _EVAL_2604;
  wire  _EVAL_2437;
  wire  _EVAL_3904;
  wire  _EVAL_2478;
  wire  _EVAL_3019;
  wire  _EVAL_463;
  wire  _EVAL_1493;
  wire  _EVAL_156;
  wire  _EVAL_3341;
  wire  _EVAL_2239;
  wire  _EVAL_3237;
  wire  _EVAL_3506;
  wire  _EVAL_924;
  wire  _EVAL_506;
  wire  _EVAL_305;
  wire  _EVAL_3132;
  wire  _EVAL_1900;
  wire  _EVAL_3346;
  wire  _EVAL_1334;
  wire  _EVAL_3668;
  wire  _EVAL_1719;
  wire  _EVAL_482;
  wire  _EVAL_3399;
  wire  _EVAL_1622;
  wire  _EVAL_2880;
  wire  _EVAL_2010;
  wire  _EVAL_3201;
  wire  _EVAL_3389;
  wire  _EVAL_2479;
  wire  _EVAL_2602;
  wire  _EVAL_2329;
  wire  _EVAL_3955;
  wire  _EVAL_426;
  wire [6:0] _EVAL_3365;
  wire  _EVAL_1074;
  wire  _EVAL_3422;
  wire  _EVAL_563;
  wire  _EVAL_855;
  wire  _EVAL_2313;
  wire  _EVAL_1361;
  wire  _EVAL_2930;
  wire  _EVAL_3929;
  wire  _EVAL_1767;
  wire  _EVAL_2392;
  wire  _EVAL_3355;
  wire  _EVAL_3592;
  wire [126:0] _EVAL_3080;
  wire [126:0] _EVAL_2719;
  wire [126:0] _EVAL_1619;
  wire [126:0] _EVAL_1373;
  wire  _EVAL_2085;
  wire  _EVAL_2367;
  wire  _EVAL_1916;
  wire  _EVAL_3666;
  wire  _EVAL_272;
  wire  _EVAL_4072;
  wire  _EVAL_627;
  wire  _EVAL_3457;
  wire [28:0] _EVAL_2738;
  wire  _EVAL_1878;
  wire  _EVAL_2894;
  wire  _EVAL_2752;
  wire  _EVAL_2799;
  wire  _EVAL_961;
  wire  _EVAL_172;
  wire  _EVAL_3309;
  wire  _EVAL_1760;
  wire  _EVAL_1687;
  wire  _EVAL_1118;
  wire  _EVAL_1844;
  wire  _EVAL_3585;
  wire  _EVAL_1058;
  wire  _EVAL_2529;
  wire  _EVAL_312;
  wire  _EVAL_1700;
  wire  _EVAL_3123;
  wire  _EVAL_2177;
  wire  _EVAL_802;
  wire  _EVAL_1056;
  wire  _EVAL_906;
  wire  _EVAL_3886;
  wire  _EVAL_3753;
  wire  _EVAL_1904;
  wire  _EVAL_2673;
  wire  _EVAL_1451;
  wire  _EVAL_1826;
  wire  _EVAL_1808;
  wire  _EVAL_2338;
  wire  _EVAL_1117;
  wire  _EVAL_2784;
  wire  _EVAL_2550;
  wire  _EVAL_1474;
  wire  _EVAL_659;
  wire  _EVAL_672;
  wire  _EVAL_2946;
  wire  _EVAL_2165;
  wire  _EVAL_3577;
  wire  _EVAL_296;
  wire  _EVAL_3076;
  wire  _EVAL_1696;
  wire  _EVAL_1007;
  wire  _EVAL_3858;
  wire  _EVAL_3778;
  wire  _EVAL_677;
  wire  _EVAL_2374;
  wire [7:0] _EVAL_3975;
  wire  _EVAL_996;
  wire  _EVAL_4051;
  wire  _EVAL_2458;
  wire  _EVAL_578;
  wire  _EVAL_2032;
  wire  _EVAL_4002;
  wire  _EVAL_2734;
  wire  _EVAL_2473;
  wire  _EVAL_407;
  wire  _EVAL_1008;
  wire  _EVAL_2905;
  wire  _EVAL_1199;
  wire  _EVAL_3792;
  wire  _EVAL_2071;
  wire  _EVAL_955;
  wire  _EVAL_1978;
  wire  _EVAL_1902;
  wire  _EVAL_1419;
  wire  _EVAL_4007;
  wire  _EVAL_3942;
  wire  _EVAL_3747;
  wire  _EVAL_1087;
  wire  _EVAL_831;
  wire  _EVAL_4030;
  wire  _EVAL_2089;
  wire  _EVAL_1604;
  wire  _EVAL_209;
  wire  _EVAL_589;
  wire  _EVAL_2476;
  wire  _EVAL_2921;
  wire  _EVAL_1684;
  wire  _EVAL_2890;
  wire  _EVAL_1908;
  wire  _EVAL_3357;
  wire  _EVAL_805;
  wire  _EVAL_2709;
  wire  _EVAL_1353;
  wire  _EVAL_3444;
  wire  _EVAL_2046;
  wire  _EVAL_3090;
  wire  _EVAL_1668;
  wire  _EVAL_838;
  wire  _EVAL_1570;
  wire  _EVAL_4057;
  wire  _EVAL_3160;
  wire  _EVAL_467;
  wire  _EVAL_3126;
  wire  _EVAL_1905;
  wire  _EVAL_1238;
  wire  _EVAL_577;
  wire  _EVAL_3703;
  wire  _EVAL_1090;
  wire  _EVAL_3854;
  wire  _EVAL_2235;
  wire  _EVAL_3386;
  wire  _EVAL_3003;
  wire  _EVAL_3349;
  wire  _EVAL_817;
  wire  _EVAL_3714;
  wire  _EVAL_1344;
  wire  _EVAL_2298;
  wire  _EVAL_2350;
  wire  _EVAL_1304;
  wire  _EVAL_1342;
  wire  _EVAL_1050;
  wire  _EVAL_860;
  wire  _EVAL_689;
  wire  _EVAL_962;
  wire  _EVAL_2077;
  wire  _EVAL_244;
  wire  _EVAL_1610;
  wire  _EVAL_3324;
  wire  _EVAL_2377;
  wire  _EVAL_528;
  wire  _EVAL_3316;
  wire  _EVAL_545;
  wire  _EVAL_486;
  wire [126:0] _EVAL_2549;
  wire  _EVAL_3340;
  wire  _EVAL_3640;
  wire  _EVAL_301;
  wire  _EVAL_3465;
  wire  _EVAL_150;
  wire  _EVAL_1214;
  wire  _EVAL_361;
  wire  _EVAL_3723;
  wire  _EVAL_3106;
  wire  _EVAL_2652;
  wire  _EVAL_2509;
  wire  _EVAL_641;
  wire  _EVAL_1268;
  wire  _EVAL_634;
  wire  _EVAL_1714;
  wire  _EVAL_3437;
  wire  _EVAL_2537;
  wire  _EVAL_3010;
  wire  _EVAL_3277;
  wire  _EVAL_162;
  wire  _EVAL_430;
  wire  _EVAL_1600;
  wire  _EVAL_1223;
  wire  _EVAL_3794;
  wire  _EVAL_1807;
  wire  _EVAL_2207;
  wire  _EVAL_3447;
  wire  _EVAL_2839;
  wire  _EVAL_2414;
  wire  _EVAL_2518;
  wire  _EVAL_307;
  wire  _EVAL_1320;
  wire  _EVAL_4045;
  wire  _EVAL_893;
  wire  _EVAL_2849;
  wire  _EVAL_3686;
  wire  _EVAL_900;
  wire  _EVAL_1138;
  wire  _EVAL_1391;
  wire  _EVAL_1033;
  wire  _EVAL_2772;
  wire  _EVAL_1953;
  wire  _EVAL_2916;
  wire  _EVAL_1693;
  wire  _EVAL_644;
  wire  _EVAL_180;
  wire  _EVAL_201;
  wire  _EVAL_158;
  wire  _EVAL_2216;
  wire  _EVAL_2472;
  wire  _EVAL_1112;
  wire  _EVAL_228;
  wire  _EVAL_601;
  wire  _EVAL_1830;
  wire  _EVAL_2186;
  wire  _EVAL_674;
  wire  _EVAL_1501;
  wire  _EVAL_3155;
  wire  _EVAL_3813;
  wire  _EVAL_3660;
  wire  _EVAL_4067;
  wire  _EVAL_2364;
  wire  _EVAL_2427;
  wire  _EVAL_2418;
  wire  _EVAL_3862;
  wire  _EVAL_628;
  wire  _EVAL_1720;
  wire  _EVAL_161;
  wire  _EVAL_3541;
  wire  _EVAL_1678;
  wire  _EVAL_842;
  wire  _EVAL_2773;
  wire  _EVAL_1255;
  wire  _EVAL_1971;
  wire  _EVAL_2327;
  wire  _EVAL_1789;
  wire  _EVAL_3086;
  wire  _EVAL_1988;
  wire  _EVAL_3435;
  wire  _EVAL_1984;
  wire  _EVAL_1675;
  wire  _EVAL_2049;
  wire  _EVAL_1615;
  wire  _EVAL_2957;
  wire  _EVAL_2268;
  wire  _EVAL_1234;
  wire  _EVAL_3947;
  wire  _EVAL_186;
  wire  _EVAL_2714;
  wire  _EVAL_1217;
  wire  _EVAL_2321;
  wire  _EVAL_2185;
  wire  _EVAL_619;
  wire  _EVAL_885;
  wire  _EVAL_3604;
  wire  _EVAL_3321;
  wire  _EVAL_3133;
  wire  _EVAL_3049;
  wire  _EVAL_281;
  wire  _EVAL_3538;
  wire  _EVAL_2542;
  wire  _EVAL_3046;
  wire  _EVAL_3227;
  wire  _EVAL_3161;
  wire  _EVAL_493;
  wire  _EVAL_3700;
  wire  _EVAL_2002;
  wire  _EVAL_239;
  wire  _EVAL_1422;
  wire  _EVAL_1606;
  wire  _EVAL_1356;
  wire  _EVAL_1336;
  wire  _EVAL_3260;
  wire  _EVAL_154;
  wire  _EVAL_1037;
  wire  _EVAL_1924;
  wire  _EVAL_1498;
  wire  _EVAL_3149;
  wire  _EVAL_2324;
  wire  _EVAL_3545;
  wire  _EVAL_160;
  wire  _EVAL_1662;
  wire  _EVAL_3658;
  wire  _EVAL_2789;
  wire  _EVAL_3193;
  wire  _EVAL_1071;
  wire  _EVAL_1146;
  wire  _EVAL_2022;
  wire  _EVAL_1411;
  wire  _EVAL_3893;
  wire  _EVAL_3040;
  wire  _EVAL_4058;
  wire  _EVAL_408;
  wire  _EVAL_2517;
  wire  _EVAL_3398;
  wire  _EVAL_1865;
  wire  _EVAL_3984;
  wire  _EVAL_3846;
  wire  _EVAL_2908;
  wire  _EVAL_2895;
  wire  _EVAL_2768;
  wire  _EVAL_2417;
  wire  _EVAL_273;
  wire  _EVAL_602;
  wire  _EVAL_2758;
  wire  _EVAL_1803;
  wire  _EVAL_3569;
  wire  _EVAL_3741;
  wire  _EVAL_3536;
  wire  _EVAL_1679;
  wire  _EVAL_322;
  wire  _EVAL_2708;
  wire  _EVAL_2328;
  wire  _EVAL_2722;
  wire  _EVAL_3302;
  wire  _EVAL_2700;
  wire  _EVAL_2213;
  wire  _EVAL_3507;
  wire  _EVAL_2586;
  wire  _EVAL_676;
  wire  _EVAL_406;
  wire  _EVAL_983;
  wire  _EVAL_3115;
  wire  _EVAL_951;
  wire  _EVAL_1254;
  wire  _EVAL_1123;
  wire  _EVAL_3058;
  wire  _EVAL_2897;
  wire  _EVAL_2934;
  wire  _EVAL_3612;
  wire  _EVAL_417;
  wire  _EVAL_3651;
  wire  _EVAL_1442;
  wire  _EVAL_3859;
  wire  _EVAL_2353;
  wire  _EVAL_3373;
  wire  _EVAL_621;
  wire  _EVAL_1256;
  wire  _EVAL_1341;
  wire  _EVAL_1539;
  wire  _EVAL_1551;
  wire  _EVAL_2813;
  wire  _EVAL_434;
  wire  _EVAL_3303;
  wire  _EVAL_1406;
  wire  _EVAL_3922;
  wire  _EVAL_2038;
  wire  _EVAL_862;
  wire  _EVAL_1798;
  wire  _EVAL_3224;
  wire  _EVAL_185;
  wire  _EVAL_3704;
  wire  _EVAL_1003;
  wire  _EVAL_2787;
  wire  _EVAL_3009;
  wire  _EVAL_2552;
  wire  _EVAL_1126;
  wire  _EVAL_2635;
  wire  _EVAL_681;
  wire  _EVAL_261;
  wire  _EVAL_908;
  wire  _EVAL_1685;
  wire  _EVAL_2045;
  wire  _EVAL_3637;
  wire  _EVAL_950;
  wire  _EVAL_2707;
  wire  _EVAL_2475;
  wire  _EVAL_749;
  wire  _EVAL_643;
  wire  _EVAL_2245;
  wire  _EVAL_3951;
  wire  _EVAL_3824;
  wire  _EVAL_3396;
  wire  _EVAL_2093;
  wire  _EVAL_1703;
  wire  _EVAL_213;
  wire  _EVAL_1832;
  wire  _EVAL_937;
  wire  _EVAL_3544;
  wire  _EVAL_3785;
  wire  _EVAL_1482;
  wire  _EVAL_3288;
  wire  _EVAL_192;
  wire  _EVAL_1363;
  wire  _EVAL_3916;
  wire  _EVAL_2967;
  wire  _EVAL_1513;
  wire  _EVAL_972;
  wire  _EVAL_3521;
  wire  _EVAL_3131;
  wire  _EVAL_2994;
  wire  _EVAL_235;
  wire  _EVAL_1165;
  wire  _EVAL_2661;
  wire  _EVAL_1011;
  wire  _EVAL_3129;
  wire  _EVAL_1348;
  wire  _EVAL_2149;
  wire  _EVAL_746;
  wire  _EVAL_1733;
  wire  _EVAL_2964;
  wire  _EVAL_2598;
  wire  _EVAL_3077;
  wire  _EVAL_850;
  wire  _EVAL_1028;
  wire  _EVAL_2028;
  wire  _EVAL_993;
  wire  _EVAL_645;
  wire  _EVAL_1770;
  wire  _EVAL_3452;
  wire  _EVAL_3178;
  wire  _EVAL_2878;
  wire  _EVAL_2626;
  wire  _EVAL_1193;
  wire  _EVAL_2727;
  wire  _EVAL_1974;
  wire  _EVAL_2238;
  wire  _EVAL_1147;
  wire  _EVAL_1712;
  wire  _EVAL_3956;
  wire  _EVAL_3559;
  wire  _EVAL_1030;
  wire  _EVAL_650;
  wire  _EVAL_1367;
  wire  _EVAL_1299;
  wire  _EVAL_2343;
  wire  _EVAL_3727;
  wire  _EVAL_1739;
  wire  _EVAL_1607;
  wire  _EVAL_2405;
  wire  _EVAL_1673;
  wire  _EVAL_3840;
  wire  _EVAL_3748;
  wire  _EVAL_3626;
  wire  _EVAL_1359;
  wire  _EVAL_798;
  wire  _EVAL_3276;
  wire  _EVAL_370;
  wire  _EVAL_2892;
  wire  _EVAL_593;
  wire  _EVAL_701;
  wire  _EVAL_3786;
  wire  _EVAL_2075;
  wire  _EVAL_3175;
  wire  _EVAL_3448;
  wire  _EVAL_2717;
  wire  _EVAL_588;
  wire  _EVAL_2562;
  wire  _EVAL_2223;
  wire  _EVAL_3414;
  wire  _EVAL_1573;
  wire  _EVAL_1302;
  wire  _EVAL_1101;
  wire  _EVAL_2385;
  wire  _EVAL_2152;
  wire  _EVAL_2461;
  wire  _EVAL_799;
  wire  _EVAL_636;
  wire  _EVAL_1928;
  wire  _EVAL_2819;
  wire  _EVAL_1374;
  wire  _EVAL_1508;
  wire  _EVAL_1520;
  wire  _EVAL_1518;
  wire  _EVAL_754;
  wire  _EVAL_2244;
  wire  _EVAL_2592;
  wire  _EVAL_2927;
  wire  _EVAL_3183;
  wire  _EVAL_1968;
  wire  _EVAL_3475;
  wire  _EVAL_713;
  wire  _EVAL_620;
  wire  _EVAL_1665;
  wire  _EVAL_572;
  wire  _EVAL_3223;
  wire  _EVAL_3576;
  wire  _EVAL_2271;
  wire  _EVAL_3915;
  wire  _EVAL_2224;
  wire  _EVAL_513;
  wire  _EVAL_1285;
  wire  _EVAL_2935;
  wire  _EVAL_729;
  wire  _EVAL_317;
  wire  _EVAL_2384;
  wire  _EVAL_3578;
  wire  _EVAL_2175;
  wire  _EVAL_2988;
  wire  _EVAL_2296;
  wire  _EVAL_1593;
  wire  _EVAL_3084;
  wire  _EVAL_1247;
  wire  _EVAL_647;
  wire  _EVAL_3420;
  wire  _EVAL_3474;
  wire  _EVAL_1994;
  wire  _EVAL_3622;
  wire  _EVAL_3430;
  wire  _EVAL_1898;
  wire  _EVAL_422;
  wire  _EVAL_932;
  wire  _EVAL_1149;
  wire  _EVAL_944;
  wire  _EVAL_3624;
  wire  _EVAL_3926;
  wire  _EVAL_3268;
  wire  _EVAL_3533;
  wire  _EVAL_2098;
  wire  _EVAL_3168;
  wire  _EVAL_3752;
  wire  _EVAL_1851;
  wire  _EVAL_2821;
  wire  _EVAL_625;
  wire  _EVAL_338;
  wire  _EVAL_2538;
  wire  _EVAL_2371;
  wire  _EVAL_587;
  wire  _EVAL_3826;
  wire  _EVAL_2876;
  wire  _EVAL_3130;
  wire  _EVAL_414;
  wire  _EVAL_861;
  wire  _EVAL_3250;
  wire  _EVAL_596;
  wire  _EVAL_2842;
  wire  _EVAL_708;
  wire  _EVAL_3307;
  wire  _EVAL_3979;
  wire  _EVAL_2315;
  wire  _EVAL_2274;
  wire  _EVAL_173;
  wire  _EVAL_230;
  wire  _EVAL_2381;
  wire  _EVAL_1150;
  wire  _EVAL_3732;
  wire  _EVAL_2394;
  wire  _EVAL_1494;
  wire  _EVAL_2368;
  wire  _EVAL_2116;
  wire  _EVAL_1276;
  wire  _EVAL_351;
  wire  _EVAL_2487;
  wire  _EVAL_259;
  wire  _EVAL_4018;
  wire  _EVAL_2987;
  wire  _EVAL_2132;
  wire  _EVAL_2495;
  wire  _EVAL_2255;
  wire  _EVAL_782;
  wire  _EVAL_3360;
  wire  _EVAL_1412;
  wire  _EVAL_560;
  wire  _EVAL_1413;
  wire  _EVAL_1649;
  wire  _EVAL_1463;
  wire  _EVAL_2735;
  wire  _EVAL_394;
  wire  _EVAL_2297;
  wire  _EVAL_382;
  wire  _EVAL_3073;
  wire  _EVAL_3855;
  wire  _EVAL_624;
  wire  _EVAL_1568;
  wire  _EVAL_580;
  wire  _EVAL_174;
  wire  _EVAL_3251;
  wire  _EVAL_3484;
  wire  _EVAL_2811;
  wire  _EVAL_3343;
  wire  _EVAL_288;
  wire  _EVAL_1346;
  wire  _EVAL_1154;
  wire  _EVAL_280;
  wire  _EVAL_2471;
  wire  _EVAL_3271;
  wire  _EVAL_3477;
  wire  _EVAL_3105;
  wire  _EVAL_2270;
  wire  _EVAL_737;
  wire  _EVAL_664;
  wire  _EVAL_1389;
  wire  _EVAL_1796;
  wire  _EVAL_2925;
  wire  _EVAL_769;
  wire  _EVAL_1115;
  wire  _EVAL_2814;
  wire  _EVAL_531;
  wire  _EVAL_1656;
  wire  _EVAL_970;
  wire  _EVAL_1569;
  wire  _EVAL_2036;
  wire  _EVAL_2833;
  wire  _EVAL_253;
  wire  _EVAL_3548;
  wire  _EVAL_1546;
  wire  _EVAL_2349;
  wire  _EVAL_3007;
  wire  _EVAL_844;
  wire  _EVAL_1657;
  wire  _EVAL_3630;
  wire  _EVAL_901;
  wire  _EVAL_278;
  wire  _EVAL_2178;
  wire  _EVAL_2997;
  wire  _EVAL_771;
  wire  _EVAL_3787;
  wire  _EVAL_2888;
  wire  _EVAL_314;
  wire  _EVAL_2409;
  wire  _EVAL_1732;
  wire  _EVAL_3900;
  wire  _EVAL_2920;
  wire  _EVAL_1797;
  wire  _EVAL_4014;
  wire  _EVAL_2345;
  wire  _EVAL_437;
  wire  _EVAL_3609;
  wire  _EVAL_976;
  wire  _EVAL_2723;
  wire  _EVAL_2896;
  wire  _EVAL_3912;
  wire  _EVAL_3114;
  wire  _EVAL_495;
  wire  _EVAL_751;
  wire  _EVAL_3518;
  wire  _EVAL_282;
  wire  _EVAL_3478;
  wire  _EVAL_3905;
  wire  _EVAL_2424;
  wire  _EVAL_2523;
  wire  _EVAL_1762;
  wire  _EVAL_1893;
  wire  _EVAL_2422;
  wire  _EVAL_2243;
  wire  _EVAL_1794;
  wire  _EVAL_2875;
  wire  _EVAL_1260;
  wire  _EVAL_3647;
  wire  _EVAL_1269;
  wire  _EVAL_2490;
  wire  _EVAL_745;
  wire  _EVAL_503;
  wire  _EVAL_918;
  wire  _EVAL_1495;
  wire  _EVAL_3425;
  wire  _EVAL_3393;
  wire  _EVAL_3938;
  wire  _EVAL_4047;
  wire  _EVAL_3254;
  wire  _EVAL_2462;
  wire  _EVAL_1954;
  wire  _EVAL_2135;
  wire  _EVAL_1909;
  wire  _EVAL_1020;
  wire  _EVAL_425;
  wire  _EVAL_2164;
  wire  _EVAL_1443;
  wire  _EVAL_3492;
  wire  _EVAL_3971;
  wire  _EVAL_1394;
  wire  _EVAL_191;
  wire  _EVAL_698;
  wire  _EVAL_3775;
  wire  _EVAL_3560;
  wire  _EVAL_1347;
  wire  _EVAL_3570;
  wire  _EVAL_2973;
  wire  _EVAL_487;
  wire  _EVAL_2351;
  wire  _EVAL_3793;
  wire  _EVAL_3473;
  wire  _EVAL_2227;
  wire  _EVAL_3205;
  wire  _EVAL_761;
  wire  _EVAL_3712;
  wire  _EVAL_2857;
  wire  _EVAL_1467;
  wire  _EVAL_3745;
  wire  _EVAL_2286;
  wire  _EVAL_1272;
  wire  _EVAL_3502;
  wire  _EVAL_2687;
  wire  _EVAL_871;
  wire  _EVAL_1184;
  wire  _EVAL_386;
  wire  _EVAL_3808;
  wire  _EVAL_2710;
  wire  _EVAL_1824;
  wire  _EVAL_3875;
  wire  _EVAL_3362;
  wire  _EVAL_2295;
  wire  _EVAL_786;
  wire  _EVAL_419;
  wire  _EVAL_616;
  wire  _EVAL_2918;
  wire  _EVAL_1981;
  wire  _EVAL_206;
  wire  _EVAL_4042;
  wire  _EVAL_1436;
  wire  _EVAL_2680;
  wire  _EVAL_1864;
  wire  _EVAL_1993;
  wire  _EVAL_1579;
  wire  _EVAL_3138;
  wire  _EVAL_1262;
  wire  _EVAL_177;
  wire  _EVAL_726;
  wire  _EVAL_3925;
  wire  _EVAL_1972;
  wire  _EVAL_2840;
  wire  _EVAL_3108;
  wire  _EVAL_2193;
  wire  _EVAL_3311;
  wire  _EVAL_3187;
  wire  _EVAL_3034;
  wire  _EVAL_3289;
  wire  _EVAL_2431;
  wire  _EVAL_839;
  wire  _EVAL_1627;
  wire  _EVAL_2282;
  wire  _EVAL_2217;
  wire  _EVAL_1349;
  wire  _EVAL_1038;
  wire  _EVAL_2019;
  wire  _EVAL_3607;
  wire  _EVAL_4036;
  wire  _EVAL_1303;
  wire  _EVAL_1623;
  wire  _EVAL_1435;
  wire  _EVAL_1478;
  wire  _EVAL_2074;
  wire  _EVAL_3483;
  wire  _EVAL_1385;
  wire  _EVAL_3182;
  wire  _EVAL_3706;
  wire  _EVAL_3902;
  wire  _EVAL_2370;
  wire  _EVAL_1757;
  wire  _EVAL_1288;
  wire  _EVAL_1529;
  wire  _EVAL_3830;
  wire  _EVAL_151;
  wire  _EVAL_3948;
  wire  _EVAL_1932;
  wire  _EVAL_3297;
  wire  _EVAL_1308;
  wire  _EVAL_3698;
  wire  _EVAL_2655;
  wire  _EVAL_2521;
  wire  _EVAL_2360;
  wire  _EVAL_227;
  wire  _EVAL_1290;
  wire  _EVAL_1896;
  wire  _EVAL_490;
  wire  _EVAL_2936;
  wire  _EVAL_4008;
  wire  _EVAL_3695;
  wire  _EVAL_3403;
  wire  _EVAL_3814;
  wire  _EVAL_292;
  wire  _EVAL_549;
  wire  _EVAL_1095;
  wire  _EVAL_1641;
  wire  _EVAL_3202;
  wire  _EVAL_3711;
  wire  _EVAL_157;
  wire  _EVAL_671;
  wire  _EVAL_2474;
  wire  _EVAL_1850;
  wire  _EVAL_2170;
  wire  _EVAL_3657;
  wire  _EVAL_2761;
  wire  _EVAL_4055;
  wire  _EVAL_2998;
  wire  _EVAL_3874;
  wire  _EVAL_610;
  wire  _EVAL_376;
  wire  _EVAL_2390;
  wire  _EVAL_2453;
  wire  _EVAL_240;
  wire  _EVAL_852;
  wire  _EVAL_1586;
  wire  _EVAL_1882;
  wire  _EVAL_383;
  wire  _EVAL_579;
  wire  _EVAL_613;
  wire  _EVAL_3978;
  wire  _EVAL_1317;
  wire  _EVAL_582;
  wire  _EVAL_1046;
  wire  _EVAL_2564;
  wire  _EVAL_714;
  wire  _EVAL_913;
  wire  _EVAL_3004;
  wire  _EVAL_3066;
  wire  _EVAL_2926;
  wire  _EVAL_1219;
  wire  _EVAL_452;
  wire  _EVAL_683;
  wire  _EVAL_1111;
  wire  _EVAL_1284;
  wire  _EVAL_224;
  wire  _EVAL_3990;
  wire  _EVAL_1006;
  wire  _EVAL_233;
  wire  _EVAL_2123;
  wire  _EVAL_787;
  wire  _EVAL_1825;
  wire  _EVAL_995;
  wire  _EVAL_3354;
  wire  _EVAL_1388;
  wire  _EVAL_1995;
  wire  _EVAL_733;
  wire  _EVAL_2262;
  wire  _EVAL_1772;
  wire  _EVAL_2067;
  wire  _EVAL_2703;
  wire  _EVAL_3739;
  wire  _EVAL_1517;
  wire  _EVAL_2519;
  wire  _EVAL_3211;
  wire  _EVAL_3111;
  wire  _EVAL_1592;
  wire  _EVAL_2466;
  wire  _EVAL_1220;
  wire  _EVAL_2168;
  wire  _EVAL_3033;
  wire  _EVAL_2246;
  wire  _EVAL_3708;
  wire  _EVAL_510;
  wire  _EVAL_433;
  wire  _EVAL_3200;
  SiFive__EVAL_181_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  assign _EVAL_2645 = Queue__EVAL_5;
  assign _EVAL_929 = _EVAL_131 & _EVAL_2645;
  assign _EVAL_534 = _EVAL_86 == 3'h4;
  assign _EVAL_3781 = _EVAL_929 & _EVAL_534;
  assign _EVAL_2747 = _EVAL_910[23:0];
  assign _EVAL_1249 = _EVAL_2747[19];
  assign _EVAL_2976 = _EVAL_2747[11];
  assign _EVAL_1925 = _EVAL_2747[10];
  assign _EVAL_2558 = _EVAL_2747[6];
  assign _EVAL_1749 = _EVAL_2747[5];
  assign _EVAL_843 = _EVAL_2747[4];
  assign _EVAL_3057 = _EVAL_2747[3];
  assign _EVAL_367 = _EVAL_2747[2];
  assign _EVAL_1519 = _EVAL_2747[1];
  assign _EVAL_974 = _EVAL_2747[0];
  assign _EVAL_2638 = {_EVAL_1249,_EVAL_2976,_EVAL_1925,_EVAL_2558,_EVAL_1749,_EVAL_843,_EVAL_3057,_EVAL_367,_EVAL_1519,_EVAL_974};
  assign _EVAL_1942 = 1024'h1 << _EVAL_2638;
  assign _EVAL_2990 = _EVAL_1942[96];
  assign _EVAL_758 = _EVAL_3781 & _EVAL_2990;
  assign _EVAL_1381 = _EVAL_1942[68];
  assign _EVAL_599 = _EVAL_3781 & _EVAL_1381;
  assign _EVAL_3143 = _EVAL_2747 & 24'hf7f380;
  assign _EVAL_246 = _EVAL_3143 == 24'h0;
  assign _EVAL_1588 = _EVAL_599 & _EVAL_246;
  assign _EVAL_1647 = _EVAL_534 == 1'h0;
  assign _EVAL_3402 = _EVAL_929 & _EVAL_1647;
  assign _EVAL_3188 = _EVAL_1942[79];
  assign _EVAL_1300 = _EVAL_3402 & _EVAL_3188;
  assign _EVAL_2191 = _EVAL_1300 & _EVAL_246;
  assign _EVAL_3225 = _EVAL_69[3];
  assign _EVAL_1726 = _EVAL_3225 ? 8'hff : 8'h0;
  assign _EVAL_2817 = _EVAL_69[2];
  assign _EVAL_3261 = _EVAL_2817 ? 8'hff : 8'h0;
  assign _EVAL_1754 = _EVAL_69[1];
  assign _EVAL_3977 = _EVAL_1754 ? 8'hff : 8'h0;
  assign _EVAL_779 = _EVAL_69[0];
  assign _EVAL_1379 = _EVAL_779 ? 8'hff : 8'h0;
  assign _EVAL_1377 = {_EVAL_1726,_EVAL_3261,_EVAL_3977,_EVAL_1379};
  assign _EVAL_347 = _EVAL_1377[2:0];
  assign _EVAL_1996 = _EVAL_347 == 3'h7;
  assign _EVAL_458 = _EVAL_2191 & _EVAL_1996;
  assign _EVAL_3286 = _EVAL_1942[18];
  assign _EVAL_402 = _EVAL_1942[128];
  assign _EVAL_2995 = _EVAL_3402 & _EVAL_402;
  assign _EVAL_1545 = _EVAL_2995 & _EVAL_246;
  assign _EVAL_3954 = _EVAL_1377[2];
  assign _EVAL_948 = _EVAL_1545 & _EVAL_3954;
  assign _EVAL_3110 = _EVAL_3059 & _EVAL_2184;
  assign _EVAL_911 = _EVAL_3059 & _EVAL_429;
  assign _EVAL_1778 = _EVAL_1942[32];
  assign _EVAL_3790 = _EVAL_1942[44];
  assign _EVAL_2551 = _EVAL_3781 & _EVAL_3790;
  assign _EVAL_1129 = _EVAL_2551 & _EVAL_246;
  assign _EVAL_889 = _EVAL_1942[41];
  assign _EVAL_1831 = _EVAL_3402 & _EVAL_889;
  assign _EVAL_1324 = _EVAL_1377[25];
  assign _EVAL_859 = _EVAL_1545 & _EVAL_1324;
  assign _EVAL_1278 = _EVAL_2999[131];
  assign _EVAL_3154 = _EVAL_3059 & _EVAL_1278;
  assign _EVAL_3075 = _EVAL_3154 & _EVAL_2267;
  assign _EVAL_3471 = _EVAL_2124[25];
  assign _EVAL_1252 = _EVAL_3075 & _EVAL_3471;
  assign _EVAL_2812 = _EVAL_3059 & _EVAL_1531;
  assign _EVAL_3446 = _EVAL_3059 & _EVAL_1886;
  assign _EVAL_958 = _EVAL_3446 & _EVAL_2267;
  assign _EVAL_3596 = _EVAL_2124[24];
  assign _EVAL_1806 = _EVAL_3075 & _EVAL_3596;
  assign _EVAL_2497 = _EVAL_1942[99];
  assign _EVAL_905 = _EVAL_3402 & _EVAL_2497;
  assign _EVAL_747 = _EVAL_905 & _EVAL_246;
  assign _EVAL_1307 = _EVAL_2999[130];
  assign _EVAL_2101 = _EVAL_3673 & _EVAL_1307;
  assign _EVAL_1279 = _EVAL_2101 & _EVAL_2267;
  assign _EVAL_3194 = _EVAL_2124[11];
  assign _EVAL_1507 = _EVAL_1279 & _EVAL_3194;
  assign _EVAL_3906 = _EVAL_1942[78];
  assign _EVAL_399 = _EVAL_3059 & _EVAL_2610;
  assign _EVAL_1543 = _EVAL_399 & _EVAL_2267;
  assign _EVAL_2961 = _EVAL_2124[22];
  assign _EVAL_4059 = _EVAL_3075 & _EVAL_2961;
  assign _EVAL_3022 = _EVAL_2999[129];
  assign _EVAL_1605 = _EVAL_3673 & _EVAL_3022;
  assign _EVAL_2112 = _EVAL_1605 & _EVAL_2267;
  assign _EVAL_806 = _EVAL_2124[18];
  assign _EVAL_454 = _EVAL_2112 & _EVAL_806;
  assign _EVAL_204 = _EVAL_1942[40];
  assign _EVAL_1024 = _EVAL_1942[131];
  assign _EVAL_1275 = _EVAL_3781 & _EVAL_1024;
  assign _EVAL_1857 = _EVAL_1275 & _EVAL_246;
  assign _EVAL_3470 = _EVAL_1377[28];
  assign _EVAL_2674 = _EVAL_1857 & _EVAL_3470;
  assign _EVAL_3568 = _EVAL_3059 & _EVAL_822;
  assign _EVAL_3330 = _EVAL_3781 & _EVAL_402;
  assign _EVAL_1470 = _EVAL_3330 & _EVAL_246;
  assign _EVAL_2020 = _EVAL_1377[20];
  assign _EVAL_2180 = _EVAL_1470 & _EVAL_2020;
  assign _EVAL_3652 = _EVAL_1942[88];
  assign _EVAL_3987 = _EVAL_3402 & _EVAL_3652;
  assign _EVAL_2585 = _EVAL_3987 & _EVAL_246;
  assign _EVAL_3901 = _EVAL_2585 & _EVAL_1996;
  assign _EVAL_2594 = _EVAL_1377[31];
  assign _EVAL_2591 = _EVAL_1857 & _EVAL_2594;
  assign _EVAL_2219 = _EVAL_3059 & _EVAL_1307;
  assign _EVAL_2986 = _EVAL_2219 & _EVAL_2267;
  assign _EVAL_1889 = _EVAL_2124[9];
  assign _EVAL_680 = _EVAL_2986 & _EVAL_1889;
  assign _EVAL_4031 = _EVAL_2124[14];
  assign _EVAL_3812 = _EVAL_3075 & _EVAL_4031;
  assign _EVAL_1209 = _EVAL_1847 - 1'h1;
  assign _EVAL_998 = _EVAL_1847 & _EVAL_1209;
  assign _EVAL_258 = _EVAL_998 == 1'h0;
  assign _EVAL_3238 = _EVAL_258 | _EVAL_105;
  assign _EVAL_2380 = _EVAL_1942[98];
  assign _EVAL_827 = _EVAL_3402 & _EVAL_2380;
  assign _EVAL_309 = _EVAL_827 & _EVAL_246;
  assign _EVAL_3558 = _EVAL_309 & _EVAL_1996;
  assign _EVAL_2676 = _EVAL_1942[50];
  assign _EVAL_1566 = _EVAL_3402 & _EVAL_2676;
  assign _EVAL_3207 = _EVAL_1942[100];
  assign _EVAL_3206 = _EVAL_3781 & _EVAL_3207;
  assign _EVAL_1174 = _EVAL_3206 & _EVAL_246;
  assign _EVAL_1643 = _EVAL_1942[123];
  assign _EVAL_1057 = _EVAL_3781 & _EVAL_1643;
  assign _EVAL_1742 = _EVAL_1057 & _EVAL_246;
  assign _EVAL_1417 = _EVAL_347 != 3'h0;
  assign _EVAL_1505 = _EVAL_1742 & _EVAL_1417;
  assign _EVAL_1010 = _EVAL_3059 & _EVAL_2122;
  assign _EVAL_3048 = _EVAL_1942[92];
  assign _EVAL_379 = _EVAL_3402 & _EVAL_3048;
  assign _EVAL_3377 = _EVAL_379 & _EVAL_246;
  assign _EVAL_496 = _EVAL_1942[23];
  assign _EVAL_3889 = _EVAL_3781 & _EVAL_496;
  assign _EVAL_3485 = _EVAL_3889 & _EVAL_246;
  assign _EVAL_2671 = _EVAL_3485 & _EVAL_1417;
  assign _EVAL_2650 = _EVAL_1942[67];
  assign _EVAL_3148 = _EVAL_1377[21];
  assign _EVAL_3461 = _EVAL_1545 & _EVAL_3148;
  assign _EVAL_1497 = _EVAL_911 & _EVAL_2267;
  assign _EVAL_1910 = _EVAL_3165 != 3'h0;
  assign _EVAL_508 = _EVAL_1497 & _EVAL_1910;
  assign _EVAL_3280 = _EVAL_1942[89];
  assign _EVAL_2211 = _EVAL_3781 & _EVAL_3280;
  assign _EVAL_1681 = _EVAL_2211 & _EVAL_246;
  assign _EVAL_694 = _EVAL_3059 & _EVAL_1907;
  assign _EVAL_1180 = _EVAL_3402 & _EVAL_3280;
  assign _EVAL_3029 = _EVAL_1180 & _EVAL_246;
  assign _EVAL_183 = _EVAL_3059 & _EVAL_1328;
  assign _EVAL_2041 = _EVAL_183 & _EVAL_2267;
  assign _EVAL_1221 = _EVAL_1332 != 7'h0;
  assign _EVAL_609 = _EVAL_2041 & _EVAL_1221;
  assign _EVAL_2062 = _EVAL_1942[121];
  assign _EVAL_3621 = _EVAL_3402 & _EVAL_2062;
  assign _EVAL_2733 = _EVAL_3621 & _EVAL_246;
  assign _EVAL_1145 = _EVAL_1377[27];
  assign _EVAL_2583 = _EVAL_1857 & _EVAL_1145;
  assign _EVAL_2941 = _EVAL_1942[257];
  assign _EVAL_2991 = _EVAL_3402 & _EVAL_2941;
  assign _EVAL_933 = _EVAL_2991 & _EVAL_246;
  assign _EVAL_692 = _EVAL_1831 & _EVAL_246;
  assign _EVAL_3295 = _EVAL_1942[82];
  assign _EVAL_2525 = _EVAL_3402 & _EVAL_3295;
  assign _EVAL_1638 = _EVAL_3059 & _EVAL_873;
  assign _EVAL_3228 = _EVAL_3059 & _EVAL_1201;
  assign _EVAL_3736 = _EVAL_3228 & _EVAL_2267;
  assign _EVAL_2319 = _EVAL_638 != 8'h0;
  assign _EVAL_2199 = _EVAL_3736 & _EVAL_2319;
  assign _EVAL_743 = _EVAL_3781 & _EVAL_2062;
  assign _EVAL_2166 = _EVAL_743 & _EVAL_246;
  assign _EVAL_1951 = _EVAL_3059 & _EVAL_1515;
  assign _EVAL_2685 = _EVAL_1951 & _EVAL_2267;
  assign _EVAL_1960 = _EVAL_2685 & _EVAL_1910;
  assign _EVAL_3063 = _EVAL_1942[258];
  assign _EVAL_250 = _EVAL_3781 & _EVAL_3063;
  assign _EVAL_1398 = _EVAL_250 & _EVAL_246;
  assign _EVAL_2699 = _EVAL_3059 & _EVAL_824;
  assign _EVAL_469 = _EVAL_2699 & _EVAL_2267;
  assign _EVAL_3562 = _EVAL_2999[128];
  assign _EVAL_3450 = _EVAL_3059 & _EVAL_3562;
  assign _EVAL_431 = _EVAL_3450 & _EVAL_2267;
  assign _EVAL_4006 = _EVAL_2124[21];
  assign _EVAL_804 = _EVAL_431 & _EVAL_4006;
  assign _EVAL_2984 = _EVAL_1377[6];
  assign _EVAL_2800 = _EVAL_1470 & _EVAL_2984;
  assign _EVAL_2091 = _EVAL_3059 & _EVAL_1475;
  assign _EVAL_1702 = _EVAL_2091 & _EVAL_2267;
  assign _EVAL_2004 = _EVAL_1702 & _EVAL_1910;
  assign _EVAL_3272 = _EVAL_1942[2];
  assign _EVAL_1092 = _EVAL_3402 & _EVAL_3272;
  assign _EVAL_3966 = _EVAL_1092 & _EVAL_246;
  assign _EVAL_717 = _EVAL_3966 & _EVAL_1996;
  assign _EVAL_3381 = _EVAL_3235 > 7'h0;
  assign _EVAL_3856 = _EVAL_1847 & _EVAL_3381;
  assign _EVAL_520 = _EVAL_1377[26];
  assign _EVAL_2794 = _EVAL_1470 & _EVAL_520;
  assign _EVAL_2042 = _EVAL_1942[22];
  assign _EVAL_1053 = _EVAL_1942[10];
  assign _EVAL_1383 = _EVAL_1942[47];
  assign _EVAL_3973 = _EVAL_3781 & _EVAL_1383;
  assign _EVAL_1818 = _EVAL_1942[124];
  assign _EVAL_2501 = _EVAL_3402 & _EVAL_1818;
  assign _EVAL_2609 = _EVAL_2501 & _EVAL_246;
  assign _EVAL_3701 = _EVAL_2124[12];
  assign _EVAL_3196 = _EVAL_3075 & _EVAL_3701;
  assign _EVAL_2340 = _EVAL_3059 & _EVAL_2835;
  assign _EVAL_3413 = _EVAL_2340 & _EVAL_2267;
  assign _EVAL_2978 = _EVAL_1942[55];
  assign _EVAL_1821 = _EVAL_3402 & _EVAL_2978;
  assign _EVAL_2397 = _EVAL_3402 & _EVAL_1024;
  assign _EVAL_3897 = _EVAL_2397 & _EVAL_246;
  assign _EVAL_1868 = _EVAL_1377[14];
  assign _EVAL_649 = _EVAL_3897 & _EVAL_1868;
  assign _EVAL_3180 = _EVAL_2124[27];
  assign _EVAL_3865 = _EVAL_431 & _EVAL_3180;
  assign _EVAL_834 = _EVAL_1942[129];
  assign _EVAL_3445 = _EVAL_3402 & _EVAL_834;
  assign _EVAL_3458 = _EVAL_3445 & _EVAL_246;
  assign _EVAL_3397 = _EVAL_1942[20];
  assign _EVAL_2732 = _EVAL_3781 & _EVAL_3397;
  assign _EVAL_1744 = _EVAL_2732 & _EVAL_246;
  assign _EVAL_1172 = _EVAL_1942[26];
  assign _EVAL_3363 = _EVAL_2124[23];
  assign _EVAL_2263 = _EVAL_1279 & _EVAL_3363;
  assign _EVAL_629 = _EVAL_1942[65];
  assign _EVAL_311 = _EVAL_3402 & _EVAL_629;
  assign _EVAL_266 = _EVAL_311 & _EVAL_246;
  assign _EVAL_215 = _EVAL_2124[0];
  assign _EVAL_1695 = _EVAL_2112 & _EVAL_215;
  assign _EVAL_3810 = _EVAL_1942[130];
  assign _EVAL_4048 = _EVAL_3402 & _EVAL_3810;
  assign _EVAL_1724 = _EVAL_4048 & _EVAL_246;
  assign _EVAL_2375 = _EVAL_1377[10];
  assign _EVAL_3264 = _EVAL_1724 & _EVAL_2375;
  assign _EVAL_2339 = _EVAL_2124[19];
  assign _EVAL_3976 = _EVAL_3075 & _EVAL_2339;
  assign _EVAL_1911 = _EVAL_1857 & _EVAL_520;
  assign _EVAL_1335 = _EVAL_1942[120];
  assign _EVAL_894 = _EVAL_3781 & _EVAL_1335;
  assign _EVAL_1862 = _EVAL_894 & _EVAL_246;
  assign _EVAL_543 = _EVAL_1377[9];
  assign _EVAL_2266 = _EVAL_3897 & _EVAL_543;
  assign _EVAL_3035 = _EVAL_3673 & _EVAL_3562;
  assign _EVAL_1553 = _EVAL_3035 & _EVAL_2267;
  assign _EVAL_3779 = _EVAL_2124[10];
  assign _EVAL_2668 = _EVAL_1553 & _EVAL_3779;
  assign _EVAL_3869 = _EVAL_3059 & _EVAL_979;
  assign _EVAL_1894 = _EVAL_3781 & _EVAL_3188;
  assign _EVAL_1504 = _EVAL_1894 & _EVAL_246;
  assign _EVAL_2053 = _EVAL_1504 & _EVAL_1417;
  assign _EVAL_1476 = _EVAL_1942[101];
  assign _EVAL_1689 = _EVAL_3781 & _EVAL_1476;
  assign _EVAL_356 = _EVAL_1942[115];
  assign _EVAL_699 = _EVAL_3781 & _EVAL_356;
  assign _EVAL_2445 = _EVAL_699 & _EVAL_246;
  assign _EVAL_2798 = _EVAL_2445 & _EVAL_1417;
  assign _EVAL_1245 = _EVAL_2124[4];
  assign _EVAL_1775 = _EVAL_1279 & _EVAL_1245;
  assign _EVAL_2105 = _EVAL_3781 & _EVAL_889;
  assign _EVAL_3664 = _EVAL_1942[109];
  assign _EVAL_1666 = _EVAL_3781 & _EVAL_3664;
  assign _EVAL_1045 = _EVAL_1377[31:24];
  assign _EVAL_2544 = _EVAL_1045 == 8'hff;
  assign _EVAL_1047 = _EVAL_3781 & _EVAL_834;
  assign _EVAL_1040 = _EVAL_1047 & _EVAL_246;
  assign _EVAL_1567 = _EVAL_1040 & _EVAL_1868;
  assign _EVAL_2712 = _EVAL_1942[13];
  assign _EVAL_2560 = _EVAL_3402 & _EVAL_2712;
  assign _EVAL_2649 = _EVAL_2560 & _EVAL_246;
  assign _EVAL_2423 = _EVAL_2649 & _EVAL_1996;
  assign _EVAL_3104 = _EVAL_3973 & _EVAL_246;
  assign _EVAL_3557 = _EVAL_3402 & _EVAL_3063;
  assign _EVAL_2173 = _EVAL_3557 & _EVAL_246;
  assign _EVAL_1371 = _EVAL_1377[7:0];
  assign _EVAL_2283 = _EVAL_1371 == 8'hff;
  assign _EVAL_1459 = _EVAL_2173 & _EVAL_2283;
  assign _EVAL_1179 = _EVAL_758 & _EVAL_246;
  assign _EVAL_321 = _EVAL_1179 & _EVAL_1417;
  assign _EVAL_3298 = _EVAL_3458 & _EVAL_1868;
  assign _EVAL_818 = _EVAL_3059 & _EVAL_4054;
  assign _EVAL_637 = _EVAL_1942[259];
  assign _EVAL_2151 = _EVAL_1942[8];
  assign _EVAL_1207 = _EVAL_3402 & _EVAL_2151;
  assign _EVAL_3376 = _EVAL_1207 & _EVAL_246;
  assign _EVAL_1228 = _EVAL_3376 & _EVAL_1996;
  assign _EVAL_4049 = _EVAL_3059 & _EVAL_1944;
  assign _EVAL_3093 = _EVAL_4049 & _EVAL_2267;
  assign _EVAL_2824 = _EVAL_1377[13];
  assign _EVAL_721 = _EVAL_1857 & _EVAL_2824;
  assign _EVAL_1903 = _EVAL_1942[76];
  assign _EVAL_2815 = _EVAL_3402 & _EVAL_1903;
  assign _EVAL_897 = _EVAL_2815 & _EVAL_246;
  assign _EVAL_611 = _EVAL_3059 & _EVAL_1533;
  assign _EVAL_2027 = _EVAL_611 & _EVAL_2267;
  assign _EVAL_1354 = _EVAL_1377[12];
  assign _EVAL_327 = _EVAL_1040 & _EVAL_1354;
  assign _EVAL_3516 = _EVAL_3059 & _EVAL_3520;
  assign _EVAL_2179 = _EVAL_3673 & _EVAL_1278;
  assign _EVAL_1034 = _EVAL_2179 & _EVAL_2267;
  assign _EVAL_1224 = _EVAL_2124[28];
  assign _EVAL_471 = _EVAL_1034 & _EVAL_1224;
  assign _EVAL_2621 = _EVAL_3781 & _EVAL_3810;
  assign _EVAL_1522 = _EVAL_2621 & _EVAL_246;
  assign _EVAL_2691 = _EVAL_1377[4];
  assign _EVAL_1012 = _EVAL_1522 & _EVAL_2691;
  assign _EVAL_914 = _EVAL_1040 & _EVAL_2984;
  assign _EVAL_3270 = _EVAL_3059 & _EVAL_3908;
  assign _EVAL_3000 = _EVAL_1377[23];
  assign _EVAL_2617 = _EVAL_1942[91];
  assign _EVAL_966 = _EVAL_3402 & _EVAL_2617;
  assign _EVAL_1901 = _EVAL_966 & _EVAL_246;
  assign _EVAL_477 = _EVAL_1901 & _EVAL_1996;
  assign _EVAL_1005 = _EVAL_3059 & _EVAL_1107;
  assign _EVAL_3503 = _EVAL_1005 & _EVAL_2267;
  assign _EVAL_1078 = _EVAL_3781 & _EVAL_2151;
  assign _EVAL_3693 = _EVAL_1377[5];
  assign _EVAL_980 = _EVAL_1040 & _EVAL_3693;
  assign _EVAL_3347 = _EVAL_1942[126];
  assign _EVAL_919 = _EVAL_3402 & _EVAL_3347;
  assign _EVAL_756 = _EVAL_919 & _EVAL_246;
  assign _EVAL_4019 = _EVAL_1942[4];
  assign _EVAL_403 = _EVAL_3402 & _EVAL_4019;
  assign _EVAL_530 = _EVAL_3059 & _EVAL_3018;
  assign _EVAL_2775 = _EVAL_530 & _EVAL_2267;
  assign _EVAL_3795 = _EVAL_2775 & _EVAL_1910;
  assign _EVAL_825 = _EVAL_2112 & _EVAL_3194;
  assign _EVAL_1079 = _EVAL_2609 & _EVAL_1996;
  assign _EVAL_4016 = _EVAL_2124[5];
  assign _EVAL_1041 = _EVAL_3075 & _EVAL_4016;
  assign _EVAL_152 = _EVAL_1942[512];
  assign _EVAL_3391 = _EVAL_3781 & _EVAL_152;
  assign _EVAL_1735 = _EVAL_3391 & _EVAL_246;
  assign _EVAL_1295 = _EVAL_1735 & _EVAL_1417;
  assign _EVAL_4069 = _EVAL_1942[127];
  assign _EVAL_1701 = _EVAL_3781 & _EVAL_4069;
  assign _EVAL_790 = _EVAL_1701 & _EVAL_246;
  assign _EVAL_957 = _EVAL_3059 & _EVAL_3022;
  assign _EVAL_2804 = _EVAL_957 & _EVAL_2267;
  assign _EVAL_2072 = _EVAL_2124[2];
  assign _EVAL_3322 = _EVAL_2804 & _EVAL_2072;
  assign _EVAL_1989 = _EVAL_1942[37];
  assign _EVAL_669 = _EVAL_1942[54];
  assign _EVAL_3248 = _EVAL_3869 & _EVAL_2267;
  assign _EVAL_868 = _EVAL_3248 & _EVAL_1910;
  assign _EVAL_3218 = _EVAL_1942[81];
  assign _EVAL_2369 = _EVAL_3781 & _EVAL_3218;
  assign _EVAL_1372 = _EVAL_1942[256];
  assign _EVAL_1834 = _EVAL_3781 & _EVAL_1372;
  assign _EVAL_3140 = _EVAL_1834 & _EVAL_246;
  assign _EVAL_2756 = _EVAL_1377[0];
  assign _EVAL_3561 = _EVAL_3140 & _EVAL_2756;
  assign _EVAL_2083 = _EVAL_3059 & _EVAL_2940;
  assign _EVAL_535 = _EVAL_2083 & _EVAL_2267;
  assign _EVAL_1048 = _EVAL_2124[26];
  assign _EVAL_1044 = _EVAL_1553 & _EVAL_1048;
  assign _EVAL_3246 = _EVAL_3059 & _EVAL_845;
  assign _EVAL_2996 = _EVAL_3246 & _EVAL_2267;
  assign _EVAL_518 = _EVAL_2996 & _EVAL_1910;
  assign _EVAL_3163 = _EVAL_3059 & _EVAL_3884;
  assign _EVAL_3472 = _EVAL_1857 & _EVAL_3148;
  assign _EVAL_3285 = _EVAL_1377[7];
  assign _EVAL_3455 = _EVAL_1545 & _EVAL_3285;
  assign _EVAL_662 = _EVAL_1377[19];
  assign _EVAL_3914 = _EVAL_3458 & _EVAL_662;
  assign _EVAL_884 = _EVAL_1857 & _EVAL_1354;
  assign _EVAL_2241 = _EVAL_1034 & _EVAL_215;
  assign _EVAL_2556 = _EVAL_1470 & _EVAL_3693;
  assign _EVAL_392 = _EVAL_1724 & _EVAL_1354;
  assign _EVAL_1621 = _EVAL_1377[11];
  assign _EVAL_1396 = _EVAL_1724 & _EVAL_1621;
  assign _EVAL_3468 = _EVAL_1942[64];
  assign _EVAL_2683 = _EVAL_3781 & _EVAL_3468;
  assign _EVAL_2043 = _EVAL_2124[13];
  assign _EVAL_3988 = _EVAL_431 & _EVAL_2043;
  assign _EVAL_3278 = _EVAL_3059 & _EVAL_1326;
  assign _EVAL_551 = _EVAL_3278 & _EVAL_2267;
  assign _EVAL_2736 = _EVAL_551 & _EVAL_1910;
  assign _EVAL_858 = _EVAL_3402 & _EVAL_2650;
  assign _EVAL_1277 = _EVAL_858 & _EVAL_246;
  assign _EVAL_755 = _EVAL_1277 & _EVAL_1996;
  assign _EVAL_2962 = _EVAL_431 & _EVAL_4031;
  assign _EVAL_2305 = _EVAL_1942[73];
  assign _EVAL_3927 = _EVAL_3402 & _EVAL_2305;
  assign _EVAL_916 = _EVAL_1942[85];
  assign _EVAL_1645 = _EVAL_3402 & _EVAL_916;
  assign _EVAL_4033 = _EVAL_1645 & _EVAL_246;
  assign _EVAL_2614 = _EVAL_4033 & _EVAL_1996;
  assign _EVAL_3770 = _EVAL_3059 & _EVAL_2252;
  assign _EVAL_3229 = _EVAL_1545 & _EVAL_2375;
  assign _EVAL_3241 = _EVAL_2124[8];
  assign _EVAL_3537 = _EVAL_2804 & _EVAL_3241;
  assign _EVAL_3051 = _EVAL_3075 & _EVAL_3779;
  assign _EVAL_3575 = _EVAL_3402 & _EVAL_1383;
  assign _EVAL_1629 = _EVAL_3575 & _EVAL_246;
  assign _EVAL_1166 = _EVAL_1034 & _EVAL_2339;
  assign _EVAL_3062 = _EVAL_3059 & _EVAL_2528;
  assign _EVAL_2273 = _EVAL_3062 & _EVAL_2267;
  assign _EVAL_2450 = _EVAL_2273 & _EVAL_1910;
  assign _EVAL_302 = _EVAL_1942[117];
  assign _EVAL_2914 = _EVAL_3402 & _EVAL_302;
  assign _EVAL_1542 = _EVAL_2914 & _EVAL_246;
  assign _EVAL_2980 = _EVAL_1542 & _EVAL_1996;
  assign _EVAL_3767 = _EVAL_1724 & _EVAL_1145;
  assign _EVAL_3821 = _EVAL_1942[69];
  assign _EVAL_3352 = _EVAL_3402 & _EVAL_3821;
  assign _EVAL_655 = _EVAL_2124[15];
  assign _EVAL_3937 = _EVAL_1279 & _EVAL_655;
  assign _EVAL_400 = _EVAL_2986 & _EVAL_2961;
  assign _EVAL_1490 = _EVAL_1377[18];
  assign _EVAL_764 = _EVAL_1470 & _EVAL_1490;
  assign _EVAL_2195 = _EVAL_1942[102];
  assign _EVAL_801 = _EVAL_3402 & _EVAL_2195;
  assign _EVAL_1143 = _EVAL_3402 & _EVAL_1476;
  assign _EVAL_2012 = _EVAL_1942[16];
  assign _EVAL_2108 = _EVAL_3781 & _EVAL_2012;
  assign _EVAL_2808 = _EVAL_1942[15];
  assign _EVAL_2442 = _EVAL_3059 & _EVAL_353;
  assign _EVAL_3405 = _EVAL_2442 & _EVAL_2267;
  assign _EVAL_2943 = _EVAL_3781 & _EVAL_3347;
  assign _EVAL_411 = _EVAL_1942[104];
  assign _EVAL_3394 = _EVAL_3402 & _EVAL_411;
  assign _EVAL_3678 = _EVAL_3394 & _EVAL_246;
  assign _EVAL_2665 = _EVAL_3059 & _EVAL_2947;
  assign _EVAL_3974 = _EVAL_2665 & _EVAL_2267;
  assign _EVAL_3969 = _EVAL_3974 & _EVAL_1910;
  assign _EVAL_2078 = _EVAL_3059 & _EVAL_3628;
  assign _EVAL_941 = _EVAL_3402 & _EVAL_637;
  assign _EVAL_2874 = _EVAL_941 & _EVAL_246;
  assign _EVAL_3249 = _EVAL_2874 & _EVAL_2544;
  assign _EVAL_2613 = _EVAL_3059 & _EVAL_1613;
  assign _EVAL_264 = _EVAL_2613 & _EVAL_2267;
  assign _EVAL_1940 = _EVAL_1942[118];
  assign _EVAL_1947 = _EVAL_1942[74];
  assign _EVAL_3145 = _EVAL_2124[20];
  assign _EVAL_1670 = _EVAL_2112 & _EVAL_3145;
  assign _EVAL_1823 = _EVAL_1942[57];
  assign _EVAL_2249 = _EVAL_3402 & _EVAL_1823;
  assign _EVAL_1524 = _EVAL_2249 & _EVAL_246;
  assign _EVAL_2285 = _EVAL_933 & _EVAL_2544;
  assign _EVAL_424 = _EVAL_1377[16];
  assign _EVAL_646 = _EVAL_3897 & _EVAL_424;
  assign _EVAL_2830 = _EVAL_1377[29];
  assign _EVAL_984 = _EVAL_1470 & _EVAL_2830;
  assign _EVAL_3746 = _EVAL_3235 > 7'h8;
  assign _EVAL_2960 = _EVAL_3402 & _EVAL_356;
  assign _EVAL_1054 = _EVAL_2960 & _EVAL_246;
  assign _EVAL_4012 = _EVAL_2124[1];
  assign _EVAL_3369 = _EVAL_1279 & _EVAL_4012;
  assign _EVAL_1885 = _EVAL_1377 != 32'h0;
  assign _EVAL_639 = _EVAL_1377[31:3];
  assign _EVAL_2470 = _EVAL_1942[125];
  assign _EVAL_1631 = _EVAL_3781 & _EVAL_2470;
  assign _EVAL_1423 = _EVAL_1631 & _EVAL_246;
  assign _EVAL_856 = _EVAL_1423 & _EVAL_1417;
  assign _EVAL_819 = _EVAL_1857 & _EVAL_3285;
  assign _EVAL_289 = _EVAL_1942[21];
  assign _EVAL_2605 = _EVAL_3402 & _EVAL_289;
  assign _EVAL_405 = _EVAL_2605 & _EVAL_246;
  assign _EVAL_1860 = _EVAL_405 & _EVAL_1996;
  assign _EVAL_2489 = _EVAL_1942[58];
  assign _EVAL_2702 = _EVAL_1942[513];
  assign _EVAL_3835 = _EVAL_3781 & _EVAL_2702;
  assign _EVAL_1969 = _EVAL_3835 & _EVAL_246;
  assign _EVAL_1982 = _EVAL_1545 & _EVAL_3470;
  assign _EVAL_1102 = _EVAL_1942[70];
  assign _EVAL_2465 = _EVAL_1942[111];
  assign _EVAL_909 = _EVAL_3402 & _EVAL_2465;
  assign _EVAL_1686 = _EVAL_909 & _EVAL_246;
  assign _EVAL_1854 = _EVAL_1686 & _EVAL_1996;
  assign _EVAL_478 = _EVAL_1942[107];
  assign _EVAL_1258 = _EVAL_1942[12];
  assign _EVAL_546 = _EVAL_3059 & _EVAL_3489;
  assign _EVAL_1017 = _EVAL_546 & _EVAL_2267;
  assign _EVAL_3171 = _EVAL_1017 & _EVAL_1910;
  assign _EVAL_3054 = _EVAL_1942[110];
  assign _EVAL_633 = _EVAL_3402 & _EVAL_3054;
  assign _EVAL_3818 = _EVAL_3059 & _EVAL_851;
  assign _EVAL_234 = _EVAL_3818 & _EVAL_2267;
  assign _EVAL_202 = _EVAL_234 & _EVAL_1910;
  assign _EVAL_2398 = _EVAL_3059 & _EVAL_455;
  assign _EVAL_3001 = _EVAL_2398 & _EVAL_2267;
  assign _EVAL_876 = _EVAL_3001 & _EVAL_1910;
  assign _EVAL_2873 = _EVAL_105 == 1'h0;
  assign _EVAL_2383 = _EVAL_3781 & _EVAL_3652;
  assign _EVAL_2276 = _EVAL_2383 & _EVAL_246;
  assign _EVAL_2030 = _EVAL_2276 & _EVAL_1417;
  assign _EVAL_1119 = _EVAL_1377[7:1];
  assign _EVAL_3953 = _EVAL_1119 != 7'h0;
  assign _EVAL_3716 = _EVAL_3140 & _EVAL_3953;
  assign _EVAL_1404 = _EVAL_801 & _EVAL_246;
  assign _EVAL_2433 = _EVAL_1942[1];
  assign _EVAL_3230 = _EVAL_3402 & _EVAL_2433;
  assign _EVAL_3782 = _EVAL_3230 & _EVAL_246;
  assign _EVAL_2009 = _EVAL_3782 & _EVAL_1996;
  assign _EVAL_3619 = _EVAL_1279 & _EVAL_1048;
  assign _EVAL_1481 = _EVAL_1942[59];
  assign _EVAL_522 = _EVAL_3059 & _EVAL_1880;
  assign _EVAL_1642 = _EVAL_1143 & _EVAL_246;
  assign _EVAL_1595 = _EVAL_1642 & _EVAL_1996;
  assign _EVAL_1809 = _EVAL_1942[90];
  assign _EVAL_969 = _EVAL_3402 & _EVAL_1809;
  assign _EVAL_661 = _EVAL_969 & _EVAL_246;
  assign _EVAL_1026 = _EVAL_1942[27];
  assign _EVAL_848 = _EVAL_3781 & _EVAL_1026;
  assign _EVAL_2724 = _EVAL_848 & _EVAL_246;
  assign _EVAL_2541 = _EVAL_3059 & _EVAL_3069;
  assign _EVAL_523 = _EVAL_2541 & _EVAL_2267;
  assign _EVAL_2622 = _EVAL_2804 & _EVAL_3180;
  assign _EVAL_2693 = _EVAL_1470 & _EVAL_2375;
  assign _EVAL_2993 = _EVAL_1470 & _EVAL_1621;
  assign _EVAL_169 = _EVAL_1377[17];
  assign _EVAL_2201 = _EVAL_3458 & _EVAL_169;
  assign _EVAL_554 = _EVAL_2112 & _EVAL_3596;
  assign _EVAL_3616 = _EVAL_3059 & _EVAL_2543;
  assign _EVAL_3528 = _EVAL_3402 & _EVAL_2012;
  assign _EVAL_465 = _EVAL_3528 & _EVAL_246;
  assign _EVAL_2401 = _EVAL_3458 & _EVAL_543;
  assign _EVAL_978 = _EVAL_1942[63];
  assign _EVAL_3190 = _EVAL_3402 & _EVAL_978;
  assign _EVAL_3653 = _EVAL_3190 & _EVAL_246;
  assign _EVAL_3119 = _EVAL_3653 & _EVAL_1996;
  assign _EVAL_1781 = _EVAL_3059 & _EVAL_926;
  assign _EVAL_598 = _EVAL_1781 & _EVAL_2267;
  assign _EVAL_3699 = _EVAL_3781 & _EVAL_1172;
  assign _EVAL_2954 = _EVAL_3402 & _EVAL_2702;
  assign _EVAL_2611 = _EVAL_3059 & _EVAL_3043;
  assign _EVAL_3807 = _EVAL_3059 & _EVAL_415;
  assign _EVAL_3052 = _EVAL_3402 & _EVAL_3664;
  assign _EVAL_1203 = _EVAL_2804 & _EVAL_1224;
  assign _EVAL_1761 = _EVAL_1942[52];
  assign _EVAL_1620 = _EVAL_3781 & _EVAL_1761;
  assign _EVAL_1103 = _EVAL_1620 & _EVAL_246;
  assign _EVAL_3648 = _EVAL_1103 & _EVAL_1417;
  assign _EVAL_2658 = _EVAL_3781 & _EVAL_2676;
  assign _EVAL_1004 = _EVAL_2658 & _EVAL_246;
  assign _EVAL_3328 = _EVAL_1004 & _EVAL_1417;
  assign _EVAL_2194 = _EVAL_3059 & _EVAL_3318;
  assign _EVAL_536 = _EVAL_1942[71];
  assign _EVAL_3462 = _EVAL_3402 & _EVAL_536;
  assign _EVAL_241 = _EVAL_3462 & _EVAL_246;
  assign _EVAL_724 = _EVAL_1377[3];
  assign _EVAL_3481 = _EVAL_3897 & _EVAL_724;
  assign _EVAL_3574 = _EVAL_3405 & _EVAL_1910;
  assign _EVAL_418 = _EVAL_3059 & _EVAL_318;
  assign _EVAL_2985 = _EVAL_418 & _EVAL_2267;
  assign _EVAL_3071 = _EVAL_1942[106];
  assign _EVAL_2741 = _EVAL_3402 & _EVAL_3071;
  assign _EVAL_3320 = _EVAL_2741 & _EVAL_246;
  assign _EVAL_1534 = _EVAL_431 & _EVAL_3363;
  assign _EVAL_2420 = _EVAL_1942[66];
  assign _EVAL_1923 = _EVAL_3402 & _EVAL_2420;
  assign _EVAL_1128 = _EVAL_1923 & _EVAL_246;
  assign _EVAL_3411 = _EVAL_1128 & _EVAL_1996;
  assign _EVAL_1950 = _EVAL_3781 & _EVAL_1102;
  assign _EVAL_1106 = _EVAL_1950 & _EVAL_246;
  assign _EVAL_1431 = _EVAL_1470 & _EVAL_3000;
  assign _EVAL_168 = _EVAL_1040 & _EVAL_2691;
  assign _EVAL_3613 = _EVAL_1942[75];
  assign _EVAL_3827 = _EVAL_3402 & _EVAL_3613;
  assign _EVAL_336 = _EVAL_3827 & _EVAL_246;
  assign _EVAL_3933 = _EVAL_3059 & _EVAL_1820;
  assign _EVAL_2805 = _EVAL_3933 & _EVAL_2267;
  assign _EVAL_1405 = _EVAL_3059 & _EVAL_1648;
  assign _EVAL_1099 = _EVAL_1405 & _EVAL_2267;
  assign _EVAL_2176 = _EVAL_1034 & _EVAL_3701;
  assign _EVAL_2979 = _EVAL_3059 & _EVAL_1230;
  assign _EVAL_3960 = _EVAL_2979 & _EVAL_2267;
  assign _EVAL_2181 = _EVAL_3059 & _EVAL_985;
  assign _EVAL_181 = _EVAL_2181 & _EVAL_2267;
  assign _EVAL_1884 = _EVAL_639 != 29'h0;
  assign _EVAL_2647 = _EVAL_1857 & _EVAL_2984;
  assign _EVAL_2386 = _EVAL_3781 & _EVAL_2305;
  assign _EVAL_2951 = _EVAL_2386 & _EVAL_246;
  assign _EVAL_872 = _EVAL_2951 & _EVAL_1417;
  assign _EVAL_3345 = _EVAL_1279 & _EVAL_4016;
  assign _EVAL_1369 = _EVAL_1942[38];
  assign _EVAL_772 = _EVAL_3781 & _EVAL_1369;
  assign _EVAL_1920 = _EVAL_772 & _EVAL_246;
  assign _EVAL_778 = _EVAL_1942[114];
  assign _EVAL_1872 = _EVAL_1666 & _EVAL_246;
  assign _EVAL_3789 = _EVAL_3781 & _EVAL_2650;
  assign _EVAL_3151 = _EVAL_3789 & _EVAL_246;
  assign _EVAL_3406 = {1'h1,_EVAL_663};
  assign _EVAL_813 = _EVAL_3402 & _EVAL_1989;
  assign _EVAL_1791 = _EVAL_1942[108];
  assign _EVAL_357 = _EVAL_3781 & _EVAL_1791;
  assign _EVAL_365 = _EVAL_790 & _EVAL_1417;
  assign _EVAL_814 = _EVAL_2525 & _EVAL_246;
  assign _EVAL_935 = _EVAL_3059 & _EVAL_886;
  assign _EVAL_2182 = _EVAL_1545 & _EVAL_1145;
  assign _EVAL_2016 = _EVAL_3781 & _EVAL_1823;
  assign _EVAL_3438 = _EVAL_2016 & _EVAL_246;
  assign _EVAL_2373 = _EVAL_3377 & _EVAL_1996;
  assign _EVAL_2284 = _EVAL_1040 & _EVAL_1145;
  assign _EVAL_145 = _EVAL_3781 & _EVAL_2978;
  assign _EVAL_992 = _EVAL_1034 & _EVAL_3471;
  assign _EVAL_977 = _EVAL_3781 & _EVAL_289;
  assign _EVAL_255 = _EVAL_3402 & _EVAL_3218;
  assign _EVAL_2778 = _EVAL_255 & _EVAL_246;
  assign _EVAL_2259 = _EVAL_1942[93];
  assign _EVAL_3848 = _EVAL_3402 & _EVAL_2259;
  assign _EVAL_297 = _EVAL_1942[62];
  assign _EVAL_2205 = _EVAL_1942[122];
  assign _EVAL_2342 = _EVAL_3402 & _EVAL_2205;
  assign _EVAL_475 = _EVAL_814 & _EVAL_1996;
  assign _EVAL_1581 = _EVAL_2112 & _EVAL_2072;
  assign _EVAL_2587 = _EVAL_2124[30];
  assign _EVAL_404 = _EVAL_2804 & _EVAL_2587;
  assign _EVAL_3210 = _EVAL_3781 & _EVAL_2195;
  assign _EVAL_3087 = _EVAL_2124[3];
  assign _EVAL_3656 = _EVAL_2112 & _EVAL_3087;
  assign _EVAL_3565 = _EVAL_3402 & _EVAL_1369;
  assign _EVAL_1140 = _EVAL_1724 & _EVAL_169;
  assign _EVAL_2253 = _EVAL_3402 & _EVAL_1026;
  assign _EVAL_1110 = _EVAL_2253 & _EVAL_246;
  assign _EVAL_3511 = _EVAL_1110 & _EVAL_1996;
  assign _EVAL_949 = _EVAL_431 & _EVAL_1224;
  assign _EVAL_2923 = _EVAL_3059 & _EVAL_4041;
  assign _EVAL_2376 = _EVAL_2923 & _EVAL_2267;
  assign _EVAL_2506 = _EVAL_1119 == 7'h7f;
  assign _EVAL_3514 = _EVAL_1942[86];
  assign _EVAL_567 = _EVAL_3781 & _EVAL_3514;
  assign _EVAL_2831 = _EVAL_567 & _EVAL_246;
  assign _EVAL_3829 = _EVAL_3059 & _EVAL_4040;
  assign _EVAL_3120 = _EVAL_3829 & _EVAL_2267;
  assign _EVAL_697 = _EVAL_3120 & _EVAL_1910;
  assign _EVAL_1976 = _EVAL_3059 & _EVAL_2731;
  assign _EVAL_1544 = _EVAL_1106 & _EVAL_1417;
  assign _EVAL_4023 = _EVAL_1522 & _EVAL_424;
  assign _EVAL_384 = _EVAL_3781 & _EVAL_3272;
  assign _EVAL_1192 = _EVAL_384 & _EVAL_246;
  assign _EVAL_210 = _EVAL_3781 & _EVAL_204;
  assign _EVAL_3016 = _EVAL_210 & _EVAL_246;
  assign _EVAL_863 = _EVAL_3016 & _EVAL_1417;
  assign _EVAL_300 = _EVAL_1942[29];
  assign _EVAL_1921 = _EVAL_3402 & _EVAL_300;
  assign _EVAL_3067 = _EVAL_1522 & _EVAL_2984;
  assign _EVAL_3173 = _EVAL_1942[19];
  assign _EVAL_3717 = _EVAL_3781 & _EVAL_3173;
  assign _EVAL_3542 = _EVAL_3402 & _EVAL_3397;
  assign _EVAL_2780 = _EVAL_3542 & _EVAL_246;
  assign _EVAL_568 = _EVAL_2780 & _EVAL_1996;
  assign _EVAL_3332 = _EVAL_1689 & _EVAL_246;
  assign _EVAL_2755 = _EVAL_3332 & _EVAL_1417;
  assign _EVAL_2294 = _EVAL_3059 & _EVAL_1502;
  assign _EVAL_1420 = _EVAL_2294 & _EVAL_2267;
  assign _EVAL_3036 = _EVAL_1942[53];
  assign _EVAL_2332 = _EVAL_1522 & _EVAL_1490;
  assign _EVAL_2922 = _EVAL_3059 & _EVAL_226;
  assign _EVAL_2322 = _EVAL_2922 & _EVAL_2267;
  assign _EVAL_953 = _EVAL_3516 & _EVAL_2267;
  assign _EVAL_2413 = _EVAL_953 & _EVAL_1910;
  assign _EVAL_2657 = _EVAL_2986 & _EVAL_1048;
  assign _EVAL_1867 = _EVAL_3059 & _EVAL_3981;
  assign _EVAL_3894 = _EVAL_3402 & _EVAL_1102;
  assign _EVAL_1514 = _EVAL_1470 & _EVAL_2594;
  assign _EVAL_3611 = _EVAL_3059 & _EVAL_3094;
  assign _EVAL_3387 = _EVAL_357 & _EVAL_246;
  assign _EVAL_2620 = _EVAL_3387 & _EVAL_1417;
  assign _EVAL_1963 = _EVAL_2124[16];
  assign _EVAL_2829 = _EVAL_2986 & _EVAL_1963;
  assign _EVAL_1897 = _EVAL_3059 & _EVAL_3873;
  assign _EVAL_3079 = _EVAL_1897 & _EVAL_2267;
  assign _EVAL_2395 = _EVAL_3079 & _EVAL_1910;
  assign _EVAL_2337 = _EVAL_1553 & _EVAL_3596;
  assign _EVAL_3530 = _EVAL_3059 & _EVAL_1634;
  assign _EVAL_3306 = _EVAL_1942[45];
  assign _EVAL_3451 = _EVAL_3402 & _EVAL_3306;
  assign _EVAL_2258 = _EVAL_3451 & _EVAL_246;
  assign _EVAL_2162 = _EVAL_3568 & _EVAL_2267;
  assign _EVAL_2402 = _EVAL_2162 & _EVAL_1910;
  assign _EVAL_3949 = _EVAL_3402 & _EVAL_1053;
  assign _EVAL_3378 = _EVAL_3949 & _EVAL_246;
  assign _EVAL_3725 = _EVAL_3378 & _EVAL_1996;
  assign _EVAL_1191 = _EVAL_3059 & _EVAL_3882;
  assign _EVAL_2694 = _EVAL_1191 & _EVAL_2267;
  assign _EVAL_2498 = _EVAL_3402 & _EVAL_1481;
  assign _EVAL_3339 = _EVAL_2498 & _EVAL_246;
  assign _EVAL_330 = _EVAL_3339 & _EVAL_1996;
  assign _EVAL_2906 = _EVAL_3458 & _EVAL_1324;
  assign _EVAL_3038 = _EVAL_1377[22];
  assign _EVAL_2632 = _EVAL_1040 & _EVAL_3038;
  assign _EVAL_1683 = _EVAL_1553 & _EVAL_1224;
  assign _EVAL_3599 = _EVAL_2986 & _EVAL_4031;
  assign _EVAL_3934 = _EVAL_1942[112];
  assign _EVAL_2293 = _EVAL_3781 & _EVAL_3934;
  assign _EVAL_728 = _EVAL_3059 & _EVAL_3707;
  assign _EVAL_2580 = _EVAL_728 & _EVAL_2267;
  assign _EVAL_767 = _EVAL_2580 & _EVAL_1910;
  assign _EVAL_1575 = _EVAL_1942[87];
  assign _EVAL_1312 = _EVAL_3402 & _EVAL_1575;
  assign _EVAL_504 = _EVAL_3781 & _EVAL_536;
  assign _EVAL_883 = _EVAL_1942[43];
  assign _EVAL_2530 = _EVAL_1545 & _EVAL_2756;
  assign _EVAL_1745 = _EVAL_3781 & _EVAL_3906;
  assign _EVAL_1836 = _EVAL_1745 & _EVAL_246;
  assign _EVAL_3208 = _EVAL_1836 & _EVAL_1417;
  assign _EVAL_960 = _EVAL_3059 & _EVAL_1432;
  assign _EVAL_243 = _EVAL_960 & _EVAL_2267;
  assign _EVAL_358 = _EVAL_3059 & _EVAL_3679;
  assign _EVAL_3141 = _EVAL_358 & _EVAL_2267;
  assign _EVAL_2444 = _EVAL_3781 & _EVAL_2497;
  assign _EVAL_2792 = _EVAL_1942[46];
  assign _EVAL_2061 = _EVAL_1942[11];
  assign _EVAL_2516 = _EVAL_3781 & _EVAL_2061;
  assign _EVAL_3095 = _EVAL_1942[103];
  assign _EVAL_474 = _EVAL_3402 & _EVAL_3095;
  assign _EVAL_2711 = _EVAL_474 & _EVAL_246;
  assign _EVAL_1609 = _EVAL_1942[6];
  assign _EVAL_2576 = _EVAL_3402 & _EVAL_1609;
  assign _EVAL_547 = _EVAL_2576 & _EVAL_246;
  assign _EVAL_1937 = _EVAL_547 & _EVAL_1996;
  assign _EVAL_3806 = _EVAL_3270 & _EVAL_2267;
  assign _EVAL_470 = _EVAL_3806 & _EVAL_1910;
  assign _EVAL_685 = _EVAL_1034 & _EVAL_4012;
  assign _EVAL_3836 = _EVAL_3059 & _EVAL_2189;
  assign _EVAL_566 = _EVAL_1942[105];
  assign _EVAL_784 = _EVAL_1040 & _EVAL_2594;
  assign _EVAL_3319 = _EVAL_1942[77];
  assign _EVAL_1491 = _EVAL_3402 & _EVAL_3319;
  assign _EVAL_279 = _EVAL_1491 & _EVAL_246;
  assign _EVAL_656 = _EVAL_279 & _EVAL_1996;
  assign _EVAL_4065 = _EVAL_1942[84];
  assign _EVAL_2667 = _EVAL_3781 & _EVAL_4065;
  assign _EVAL_2636 = _EVAL_2667 & _EVAL_246;
  assign _EVAL_3735 = _EVAL_3402 & _EVAL_3036;
  assign _EVAL_696 = _EVAL_2124[29];
  assign _EVAL_1484 = _EVAL_1279 & _EVAL_696;
  assign _EVAL_2331 = _EVAL_3059 & _EVAL_1922;
  assign _EVAL_2196 = _EVAL_2331 & _EVAL_2267;
  assign _EVAL_3737 = _EVAL_1976 & _EVAL_2267;
  assign _EVAL_1322 = _EVAL_3402 & _EVAL_2042;
  assign _EVAL_3440 = _EVAL_1322 & _EVAL_246;
  assign _EVAL_657 = _EVAL_3781 & _EVAL_669;
  assign _EVAL_1618 = _EVAL_657 & _EVAL_246;
  assign _EVAL_1800 = _EVAL_1942[48];
  assign _EVAL_2040 = _EVAL_3402 & _EVAL_1800;
  assign _EVAL_3441 = _EVAL_3781 & _EVAL_3821;
  assign _EVAL_1016 = _EVAL_3441 & _EVAL_246;
  assign _EVAL_686 = _EVAL_465 & _EVAL_1996;
  assign _EVAL_1895 = _EVAL_3807 & _EVAL_2267;
  assign _EVAL_3408 = _EVAL_3372 != 8'h0;
  assign _EVAL_1766 = _EVAL_1895 & _EVAL_3408;
  assign _EVAL_887 = _EVAL_1377[1];
  assign _EVAL_2087 = _EVAL_3897 & _EVAL_887;
  assign _EVAL_849 = _EVAL_1942[28];
  assign _EVAL_2726 = _EVAL_3402 & _EVAL_849;
  assign _EVAL_3968 = _EVAL_2726 & _EVAL_246;
  assign _EVAL_498 = _EVAL_3968 & _EVAL_1996;
  assign _EVAL_3982 = _EVAL_2112 & _EVAL_2043;
  assign _EVAL_1415 = _EVAL_3059 & _EVAL_260;
  assign _EVAL_1817 = _EVAL_1415 & _EVAL_2267;
  assign _EVAL_3480 = _EVAL_1817 & _EVAL_1910;
  assign _EVAL_3771 = _EVAL_3059 & _EVAL_515;
  assign _EVAL_2044 = _EVAL_3771 & _EVAL_2267;
  assign _EVAL_3845 = _EVAL_933 & _EVAL_2283;
  assign _EVAL_2326 = _EVAL_2804 & _EVAL_3701;
  assign _EVAL_1426 = _EVAL_3781 & _EVAL_300;
  assign _EVAL_1310 = _EVAL_1629 & _EVAL_1996;
  assign _EVAL_1949 = _EVAL_2322 & _EVAL_1910;
  assign _EVAL_2757 = _EVAL_3059 & _EVAL_2743;
  assign _EVAL_1636 = _EVAL_1724 & _EVAL_3954;
  assign _EVAL_763 = _EVAL_2943 & _EVAL_246;
  assign _EVAL_999 = _EVAL_1942[49];
  assign _EVAL_3326 = _EVAL_1942[17];
  assign _EVAL_869 = _EVAL_3781 & _EVAL_3326;
  assign _EVAL_3162 = _EVAL_869 & _EVAL_246;
  assign _EVAL_1263 = _EVAL_3894 & _EVAL_246;
  assign _EVAL_3366 = _EVAL_1263 & _EVAL_1996;
  assign _EVAL_2348 = _EVAL_1034 & _EVAL_3241;
  assign _EVAL_2379 = _EVAL_1942[83];
  assign _EVAL_332 = _EVAL_3781 & _EVAL_2379;
  assign _EVAL_499 = _EVAL_332 & _EVAL_246;
  assign _EVAL_1538 = _EVAL_3059 & _EVAL_1439;
  assign _EVAL_3257 = _EVAL_1522 & _EVAL_2830;
  assign _EVAL_3209 = _EVAL_2124[7];
  assign _EVAL_2740 = _EVAL_2986 & _EVAL_3209;
  assign _EVAL_1705 = _EVAL_694 & _EVAL_2267;
  assign _EVAL_2396 = _EVAL_1705 & _EVAL_1910;
  assign _EVAL_494 = _EVAL_3402 & _EVAL_1940;
  assign _EVAL_3805 = _EVAL_494 & _EVAL_246;
  assign _EVAL_1829 = _EVAL_2986 & _EVAL_2339;
  assign _EVAL_3730 = _EVAL_1681 & _EVAL_1417;
  assign _EVAL_2706 = _EVAL_3059 & _EVAL_1216;
  assign _EVAL_501 = _EVAL_2706 & _EVAL_2267;
  assign _EVAL_2820 = _EVAL_3402 & _EVAL_2990;
  assign _EVAL_3582 = _EVAL_3059 & _EVAL_2644;
  assign _EVAL_1748 = _EVAL_3402 & _EVAL_1643;
  assign _EVAL_550 = _EVAL_1748 & _EVAL_246;
  assign _EVAL_432 = _EVAL_550 & _EVAL_1996;
  assign _EVAL_179 = _EVAL_1470 & _EVAL_887;
  assign _EVAL_198 = _EVAL_3059 & _EVAL_3101;
  assign _EVAL_1577 = _EVAL_198 & _EVAL_2267;
  assign _EVAL_3876 = _EVAL_1553 & _EVAL_3145;
  assign _EVAL_398 = _EVAL_2124[17];
  assign _EVAL_3368 = _EVAL_1553 & _EVAL_398;
  assign _EVAL_324 = _EVAL_1942[36];
  assign _EVAL_3791 = _EVAL_3781 & _EVAL_324;
  assign _EVAL_4035 = _EVAL_3791 & _EVAL_246;
  assign _EVAL_284 = _EVAL_3059 & _EVAL_1325;
  assign _EVAL_2928 = _EVAL_284 & _EVAL_2267;
  assign _EVAL_2221 = _EVAL_3059 & _EVAL_3350;
  assign _EVAL_1883 = _EVAL_2221 & _EVAL_2267;
  assign _EVAL_904 = _EVAL_1724 & _EVAL_1868;
  assign _EVAL_340 = _EVAL_2078 & _EVAL_2267;
  assign _EVAL_2145 = _EVAL_3059 & _EVAL_2567;
  assign _EVAL_3631 = _EVAL_3781 & _EVAL_2489;
  assign _EVAL_3697 = _EVAL_3631 & _EVAL_246;
  assign _EVAL_440 = _EVAL_1724 & _EVAL_3285;
  assign _EVAL_687 = _EVAL_3059 & _EVAL_3088;
  assign _EVAL_635 = _EVAL_3897 & _EVAL_1354;
  assign _EVAL_2236 = _EVAL_3897 & _EVAL_1324;
  assign _EVAL_2508 = _EVAL_3059 & _EVAL_938;
  assign _EVAL_2363 = _EVAL_2508 & _EVAL_2267;
  assign _EVAL_3189 = _EVAL_2363 & _EVAL_1910;
  assign _EVAL_3633 = _EVAL_2196 & _EVAL_1910;
  assign _EVAL_931 = _EVAL_3735 & _EVAL_246;
  assign _EVAL_442 = _EVAL_3402 & _EVAL_1381;
  assign _EVAL_1455 = _EVAL_3781 & _EVAL_1940;
  assign _EVAL_319 = _EVAL_3075 & _EVAL_4012;
  assign _EVAL_538 = _EVAL_2040 & _EVAL_246;
  assign _EVAL_2540 = _EVAL_538 & _EVAL_1996;
  assign _EVAL_1792 = _EVAL_3402 & _EVAL_204;
  assign _EVAL_3294 = _EVAL_1942[24];
  assign _EVAL_2407 = _EVAL_3781 & _EVAL_3294;
  assign _EVAL_1983 = _EVAL_2407 & _EVAL_246;
  assign _EVAL_719 = _EVAL_1983 & _EVAL_1417;
  assign _EVAL_564 = _EVAL_2986 & _EVAL_3701;
  assign _EVAL_1155 = _EVAL_1078 & _EVAL_246;
  assign _EVAL_1248 = _EVAL_3402 & _EVAL_1258;
  assign _EVAL_2403 = _EVAL_1248 & _EVAL_246;
  assign _EVAL_1935 = _EVAL_3402 & _EVAL_3790;
  assign _EVAL_232 = _EVAL_1935 & _EVAL_246;
  assign _EVAL_3872 = _EVAL_1942[116];
  assign _EVAL_2203 = _EVAL_3402 & _EVAL_3872;
  assign _EVAL_2086 = _EVAL_2203 & _EVAL_246;
  assign _EVAL_2534 = _EVAL_2086 & _EVAL_1996;
  assign _EVAL_2836 = _EVAL_2293 & _EVAL_246;
  assign _EVAL_2679 = _EVAL_1279 & _EVAL_4031;
  assign _EVAL_920 = _EVAL_3055 != 8'h0;
  assign _EVAL_2412 = _EVAL_1377[30];
  assign _EVAL_1715 = _EVAL_3458 & _EVAL_2412;
  assign _EVAL_3742 = _EVAL_1857 & _EVAL_887;
  assign _EVAL_1089 = _EVAL_3075 & _EVAL_696;
  assign _EVAL_752 = _EVAL_1040 & _EVAL_2756;
  assign _EVAL_3217 = _EVAL_1371 != 8'h0;
  assign _EVAL_2428 = _EVAL_1398 & _EVAL_3217;
  assign _EVAL_2522 = _EVAL_3059 & _EVAL_1948;
  assign _EVAL_3702 = _EVAL_2522 & _EVAL_2267;
  assign _EVAL_2859 = _EVAL_3059 & _EVAL_3287;
  assign _EVAL_1814 = _EVAL_2859 & _EVAL_2267;
  assign _EVAL_2783 = _EVAL_1814 & _EVAL_1910;
  assign _EVAL_2547 = _EVAL_1857 & _EVAL_2412;
  assign _EVAL_328 = _EVAL_598 & _EVAL_1910;
  assign _EVAL_3819 = _EVAL_1990 & _EVAL_3861;
  assign _EVAL_1437 = _EVAL_3402 & _EVAL_3468;
  assign _EVAL_3089 = _EVAL_1279 & _EVAL_3087;
  assign _EVAL_500 = _EVAL_1522 & _EVAL_2412;
  assign _EVAL_1926 = _EVAL_3059 & _EVAL_3847;
  assign _EVAL_211 = _EVAL_1942[80];
  assign _EVAL_2721 = _EVAL_3781 & _EVAL_211;
  assign _EVAL_823 = _EVAL_2721 & _EVAL_246;
  assign _EVAL_1274 = _EVAL_3781 & _EVAL_3295;
  assign _EVAL_1813 = _EVAL_1942[51];
  assign _EVAL_3290 = _EVAL_3781 & _EVAL_1813;
  assign _EVAL_388 = _EVAL_695 != 8'h0;
  assign _EVAL_2577 = _EVAL_3736 & _EVAL_388;
  assign _EVAL_3467 = _EVAL_2145 & _EVAL_2267;
  assign _EVAL_1188 = _EVAL_3467 & _EVAL_1910;
  assign _EVAL_2029 = _EVAL_3052 & _EVAL_246;
  assign _EVAL_1314 = _EVAL_2029 & _EVAL_1996;
  assign _EVAL_892 = _EVAL_181 & _EVAL_1910;
  assign _EVAL_2021 = _EVAL_3402 & _EVAL_778;
  assign _EVAL_446 = _EVAL_2021 & _EVAL_246;
  assign _EVAL_2323 = _EVAL_446 & _EVAL_1996;
  assign _EVAL_3935 = _EVAL_1034 & _EVAL_806;
  assign _EVAL_1612 = _EVAL_3582 & _EVAL_2267;
  assign _EVAL_413 = _EVAL_1612 & _EVAL_1910;
  assign _EVAL_2919 = _EVAL_1942[95];
  assign _EVAL_2793 = _EVAL_3781 & _EVAL_2712;
  assign _EVAL_2884 = _EVAL_2793 & _EVAL_246;
  assign _EVAL_2795 = _EVAL_3238 == 1'h0;
  assign _EVAL_1561 = _EVAL_3059 & _EVAL_3932;
  assign _EVAL_2643 = _EVAL_431 & _EVAL_3209;
  assign _EVAL_3863 = _EVAL_1545 & _EVAL_1868;
  assign _EVAL_3962 = _EVAL_3402 & _EVAL_883;
  assign _EVAL_3643 = _EVAL_3962 & _EVAL_246;
  assign _EVAL_3501 = _EVAL_1553 & _EVAL_215;
  assign _EVAL_3684 = _EVAL_3781 & _EVAL_1609;
  assign _EVAL_575 = _EVAL_3684 & _EVAL_246;
  assign _EVAL_1464 = _EVAL_575 & _EVAL_1417;
  assign _EVAL_3797 = _EVAL_3059 & _EVAL_1833;
  assign _EVAL_1409 = _EVAL_3797 & _EVAL_2267;
  assign _EVAL_2419 = _EVAL_1409 & _EVAL_1910;
  assign _EVAL_3634 = _EVAL_3059 & _EVAL_939;
  assign _EVAL_333 = _EVAL_1744 & _EVAL_1417;
  assign _EVAL_2080 = _EVAL_3059 & _EVAL_308;
  assign _EVAL_1743 = _EVAL_431 & _EVAL_1889;
  assign _EVAL_3809 = _EVAL_3781 & _EVAL_2433;
  assign _EVAL_1729 = _EVAL_3809 & _EVAL_246;
  assign _EVAL_2393 = _EVAL_1729 & _EVAL_1417;
  assign _EVAL_1480 = _EVAL_3059 & _EVAL_2742;
  assign _EVAL_1616 = _EVAL_241 & _EVAL_1996;
  assign _EVAL_3512 = _EVAL_2812 & _EVAL_2267;
  assign _EVAL_1029 = _EVAL_3402 & _EVAL_1172;
  assign _EVAL_451 = _EVAL_2928 & _EVAL_1910;
  assign _EVAL_2846 = _EVAL_2986 & _EVAL_806;
  assign _EVAL_1554 = _EVAL_1942[7];
  assign _EVAL_705 = _EVAL_3781 & _EVAL_1554;
  assign _EVAL_2357 = _EVAL_705 & _EVAL_246;
  assign _EVAL_1169 = _EVAL_3402 & _EVAL_152;
  assign _EVAL_882 = _EVAL_1169 & _EVAL_246;
  assign _EVAL_2260 = _EVAL_639 == 29'h1fffffff;
  assign _EVAL_1560 = _EVAL_882 & _EVAL_2260;
  assign _EVAL_1646 = _EVAL_1942[35];
  assign _EVAL_3696 = _EVAL_3781 & _EVAL_1646;
  assign _EVAL_3833 = _EVAL_882 & _EVAL_1996;
  assign _EVAL_2344 = _EVAL_2124[31];
  assign _EVAL_1563 = _EVAL_431 & _EVAL_2344;
  assign _EVAL_2933 = _EVAL_3059 & _EVAL_3682;
  assign _EVAL_1869 = _EVAL_2933 & _EVAL_2267;
  assign _EVAL_1340 = _EVAL_504 & _EVAL_246;
  assign _EVAL_1395 = _EVAL_2112 & _EVAL_3363;
  assign _EVAL_597 = _EVAL_3781 & _EVAL_3095;
  assign _EVAL_934 = _EVAL_597 & _EVAL_246;
  assign _EVAL_3449 = _EVAL_934 & _EVAL_1417;
  assign _EVAL_3427 = _EVAL_2831 & _EVAL_1417;
  assign _EVAL_1846 = _EVAL_2820 & _EVAL_246;
  assign _EVAL_2469 = _EVAL_1522 & _EVAL_520;
  assign _EVAL_776 = _EVAL_1942[14];
  assign _EVAL_1782 = _EVAL_3781 & _EVAL_776;
  assign _EVAL_3761 = _EVAL_1942[34];
  assign _EVAL_2452 = _EVAL_3781 & _EVAL_3761;
  assign _EVAL_2949 = _EVAL_2041 & _EVAL_388;
  assign _EVAL_1523 = _EVAL_3781 & _EVAL_297;
  assign _EVAL_468 = _EVAL_1523 & _EVAL_246;
  assign _EVAL_1331 = _EVAL_468 & _EVAL_1417;
  assign _EVAL_2901 = _EVAL_1942[60];
  assign _EVAL_1183 = _EVAL_2986 & _EVAL_1245;
  assign _EVAL_997 = _EVAL_3059 & _EVAL_1013;
  assign _EVAL_3849 = _EVAL_997 & _EVAL_2267;
  assign _EVAL_3333 = _EVAL_1942[72];
  assign _EVAL_3685 = _EVAL_3402 & _EVAL_3333;
  assign _EVAL_435 = _EVAL_1942[31];
  assign _EVAL_1688 = _EVAL_3402 & _EVAL_435;
  assign _EVAL_3032 = _EVAL_1688 & _EVAL_246;
  assign _EVAL_740 = _EVAL_3032 & _EVAL_1996;
  assign _EVAL_2871 = _EVAL_3781 & _EVAL_3319;
  assign _EVAL_1812 = _EVAL_2871 & _EVAL_246;
  assign _EVAL_1787 = _EVAL_3059 & _EVAL_1182;
  assign _EVAL_3980 = _EVAL_1787 & _EVAL_2267;
  assign _EVAL_2689 = _EVAL_935 & _EVAL_2267;
  assign _EVAL_1152 = _EVAL_2689 & _EVAL_1910;
  assign _EVAL_1871 = _EVAL_3781 & _EVAL_3048;
  assign _EVAL_2247 = _EVAL_1871 & _EVAL_246;
  assign _EVAL_3128 = _EVAL_2247 & _EVAL_1417;
  assign _EVAL_2641 = _EVAL_3781 & _EVAL_3872;
  assign _EVAL_1589 = _EVAL_2641 & _EVAL_246;
  assign _EVAL_1691 = _EVAL_2112 & _EVAL_4031;
  assign _EVAL_2900 = _EVAL_1377[15:8];
  assign _EVAL_2456 = _EVAL_2900 == 8'hff;
  assign _EVAL_1296 = _EVAL_3458 & _EVAL_2594;
  assign _EVAL_1158 = _EVAL_3402 & _EVAL_2061;
  assign _EVAL_2240 = _EVAL_1638 & _EVAL_2267;
  assign _EVAL_2891 = _EVAL_1792 & _EVAL_246;
  assign _EVAL_1457 = _EVAL_2891 & _EVAL_1996;
  assign _EVAL_1153 = _EVAL_3736 & _EVAL_920;
  assign _EVAL_526 = _EVAL_2874 & _EVAL_2456;
  assign _EVAL_2457 = _EVAL_2804 & _EVAL_4031;
  assign _EVAL_2606 = _EVAL_3781 & _EVAL_778;
  assign _EVAL_1084 = _EVAL_3320 & _EVAL_1996;
  assign _EVAL_3691 = _EVAL_1990 - 1'h1;
  assign _EVAL_3920 = _EVAL_1377[24];
  assign _EVAL_4000 = _EVAL_3402 & _EVAL_1778;
  assign _EVAL_1603 = _EVAL_4000 & _EVAL_246;
  assign _EVAL_3153 = _EVAL_1603 & _EVAL_1996;
  assign _EVAL_1630 = _EVAL_3059 & _EVAL_3844;
  assign _EVAL_3963 = _EVAL_3781 & _EVAL_3054;
  assign _EVAL_1330 = _EVAL_3963 & _EVAL_246;
  assign _EVAL_1281 = _EVAL_431 & _EVAL_3145;
  assign _EVAL_393 = _EVAL_3402 & _EVAL_2792;
  assign _EVAL_3417 = _EVAL_393 & _EVAL_246;
  assign _EVAL_1576 = _EVAL_1553 & _EVAL_1889;
  assign _EVAL_4060 = _EVAL_3059 & _EVAL_3213;
  assign _EVAL_3524 = _EVAL_4060 & _EVAL_2267;
  assign _EVAL_3395 = _EVAL_3524 & _EVAL_1910;
  assign _EVAL_3635 = _EVAL_1522 & _EVAL_3920;
  assign _EVAL_678 = _EVAL_1724 & _EVAL_2594;
  assign _EVAL_166 = _EVAL_818 & _EVAL_2267;
  assign _EVAL_184 = _EVAL_166 & _EVAL_1910;
  assign _EVAL_803 = _EVAL_2124[6];
  assign _EVAL_2618 = _EVAL_1279 & _EVAL_803;
  assign _EVAL_965 = _EVAL_2804 & _EVAL_2043;
  assign _EVAL_175 = _EVAL_2683 & _EVAL_246;
  assign _EVAL_3986 = _EVAL_175 & _EVAL_1417;
  assign _EVAL_1091 = _EVAL_1857 & _EVAL_1621;
  assign _EVAL_1694 = _EVAL_431 & _EVAL_1963;
  assign _EVAL_2945 = _EVAL_431 & _EVAL_4012;
  assign _EVAL_3600 = _EVAL_1274 & _EVAL_246;
  assign _EVAL_1445 = _EVAL_3075 & _EVAL_655;
  assign _EVAL_2483 = _EVAL_3781 & _EVAL_2259;
  assign _EVAL_1624 = _EVAL_2483 & _EVAL_246;
  assign _EVAL_3654 = _EVAL_1624 & _EVAL_1417;
  assign _EVAL_2280 = _EVAL_2444 & _EVAL_246;
  assign _EVAL_2161 = _EVAL_2778 & _EVAL_1996;
  assign _EVAL_810 = _EVAL_3781 & _EVAL_849;
  assign _EVAL_2765 = _EVAL_810 & _EVAL_246;
  assign _EVAL_3116 = _EVAL_2765 & _EVAL_1417;
  assign _EVAL_2862 = _EVAL_1522 & _EVAL_2824;
  assign _EVAL_1086 = _EVAL_2105 & _EVAL_246;
  assign _EVAL_3068 = _EVAL_1086 & _EVAL_1417;
  assign _EVAL_3342 = _EVAL_2804 & _EVAL_3471;
  assign _EVAL_2983 = _EVAL_1942[113];
  assign _EVAL_952 = _EVAL_3781 & _EVAL_2983;
  assign _EVAL_3310 = _EVAL_952 & _EVAL_246;
  assign _EVAL_3754 = _EVAL_3310 & _EVAL_1417;
  assign _EVAL_3304 = _EVAL_3059 & _EVAL_4062;
  assign _EVAL_205 = _EVAL_3304 & _EVAL_2267;
  assign _EVAL_3924 = _EVAL_205 & _EVAL_1910;
  assign _EVAL_3532 = _EVAL_2804 & _EVAL_1963;
  assign _EVAL_385 = _EVAL_3059 & _EVAL_847;
  assign _EVAL_502 = _EVAL_2986 & _EVAL_3241;
  assign _EVAL_4024 = _EVAL_1034 & _EVAL_803;
  assign _EVAL_1967 = _EVAL_3781 & _EVAL_1053;
  assign _EVAL_2904 = _EVAL_1967 & _EVAL_246;
  assign _EVAL_3027 = _EVAL_3059 & _EVAL_1650;
  assign _EVAL_1661 = _EVAL_3027 & _EVAL_2267;
  assign _EVAL_670 = _EVAL_1942[3];
  assign _EVAL_2372 = _EVAL_3781 & _EVAL_670;
  assign _EVAL_223 = _EVAL_3402 & _EVAL_2379;
  assign _EVAL_256 = _EVAL_223 & _EVAL_246;
  assign _EVAL_2272 = _EVAL_1522 & _EVAL_3954;
  assign _EVAL_2127 = _EVAL_3458 & _EVAL_2375;
  assign _EVAL_216 = _EVAL_3402 & _EVAL_669;
  assign _EVAL_3958 = _EVAL_2376 & _EVAL_1910;
  assign _EVAL_3164 = _EVAL_3402 & _EVAL_566;
  assign _EVAL_3985 = _EVAL_3164 & _EVAL_246;
  assign _EVAL_3877 = _EVAL_3985 & _EVAL_1996;
  assign _EVAL_2566 = _EVAL_1724 & _EVAL_3693;
  assign _EVAL_2599 = _EVAL_2804 & _EVAL_3363;
  assign _EVAL_1692 = _EVAL_3458 & _EVAL_1621;
  assign _EVAL_4046 = _EVAL_2986 & _EVAL_398;
  assign _EVAL_744 = _EVAL_1857 & _EVAL_2020;
  assign _EVAL_2974 = _EVAL_3634 & _EVAL_2267;
  assign _EVAL_441 = _EVAL_2974 & _EVAL_1910;
  assign _EVAL_1840 = _EVAL_3075 & _EVAL_3180;
  assign _EVAL_1382 = _EVAL_1522 & _EVAL_2594;
  assign _EVAL_1083 = _EVAL_2900 != 8'h0;
  assign _EVAL_3763 = _EVAL_1553 & _EVAL_2043;
  assign _EVAL_1125 = _EVAL_2804 & _EVAL_3087;
  assign _EVAL_3597 = _EVAL_3781 & _EVAL_302;
  assign _EVAL_3121 = _EVAL_3597 & _EVAL_246;
  assign _EVAL_2879 = _EVAL_1279 & _EVAL_806;
  assign _EVAL_3555 = _EVAL_2804 & _EVAL_3194;
  assign _EVAL_3487 = _EVAL_2757 & _EVAL_2267;
  assign _EVAL_2692 = _EVAL_1942[61];
  assign _EVAL_290 = _EVAL_3781 & _EVAL_2692;
  assign _EVAL_344 = _EVAL_290 & _EVAL_246;
  assign _EVAL_2505 = _EVAL_344 & _EVAL_1417;
  assign _EVAL_1664 = _EVAL_2954 & _EVAL_246;
  assign _EVAL_2034 = _EVAL_1377 == 32'hffffffff;
  assign _EVAL_967 = _EVAL_1664 & _EVAL_2034;
  assign _EVAL_2637 = _EVAL_1942[56];
  assign _EVAL_1530 = _EVAL_3781 & _EVAL_2637;
  assign _EVAL_1043 = _EVAL_1530 & _EVAL_246;
  assign _EVAL_2230 = _EVAL_2804 & _EVAL_4012;
  assign _EVAL_3479 = _EVAL_1553 & _EVAL_1963;
  assign _EVAL_3989 = _EVAL_1377[15];
  assign _EVAL_2493 = _EVAL_1857 & _EVAL_3989;
  assign _EVAL_665 = _EVAL_3781 & _EVAL_2465;
  assign _EVAL_3601 = _EVAL_665 & _EVAL_246;
  assign _EVAL_1499 = _EVAL_3402 & _EVAL_3514;
  assign _EVAL_874 = _EVAL_1499 & _EVAL_246;
  assign _EVAL_857 = _EVAL_874 & _EVAL_1996;
  assign _EVAL_877 = _EVAL_1420 & _EVAL_2319;
  assign _EVAL_1060 = _EVAL_3402 & _EVAL_4065;
  assign _EVAL_3838 = _EVAL_1060 & _EVAL_246;
  assign _EVAL_483 = _EVAL_431 & _EVAL_2587;
  assign _EVAL_936 = _EVAL_2108 & _EVAL_246;
  assign _EVAL_1316 = _EVAL_1883 & _EVAL_1910;
  assign _EVAL_4071 = _EVAL_2724 & _EVAL_1417;
  assign _EVAL_4004 = _EVAL_633 & _EVAL_246;
  assign _EVAL_777 = _EVAL_4004 & _EVAL_1996;
  assign _EVAL_3676 = _EVAL_3781 & _EVAL_3613;
  assign _EVAL_2725 = _EVAL_1040 & _EVAL_724;
  assign _EVAL_1447 = _EVAL_3781 & _EVAL_3306;
  assign _EVAL_1000 = _EVAL_1447 & _EVAL_246;
  assign _EVAL_2837 = _EVAL_3402 & _EVAL_1813;
  assign _EVAL_982 = _EVAL_2837 & _EVAL_246;
  assign _EVAL_2834 = _EVAL_982 & _EVAL_1996;
  assign _EVAL_1532 = _EVAL_1034 & _EVAL_3363;
  assign _EVAL_3639 = _EVAL_3503 & _EVAL_1910;
  assign _EVAL_3176 = _EVAL_1857 & _EVAL_1324;
  assign _EVAL_1375 = _EVAL_3075 & _EVAL_3363;
  assign _EVAL_3144 = _EVAL_1099 & _EVAL_1910;
  assign _EVAL_3891 = _EVAL_3402 & _EVAL_1372;
  assign _EVAL_1822 = _EVAL_3891 & _EVAL_246;
  assign _EVAL_4022 = _EVAL_3059 & _EVAL_3508;
  assign _EVAL_2138 = _EVAL_4022 & _EVAL_2267;
  assign _EVAL_3694 = _EVAL_1857 & _EVAL_3920;
  assign _EVAL_2014 = _EVAL_1618 & _EVAL_1417;
  assign _EVAL_668 = _EVAL_3781 & _EVAL_1481;
  assign _EVAL_3871 = _EVAL_3059 & _EVAL_3423;
  assign _EVAL_3917 = _EVAL_3871 & _EVAL_2267;
  assign _EVAL_164 = _EVAL_3917 & _EVAL_1910;
  assign _EVAL_3367 = _EVAL_522 & _EVAL_2267;
  assign _EVAL_766 = _EVAL_3367 & _EVAL_1910;
  assign _EVAL_2596 = _EVAL_3565 & _EVAL_246;
  assign _EVAL_2359 = _EVAL_2596 & _EVAL_1996;
  assign _EVAL_1364 = _EVAL_3059 & _EVAL_2823;
  assign _EVAL_3482 = _EVAL_431 & _EVAL_3241;
  assign _EVAL_1401 = _EVAL_1279 & _EVAL_2961;
  assign _EVAL_2681 = _EVAL_1420 & _EVAL_3408;
  assign _EVAL_3092 = _EVAL_3530 & _EVAL_2267;
  assign _EVAL_702 = _EVAL_3402 & _EVAL_2470;
  assign _EVAL_2400 = _EVAL_702 & _EVAL_246;
  assign _EVAL_196 = _EVAL_3059 & _EVAL_1113;
  assign _EVAL_3692 = _EVAL_3402 & _EVAL_3294;
  assign _EVAL_1358 = _EVAL_3692 & _EVAL_246;
  assign _EVAL_275 = _EVAL_1867 & _EVAL_2267;
  assign _EVAL_1022 = _EVAL_275 & _EVAL_1910;
  assign _EVAL_4037 = _EVAL_958 & _EVAL_1910;
  assign _EVAL_1116 = _EVAL_2804 & _EVAL_655;
  assign _EVAL_1319 = _EVAL_3781 & _EVAL_2617;
  assign _EVAL_2312 = _EVAL_1319 & _EVAL_246;
  assign _EVAL_3517 = _EVAL_2312 & _EVAL_1417;
  assign _EVAL_1049 = _EVAL_3781 & _EVAL_629;
  assign _EVAL_1031 = _EVAL_2804 & _EVAL_2339;
  assign _EVAL_153 = _EVAL_3927 & _EVAL_246;
  assign _EVAL_2264 = _EVAL_153 & _EVAL_1996;
  assign _EVAL_3610 = _EVAL_3856 | _EVAL_1990;
  assign _EVAL_2769 = _EVAL_1377[8];
  assign _EVAL_337 = _EVAL_1724 & _EVAL_2769;
  assign _EVAL_2569 = _EVAL_1279 & _EVAL_215;
  assign _EVAL_2759 = _EVAL_2804 & _EVAL_215;
  assign _EVAL_484 = _EVAL_1040 & _EVAL_2830;
  assign _EVAL_3885 = _EVAL_3781 & _EVAL_411;
  assign _EVAL_1653 = _EVAL_431 & _EVAL_3779;
  assign _EVAL_3834 = _EVAL_3029 & _EVAL_1996;
  assign _EVAL_1755 = _EVAL_2044 & _EVAL_1910;
  assign _EVAL_558 = _EVAL_3781 & _EVAL_883;
  assign _EVAL_1912 = _EVAL_558 & _EVAL_246;
  assign _EVAL_2250 = _EVAL_1912 & _EVAL_1417;
  assign _EVAL_1384 = _EVAL_2516 & _EVAL_246;
  assign _EVAL_1065 = _EVAL_1545 & _EVAL_2769;
  assign _EVAL_1997 = _EVAL_1942[25];
  assign _EVAL_544 = _EVAL_3781 & _EVAL_1997;
  assign _EVAL_2275 = _EVAL_544 & _EVAL_246;
  assign _EVAL_991 = _EVAL_3121 & _EVAL_1417;
  assign _EVAL_903 = _EVAL_3781 & _EVAL_637;
  assign _EVAL_3496 = _EVAL_903 & _EVAL_246;
  assign _EVAL_1098 = _EVAL_1045 != 8'h0;
  assign _EVAL_3313 = _EVAL_3496 & _EVAL_1098;
  assign _EVAL_1961 = _EVAL_747 & _EVAL_1996;
  assign _EVAL_3327 = _EVAL_2080 & _EVAL_2267;
  assign _EVAL_1652 = _EVAL_3781 & _EVAL_2808;
  assign _EVAL_1659 = _EVAL_3402 & _EVAL_3173;
  assign _EVAL_3375 = _EVAL_3697 & _EVAL_1417;
  assign _EVAL_3777 = _EVAL_1821 & _EVAL_246;
  assign _EVAL_2855 = _EVAL_3777 & _EVAL_1996;
  assign _EVAL_1001 = _EVAL_3496 & _EVAL_3217;
  assign _EVAL_2678 = _EVAL_1470 & _EVAL_1868;
  assign _EVAL_2630 = _EVAL_3075 & _EVAL_1048;
  assign _EVAL_2488 = _EVAL_3059 & _EVAL_236;
  assign _EVAL_1941 = _EVAL_2488 & _EVAL_2267;
  assign _EVAL_2753 = _EVAL_1941 & _EVAL_1910;
  assign _EVAL_3931 = _EVAL_3402 & _EVAL_776;
  assign _EVAL_456 = _EVAL_3931 & _EVAL_246;
  assign _EVAL_654 = _EVAL_3512 & _EVAL_1910;
  assign _EVAL_785 = _EVAL_3059 & _EVAL_2302;
  assign _EVAL_2154 = _EVAL_785 & _EVAL_2267;
  assign _EVAL_2992 = _EVAL_2154 & _EVAL_1910;
  assign _EVAL_1759 = _EVAL_3402 & _EVAL_2808;
  assign _EVAL_3580 = _EVAL_1759 & _EVAL_246;
  assign _EVAL_3392 = _EVAL_3059 & _EVAL_1706;
  assign _EVAL_2212 = _EVAL_2636 & _EVAL_1417;
  assign _EVAL_789 = _EVAL_1942[94];
  assign _EVAL_3085 = _EVAL_3402 & _EVAL_789;
  assign _EVAL_783 = _EVAL_3897 & _EVAL_3285;
  assign _EVAL_2546 = _EVAL_3110 & _EVAL_2267;
  assign _EVAL_3197 = _EVAL_431 & _EVAL_803;
  assign _EVAL_2039 = _EVAL_3402 & _EVAL_1761;
  assign _EVAL_2387 = _EVAL_2039 & _EVAL_246;
  assign _EVAL_2816 = _EVAL_3059 & _EVAL_268;
  assign _EVAL_2069 = _EVAL_2816 & _EVAL_2267;
  assign _EVAL_3598 = _EVAL_3458 & _EVAL_3285;
  assign _EVAL_2570 = _EVAL_1942[97];
  assign _EVAL_3212 = _EVAL_3402 & _EVAL_2570;
  assign _EVAL_3253 = _EVAL_3212 & _EVAL_246;
  assign _EVAL_2352 = _EVAL_3836 & _EVAL_2267;
  assign _EVAL_1428 = _EVAL_2352 & _EVAL_1910;
  assign _EVAL_3124 = _EVAL_3059 & _EVAL_3642;
  assign _EVAL_3672 = _EVAL_3770 & _EVAL_2267;
  assign _EVAL_1964 = _EVAL_3672 & _EVAL_1910;
  assign _EVAL_1747 = _EVAL_3402 & _EVAL_496;
  assign _EVAL_1039 = _EVAL_1747 & _EVAL_246;
  assign _EVAL_642 = _EVAL_2986 & _EVAL_2587;
  assign _EVAL_2672 = _EVAL_3897 & _EVAL_2756;
  assign _EVAL_3567 = _EVAL_1553 & _EVAL_696;
  assign _EVAL_630 = _EVAL_1942[30];
  assign _EVAL_895 = _EVAL_3781 & _EVAL_630;
  assign _EVAL_3983 = _EVAL_3781 & _EVAL_3286;
  assign _EVAL_2406 = _EVAL_3983 & _EVAL_246;
  assign _EVAL_453 = _EVAL_2406 & _EVAL_1417;
  assign _EVAL_1105 = _EVAL_3897 & _EVAL_2691;
  assign _EVAL_1828 = _EVAL_3897 & _EVAL_662;
  assign _EVAL_1233 = _EVAL_1553 & _EVAL_803;
  assign _EVAL_853 = _EVAL_3059 & _EVAL_828;
  assign _EVAL_2292 = _EVAL_853 & _EVAL_2267;
  assign _EVAL_2695 = _EVAL_1942[119];
  assign _EVAL_3255 = _EVAL_1553 & _EVAL_3180;
  assign _EVAL_2822 = _EVAL_3960 & _EVAL_1910;
  assign _EVAL_170 = _EVAL_3643 & _EVAL_1996;
  assign _EVAL_3031 = _EVAL_2112 & _EVAL_3779;
  assign _EVAL_2512 = _EVAL_1857 & _EVAL_543;
  assign _EVAL_2887 = _EVAL_3781 & _EVAL_566;
  assign _EVAL_2200 = _EVAL_1279 & _EVAL_3596;
  assign _EVAL_2222 = _EVAL_1577 & _EVAL_1910;
  assign _EVAL_2924 = _EVAL_3392 & _EVAL_2267;
  assign _EVAL_1975 = _EVAL_2924 & _EVAL_1910;
  assign _EVAL_3170 = _EVAL_3458 & _EVAL_2984;
  assign _EVAL_3967 = _EVAL_3601 & _EVAL_1417;
  assign _EVAL_738 = _EVAL_3676 & _EVAL_246;
  assign _EVAL_3498 = _EVAL_738 & _EVAL_1417;
  assign _EVAL_2604 = _EVAL_1920 & _EVAL_1417;
  assign _EVAL_2437 = _EVAL_3402 & _EVAL_211;
  assign _EVAL_3904 = _EVAL_2437 & _EVAL_246;
  assign _EVAL_2478 = _EVAL_3904 & _EVAL_1996;
  assign _EVAL_3019 = _EVAL_3253 & _EVAL_1996;
  assign _EVAL_463 = _EVAL_2804 & _EVAL_4016;
  assign _EVAL_1493 = _EVAL_2112 & _EVAL_3701;
  assign _EVAL_156 = _EVAL_2369 & _EVAL_246;
  assign _EVAL_3341 = _EVAL_1846 & _EVAL_1996;
  assign _EVAL_2239 = _EVAL_2069 & _EVAL_1910;
  assign _EVAL_3237 = _EVAL_3781 & _EVAL_2042;
  assign _EVAL_3506 = _EVAL_3487 & _EVAL_1910;
  assign _EVAL_924 = _EVAL_3059 & _EVAL_3816;
  assign _EVAL_506 = _EVAL_924 & _EVAL_2267;
  assign _EVAL_305 = _EVAL_1942[42];
  assign _EVAL_3132 = _EVAL_3781 & _EVAL_305;
  assign _EVAL_1900 = _EVAL_3132 & _EVAL_246;
  assign _EVAL_3346 = _EVAL_1279 & _EVAL_3180;
  assign _EVAL_1334 = _EVAL_1522 & _EVAL_1324;
  assign _EVAL_3668 = _EVAL_3781 & _EVAL_1258;
  assign _EVAL_1719 = _EVAL_3668 & _EVAL_246;
  assign _EVAL_482 = _EVAL_431 & _EVAL_696;
  assign _EVAL_3399 = _EVAL_3059 & _EVAL_265;
  assign _EVAL_1622 = _EVAL_3399 & _EVAL_2267;
  assign _EVAL_2880 = _EVAL_3402 & _EVAL_3761;
  assign _EVAL_2010 = _EVAL_3059 & _EVAL_1400;
  assign _EVAL_3201 = _EVAL_2010 & _EVAL_2267;
  assign _EVAL_3389 = _EVAL_3201 & _EVAL_1910;
  assign _EVAL_2479 = _EVAL_3781 & _EVAL_1989;
  assign _EVAL_2602 = _EVAL_2479 & _EVAL_246;
  assign _EVAL_2329 = _EVAL_3781 & _EVAL_3036;
  assign _EVAL_3955 = _EVAL_2329 & _EVAL_246;
  assign _EVAL_426 = _EVAL_3955 & _EVAL_1417;
  assign _EVAL_3365 = {{3'd0}, _EVAL_3406};
  assign _EVAL_1074 = _EVAL_3235 <= _EVAL_3365;
  assign _EVAL_3422 = _EVAL_3746 & _EVAL_1074;
  assign _EVAL_563 = _EVAL_3402 & _EVAL_305;
  assign _EVAL_855 = _EVAL_1630 & _EVAL_2267;
  assign _EVAL_2313 = _EVAL_232 & _EVAL_1996;
  assign _EVAL_1361 = _EVAL_1857 & _EVAL_724;
  assign _EVAL_2930 = _EVAL_823 & _EVAL_1417;
  assign _EVAL_3929 = _EVAL_3897 & _EVAL_1490;
  assign _EVAL_1767 = _EVAL_3402 & _EVAL_1997;
  assign _EVAL_2392 = _EVAL_1767 & _EVAL_246;
  assign _EVAL_3355 = _EVAL_3897 & _EVAL_2375;
  assign _EVAL_3592 = _EVAL_3781 & _EVAL_4019;
  assign _EVAL_3080 = _EVAL_2527 & _EVAL_3572;
  assign _EVAL_2719 = ~ _EVAL_3531;
  assign _EVAL_1619 = _EVAL_3080 & _EVAL_2719;
  assign _EVAL_1373 = _EVAL_1619 - 127'h1;
  assign _EVAL_2085 = _EVAL_403 & _EVAL_246;
  assign _EVAL_2367 = _EVAL_2085 & _EVAL_1996;
  assign _EVAL_1916 = _EVAL_3402 & _EVAL_2695;
  assign _EVAL_3666 = _EVAL_1916 & _EVAL_246;
  assign _EVAL_272 = _EVAL_3059 & _EVAL_3117;
  assign _EVAL_4072 = _EVAL_272 & _EVAL_2267;
  assign _EVAL_627 = _EVAL_1895 & _EVAL_920;
  assign _EVAL_3457 = _EVAL_431 & _EVAL_2072;
  assign _EVAL_2738 = _EVAL_2124[31:3];
  assign _EVAL_1878 = _EVAL_1040 & _EVAL_3954;
  assign _EVAL_2894 = _EVAL_563 & _EVAL_246;
  assign _EVAL_2752 = _EVAL_3781 & _EVAL_2695;
  assign _EVAL_2799 = _EVAL_2752 & _EVAL_246;
  assign _EVAL_961 = _EVAL_2799 & _EVAL_1417;
  assign _EVAL_172 = _EVAL_1942[5];
  assign _EVAL_3309 = _EVAL_3402 & _EVAL_172;
  assign _EVAL_1760 = _EVAL_3059 & _EVAL_2608;
  assign _EVAL_1687 = _EVAL_1760 & _EVAL_2267;
  assign _EVAL_1118 = _EVAL_1687 & _EVAL_1910;
  assign _EVAL_1844 = _EVAL_1034 & _EVAL_2344;
  assign _EVAL_3585 = _EVAL_2342 & _EVAL_246;
  assign _EVAL_1058 = _EVAL_3585 & _EVAL_1996;
  assign _EVAL_2529 = _EVAL_3327 & _EVAL_1910;
  assign _EVAL_312 = _EVAL_3075 & _EVAL_1224;
  assign _EVAL_1700 = _EVAL_3059 & _EVAL_829;
  assign _EVAL_3123 = _EVAL_1700 & _EVAL_2267;
  assign _EVAL_2177 = _EVAL_3123 & _EVAL_1910;
  assign _EVAL_802 = _EVAL_3402 & _EVAL_2983;
  assign _EVAL_1056 = _EVAL_431 & _EVAL_3701;
  assign _EVAL_906 = _EVAL_3781 & _EVAL_2570;
  assign _EVAL_3886 = _EVAL_431 & _EVAL_4016;
  assign _EVAL_3753 = _EVAL_3458 & _EVAL_3470;
  assign _EVAL_1904 = _EVAL_1522 & _EVAL_3989;
  assign _EVAL_2673 = _EVAL_3402 & _EVAL_2919;
  assign _EVAL_1451 = _EVAL_2673 & _EVAL_246;
  assign _EVAL_1826 = _EVAL_3402 & _EVAL_670;
  assign _EVAL_1808 = _EVAL_1826 & _EVAL_246;
  assign _EVAL_2338 = _EVAL_1470 & _EVAL_3989;
  assign _EVAL_1117 = _EVAL_1279 & _EVAL_3145;
  assign _EVAL_2784 = _EVAL_3210 & _EVAL_246;
  assign _EVAL_2550 = _EVAL_2784 & _EVAL_1417;
  assign _EVAL_1474 = _EVAL_3897 & _EVAL_2020;
  assign _EVAL_659 = _EVAL_3075 & _EVAL_3145;
  assign _EVAL_672 = _EVAL_1553 & _EVAL_3209;
  assign _EVAL_2946 = _EVAL_2874 & _EVAL_2283;
  assign _EVAL_2165 = _EVAL_3059 & _EVAL_2856;
  assign _EVAL_3577 = _EVAL_2165 & _EVAL_2267;
  assign _EVAL_296 = _EVAL_1857 & _EVAL_2691;
  assign _EVAL_3076 = _EVAL_3458 & _EVAL_424;
  assign _EVAL_1696 = _EVAL_2986 & _EVAL_3363;
  assign _EVAL_1007 = _EVAL_3402 & _EVAL_1554;
  assign _EVAL_3858 = _EVAL_3781 & _EVAL_2941;
  assign _EVAL_3778 = _EVAL_3858 & _EVAL_246;
  assign _EVAL_677 = _EVAL_3778 & _EVAL_1098;
  assign _EVAL_2374 = _EVAL_1398 & _EVAL_1083;
  assign _EVAL_3975 = _EVAL_1377[23:16];
  assign _EVAL_996 = _EVAL_3975 != 8'h0;
  assign _EVAL_4051 = _EVAL_3402 & _EVAL_3326;
  assign _EVAL_2458 = _EVAL_2805 & _EVAL_1910;
  assign _EVAL_578 = _EVAL_3075 & _EVAL_3194;
  assign _EVAL_2032 = _EVAL_1724 & _EVAL_3000;
  assign _EVAL_4002 = _EVAL_3781 & _EVAL_2792;
  assign _EVAL_2734 = _EVAL_4002 & _EVAL_246;
  assign _EVAL_2473 = _EVAL_3402 & _EVAL_1335;
  assign _EVAL_407 = _EVAL_2473 & _EVAL_246;
  assign _EVAL_1008 = _EVAL_407 & _EVAL_1996;
  assign _EVAL_2905 = _EVAL_1553 & _EVAL_2961;
  assign _EVAL_1199 = _EVAL_1921 & _EVAL_246;
  assign _EVAL_3792 = _EVAL_216 & _EVAL_246;
  assign _EVAL_2071 = _EVAL_3696 & _EVAL_246;
  assign _EVAL_955 = _EVAL_2071 & _EVAL_1417;
  assign _EVAL_1978 = _EVAL_3140 & _EVAL_996;
  assign _EVAL_1902 = _EVAL_2986 & _EVAL_3145;
  assign _EVAL_1419 = _EVAL_1724 & _EVAL_2020;
  assign _EVAL_4007 = _EVAL_1857 & _EVAL_1490;
  assign _EVAL_3942 = _EVAL_1545 & _EVAL_887;
  assign _EVAL_3747 = _EVAL_1545 & _EVAL_2824;
  assign _EVAL_1087 = _EVAL_2986 & _EVAL_3596;
  assign _EVAL_831 = _EVAL_3059 & _EVAL_3919;
  assign _EVAL_4030 = _EVAL_1872 & _EVAL_1417;
  assign _EVAL_2089 = _EVAL_1522 & _EVAL_1868;
  assign _EVAL_1604 = _EVAL_3402 & _EVAL_297;
  assign _EVAL_209 = _EVAL_906 & _EVAL_246;
  assign _EVAL_589 = _EVAL_3897 & _EVAL_2769;
  assign _EVAL_2476 = _EVAL_2986 & _EVAL_2344;
  assign _EVAL_2921 = _EVAL_3402 & _EVAL_4069;
  assign _EVAL_1684 = _EVAL_2921 & _EVAL_246;
  assign _EVAL_2890 = _EVAL_1684 & _EVAL_1996;
  assign _EVAL_1908 = _EVAL_1279 & _EVAL_2344;
  assign _EVAL_3357 = _EVAL_1857 & _EVAL_3038;
  assign _EVAL_805 = _EVAL_1724 & _EVAL_543;
  assign _EVAL_2709 = _EVAL_1040 & _EVAL_3285;
  assign _EVAL_1353 = _EVAL_3685 & _EVAL_246;
  assign _EVAL_3444 = _EVAL_1192 & _EVAL_1417;
  assign _EVAL_2046 = _EVAL_1034 & _EVAL_4016;
  assign _EVAL_3090 = _EVAL_1857 & _EVAL_424;
  assign _EVAL_1668 = _EVAL_1545 & _EVAL_2594;
  assign _EVAL_838 = _EVAL_1724 & _EVAL_2830;
  assign _EVAL_1570 = _EVAL_1451 & _EVAL_1996;
  assign _EVAL_4057 = _EVAL_1470 & _EVAL_3470;
  assign _EVAL_3160 = _EVAL_2880 & _EVAL_246;
  assign _EVAL_467 = _EVAL_3438 & _EVAL_1417;
  assign _EVAL_3126 = _EVAL_1659 & _EVAL_246;
  assign _EVAL_1905 = _EVAL_831 & _EVAL_2267;
  assign _EVAL_1238 = _EVAL_1905 & _EVAL_1910;
  assign _EVAL_577 = _EVAL_2804 & _EVAL_3145;
  assign _EVAL_3703 = _EVAL_1034 & _EVAL_2043;
  assign _EVAL_1090 = _EVAL_3885 & _EVAL_246;
  assign _EVAL_3854 = _EVAL_1090 & _EVAL_1417;
  assign _EVAL_2235 = _EVAL_1279 & _EVAL_3209;
  assign _EVAL_3386 = _EVAL_3151 & _EVAL_1417;
  assign _EVAL_3003 = _EVAL_3897 & _EVAL_3920;
  assign _EVAL_3349 = _EVAL_1040 & _EVAL_1490;
  assign _EVAL_817 = _EVAL_1470 & _EVAL_724;
  assign _EVAL_3714 = _EVAL_3458 & _EVAL_2824;
  assign _EVAL_1344 = _EVAL_1040 & _EVAL_887;
  assign _EVAL_2298 = _EVAL_1724 & _EVAL_1324;
  assign _EVAL_2350 = _EVAL_3075 & _EVAL_1245;
  assign _EVAL_1304 = _EVAL_2611 & _EVAL_2267;
  assign _EVAL_1342 = _EVAL_1304 & _EVAL_1910;
  assign _EVAL_1050 = _EVAL_2452 & _EVAL_246;
  assign _EVAL_860 = _EVAL_2387 & _EVAL_1996;
  assign _EVAL_689 = _EVAL_3059 & _EVAL_3325;
  assign _EVAL_962 = _EVAL_689 & _EVAL_2267;
  assign _EVAL_2077 = _EVAL_962 & _EVAL_1910;
  assign _EVAL_244 = _EVAL_3059 & _EVAL_2959;
  assign _EVAL_1610 = _EVAL_244 & _EVAL_2267;
  assign _EVAL_3324 = _EVAL_1553 & _EVAL_4016;
  assign _EVAL_2377 = _EVAL_1808 & _EVAL_1996;
  assign _EVAL_528 = _EVAL_2986 & _EVAL_4006;
  assign _EVAL_3316 = _EVAL_2112 & _EVAL_3471;
  assign _EVAL_545 = _EVAL_1822 & _EVAL_2544;
  assign _EVAL_486 = _EVAL_3085 & _EVAL_246;
  assign _EVAL_2549 = _EVAL_1619 & _EVAL_1373;
  assign _EVAL_3340 = _EVAL_3402 & _EVAL_999;
  assign _EVAL_3640 = _EVAL_3340 & _EVAL_246;
  assign _EVAL_301 = _EVAL_3640 & _EVAL_1996;
  assign _EVAL_3465 = _EVAL_431 & _EVAL_1048;
  assign _EVAL_150 = _EVAL_1942[39];
  assign _EVAL_1214 = _EVAL_3781 & _EVAL_150;
  assign _EVAL_361 = _EVAL_1214 & _EVAL_246;
  assign _EVAL_3723 = _EVAL_361 & _EVAL_1417;
  assign _EVAL_3106 = _EVAL_3402 & _EVAL_3906;
  assign _EVAL_2652 = _EVAL_1470 & _EVAL_2691;
  assign _EVAL_2509 = _EVAL_2292 & _EVAL_1910;
  assign _EVAL_641 = _EVAL_3402 & _EVAL_2489;
  assign _EVAL_1268 = _EVAL_641 & _EVAL_246;
  assign _EVAL_634 = _EVAL_1622 & _EVAL_1910;
  assign _EVAL_1714 = _EVAL_1724 & _EVAL_2691;
  assign _EVAL_3437 = _EVAL_1040 & _EVAL_520;
  assign _EVAL_2537 = _EVAL_3352 & _EVAL_246;
  assign _EVAL_3010 = _EVAL_2537 & _EVAL_1996;
  assign _EVAL_3277 = _EVAL_3402 & _EVAL_3207;
  assign _EVAL_162 = _EVAL_3736 & _EVAL_3408;
  assign _EVAL_430 = _EVAL_931 & _EVAL_1996;
  assign _EVAL_1600 = _EVAL_1610 & _EVAL_1910;
  assign _EVAL_1223 = _EVAL_3277 & _EVAL_246;
  assign _EVAL_3794 = _EVAL_3897 & _EVAL_3954;
  assign _EVAL_1807 = _EVAL_3781 & _EVAL_2919;
  assign _EVAL_2207 = _EVAL_3402 & _EVAL_630;
  assign _EVAL_3447 = _EVAL_2207 & _EVAL_246;
  assign _EVAL_2839 = _EVAL_3447 & _EVAL_1996;
  assign _EVAL_2414 = _EVAL_3458 & _EVAL_2756;
  assign _EVAL_2518 = _EVAL_2112 & _EVAL_2587;
  assign _EVAL_307 = _EVAL_3458 & _EVAL_3693;
  assign _EVAL_1320 = _EVAL_1040 & _EVAL_3920;
  assign _EVAL_4045 = _EVAL_1545 & _EVAL_2412;
  assign _EVAL_893 = _EVAL_1522 & _EVAL_1354;
  assign _EVAL_2849 = _EVAL_431 & _EVAL_398;
  assign _EVAL_3686 = _EVAL_3458 & _EVAL_2830;
  assign _EVAL_900 = _EVAL_1470 & _EVAL_424;
  assign _EVAL_1138 = _EVAL_3075 & _EVAL_2072;
  assign _EVAL_1391 = _EVAL_1034 & _EVAL_3194;
  assign _EVAL_1033 = _EVAL_1034 & _EVAL_3209;
  assign _EVAL_2772 = _EVAL_1724 & _EVAL_3148;
  assign _EVAL_1953 = _EVAL_1049 & _EVAL_246;
  assign _EVAL_2916 = _EVAL_1353 & _EVAL_1996;
  assign _EVAL_1693 = _EVAL_1040 & _EVAL_169;
  assign _EVAL_644 = _EVAL_1895 & _EVAL_388;
  assign _EVAL_180 = _EVAL_3059 & _EVAL_3215;
  assign _EVAL_201 = _EVAL_180 & _EVAL_2267;
  assign _EVAL_158 = _EVAL_201 & _EVAL_1910;
  assign _EVAL_2216 = _EVAL_1040 & _EVAL_2412;
  assign _EVAL_2472 = _EVAL_895 & _EVAL_246;
  assign _EVAL_1112 = _EVAL_2112 & _EVAL_803;
  assign _EVAL_228 = _EVAL_3059 & _EVAL_1236;
  assign _EVAL_601 = _EVAL_228 & _EVAL_2267;
  assign _EVAL_1830 = _EVAL_3124 & _EVAL_2267;
  assign _EVAL_2186 = _EVAL_3737 & _EVAL_1910;
  assign _EVAL_674 = _EVAL_336 & _EVAL_1996;
  assign _EVAL_1501 = _EVAL_2112 & _EVAL_3241;
  assign _EVAL_3155 = _EVAL_3402 & _EVAL_1947;
  assign _EVAL_3813 = _EVAL_3155 & _EVAL_246;
  assign _EVAL_3660 = _EVAL_1524 & _EVAL_1996;
  assign _EVAL_4067 = _EVAL_431 & _EVAL_806;
  assign _EVAL_2364 = _EVAL_1862 & _EVAL_1417;
  assign _EVAL_2427 = _EVAL_3781 & _EVAL_1818;
  assign _EVAL_2418 = _EVAL_2427 & _EVAL_246;
  assign _EVAL_3862 = _EVAL_2418 & _EVAL_1417;
  assign _EVAL_628 = _EVAL_1990 & _EVAL_3691;
  assign _EVAL_1720 = _EVAL_628 == 1'h0;
  assign _EVAL_161 = _EVAL_1720 | _EVAL_105;
  assign _EVAL_3541 = _EVAL_161 == 1'h0;
  assign _EVAL_1678 = _EVAL_2606 & _EVAL_246;
  assign _EVAL_842 = _EVAL_2166 & _EVAL_1417;
  assign _EVAL_2773 = _EVAL_2985 & _EVAL_1910;
  assign _EVAL_1255 = _EVAL_1279 & _EVAL_398;
  assign _EVAL_1971 = _EVAL_3458 & _EVAL_1490;
  assign _EVAL_2327 = _EVAL_1857 & _EVAL_1868;
  assign _EVAL_1789 = _EVAL_3059 & _EVAL_925;
  assign _EVAL_3086 = _EVAL_1279 & _EVAL_3701;
  assign _EVAL_1988 = _EVAL_1553 & _EVAL_3194;
  assign _EVAL_3435 = _EVAL_1857 & _EVAL_2756;
  assign _EVAL_1984 = _EVAL_666 == _EVAL_666;
  assign _EVAL_1675 = _EVAL_1984 | _EVAL_105;
  assign _EVAL_2049 = _EVAL_1675 == 1'h0;
  assign _EVAL_1615 = _EVAL_3781 & _EVAL_1800;
  assign _EVAL_2957 = _EVAL_1615 & _EVAL_246;
  assign _EVAL_2268 = _EVAL_2957 & _EVAL_1417;
  assign _EVAL_1234 = _EVAL_2041 & _EVAL_215;
  assign _EVAL_3947 = _EVAL_3059 & _EVAL_2713;
  assign _EVAL_186 = _EVAL_3947 & _EVAL_2267;
  assign _EVAL_2714 = _EVAL_2986 & _EVAL_3087;
  assign _EVAL_1217 = _EVAL_3781 & _EVAL_2205;
  assign _EVAL_2321 = _EVAL_1217 & _EVAL_246;
  assign _EVAL_2185 = _EVAL_3778 & _EVAL_1083;
  assign _EVAL_619 = _EVAL_506 & _EVAL_1910;
  assign _EVAL_885 = _EVAL_1029 & _EVAL_246;
  assign _EVAL_3604 = _EVAL_431 & _EVAL_655;
  assign _EVAL_3321 = _EVAL_1789 & _EVAL_2267;
  assign _EVAL_3133 = _EVAL_1566 & _EVAL_246;
  assign _EVAL_3049 = _EVAL_3133 & _EVAL_1996;
  assign _EVAL_281 = _EVAL_1553 & _EVAL_806;
  assign _EVAL_3538 = _EVAL_3781 & _EVAL_478;
  assign _EVAL_2542 = _EVAL_763 & _EVAL_1417;
  assign _EVAL_3046 = _EVAL_3059 & _EVAL_1064;
  assign _EVAL_3227 = _EVAL_2112 & _EVAL_4006;
  assign _EVAL_3161 = _EVAL_1724 & _EVAL_2984;
  assign _EVAL_493 = _EVAL_1470 & _EVAL_169;
  assign _EVAL_3700 = _EVAL_1279 & _EVAL_2339;
  assign _EVAL_2002 = _EVAL_3458 & _EVAL_1354;
  assign _EVAL_239 = _EVAL_2986 & _EVAL_3180;
  assign _EVAL_1422 = _EVAL_3458 & _EVAL_2769;
  assign _EVAL_1606 = _EVAL_802 & _EVAL_246;
  assign _EVAL_1356 = _EVAL_3413 & _EVAL_1910;
  assign _EVAL_1336 = _EVAL_2986 & _EVAL_215;
  assign _EVAL_3260 = _EVAL_2372 & _EVAL_246;
  assign _EVAL_154 = _EVAL_3260 & _EVAL_1417;
  assign _EVAL_1037 = _EVAL_3781 & _EVAL_1903;
  assign _EVAL_1924 = _EVAL_3141 & _EVAL_1910;
  assign _EVAL_1498 = _EVAL_2112 & _EVAL_1963;
  assign _EVAL_3149 = _EVAL_3702 & _EVAL_1910;
  assign _EVAL_2324 = _EVAL_3897 & _EVAL_2412;
  assign _EVAL_3545 = _EVAL_2694 & _EVAL_1910;
  assign _EVAL_160 = _EVAL_209 & _EVAL_1417;
  assign _EVAL_1662 = _EVAL_1724 & _EVAL_520;
  assign _EVAL_3658 = _EVAL_186 & _EVAL_1910;
  assign _EVAL_2789 = _EVAL_3980 & _EVAL_1910;
  assign _EVAL_3193 = _EVAL_3856 & _EVAL_1327;
  assign _EVAL_1071 = _EVAL_2734 & _EVAL_1417;
  assign _EVAL_1146 = _EVAL_1040 & _EVAL_2769;
  assign _EVAL_2022 = _EVAL_2240 & _EVAL_1910;
  assign _EVAL_1411 = _EVAL_3106 & _EVAL_246;
  assign _EVAL_3893 = _EVAL_885 & _EVAL_1996;
  assign _EVAL_3040 = _EVAL_1942[33];
  assign _EVAL_4058 = _EVAL_3402 & _EVAL_3040;
  assign _EVAL_408 = _EVAL_3458 & _EVAL_724;
  assign _EVAL_2517 = _EVAL_2986 & _EVAL_3779;
  assign _EVAL_3398 = _EVAL_1455 & _EVAL_246;
  assign _EVAL_1865 = _EVAL_3237 & _EVAL_246;
  assign _EVAL_3984 = _EVAL_3059 & _EVAL_1235;
  assign _EVAL_3846 = _EVAL_3984 & _EVAL_2267;
  assign _EVAL_2908 = _EVAL_3846 & _EVAL_1910;
  assign _EVAL_2895 = _EVAL_977 & _EVAL_246;
  assign _EVAL_2768 = _EVAL_3781 & _EVAL_978;
  assign _EVAL_2417 = _EVAL_2768 & _EVAL_246;
  assign _EVAL_273 = _EVAL_1857 & _EVAL_2769;
  assign _EVAL_602 = _EVAL_1404 & _EVAL_1996;
  assign _EVAL_2758 = _EVAL_3975 == 8'hff;
  assign _EVAL_1803 = _EVAL_2173 & _EVAL_2758;
  assign _EVAL_3569 = _EVAL_3580 & _EVAL_1996;
  assign _EVAL_3741 = _EVAL_2546 & _EVAL_1910;
  assign _EVAL_3536 = _EVAL_431 & _EVAL_1245;
  assign _EVAL_1679 = _EVAL_1279 & _EVAL_1963;
  assign _EVAL_322 = _EVAL_2804 & _EVAL_3209;
  assign _EVAL_2708 = _EVAL_3781 & _EVAL_1809;
  assign _EVAL_2328 = _EVAL_2708 & _EVAL_246;
  assign _EVAL_2722 = _EVAL_2328 & _EVAL_1417;
  assign _EVAL_3302 = _EVAL_1470 & _EVAL_3954;
  assign _EVAL_2700 = _EVAL_3402 & _EVAL_150;
  assign _EVAL_2213 = _EVAL_1199 & _EVAL_1996;
  assign _EVAL_3507 = _EVAL_3059 & _EVAL_295;
  assign _EVAL_2586 = _EVAL_3507 & _EVAL_2267;
  assign _EVAL_676 = _EVAL_2586 & _EVAL_1910;
  assign _EVAL_406 = _EVAL_601 & _EVAL_1910;
  assign _EVAL_983 = _EVAL_3059 & _EVAL_2054;
  assign _EVAL_3115 = _EVAL_3290 & _EVAL_246;
  assign _EVAL_951 = _EVAL_3115 & _EVAL_1417;
  assign _EVAL_1254 = _EVAL_1437 & _EVAL_246;
  assign _EVAL_1123 = _EVAL_3059 & _EVAL_2866;
  assign _EVAL_3058 = _EVAL_1123 & _EVAL_2267;
  assign _EVAL_2897 = _EVAL_3699 & _EVAL_246;
  assign _EVAL_2934 = _EVAL_3600 & _EVAL_1417;
  assign _EVAL_3612 = _EVAL_3059 & _EVAL_2520;
  assign _EVAL_417 = _EVAL_3781 & _EVAL_2420;
  assign _EVAL_3651 = _EVAL_417 & _EVAL_246;
  assign _EVAL_1442 = _EVAL_3781 & _EVAL_172;
  assign _EVAL_3859 = _EVAL_1942[9];
  assign _EVAL_2353 = _EVAL_3402 & _EVAL_3859;
  assign _EVAL_3373 = _EVAL_2353 & _EVAL_246;
  assign _EVAL_621 = _EVAL_3373 & _EVAL_1996;
  assign _EVAL_1256 = _EVAL_3059 & _EVAL_927;
  assign _EVAL_1341 = _EVAL_1256 & _EVAL_2267;
  assign _EVAL_1539 = _EVAL_1341 & _EVAL_1910;
  assign _EVAL_1551 = _EVAL_1807 & _EVAL_246;
  assign _EVAL_2813 = _EVAL_1442 & _EVAL_246;
  assign _EVAL_434 = _EVAL_1155 & _EVAL_1417;
  assign _EVAL_3303 = _EVAL_3402 & _EVAL_2637;
  assign _EVAL_1406 = _EVAL_3303 & _EVAL_246;
  assign _EVAL_3922 = _EVAL_1522 & _EVAL_3038;
  assign _EVAL_2038 = _EVAL_2258 & _EVAL_1996;
  assign _EVAL_862 = _EVAL_1522 & _EVAL_2375;
  assign _EVAL_1798 = _EVAL_1040 & _EVAL_3000;
  assign _EVAL_3224 = _EVAL_3611 & _EVAL_2267;
  assign _EVAL_185 = _EVAL_3781 & _EVAL_3071;
  assign _EVAL_3704 = _EVAL_185 & _EVAL_246;
  assign _EVAL_1003 = _EVAL_1522 & _EVAL_3470;
  assign _EVAL_2787 = _EVAL_3458 & _EVAL_520;
  assign _EVAL_3009 = _EVAL_3059 & _EVAL_2571;
  assign _EVAL_2552 = _EVAL_3009 & _EVAL_2267;
  assign _EVAL_1126 = _EVAL_2552 & _EVAL_1910;
  assign _EVAL_2635 = _EVAL_1470 & _EVAL_662;
  assign _EVAL_681 = _EVAL_1254 & _EVAL_1996;
  assign _EVAL_261 = _EVAL_1398 & _EVAL_996;
  assign _EVAL_908 = _EVAL_3309 & _EVAL_246;
  assign _EVAL_1685 = _EVAL_3402 & _EVAL_324;
  assign _EVAL_2045 = _EVAL_1685 & _EVAL_246;
  assign _EVAL_3637 = _EVAL_2045 & _EVAL_1996;
  assign _EVAL_950 = _EVAL_3897 & _EVAL_2830;
  assign _EVAL_2707 = _EVAL_3059 & _EVAL_2052;
  assign _EVAL_2475 = _EVAL_2707 & _EVAL_2267;
  assign _EVAL_749 = _EVAL_2475 & _EVAL_1910;
  assign _EVAL_643 = _EVAL_1545 & _EVAL_3693;
  assign _EVAL_2245 = _EVAL_3781 & _EVAL_3040;
  assign _EVAL_3951 = _EVAL_3059 & _EVAL_3820;
  assign _EVAL_3824 = _EVAL_2874 & _EVAL_2758;
  assign _EVAL_3396 = _EVAL_668 & _EVAL_246;
  assign _EVAL_2093 = _EVAL_2549 != 127'h0;
  assign _EVAL_1703 = _EVAL_1522 & _EVAL_169;
  assign _EVAL_213 = _EVAL_1034 & _EVAL_3180;
  assign _EVAL_1832 = _EVAL_1545 & _EVAL_543;
  assign _EVAL_937 = _EVAL_1522 & _EVAL_887;
  assign _EVAL_3544 = _EVAL_1522 & _EVAL_543;
  assign _EVAL_3785 = _EVAL_1470 & _EVAL_1145;
  assign _EVAL_1482 = _EVAL_1420 & _EVAL_920;
  assign _EVAL_3288 = _EVAL_3458 & _EVAL_3148;
  assign _EVAL_192 = _EVAL_2804 & _EVAL_803;
  assign _EVAL_1363 = _EVAL_1553 & _EVAL_1245;
  assign _EVAL_3916 = _EVAL_1553 & _EVAL_655;
  assign _EVAL_2967 = _EVAL_3781 & _EVAL_916;
  assign _EVAL_1513 = _EVAL_2967 & _EVAL_246;
  assign _EVAL_972 = _EVAL_1513 & _EVAL_1417;
  assign _EVAL_3521 = _EVAL_1545 & _EVAL_3920;
  assign _EVAL_3131 = _EVAL_1040 & _EVAL_1324;
  assign _EVAL_2994 = _EVAL_4058 & _EVAL_246;
  assign _EVAL_235 = _EVAL_1553 & _EVAL_4006;
  assign _EVAL_1165 = _EVAL_442 & _EVAL_246;
  assign _EVAL_2661 = _EVAL_1165 & _EVAL_1996;
  assign _EVAL_1011 = _EVAL_1545 & _EVAL_3989;
  assign _EVAL_3129 = _EVAL_1426 & _EVAL_246;
  assign _EVAL_1348 = _EVAL_3059 & _EVAL_1240;
  assign _EVAL_2149 = _EVAL_1348 & _EVAL_2267;
  assign _EVAL_746 = _EVAL_2149 & _EVAL_1910;
  assign _EVAL_1733 = _EVAL_1545 & _EVAL_1621;
  assign _EVAL_2964 = _EVAL_1822 & _EVAL_2456;
  assign _EVAL_2598 = _EVAL_3058 & _EVAL_1910;
  assign _EVAL_3077 = _EVAL_3849 & _EVAL_1910;
  assign _EVAL_850 = _EVAL_3402 & _EVAL_1646;
  assign _EVAL_1028 = _EVAL_850 & _EVAL_246;
  assign _EVAL_2028 = _EVAL_2804 & _EVAL_806;
  assign _EVAL_993 = _EVAL_1034 & _EVAL_696;
  assign _EVAL_645 = _EVAL_3778 & _EVAL_996;
  assign _EVAL_1770 = _EVAL_1735 & _EVAL_1884;
  assign _EVAL_3452 = _EVAL_1480 & _EVAL_2267;
  assign _EVAL_3178 = _EVAL_3162 & _EVAL_1417;
  assign _EVAL_2878 = _EVAL_3104 & _EVAL_1417;
  assign _EVAL_2626 = _EVAL_3075 & _EVAL_2344;
  assign _EVAL_1193 = _EVAL_3717 & _EVAL_246;
  assign _EVAL_2727 = _EVAL_2275 & _EVAL_1417;
  assign _EVAL_1974 = _EVAL_1279 & _EVAL_2587;
  assign _EVAL_2238 = _EVAL_1279 & _EVAL_1889;
  assign _EVAL_1147 = _EVAL_3897 & _EVAL_2824;
  assign _EVAL_1712 = _EVAL_1158 & _EVAL_246;
  assign _EVAL_3956 = _EVAL_1712 & _EVAL_1996;
  assign _EVAL_3559 = _EVAL_1678 & _EVAL_1417;
  assign _EVAL_1030 = _EVAL_1223 & _EVAL_1996;
  assign _EVAL_650 = _EVAL_1129 & _EVAL_1417;
  assign _EVAL_1367 = _EVAL_1034 & _EVAL_4031;
  assign _EVAL_1299 = _EVAL_1312 & _EVAL_246;
  assign _EVAL_2343 = _EVAL_3496 & _EVAL_996;
  assign _EVAL_3727 = _EVAL_3538 & _EVAL_246;
  assign _EVAL_1739 = _EVAL_3727 & _EVAL_1417;
  assign _EVAL_1607 = _EVAL_3075 & _EVAL_3209;
  assign _EVAL_2405 = _EVAL_2472 & _EVAL_1417;
  assign _EVAL_1673 = _EVAL_2894 & _EVAL_1996;
  assign _EVAL_3840 = _EVAL_2112 & _EVAL_4012;
  assign _EVAL_3748 = _EVAL_431 & _EVAL_2961;
  assign _EVAL_3626 = _EVAL_3075 & _EVAL_1889;
  assign _EVAL_1359 = _EVAL_3321 & _EVAL_1910;
  assign _EVAL_798 = _EVAL_2112 & _EVAL_3209;
  assign _EVAL_3276 = _EVAL_3781 & _EVAL_1947;
  assign _EVAL_370 = _EVAL_3276 & _EVAL_246;
  assign _EVAL_2892 = _EVAL_3075 & _EVAL_3241;
  assign _EVAL_593 = _EVAL_2403 & _EVAL_1996;
  assign _EVAL_701 = _EVAL_2733 & _EVAL_1996;
  assign _EVAL_3786 = _EVAL_1470 & _EVAL_1354;
  assign _EVAL_2075 = _EVAL_1926 & _EVAL_2267;
  assign _EVAL_3175 = _EVAL_2075 & _EVAL_1910;
  assign _EVAL_3448 = _EVAL_3402 & _EVAL_3934;
  assign _EVAL_2717 = _EVAL_3448 & _EVAL_246;
  assign _EVAL_588 = _EVAL_2717 & _EVAL_1996;
  assign _EVAL_2562 = _EVAL_1007 & _EVAL_246;
  assign _EVAL_2223 = _EVAL_2562 & _EVAL_1996;
  assign _EVAL_3414 = _EVAL_1553 & _EVAL_2344;
  assign _EVAL_1573 = _EVAL_145 & _EVAL_246;
  assign _EVAL_1302 = _EVAL_3059 & _EVAL_2303;
  assign _EVAL_1101 = _EVAL_1561 & _EVAL_2267;
  assign _EVAL_2385 = _EVAL_1101 & _EVAL_1910;
  assign _EVAL_2152 = _EVAL_3897 & _EVAL_3693;
  assign _EVAL_2461 = _EVAL_3781 & _EVAL_2380;
  assign _EVAL_799 = _EVAL_2461 & _EVAL_246;
  assign _EVAL_636 = _EVAL_2027 & _EVAL_1910;
  assign _EVAL_1928 = _EVAL_3075 & _EVAL_1963;
  assign _EVAL_2819 = _EVAL_1470 & _EVAL_2756;
  assign _EVAL_1374 = _EVAL_2738 != 29'h0;
  assign _EVAL_1508 = _EVAL_3126 & _EVAL_1996;
  assign _EVAL_1520 = _EVAL_2887 & _EVAL_246;
  assign _EVAL_1518 = _EVAL_1520 & _EVAL_1417;
  assign _EVAL_754 = _EVAL_1719 & _EVAL_1417;
  assign _EVAL_2244 = _EVAL_855 & _EVAL_1910;
  assign _EVAL_2592 = _EVAL_3781 & _EVAL_789;
  assign _EVAL_2927 = _EVAL_2592 & _EVAL_246;
  assign _EVAL_3183 = _EVAL_2927 & _EVAL_1417;
  assign _EVAL_1968 = _EVAL_1538 & _EVAL_2267;
  assign _EVAL_3475 = _EVAL_1968 & _EVAL_1910;
  assign _EVAL_713 = _EVAL_3592 & _EVAL_246;
  assign _EVAL_620 = _EVAL_3781 & _EVAL_999;
  assign _EVAL_1665 = _EVAL_2112 & _EVAL_2961;
  assign _EVAL_572 = _EVAL_1553 & _EVAL_3087;
  assign _EVAL_3223 = _EVAL_340 & _EVAL_1910;
  assign _EVAL_3576 = _EVAL_3402 & _EVAL_3286;
  assign _EVAL_2271 = _EVAL_3576 & _EVAL_246;
  assign _EVAL_3915 = _EVAL_1724 & _EVAL_662;
  assign _EVAL_2224 = _EVAL_1543 & _EVAL_1910;
  assign _EVAL_513 = _EVAL_1573 & _EVAL_1417;
  assign _EVAL_1285 = _EVAL_1470 & _EVAL_3920;
  assign _EVAL_2935 = _EVAL_1340 & _EVAL_1417;
  assign _EVAL_729 = _EVAL_3951 & _EVAL_2267;
  assign _EVAL_317 = _EVAL_729 & _EVAL_1910;
  assign _EVAL_2384 = _EVAL_3897 & _EVAL_1145;
  assign _EVAL_3578 = _EVAL_1545 & _EVAL_520;
  assign _EVAL_2175 = _EVAL_2357 & _EVAL_1417;
  assign _EVAL_2988 = _EVAL_1470 & _EVAL_2769;
  assign _EVAL_2296 = _EVAL_3612 & _EVAL_2267;
  assign _EVAL_1593 = _EVAL_1553 & _EVAL_2339;
  assign _EVAL_3084 = _EVAL_3781 & _EVAL_1778;
  assign _EVAL_1247 = _EVAL_3084 & _EVAL_246;
  assign _EVAL_647 = _EVAL_1279 & _EVAL_2072;
  assign _EVAL_3420 = _EVAL_1522 & _EVAL_3148;
  assign _EVAL_3474 = _EVAL_1588 & _EVAL_1417;
  assign _EVAL_1994 = _EVAL_1470 & _EVAL_3148;
  assign _EVAL_3622 = _EVAL_3075 & _EVAL_803;
  assign _EVAL_3430 = _EVAL_3897 & _EVAL_3470;
  assign _EVAL_1898 = _EVAL_3458 & _EVAL_2691;
  assign _EVAL_422 = _EVAL_3781 & _EVAL_435;
  assign _EVAL_932 = _EVAL_422 & _EVAL_246;
  assign _EVAL_1149 = _EVAL_2112 & _EVAL_1224;
  assign _EVAL_944 = _EVAL_1545 & _EVAL_2984;
  assign _EVAL_3624 = _EVAL_1553 & _EVAL_2072;
  assign _EVAL_3926 = _EVAL_756 & _EVAL_1996;
  assign _EVAL_3268 = _EVAL_3402 & _EVAL_1791;
  assign _EVAL_3533 = _EVAL_2804 & _EVAL_2344;
  assign _EVAL_2098 = _EVAL_1040 & _EVAL_2020;
  assign _EVAL_3168 = _EVAL_501 & _EVAL_1910;
  assign _EVAL_3752 = _EVAL_3140 & _EVAL_1098;
  assign _EVAL_1851 = _EVAL_1724 & _EVAL_424;
  assign _EVAL_2821 = _EVAL_1606 & _EVAL_1996;
  assign _EVAL_625 = _EVAL_3075 & _EVAL_806;
  assign _EVAL_338 = _EVAL_2400 & _EVAL_1996;
  assign _EVAL_2538 = _EVAL_266 & _EVAL_1996;
  assign _EVAL_2371 = _EVAL_2711 & _EVAL_1996;
  assign _EVAL_587 = _EVAL_933 & _EVAL_2456;
  assign _EVAL_3826 = _EVAL_1279 & _EVAL_3779;
  assign _EVAL_2876 = _EVAL_3458 & _EVAL_1145;
  assign _EVAL_3130 = _EVAL_431 & _EVAL_3194;
  assign _EVAL_414 = _EVAL_3059 & _EVAL_1213;
  assign _EVAL_861 = _EVAL_414 & _EVAL_2267;
  assign _EVAL_3250 = _EVAL_861 & _EVAL_1910;
  assign _EVAL_596 = _EVAL_2986 & _EVAL_3471;
  assign _EVAL_2842 = _EVAL_2700 & _EVAL_246;
  assign _EVAL_708 = _EVAL_2842 & _EVAL_1996;
  assign _EVAL_3307 = _EVAL_1553 & _EVAL_2587;
  assign _EVAL_3979 = _EVAL_2804 & _EVAL_2961;
  assign _EVAL_2315 = _EVAL_3781 & _EVAL_1575;
  assign _EVAL_2274 = _EVAL_1279 & _EVAL_4006;
  assign _EVAL_173 = _EVAL_3848 & _EVAL_246;
  assign _EVAL_230 = _EVAL_3781 & _EVAL_2901;
  assign _EVAL_2381 = _EVAL_230 & _EVAL_246;
  assign _EVAL_1150 = _EVAL_2381 & _EVAL_1417;
  assign _EVAL_3732 = _EVAL_1812 & _EVAL_1417;
  assign _EVAL_2394 = _EVAL_196 & _EVAL_2267;
  assign _EVAL_1494 = _EVAL_3059 & _EVAL_3454;
  assign _EVAL_2368 = _EVAL_1494 & _EVAL_2267;
  assign _EVAL_2116 = _EVAL_2368 & _EVAL_1910;
  assign _EVAL_1276 = _EVAL_3805 & _EVAL_1996;
  assign _EVAL_351 = _EVAL_2986 & _EVAL_1224;
  assign _EVAL_2487 = _EVAL_3402 & _EVAL_2692;
  assign _EVAL_259 = _EVAL_2487 & _EVAL_246;
  assign _EVAL_4018 = _EVAL_259 & _EVAL_1996;
  assign _EVAL_2987 = _EVAL_1034 & _EVAL_3145;
  assign _EVAL_2132 = _EVAL_2296 & _EVAL_1910;
  assign _EVAL_2495 = _EVAL_1039 & _EVAL_1996;
  assign _EVAL_2255 = _EVAL_3577 & _EVAL_1910;
  assign _EVAL_782 = _EVAL_1545 & _EVAL_3000;
  assign _EVAL_3360 = _EVAL_3129 & _EVAL_1417;
  assign _EVAL_1412 = _EVAL_1034 & _EVAL_2587;
  assign _EVAL_560 = _EVAL_1652 & _EVAL_246;
  assign _EVAL_1413 = _EVAL_1724 & _EVAL_2824;
  assign _EVAL_1649 = _EVAL_3059 & _EVAL_2234;
  assign _EVAL_1463 = _EVAL_1649 & _EVAL_2267;
  assign _EVAL_2735 = _EVAL_1463 & _EVAL_1910;
  assign _EVAL_394 = _EVAL_2417 & _EVAL_1417;
  assign _EVAL_2297 = _EVAL_2804 & _EVAL_1889;
  assign _EVAL_382 = _EVAL_1034 & _EVAL_1048;
  assign _EVAL_3073 = _EVAL_1545 & _EVAL_2020;
  assign _EVAL_3855 = _EVAL_1545 & _EVAL_724;
  assign _EVAL_624 = _EVAL_3813 & _EVAL_1996;
  assign _EVAL_1568 = _EVAL_1724 & _EVAL_3920;
  assign _EVAL_580 = _EVAL_2738 == 29'h1fffffff;
  assign _EVAL_174 = _EVAL_3669 & _EVAL_580;
  assign _EVAL_3251 = _EVAL_243 & _EVAL_1910;
  assign _EVAL_3484 = _EVAL_3781 & _EVAL_3333;
  assign _EVAL_2811 = _EVAL_3484 & _EVAL_246;
  assign _EVAL_3343 = _EVAL_2811 & _EVAL_1417;
  assign _EVAL_288 = _EVAL_1470 & _EVAL_543;
  assign _EVAL_1346 = _EVAL_3458 & _EVAL_3920;
  assign _EVAL_1154 = _EVAL_1010 & _EVAL_2267;
  assign _EVAL_280 = _EVAL_1154 & _EVAL_1910;
  assign _EVAL_2471 = _EVAL_2804 & _EVAL_1245;
  assign _EVAL_3271 = _EVAL_1040 & _EVAL_3989;
  assign _EVAL_3477 = _EVAL_3594 & _EVAL_215;
  assign _EVAL_3105 = _EVAL_1724 & _EVAL_2412;
  assign _EVAL_2270 = _EVAL_2804 & _EVAL_398;
  assign _EVAL_737 = _EVAL_1822 & _EVAL_2506;
  assign _EVAL_664 = _EVAL_1589 & _EVAL_1417;
  assign _EVAL_1389 = _EVAL_1034 & _EVAL_3779;
  assign _EVAL_1796 = _EVAL_3897 & _EVAL_1621;
  assign _EVAL_2925 = _EVAL_3046 & _EVAL_2267;
  assign _EVAL_769 = _EVAL_2925 & _EVAL_1910;
  assign _EVAL_1115 = _EVAL_3075 & _EVAL_398;
  assign _EVAL_2814 = _EVAL_385 & _EVAL_2267;
  assign _EVAL_531 = _EVAL_2814 & _EVAL_1910;
  assign _EVAL_1656 = _EVAL_1522 & _EVAL_3285;
  assign _EVAL_970 = _EVAL_897 & _EVAL_1996;
  assign _EVAL_1569 = _EVAL_456 & _EVAL_1996;
  assign _EVAL_2036 = _EVAL_2173 & _EVAL_2544;
  assign _EVAL_2833 = _EVAL_1604 & _EVAL_246;
  assign _EVAL_253 = _EVAL_1034 & _EVAL_1889;
  assign _EVAL_3548 = _EVAL_2836 & _EVAL_1417;
  assign _EVAL_1546 = _EVAL_1406 & _EVAL_1996;
  assign _EVAL_2349 = _EVAL_1724 & _EVAL_724;
  assign _EVAL_3007 = _EVAL_1724 & _EVAL_3470;
  assign _EVAL_844 = _EVAL_2112 & _EVAL_3180;
  assign _EVAL_1657 = _EVAL_1724 & _EVAL_3038;
  assign _EVAL_3630 = _EVAL_1279 & _EVAL_3471;
  assign _EVAL_901 = _EVAL_1411 & _EVAL_1996;
  assign _EVAL_278 = _EVAL_1034 & _EVAL_3087;
  assign _EVAL_2178 = _EVAL_264 & _EVAL_1910;
  assign _EVAL_2997 = _EVAL_1822 & _EVAL_2756;
  assign _EVAL_771 = _EVAL_3059 & _EVAL_3579;
  assign _EVAL_3787 = _EVAL_2986 & _EVAL_2043;
  assign _EVAL_2888 = _EVAL_3897 & _EVAL_3148;
  assign _EVAL_314 = _EVAL_620 & _EVAL_246;
  assign _EVAL_2409 = _EVAL_314 & _EVAL_1417;
  assign _EVAL_1732 = _EVAL_4035 & _EVAL_1417;
  assign _EVAL_3900 = _EVAL_469 & _EVAL_1910;
  assign _EVAL_2920 = _EVAL_1470 & _EVAL_2824;
  assign _EVAL_1797 = _EVAL_1299 & _EVAL_1996;
  assign _EVAL_4014 = _EVAL_2112 & _EVAL_655;
  assign _EVAL_2345 = _EVAL_1040 & _EVAL_662;
  assign _EVAL_437 = _EVAL_1522 & _EVAL_3000;
  assign _EVAL_3609 = _EVAL_3163 & _EVAL_2267;
  assign _EVAL_976 = _EVAL_3609 & _EVAL_1910;
  assign _EVAL_2723 = _EVAL_3792 & _EVAL_1996;
  assign _EVAL_2896 = _EVAL_932 & _EVAL_1417;
  assign _EVAL_3912 = _EVAL_3160 & _EVAL_1996;
  assign _EVAL_3114 = _EVAL_1040 & _EVAL_3470;
  assign _EVAL_495 = _EVAL_3666 & _EVAL_1996;
  assign _EVAL_751 = _EVAL_560 & _EVAL_1417;
  assign _EVAL_3518 = _EVAL_1054 & _EVAL_1996;
  assign _EVAL_282 = _EVAL_3616 & _EVAL_2267;
  assign _EVAL_3478 = _EVAL_282 & _EVAL_1910;
  assign _EVAL_3905 = _EVAL_1034 & _EVAL_398;
  assign _EVAL_2424 = _EVAL_2897 & _EVAL_1417;
  assign _EVAL_2523 = _EVAL_1000 & _EVAL_1417;
  assign _EVAL_1762 = _EVAL_1900 & _EVAL_1417;
  assign _EVAL_1893 = _EVAL_1028 & _EVAL_1996;
  assign _EVAL_2422 = _EVAL_1268 & _EVAL_1996;
  assign _EVAL_2243 = _EVAL_692 & _EVAL_1996;
  assign _EVAL_1794 = _EVAL_3897 & _EVAL_3000;
  assign _EVAL_2875 = _EVAL_1522 & _EVAL_1145;
  assign _EVAL_1260 = _EVAL_771 & _EVAL_2267;
  assign _EVAL_3647 = _EVAL_1260 & _EVAL_1910;
  assign _EVAL_1269 = _EVAL_1553 & _EVAL_3241;
  assign _EVAL_2490 = _EVAL_3075 & _EVAL_2043;
  assign _EVAL_745 = _EVAL_431 & _EVAL_3596;
  assign _EVAL_503 = _EVAL_3140 & _EVAL_1083;
  assign _EVAL_918 = _EVAL_2986 & _EVAL_4016;
  assign _EVAL_1495 = _EVAL_1522 & _EVAL_724;
  assign _EVAL_3425 = _EVAL_1545 & _EVAL_2691;
  assign _EVAL_3393 = _EVAL_713 & _EVAL_1417;
  assign _EVAL_3938 = _EVAL_1830 & _EVAL_1910;
  assign _EVAL_4047 = _EVAL_2112 & _EVAL_696;
  assign _EVAL_3254 = _EVAL_431 & _EVAL_3087;
  assign _EVAL_2462 = _EVAL_1384 & _EVAL_1417;
  assign _EVAL_1954 = _EVAL_1034 & _EVAL_4006;
  assign _EVAL_2135 = _EVAL_1857 & _EVAL_662;
  assign _EVAL_1909 = _EVAL_799 & _EVAL_1417;
  assign _EVAL_1020 = _EVAL_3496 & _EVAL_1083;
  assign _EVAL_425 = _EVAL_1822 & _EVAL_2758;
  assign _EVAL_2164 = _EVAL_3778 & _EVAL_3217;
  assign _EVAL_1443 = _EVAL_1174 & _EVAL_1417;
  assign _EVAL_3492 = _EVAL_2804 & _EVAL_3779;
  assign _EVAL_3971 = _EVAL_1247 & _EVAL_1417;
  assign _EVAL_1394 = _EVAL_2813 & _EVAL_1417;
  assign _EVAL_191 = _EVAL_1034 & _EVAL_2072;
  assign _EVAL_698 = _EVAL_1545 & _EVAL_424;
  assign _EVAL_3775 = _EVAL_4051 & _EVAL_246;
  assign _EVAL_3560 = _EVAL_3775 & _EVAL_1996;
  assign _EVAL_1347 = _EVAL_1553 & _EVAL_3363;
  assign _EVAL_3570 = _EVAL_2986 & _EVAL_3194;
  assign _EVAL_2973 = _EVAL_3458 & _EVAL_3038;
  assign _EVAL_487 = _EVAL_2884 & _EVAL_1417;
  assign _EVAL_2351 = _EVAL_1545 & _EVAL_3038;
  assign _EVAL_3793 = _EVAL_3075 & _EVAL_3087;
  assign _EVAL_3473 = _EVAL_1040 & _EVAL_424;
  assign _EVAL_2227 = _EVAL_3458 & _EVAL_3000;
  assign _EVAL_3205 = _EVAL_1398 & _EVAL_1098;
  assign _EVAL_761 = _EVAL_499 & _EVAL_1417;
  assign _EVAL_3712 = _EVAL_3458 & _EVAL_3954;
  assign _EVAL_2857 = _EVAL_1040 & _EVAL_2824;
  assign _EVAL_1467 = _EVAL_1895 & _EVAL_2319;
  assign _EVAL_3745 = _EVAL_1037 & _EVAL_246;
  assign _EVAL_2286 = _EVAL_3745 & _EVAL_1417;
  assign _EVAL_1272 = _EVAL_1193 & _EVAL_1417;
  assign _EVAL_3502 = _EVAL_983 & _EVAL_2267;
  assign _EVAL_2687 = _EVAL_1522 & _EVAL_2769;
  assign _EVAL_871 = _EVAL_3075 & _EVAL_215;
  assign _EVAL_1184 = _EVAL_1522 & _EVAL_2756;
  assign _EVAL_386 = _EVAL_1034 & _EVAL_2961;
  assign _EVAL_3808 = _EVAL_1865 & _EVAL_1417;
  assign _EVAL_2710 = _EVAL_1545 & _EVAL_1490;
  assign _EVAL_1824 = _EVAL_687 & _EVAL_2267;
  assign _EVAL_3875 = _EVAL_1724 & _EVAL_887;
  assign _EVAL_3362 = _EVAL_3402 & _EVAL_2901;
  assign _EVAL_2295 = _EVAL_2112 & _EVAL_2339;
  assign _EVAL_786 = _EVAL_431 & _EVAL_215;
  assign _EVAL_419 = _EVAL_1043 & _EVAL_1417;
  assign _EVAL_616 = _EVAL_3458 & _EVAL_2020;
  assign _EVAL_2918 = _EVAL_3268 & _EVAL_246;
  assign _EVAL_1981 = _EVAL_1470 & _EVAL_1324;
  assign _EVAL_206 = _EVAL_1857 & _EVAL_3000;
  assign _EVAL_4042 = _EVAL_2112 & _EVAL_1245;
  assign _EVAL_1436 = _EVAL_2112 & _EVAL_2344;
  assign _EVAL_2680 = _EVAL_256 & _EVAL_1996;
  assign _EVAL_1864 = _EVAL_1724 & _EVAL_2756;
  assign _EVAL_1993 = _EVAL_3362 & _EVAL_246;
  assign _EVAL_1579 = _EVAL_1302 & _EVAL_2267;
  assign _EVAL_3138 = _EVAL_1579 & _EVAL_1910;
  assign _EVAL_1262 = _EVAL_1016 & _EVAL_1417;
  assign _EVAL_177 = _EVAL_3093 & _EVAL_1910;
  assign _EVAL_726 = _EVAL_173 & _EVAL_1996;
  assign _EVAL_3925 = _EVAL_535 & _EVAL_1910;
  assign _EVAL_1972 = _EVAL_1034 & _EVAL_1963;
  assign _EVAL_2840 = _EVAL_4072 & _EVAL_1910;
  assign _EVAL_3108 = _EVAL_1969 & _EVAL_1885;
  assign _EVAL_2193 = _EVAL_1050 & _EVAL_1417;
  assign _EVAL_3311 = _EVAL_3075 & _EVAL_4006;
  assign _EVAL_3187 = _EVAL_1993 & _EVAL_1996;
  assign _EVAL_3034 = _EVAL_2041 & _EVAL_3408;
  assign _EVAL_3289 = _EVAL_3781 & _EVAL_3859;
  assign _EVAL_2431 = _EVAL_3289 & _EVAL_246;
  assign _EVAL_839 = _EVAL_2918 & _EVAL_1996;
  assign _EVAL_1627 = _EVAL_3897 & _EVAL_169;
  assign _EVAL_2282 = _EVAL_1551 & _EVAL_1417;
  assign _EVAL_2217 = _EVAL_2245 & _EVAL_246;
  assign _EVAL_1349 = _EVAL_2986 & _EVAL_696;
  assign _EVAL_1038 = _EVAL_2804 & _EVAL_4006;
  assign _EVAL_2019 = _EVAL_2804 & _EVAL_3596;
  assign _EVAL_3607 = _EVAL_1545 & _EVAL_662;
  assign _EVAL_4036 = _EVAL_1724 & _EVAL_1490;
  assign _EVAL_1303 = _EVAL_1358 & _EVAL_1996;
  assign _EVAL_1623 = _EVAL_2321 & _EVAL_1417;
  assign _EVAL_1435 = _EVAL_1782 & _EVAL_246;
  assign _EVAL_1478 = _EVAL_1034 & _EVAL_1245;
  assign _EVAL_2074 = _EVAL_1040 & _EVAL_3148;
  assign _EVAL_3483 = _EVAL_1522 & _EVAL_662;
  assign _EVAL_1385 = _EVAL_523 & _EVAL_1910;
  assign _EVAL_3182 = _EVAL_1857 & _EVAL_2830;
  assign _EVAL_3706 = _EVAL_1553 & _EVAL_3701;
  assign _EVAL_3902 = _EVAL_1034 & _EVAL_3596;
  assign _EVAL_2370 = _EVAL_1470 & _EVAL_3285;
  assign _EVAL_1757 = _EVAL_2392 & _EVAL_1996;
  assign _EVAL_1288 = _EVAL_3897 & _EVAL_3989;
  assign _EVAL_1529 = _EVAL_3224 & _EVAL_1910;
  assign _EVAL_3830 = _EVAL_2986 & _EVAL_655;
  assign _EVAL_151 = _EVAL_1857 & _EVAL_2375;
  assign _EVAL_3948 = _EVAL_2895 & _EVAL_1417;
  assign _EVAL_1932 = _EVAL_813 & _EVAL_246;
  assign _EVAL_3297 = _EVAL_1932 & _EVAL_1996;
  assign _EVAL_1308 = _EVAL_2112 & _EVAL_1889;
  assign _EVAL_3698 = _EVAL_1279 & _EVAL_3241;
  assign _EVAL_2655 = _EVAL_3838 & _EVAL_1996;
  assign _EVAL_2521 = _EVAL_1364 & _EVAL_2267;
  assign _EVAL_2360 = _EVAL_3512 & _EVAL_1374;
  assign _EVAL_227 = _EVAL_3092 & _EVAL_1910;
  assign _EVAL_1290 = _EVAL_1857 & _EVAL_3693;
  assign _EVAL_1896 = _EVAL_1470 & _EVAL_3038;
  assign _EVAL_490 = _EVAL_2041 & _EVAL_2319;
  assign _EVAL_2936 = _EVAL_3396 & _EVAL_1417;
  assign _EVAL_4008 = _EVAL_3651 & _EVAL_1417;
  assign _EVAL_3695 = _EVAL_2521 & _EVAL_1910;
  assign _EVAL_3403 = _EVAL_936 & _EVAL_1417;
  assign _EVAL_3814 = _EVAL_3458 & _EVAL_887;
  assign _EVAL_292 = _EVAL_1553 & _EVAL_4012;
  assign _EVAL_549 = _EVAL_2138 & _EVAL_1910;
  assign _EVAL_1095 = _EVAL_1869 & _EVAL_1910;
  assign _EVAL_1641 = _EVAL_3678 & _EVAL_1996;
  assign _EVAL_3202 = _EVAL_2986 & _EVAL_4012;
  assign _EVAL_3711 = _EVAL_1724 & _EVAL_3989;
  assign _EVAL_157 = _EVAL_2394 & _EVAL_1910;
  assign _EVAL_671 = _EVAL_3897 & _EVAL_2984;
  assign _EVAL_2474 = _EVAL_2173 & _EVAL_2456;
  assign _EVAL_1850 = _EVAL_1522 & _EVAL_3693;
  assign _EVAL_2170 = _EVAL_1857 & _EVAL_169;
  assign _EVAL_3657 = _EVAL_1034 & _EVAL_655;
  assign _EVAL_2761 = _EVAL_2833 & _EVAL_1996;
  assign _EVAL_4055 = _EVAL_1553 & _EVAL_4031;
  assign _EVAL_2998 = _EVAL_3417 & _EVAL_1996;
  assign _EVAL_3874 = _EVAL_1824 & _EVAL_1910;
  assign _EVAL_610 = _EVAL_3440 & _EVAL_1996;
  assign _EVAL_376 = _EVAL_2804 & _EVAL_696;
  assign _EVAL_2390 = _EVAL_1040 & _EVAL_1621;
  assign _EVAL_2453 = _EVAL_3897 & _EVAL_3038;
  assign _EVAL_240 = _EVAL_1661 & _EVAL_1910;
  assign _EVAL_852 = _EVAL_908 & _EVAL_1996;
  assign _EVAL_1586 = _EVAL_431 & _EVAL_3471;
  assign _EVAL_1882 = _EVAL_1420 & _EVAL_388;
  assign _EVAL_383 = _EVAL_1545 & _EVAL_2830;
  assign _EVAL_579 = _EVAL_2112 & _EVAL_4016;
  assign _EVAL_613 = _EVAL_1330 & _EVAL_1417;
  assign _EVAL_3978 = _EVAL_2602 & _EVAL_1417;
  assign _EVAL_1317 = _EVAL_933 & _EVAL_2758;
  assign _EVAL_582 = _EVAL_3402 & _EVAL_478;
  assign _EVAL_1046 = _EVAL_582 & _EVAL_246;
  assign _EVAL_2564 = _EVAL_1553 & _EVAL_3471;
  assign _EVAL_714 = _EVAL_3458 & _EVAL_3989;
  assign _EVAL_913 = _EVAL_2271 & _EVAL_1996;
  assign _EVAL_3004 = _EVAL_2217 & _EVAL_1417;
  assign _EVAL_3066 = _EVAL_2280 & _EVAL_1417;
  assign _EVAL_2926 = _EVAL_2431 & _EVAL_1417;
  assign _EVAL_1219 = _EVAL_1857 & _EVAL_3954;
  assign _EVAL_452 = _EVAL_1279 & _EVAL_1224;
  assign _EVAL_683 = _EVAL_2986 & _EVAL_2072;
  assign _EVAL_1111 = _EVAL_1040 & _EVAL_2375;
  assign _EVAL_1284 = _EVAL_2986 & _EVAL_803;
  assign _EVAL_224 = _EVAL_1545 & _EVAL_1354;
  assign _EVAL_3990 = _EVAL_2315 & _EVAL_246;
  assign _EVAL_1006 = _EVAL_1953 & _EVAL_1417;
  assign _EVAL_233 = _EVAL_2194 & _EVAL_2267;
  assign _EVAL_2123 = _EVAL_156 & _EVAL_1417;
  assign _EVAL_787 = _EVAL_2112 & _EVAL_1048;
  assign _EVAL_1825 = _EVAL_1470 & _EVAL_2412;
  assign _EVAL_995 = _EVAL_3398 & _EVAL_1417;
  assign _EVAL_3354 = _EVAL_431 & _EVAL_2339;
  assign _EVAL_1388 = _EVAL_2904 & _EVAL_1417;
  assign _EVAL_1995 = _EVAL_1040 & _EVAL_543;
  assign _EVAL_733 = _EVAL_233 & _EVAL_1910;
  assign _EVAL_2262 = _EVAL_3452 & _EVAL_1910;
  assign _EVAL_1772 = _EVAL_2804 & _EVAL_1048;
  assign _EVAL_2067 = _EVAL_1279 & _EVAL_2043;
  assign _EVAL_2703 = _EVAL_1435 & _EVAL_1417;
  assign _EVAL_3739 = _EVAL_3075 & _EVAL_2587;
  assign _EVAL_1517 = _EVAL_2112 & _EVAL_398;
  assign _EVAL_2519 = _EVAL_1046 & _EVAL_1996;
  assign _EVAL_3211 = _EVAL_3897 & _EVAL_520;
  assign _EVAL_3111 = _EVAL_661 & _EVAL_1996;
  assign _EVAL_1592 = _EVAL_486 & _EVAL_1996;
  assign _EVAL_2466 = _EVAL_370 & _EVAL_1417;
  assign _EVAL_1220 = _EVAL_2994 & _EVAL_1996;
  assign _EVAL_2168 = _EVAL_1522 & _EVAL_2020;
  assign _EVAL_3033 = _EVAL_1522 & _EVAL_1621;
  assign _EVAL_2246 = _EVAL_3502 & _EVAL_1910;
  assign _EVAL_3708 = _EVAL_3704 & _EVAL_1417;
  assign _EVAL_510 = _EVAL_1545 & _EVAL_169;
  assign _EVAL_433 = _EVAL_3990 & _EVAL_1417;
  assign _EVAL_3200 = _EVAL_3897 & _EVAL_2594;
  assign TLMonitor__EVAL_0 = _EVAL_86;
  assign TLMonitor__EVAL_7 = _EVAL_131;
  assign TLMonitor__EVAL_5 = _EVAL_59;
  assign TLMonitor__EVAL_2 = _EVAL_51;
  assign TLMonitor__EVAL_13 = _EVAL_20;
  assign TLMonitor__EVAL = _EVAL_143;
  assign TLMonitor__EVAL_11 = Queue__EVAL_5;
  assign TLMonitor__EVAL_12 = _EVAL_69;
  assign TLMonitor__EVAL_8 = _EVAL_79;
  assign TLMonitor__EVAL_10 = _EVAL_291[1:0];
  assign TLMonitor__EVAL_1 = _EVAL_58;
  assign TLMonitor__EVAL_4 = _EVAL_142;
  assign TLMonitor__EVAL_6 = {{2'd0}, _EVAL_815};
  assign TLMonitor__EVAL_3 = _EVAL_105;
  assign TLMonitor__EVAL_9 = Queue__EVAL_12;
  assign TLMonitor__EVAL_14 = _EVAL_291[13:2];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_1327 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {4{`RANDOM}};
  _EVAL_3531 = _RAND_1[126:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_3861 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_142) begin
    if (_EVAL_105) begin
      _EVAL_1327 <= 1'h0;
    end else begin
      if (_EVAL_3610) begin
        _EVAL_1327 <= _EVAL_3856;
      end
    end
    _EVAL_3531 <= _EVAL_2527 & _EVAL_3572;
    if (_EVAL_105) begin
      _EVAL_3861 <= 1'h0;
    end else begin
      if (_EVAL_3610) begin
        _EVAL_3861 <= _EVAL_1990;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e9aafeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3460 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b868c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3795 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c09a6e2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2175 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7b6a93d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2360 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1576 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c437cbdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2770 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25186cbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3073 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95c768e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_656 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55687607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1118 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(169f8252)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ef59654)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2888 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ff1ab89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2212 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c37d86c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_745 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d16b2174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3604 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2609f161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82eb4b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4055 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef904156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2523 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54b39e10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2014 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78779897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2787 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ebf645d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_467 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a1a4f6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3748 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d62a339a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cabbc3f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1508 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86b3dada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2216 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0662945)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3922 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f35b623f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_844 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdee35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1696 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ebac427)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3819 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b8d6055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_993 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c7c66d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bf8e537)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1928 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8583551e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3767 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1efb3e33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4da6a65f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3845 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2f939ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d8e0f5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_532 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e28c900)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3700 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d716b4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2098 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b388ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2876 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40f054f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2223 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff992dc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c375f4cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1501 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8020867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3794 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(959cc2e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3703 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23c56401)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3660 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e281e33a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_984 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee417c73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_719 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4174f04d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3430 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(768b8345)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2678 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(641b990f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_579 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7126d78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3357 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35926fb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2116 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9fc399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_995 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd93be59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2945 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14ee59cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1592 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(543a514b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2879 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d5ce771)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_970 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f0dedb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_571 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27db0bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_647 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28514c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2409 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c80dc48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3422 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d757f902)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3068 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b303b4f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1707 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(719b7c7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1041 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea102e16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1733 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f145f0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1595 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9326cba5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2896 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ebbf6c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1285 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ebb96ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2934 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b250452)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1961 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad1aa68f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3876 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(289aceb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2351 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ae07125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3185 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9de9f5eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_513 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd92fb66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1850 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69842792)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1743 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c7418e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1147 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5431db8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25d836e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2785e72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1234 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2002 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71dcb49b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2654 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b309348f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2773 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9edd4bf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3131 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25b8b137)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_744 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9beae55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2795) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78c371e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1546 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1574995)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2349 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b59e56b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1842 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c9c549a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_463 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f4d2ea2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3375 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d450d9b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3730 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ce911a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3958 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c22e49ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2538 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaacf156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2906 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3be819e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2401 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38fa64e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2053 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a83e4586)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1436 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a117b423)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_425 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9d5f9b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1772 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(986c5c8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_636 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c7fb456)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_721 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85a70697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e232ba17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1847 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fb60646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7130698)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3723 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4620b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3725 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1beffc4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_678 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4936c1f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1662 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aad7811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1efbcf46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2556 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1497dff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4042 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf3f5dc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1972 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e96ea8ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1150 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d8c4a0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1058 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c93fca77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2865 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dfebd92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1964 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a37f76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff504738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3763 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9efbf9f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4036 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(463adac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_554 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8f00e42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1403 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab5b28d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3982 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e7e8f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2262 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aefe9ee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2213 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b415faf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1445 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(332a3223)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_838 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c1f33e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_972 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeb18e39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2377 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(deed2786)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_767 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1021ad68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3478 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eb79506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3574 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1cc236f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1382 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc939bad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3411 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61f73a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2048 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf8564e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c01ad95a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918722b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1641 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc24ecc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1443 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c940c7b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3208 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b4f0e06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2087 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3c45b7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2370 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c78d9c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2393 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e930e710)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1636 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d130bd29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2074 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cf2164f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4024 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a77642ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2046 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf3f1d67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1467 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(179ff943)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_680 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de1f1b46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3456 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf05df1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3197 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(937e87ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3787 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45c42c9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3328 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a22117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1797 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13d1efe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1220 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b59481b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_893 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64301352)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3658 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8db88cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2577 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1849c78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2583 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2dec1da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_576 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81e9165f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2019 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1900ef67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3307 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7bc5583)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3152 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6a9337c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3569 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(389b1258)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1126 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ac6b11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3076 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34c306ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3657 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b91760ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1841 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c67f98d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3086 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66f6a0a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2367 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0e19313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3457 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(560c3128)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3475 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f80dbfc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2255 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aed45b43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c2b5c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1656 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(388ec326)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2598 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eb4d7b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2620 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b75b5060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_717 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f7b16b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_751 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5edad709)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2794 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(899b08ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3741 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f33a635)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_877 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(655e2f62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69704538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3138 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1c7cc3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_659 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eddc0665)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2550 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb75b94f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_609 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa808b10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1146 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(829d0984)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_819 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c79c91a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_914 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b6bf82f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2176 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b29e6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4047 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f51df37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3250 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(361380fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3739 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c10923b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2490 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8e683ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1459 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ed5b155)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3716 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f13c680)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3916 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5db64224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2233 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d521daba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2569 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b26a57e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5b5b4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1166 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef59840e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3893 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17546d57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2687 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(793a5dcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2603 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ef11262)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1116 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78378fec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4092ff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da4fc7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2930 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba83315f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3200 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d01ae6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e37a5689)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f991fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3832 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f462d30e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2246 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebb2924c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3255 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cea277a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_754 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65c1141a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_541 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(297bc069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2272 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cabb04f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1272 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce59d462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2458 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a34329f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2825 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13cdb07d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dc726b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2390 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61c4b63b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bfd1aea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2264 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9c14917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3114 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f51f13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3284 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f61ce875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_466 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c90d84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3316 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3514af93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_674 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8a37e67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2614 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6708a2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3414 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ede3ad05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_625 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16045198)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e790a448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_951 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c71f9f9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1125 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cff88408)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1474 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d78e8a25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3183 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4dfede4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1478 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b9e908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2161 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20ebaa54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2405 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e932df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_872 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2702af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e0edf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1027 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32c96848)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3234 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9959b9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2160 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(914abc25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_783 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e581d510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2359 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8491e60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1739 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0d2874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3712 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43122749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3342 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eba6a4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1388 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14e33d9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdf3e0bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1924 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d37757f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_634 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3429e78c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2297 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ea0a39f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3506 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7aec368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1507 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ca293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1518 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64ce5d11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2270 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62c75522)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1149 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72f1c782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1534 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b122877f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1378 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c505259)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3986 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34df2394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_859 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(335a9dc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3007 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(658ad808)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1284 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5a8427f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3978 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9f9c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3785 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ec6324a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1065 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a552f014)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2474 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e3c9f5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2274 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf40d54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3988 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e29ab1a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3481 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22380dcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2284 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73e71190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_868 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ca4fef2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3635 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2df556cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3925 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(286e0ba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3948 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd4df460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1898 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9d02fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2067 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8d0cc21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2343 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a259bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2424 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4d2f531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1966 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a9760e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2466 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc98c52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2926 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(738db8c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3313 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(620bf1d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3902 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2591e783)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1087 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(920bb83f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1794 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64bb3b20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2028 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c56bf47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2857 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa2cb394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3483 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb3d3ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_892 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89c9e8e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3599 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdd79cac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2639 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a71f3c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f654927c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3435 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4c18f25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3840 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b26f7c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2422 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46bab563)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4007 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1f454c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3647 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5eaca5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1937 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b12def2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_593 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2afdaca3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2714 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edf38f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1982 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689ef4e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2903 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ae2e1ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3251 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49404dda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_627 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d800dbb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2402 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f67ebcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3793 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d5895fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4030 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9a33d6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1694 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(753ed9e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2878 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25507c3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_644 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65879bb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2396 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc6fcc69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2920 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f18d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2374 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f368172a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f3c92ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2785 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d95bfed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(709f2871)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1067 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b322779c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_817 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6715b1ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2177 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb3fdbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_761 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30bb11eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4194bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bca61797)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3034 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9833c5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_500 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9d70b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2244 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c8fe930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3998 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9be76ae5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3298 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f8e52c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2540 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7e3e34b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1012 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bea31146)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3630 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b489c6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b694ff6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_400 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c56162a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3168 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f18c3c74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1309 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a6ed96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3227 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e30508d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2324 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba7db74a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1882 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7fad00b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3764 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2858b36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2618 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99cf8130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3545 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b832d0d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(555a0d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1084 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a24cffa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3698 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5113286b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3223 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7a39679)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc51e46e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_432 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b4644c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3271 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d89dfe9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2428 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b8d49f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2740 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742eecc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1262 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8260b57d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3938 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15f20ba8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2193 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f1b4247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0d3c44b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2992 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a32577d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_676 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ba2389)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3064 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6506f631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2798 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7f12700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1344 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eec7860)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3461 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb6e6c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3116 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cd2dd1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2869 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd518d49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3161 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c74384f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3031 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbcc45b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1703 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(715c8703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2783 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9043f673)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_737 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f973d2d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0631d6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3937 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6036a79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1784 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(211b913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3754 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(716bb87f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2268 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8c3f934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1111 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d22f2929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3578 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c67c43a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3912 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed746ee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_860 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e27af28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1960 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f2764de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3924 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1220f0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2729 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8595b705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86ce8a0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f71cac42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1971 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c6fddff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3198 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf2a9a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2236 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce7d1393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54d7284f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1558 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23b2f7e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2476 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a30fc107)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3877 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dd4ceb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42a2a462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2373 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(939965eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1308 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc6580a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1732 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b5bea1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3311 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9174412f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3558 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a7c5d27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2681 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0868a39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2703 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3788dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1498 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c65ca43e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3874 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fad7bc4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2755 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1218fed5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2327 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88e40b29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c13322f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2632 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aa1c5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3555 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1d14dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_683 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4eac6c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1607 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63af7a2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2004 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67275845)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3420 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17868402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_714 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee706a35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b833df00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6874ce06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1089 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21c283d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2049) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3868be7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3389 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(223e027c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_651 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1be70b1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_635 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(864933fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1623 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(573dd715)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1949 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219796b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_498 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98547657)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b23d7944)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2170 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caa85850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_545 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9252f48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2414 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe01d358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4023 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(857529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_596 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c131d5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3077 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1452200d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2323 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f682bf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1033 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9cf584a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3518 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7beabde6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3193 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aa56521)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2839 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29a08ff3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1396 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe6fb7ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1714 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2a087a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2998 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3b0d031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2890 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f10322d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(737f03f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2964 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0b1eee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3176 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d6106a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d47fed08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1773 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(661b0e47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2566 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e0669e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2130 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70ea6007)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad77a775)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2935 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f5ce52d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1904 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6050303a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1271 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69818a17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2143 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(107699ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3855 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c23b8a07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1627 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(813dd588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1238 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78cab82f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1829 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e80f44b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2109 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a03fc15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1276 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec7cce80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3637 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9c888db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_862 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dd52ac7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3826 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(912d3750)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1854 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(804fd8a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3940 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8c291e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1367 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9c697a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_610 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff0c4dc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2517 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c9ed3ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1115 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c45e264a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2840 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2329893a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2182 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d8c53db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1233 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9be1b00c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_419 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df323a7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1911 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71fa1221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9651fa1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2099 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b2d3f2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48d3bfa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1389 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5bd66ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3862 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(551e4357)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e56155e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1472 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ced6870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2630 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d994aa0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1316 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b894d35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3752 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7c75ad2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_392 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7bdceac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1008 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52009089)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1139 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa6f885)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1355 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4410704)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2776 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d6973bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1570 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c480ca0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c13031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2643 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4556106b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2647 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(449f0e71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(762af327)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2235 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a90bfeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_327 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75a3a216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2077 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(995137b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3971 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9310337c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2337 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fccfc207)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_769 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b78e230c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2671 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf7ce9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3346 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba64244e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_708 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba562fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3324 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da2a796b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_667 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7a33e98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1653 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e31f8aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3774 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c3d1f5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3202 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90f99e5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a73e90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75e40229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1798 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36740d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3544 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2549e7c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2849 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6cd7260)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1120 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a293f4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_991 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a879131b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1995 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76865716)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2819 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3409 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d151dbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_839 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a94f287a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3473 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b56a6be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3979 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73c56957)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1336 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(625c2ee4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_503 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20d644a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1510 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16b42f7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2295 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b5a916c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a7c034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_965 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae29c1a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_733 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eff14e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1431 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ebf38e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2469 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd3ec50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0423a6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1428 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7063542b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_677 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a7a75f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2009 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feeb400)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_782 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cd9fb09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2036 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93378c20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1314 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93e92463)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1529 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c8d40d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3654 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7bd4a87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2222 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(908bfddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_796 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(873e1096)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_440 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae7139c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3812 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75cda347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_937 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2739db1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_948 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(901410de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3967 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4f69134)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2679 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f6fa743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2845 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b206727)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(385ccfdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1548 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f52c2d79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_671 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(972898b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c29618a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3153 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78595d97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_430 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98f921aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3492 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be84db39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aaff4ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3171 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a4bc4a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_949 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7a69538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3830 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d047649d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2657 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74cf9a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13c23158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28ce0b6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2135 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33103382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2462 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e77726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3187 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b34eed20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_376 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c595a33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2001 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d93ce5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_518 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdbef918)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3521 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b8ae9b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1482 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b749752)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2709 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7e28e5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1082 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97b524b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_755 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67334c36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3360 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(610161af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1532 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7780dae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2515 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1c4858a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3474 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c5008f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb69e9e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2987 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9cf06c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2591 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96831010)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3511 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f4319f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2180 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b206283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3533 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d5a29a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_740 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf8c9cf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3854 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8a7dd9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1117 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a153f51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2512 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8e6b483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_686 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f1316e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2093 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38ec23e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2660 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(757d7345)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_660 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64ff547f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1517 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f35f8124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3345 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f1e9bb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3997 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f80d2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_804 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26054a65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3254 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce952057)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4045 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3f5d69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1909 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cccb03d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3366 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8515992c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7288eda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4008 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(754f2932)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2564 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbf8cc51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3842 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98617347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2326 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8142a19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1484 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b25036b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1219 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(246c6ade)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2962 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(687a2115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_649 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b27cd645)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_454 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6079d3da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2227 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ba119e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2668 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3969a91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3257 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ecd015d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3178 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeb69876)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2723 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f5a39bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2822 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dce6e87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1775 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bc4e8e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2905 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fb0443f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1184 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ddfcd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_697 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5da56a6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b0f884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3886 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc6ac260)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3288 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59b2a264)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2505 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab98eaf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_433 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5e5e5cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1006 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c73238d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2997 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cdeb206)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(948d65e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2132 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(278450d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3395 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33eeee9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3010 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6a6204)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2185 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c5ca665)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2408 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b34ed6a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1281 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8770f90d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1806 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da9f732)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3090 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b46097f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85527eae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1715 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59902093)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3956 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b65f04e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1755 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e69d04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3128 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1807f28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3465 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba029920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3915 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c0600f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1493 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bfcfdd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2200 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77cab69f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2e81fba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2152 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3205 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c67cad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_752 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dc4b1b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_564 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b565831b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3539 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade69ebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2030 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeed6087)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1178 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(539167e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3108 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0e7aa39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3900 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3981011b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1317 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a0faf12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3865 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d76dad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3901 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b14bc221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50820a74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3386 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a23a63b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2168 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f610782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1655 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6338da0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(975e9214)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2892 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(218a5b15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2946 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb5e76d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1011 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd8b2162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1095 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ce4668c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2753 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fefde68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3593 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81ee5f86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3833 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb34ce63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_528 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbbc0faf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2423 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb0d6ffe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_961 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(558f80e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1670 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf940ce9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2298 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f8eea85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3211 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(569b4f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_487 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9369059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2672 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b46a7c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3618 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d08dc4e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1461 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc7911cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3264 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69021ab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa49397e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4071 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3956936d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3368 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a7eb93f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1295 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d14dbed5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2534 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93519a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1974 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e8130c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3541) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d5c4cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2674 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ddfeb1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1056 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9235432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2285 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8fb913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3875 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d08a8e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4061 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d46add85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(178261a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3369 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43abd052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2015 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e35e256d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_484 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b478bcec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3425 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c076f2c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_568 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f9fd102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1079 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3bb5182)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_612 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be43bc74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1337 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c273ef36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfbf7e94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3532 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50359124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1691 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b388337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_701 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adadeb6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f79a023d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_619 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99f5c89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3353 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(392396b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3708 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(172ca0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2655 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecaaa4b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3427 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(891ccede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2626 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95acf987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1161 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fda113a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3650 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93e7c2ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1840 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b072819)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_479 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c344277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3119 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e293c64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2509 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c29f7322)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4018 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc88272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2426 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6032f8e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1303 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a83b4276)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1695 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d44b8efd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1762 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5325b35c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1514 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8109a88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1020 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(739b37a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3738 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2886a42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3449 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ab790e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7091d7ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2199 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3553db0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2411 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5032c0fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_746 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a42ea557)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3786 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4100740)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1766 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88b7a23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3341 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd22bc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2696 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9de67957)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2875 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f37c9dff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_901 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(571743e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1908 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(491a8d15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1419 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(551de8cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_490 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53e64fa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(effcb701)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1618c580)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1693 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7c939e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1071 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60ff089d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_426 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30b52d6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9df72bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2547 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06932ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3517 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7623fc67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c507e6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3130 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cac69e35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60e3a939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1591 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dda026ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3297 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb79605e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2313 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84b65dd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2420717f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3004 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8aa10ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1363 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea31affc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1157 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39bc7191)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2800 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(552914e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2413 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95b49dbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3622 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33562f6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2089 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a094b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2201 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76367f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1334 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a76c2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1003 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bd6a49e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1457 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(748297b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1203 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c44be8ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3808 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(653a4a4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1288 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ffe10e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(292c1bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1893 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(344b71ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2493 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad68c089)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5d6e0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1025 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38835e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1994 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c6da40f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3926 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edffa987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2338 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(231f5f5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2224 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ca0fb5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_726 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b14335e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1015 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a1ab988)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3105 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc1e606)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1395 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc8d5c82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3343 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edce4c42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4014 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdf1f9c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3337 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b787d497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2563 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8a58ca5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2829 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc1836e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3437 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41ae2315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1569 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c33379dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4207ac1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2795) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_451 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83973aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3648 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c0344f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_406 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39a22803)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3824 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ecf417e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3537 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6576754b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3444 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2ca2da9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3003 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f7aad32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3393 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d7a0b68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_876 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(add470d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2266 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1845dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_992 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98d30e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_749 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9432611b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_777 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89e2be3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3744 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487b97c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2519 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8e13476)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3929 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e608fac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3619 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53767324)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1975 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9358332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_471 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d9f618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6b05c45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1359 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2825f632)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3472 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(909c97a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2652 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ff2a178)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3536 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1204d451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_531 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e9da874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_706 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f97f158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2395 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3644903b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2345 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68aadee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1044 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(877b7f61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1346 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6cc5c34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e0f406)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_866 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b76a47e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2453 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2028723c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1042 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1aec81b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1031 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3e100e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3681 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a2f14c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3322 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a53ff0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2622 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d22cffe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1290 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3b90b6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1140 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b026c2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7be328)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3753 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4929ba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2364 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33fe48f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29c64afa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1342 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6024ea7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_950 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(958a72cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1001 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32307201)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1825 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c79bb01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1567 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0998bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2604 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57857f53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1878 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3641b81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_685 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(703c4d5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3695 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57a12214)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3598 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8f03cda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3067 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(808c54c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3191 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(895b3e16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0b3dd10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_654 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69e1379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_900 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f973db81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3742 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2ecddb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3726 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816fa2e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1228 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5cf5f33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3019 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65d01191)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_394 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b4bbd84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1187 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c849e3ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11017852)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_975 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a69bd6c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1796 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a334c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3711 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(415f5ed7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2057 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39a517fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3656 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc8d1cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2710 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(189c8e10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4057 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b89b333)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_857 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60c679d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4067 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5949271c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3714 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(908cad22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1361 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fae71bf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1347 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ca60d34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1138 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dedc94ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2529 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c968443c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3355 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a1be0c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2862 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4d91c25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1563 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a64839f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba0fef74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_863 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c454fb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3302 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(732342a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1183 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83de27b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2663 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(404240cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3229 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bad7195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1030 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a615f9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3633 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a62016)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2693 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6708bf72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2916 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb97356f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3914 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(301b94d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1844 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8abc80dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1600 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(786184b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aecf6c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3639 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2299162c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_904 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48a8f903)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2661 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5695adb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1205 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be1a358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1657 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(340f97b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2533 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4bea6a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3144 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6806a44c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1586 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba142726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3498 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fec1afd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2243 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6192faf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2973 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7767c30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6b1ce17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2450 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93aebb7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8aef796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2495 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7b6e41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3005 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d8a1875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_980 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d756aab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2123 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5390d02c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3480 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91b0c8c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3814 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62db877a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3349 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe92366c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3939 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(836178e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1957 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e710c458)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1832 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7af87ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1902 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab6de5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1954 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6805247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2371 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a680b7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_698 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1201e89a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_453 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1577ccb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2511 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(562ada94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d24299fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2635 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a222e102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2218 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4ae15e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7789836c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4001 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24f3dd35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3541) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3111 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5379d56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3976 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5211597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2178 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5f6eabe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2599 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfba3be8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1851 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a912395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3482 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e048a738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1692 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e447b17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3249 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2db54f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1356 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ca43531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2855 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9d19051)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2680 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aea6695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1a68706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1581 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18451ed4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1803 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96f99d2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3559 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99b1c640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1394 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afdb609)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1232 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92052c16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3495fbc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4046 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fece5d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3560 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(639260d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2736 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab64ec8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1112 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e582cd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1568 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(783dbc0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4009 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4973270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2908 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8265ba8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2478 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff30e79b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_664 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d96da7a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3214 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b12679e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5090d7c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1310 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(700a9526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a9813)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3049 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fdb2d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3455 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c18265a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2239 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff37e457)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_852 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7896441)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2846 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb4c431d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2735 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eccb102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2457 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f20cea9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_351 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d400cd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f95d221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3051 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f06d6ae7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccdb5835)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_437 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e317badd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3149 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f50426b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3196 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c0a1cb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2164 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62b65de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_681 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a2dde8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3182 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b6dffe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3567 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43543936)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2993 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e21cdc8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1828 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32aa7dde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2542 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e957811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3942 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c81bff3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_412 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3058d08a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2789 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85ef7e14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3686 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de3e713)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fa1421f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2759 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6b42d1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_784 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aad53b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4059 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf3b17de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d297f51b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1673 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2f90338)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2241 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40f1277a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3570 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8412a58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2949 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf543040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1544 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(940f65b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb8c72ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3066 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eac610b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1252 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24cdf61e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1981 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41ac24e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1560 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3583 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19337ec2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2697 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10f85909)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2348 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf74ac84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2384 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc60ebc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_967 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bceaa14e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1349 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(391f3e68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_825 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2be53637)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db72aad9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3561 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1682 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeed783b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2286 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f04a75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3103 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa03d1d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66f8e326)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1422 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df7a90fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3479 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dc0cfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d221e9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3175 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83e8647c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2350 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25265e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1385 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b473b335)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2518 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd1085a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2282 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2a3aaa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1153 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d027f1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b2499c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3170 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ce038)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3747 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76f05785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2722 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4614af31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(998707cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2834 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d54fe638)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2250 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24911d93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_807 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc7fa1a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3683 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a032e1c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da0759dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2821 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de017651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3935 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed0f8d09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_955 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd284f03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3024 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87fef7f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_805 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e41c0318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2727 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d77afd83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2186 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9a5a739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_954 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a42f480)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1311 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(358b158a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2263 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15a8d24f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2530 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2419 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c872bcf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2690 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85782dfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1616 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d0ebc8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1464 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ca4e3dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_913 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0543965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3089 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27c58e23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1386 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f83e7df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1446 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64fe5d92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3969 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d27c2d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1770 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3624 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3361d7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1269 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c17fba45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3863 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a50b1142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_624 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdcd1f12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3694 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef48b175)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2058 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4de705a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1860 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54d4274a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2744 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2ef95d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2127 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59943b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2332 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fb4b6a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2761 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c937c358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_856 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bcb268e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2988 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe403e2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2097 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc64ac5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_493 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1d246a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_798 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928f2509)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3905 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc50729c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2725 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1401fdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1188 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b53f4529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3403 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc49bb18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aec9186f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1593 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e79cfc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2471 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(104d4258)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1091 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a99eca22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1495 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8edda769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3626 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9b866a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2936 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffa63a44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3834 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4f7ff6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1215 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bada7aea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1978 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99434e54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2439 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ccc497d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1679 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee506067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3732 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5975ba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3033 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc8d89b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_408 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ff5adb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3189 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3851381d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1665 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e407d98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1152 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3bee3d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3706 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8201365)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3548 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c153ce79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(262ebd17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_787 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8780004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3477 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2980 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0ea081a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2772 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728b485)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1391 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(848fb226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_616 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd1de8ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1038 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5cff14e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_642 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(858bfe16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3501 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4037 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(388561b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1998 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f455322f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2049) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1331 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a27fe0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1668 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaec2fa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3354 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a261c5fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3607 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d2b4fcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2385 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca44934f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_918 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdd1a4fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_602 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27fdc6d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2238 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86db1e31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_391 & _EVAL_2873) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9682988)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
