//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_45_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [5:0]  _EVAL_3,
  input         _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [5:0]  _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_32;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_63;
  reg [31:0] _RAND_1;
  reg  _EVAL_64;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_71;
  reg [31:0] _RAND_3;
  reg [5:0] _EVAL_87;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_107;
  reg [31:0] _RAND_5;
  reg [5:0] _EVAL_110;
  reg [31:0] _RAND_6;
  reg [5:0] _EVAL_117;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_119;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_156;
  reg [31:0] _RAND_9;
  reg [32:0] _EVAL_168;
  reg [63:0] _RAND_10;
  reg [31:0] _EVAL_189;
  reg [31:0] _RAND_11;
  reg [5:0] _EVAL_198;
  reg [31:0] _RAND_12;
  reg  _EVAL_200;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_222;
  reg [31:0] _RAND_14;
  reg [5:0] _EVAL_247;
  reg [31:0] _RAND_15;
  reg [31:0] _EVAL_332;
  reg [31:0] _RAND_16;
  wire [2:0] _EVAL_39;
  wire  _EVAL_165;
  wire  _EVAL_164;
  wire  _EVAL_329;
  wire  _EVAL_158;
  wire [63:0] _EVAL_277;
  wire [63:0] _EVAL_173;
  wire [32:0] _EVAL_275;
  wire  _EVAL_344;
  wire  _EVAL_350;
  wire  _EVAL_316;
  wire  _EVAL_338;
  wire [31:0] _EVAL_31;
  wire [32:0] _EVAL_325;
  wire [32:0] _EVAL_103;
  wire [32:0] _EVAL_111;
  wire  _EVAL_278;
  wire  _EVAL_90;
  wire  _EVAL_267;
  wire [1:0] _EVAL_336;
  wire [1:0] _EVAL_206;
  wire  _EVAL_109;
  wire  _EVAL_88;
  wire  _EVAL_288;
  wire  _EVAL_327;
  wire  _EVAL_282;
  wire  _EVAL_363;
  wire  _EVAL_41;
  wire  _EVAL_78;
  wire  _EVAL_105;
  wire  _EVAL_65;
  wire  _EVAL_343;
  wire  _EVAL_331;
  wire  _EVAL_86;
  wire  _EVAL_40;
  wire [63:0] _EVAL_43;
  wire [63:0] _EVAL_213;
  wire [32:0] _EVAL_135;
  wire  _EVAL_259;
  wire  _EVAL_181;
  wire  _EVAL_280;
  wire  _EVAL_192;
  wire  _EVAL_172;
  wire  _EVAL_208;
  wire  _EVAL_294;
  wire  _EVAL_320;
  wire  _EVAL_52;
  wire  _EVAL_299;
  wire  _EVAL_93;
  wire  _EVAL_187;
  wire [32:0] _EVAL_59;
  wire  _EVAL_306;
  wire  _EVAL_229;
  wire  _EVAL_340;
  wire [32:0] _EVAL_159;
  wire [32:0] _EVAL_263;
  wire  _EVAL_139;
  wire  _EVAL_335;
  wire  _EVAL_46;
  wire [22:0] _EVAL_254;
  wire [7:0] _EVAL_230;
  wire  _EVAL_197;
  wire  _EVAL_23;
  wire  _EVAL_334;
  wire [31:0] _EVAL_261;
  wire [32:0] _EVAL_76;
  wire [32:0] _EVAL_279;
  wire [32:0] _EVAL_204;
  wire  _EVAL_104;
  wire  _EVAL_297;
  wire [31:0] _EVAL_203;
  wire [32:0] _EVAL_323;
  wire [32:0] _EVAL_157;
  wire [32:0] _EVAL_195;
  wire  _EVAL_364;
  wire [31:0] _EVAL_154;
  wire [32:0] _EVAL_322;
  wire [32:0] _EVAL_113;
  wire [32:0] _EVAL_112;
  wire  _EVAL_352;
  wire  _EVAL_270;
  wire  _EVAL_303;
  wire  _EVAL_186;
  wire  _EVAL_274;
  wire [31:0] _EVAL_174;
  wire [32:0] _EVAL_360;
  wire [32:0] _EVAL_35;
  wire [32:0] _EVAL_337;
  wire  _EVAL_155;
  wire  _EVAL_356;
  wire [31:0] _EVAL_310;
  wire [32:0] _EVAL_199;
  wire [32:0] _EVAL_142;
  wire [32:0] _EVAL_50;
  wire  _EVAL_44;
  wire  _EVAL_162;
  wire [32:0] _EVAL_219;
  wire [32:0] _EVAL_19;
  wire [32:0] _EVAL_137;
  wire  _EVAL_296;
  wire  _EVAL_144;
  wire  _EVAL_286;
  wire  _EVAL_99;
  wire  _EVAL_290;
  wire [22:0] _EVAL_268;
  wire [7:0] _EVAL_27;
  wire [7:0] _EVAL_193;
  wire  _EVAL_30;
  wire  _EVAL_167;
  wire  _EVAL_121;
  wire  _EVAL_211;
  wire  _EVAL_51;
  wire  _EVAL_345;
  wire [32:0] _EVAL_70;
  wire  _EVAL_180;
  wire  _EVAL_114;
  wire  _EVAL_77;
  wire [31:0] _EVAL_169;
  wire [32:0] _EVAL_289;
  wire  _EVAL_207;
  wire  _EVAL_161;
  wire  _EVAL_69;
  wire  _EVAL_228;
  wire  _EVAL_217;
  wire  _EVAL_129;
  wire  _EVAL_145;
  wire  _EVAL_353;
  wire  _EVAL_341;
  wire  _EVAL_238;
  wire  _EVAL_115;
  wire  _EVAL_262;
  wire  _EVAL_55;
  wire  _EVAL_300;
  wire [3:0] _EVAL_150;
  wire [3:0] _EVAL_215;
  wire [3:0] _EVAL_358;
  wire  _EVAL_20;
  wire  _EVAL_266;
  wire [7:0] _EVAL_194;
  wire [5:0] _EVAL_36;
  wire [5:0] _EVAL_237;
  wire [32:0] _EVAL_54;
  wire  _EVAL_118;
  wire  _EVAL_362;
  wire [31:0] _EVAL_185;
  wire [31:0] _EVAL_342;
  wire  _EVAL_245;
  wire  _EVAL_183;
  wire  _EVAL_61;
  wire  _EVAL_234;
  wire [2:0] _EVAL_196;
  wire  _EVAL_349;
  wire  _EVAL_317;
  wire  _EVAL_212;
  wire  _EVAL_170;
  wire  _EVAL_205;
  wire  _EVAL_138;
  wire  _EVAL_128;
  wire  _EVAL_239;
  wire  _EVAL_82;
  wire  _EVAL_253;
  wire  _EVAL_256;
  wire  _EVAL_255;
  wire  _EVAL_214;
  wire  _EVAL_178;
  wire  _EVAL_81;
  wire  _EVAL_101;
  wire  _EVAL_226;
  wire [31:0] _EVAL_120;
  wire [32:0] _EVAL_359;
  wire [32:0] _EVAL_123;
  wire [32:0] _EVAL_85;
  wire  _EVAL_285;
  wire  _EVAL_328;
  wire [32:0] _EVAL_130;
  wire  _EVAL_309;
  wire  _EVAL_302;
  wire  _EVAL_287;
  wire  _EVAL_339;
  wire  _EVAL_141;
  wire  _EVAL_311;
  wire [5:0] _EVAL_315;
  wire  _EVAL_66;
  wire  _EVAL_84;
  wire  _EVAL_240;
  wire [32:0] _EVAL_89;
  wire [32:0] _EVAL_361;
  wire [5:0] _EVAL_301;
  wire  _EVAL_218;
  wire  _EVAL_60;
  wire  _EVAL_241;
  wire  _EVAL_62;
  wire  _EVAL_106;
  wire  _EVAL_223;
  wire  _EVAL_74;
  wire  _EVAL_131;
  wire  _EVAL_73;
  wire  _EVAL_49;
  wire  _EVAL_79;
  wire  _EVAL_126;
  wire  _EVAL_134;
  wire  _EVAL_324;
  wire  _EVAL_67;
  wire  _EVAL_221;
  wire  _EVAL_25;
  wire  _EVAL_281;
  wire  _EVAL_97;
  wire  _EVAL_184;
  wire  _EVAL_140;
  wire  _EVAL_246;
  wire  _EVAL_100;
  wire  _EVAL_136;
  wire  _EVAL_313;
  wire [5:0] _EVAL_108;
  wire [5:0] _EVAL_271;
  wire [31:0] _EVAL_244;
  wire  _EVAL_95;
  wire  _EVAL_94;
  wire  _EVAL_102;
  wire  _EVAL_153;
  wire  _EVAL_116;
  wire  _EVAL_347;
  wire  _EVAL_351;
  wire  _EVAL_250;
  wire  _EVAL_326;
  wire  _EVAL_151;
  wire  _EVAL_235;
  wire  _EVAL_125;
  wire  _EVAL_312;
  wire  _EVAL_321;
  wire  _EVAL_163;
  wire  _EVAL_57;
  wire  _EVAL_355;
  wire  _EVAL_53;
  wire  _EVAL_148;
  wire  _EVAL_233;
  wire  _EVAL_92;
  wire  _EVAL_298;
  wire  _EVAL_231;
  wire  _EVAL_291;
  wire  _EVAL_22;
  wire  _EVAL_48;
  wire  _EVAL_330;
  wire  _EVAL_248;
  wire  _EVAL_179;
  wire  _EVAL_143;
  wire  _EVAL_146;
  wire  _EVAL_242;
  wire  _EVAL_293;
  wire  _EVAL_80;
  wire  _EVAL_34;
  wire  _EVAL_133;
  wire  _EVAL_160;
  wire  _EVAL_251;
  wire  _EVAL_292;
  wire  _EVAL_171;
  wire  _EVAL_249;
  wire  _EVAL_216;
  wire  _EVAL_124;
  wire  _EVAL_45;
  wire  _EVAL_269;
  wire [3:0] _EVAL_284;
  wire  _EVAL_236;
  wire  _EVAL_191;
  wire  _EVAL_225;
  wire  _EVAL_175;
  wire  _EVAL_264;
  wire  _EVAL_176;
  wire  _EVAL_210;
  wire  _EVAL_202;
  wire  _EVAL_232;
  wire  _EVAL_21;
  wire  _EVAL_68;
  wire  _EVAL_56;
  wire  _EVAL_83;
  wire  _EVAL_272;
  wire  _EVAL_209;
  wire  _EVAL_122;
  wire  _EVAL_26;
  wire  _EVAL_58;
  wire  _EVAL_29;
  wire  _EVAL_305;
  wire  _EVAL_333;
  wire  _EVAL_265;
  wire  _EVAL_38;
  wire  _EVAL_354;
  wire  _EVAL_258;
  wire  _EVAL_24;
  wire  _EVAL_28;
  wire  _EVAL_98;
  wire  _EVAL_224;
  wire  _EVAL_33;
  wire  _EVAL_47;
  wire  _EVAL_257;
  wire  _EVAL_72;
  wire  _EVAL_273;
  wire  _EVAL_304;
  wire  _EVAL_188;
  wire  _EVAL_308;
  wire  _EVAL_295;
  wire  _EVAL_252;
  wire  _EVAL_91;
  wire  _EVAL_346;
  wire  _EVAL_42;
  wire  _EVAL_96;
  wire  _EVAL_319;
  wire  _EVAL_227;
  wire  _EVAL_182;
  wire  _EVAL_127;
  wire  _EVAL_283;
  wire  _EVAL_75;
  wire  _EVAL_147;
  wire  _EVAL_152;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_39 = _EVAL_6[5:3];
  assign _EVAL_165 = _EVAL_12 == _EVAL_71;
  assign _EVAL_164 = _EVAL_13 & _EVAL_10;
  assign _EVAL_329 = _EVAL_156 == 6'h0;
  assign _EVAL_158 = _EVAL_164 & _EVAL_329;
  assign _EVAL_277 = 64'h1 << _EVAL_6;
  assign _EVAL_173 = _EVAL_158 ? _EVAL_277 : 64'h0;
  assign _EVAL_275 = _EVAL_173[32:0];
  assign _EVAL_344 = _EVAL_16 == _EVAL_222;
  assign _EVAL_350 = _EVAL_344 | _EVAL_4;
  assign _EVAL_316 = _EVAL_350 == 1'h0;
  assign _EVAL_338 = _EVAL_2 == _EVAL_200;
  assign _EVAL_31 = _EVAL_14 ^ 32'h1800000;
  assign _EVAL_325 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_103 = $signed(_EVAL_325) & $signed(-33'sh8000);
  assign _EVAL_111 = $signed(_EVAL_103);
  assign _EVAL_278 = $signed(_EVAL_111) == $signed(33'sh0);
  assign _EVAL_90 = _EVAL_332 < plusarg_reader_out;
  assign _EVAL_267 = _EVAL_18[0];
  assign _EVAL_336 = 2'h1 << _EVAL_267;
  assign _EVAL_206 = _EVAL_336 | 2'h1;
  assign _EVAL_109 = _EVAL_206[0];
  assign _EVAL_88 = _EVAL_14[1];
  assign _EVAL_288 = _EVAL_14[0];
  assign _EVAL_327 = _EVAL_88 & _EVAL_288;
  assign _EVAL_282 = _EVAL_109 & _EVAL_327;
  assign _EVAL_363 = _EVAL <= 3'h3;
  assign _EVAL_41 = _EVAL_363 | _EVAL_4;
  assign _EVAL_78 = _EVAL_41 == 1'h0;
  assign _EVAL_105 = _EVAL_15 & _EVAL_17;
  assign _EVAL_65 = _EVAL_117 == 6'h0;
  assign _EVAL_343 = _EVAL_105 & _EVAL_65;
  assign _EVAL_331 = _EVAL_1 == 3'h6;
  assign _EVAL_86 = _EVAL_331 == 1'h0;
  assign _EVAL_40 = _EVAL_343 & _EVAL_86;
  assign _EVAL_43 = 64'h1 << _EVAL_3;
  assign _EVAL_213 = _EVAL_40 ? _EVAL_43 : 64'h0;
  assign _EVAL_135 = _EVAL_213[32:0];
  assign _EVAL_259 = _EVAL_275 != _EVAL_135;
  assign _EVAL_181 = _EVAL_275 != 33'h0;
  assign _EVAL_280 = _EVAL_181 == 1'h0;
  assign _EVAL_192 = _EVAL_259 | _EVAL_280;
  assign _EVAL_172 = _EVAL == 3'h0;
  assign _EVAL_208 = _EVAL_8[2];
  assign _EVAL_294 = _EVAL_208 == 1'h0;
  assign _EVAL_320 = _EVAL_3 == 6'h20;
  assign _EVAL_52 = _EVAL_39 == 3'h1;
  assign _EVAL_299 = _EVAL_12 == 2'h0;
  assign _EVAL_93 = _EVAL_299 | _EVAL_4;
  assign _EVAL_187 = _EVAL_93 == 1'h0;
  assign _EVAL_59 = _EVAL_168 >> _EVAL_6;
  assign _EVAL_306 = _EVAL_59[0];
  assign _EVAL_229 = _EVAL_306 == 1'h0;
  assign _EVAL_340 = _EVAL_229 | _EVAL_4;
  assign _EVAL_159 = _EVAL_275 | _EVAL_168;
  assign _EVAL_263 = _EVAL_159 >> _EVAL_3;
  assign _EVAL_139 = _EVAL_1 == 3'h2;
  assign _EVAL_335 = _EVAL_17 & _EVAL_139;
  assign _EVAL_46 = _EVAL_8 == 3'h3;
  assign _EVAL_254 = 23'hff << _EVAL_16;
  assign _EVAL_230 = _EVAL_254[7:0];
  assign _EVAL_197 = _EVAL_1 == 3'h4;
  assign _EVAL_23 = _EVAL_17 & _EVAL_197;
  assign _EVAL_334 = _EVAL_18 <= 4'h8;
  assign _EVAL_261 = _EVAL_14 ^ 32'h3000;
  assign _EVAL_76 = {1'b0,$signed(_EVAL_261)};
  assign _EVAL_279 = $signed(_EVAL_76) & $signed(-33'sh1000);
  assign _EVAL_204 = $signed(_EVAL_279);
  assign _EVAL_104 = $signed(_EVAL_204) == $signed(33'sh0);
  assign _EVAL_297 = _EVAL_334 & _EVAL_104;
  assign _EVAL_203 = _EVAL_14 ^ 32'h40000000;
  assign _EVAL_323 = {1'b0,$signed(_EVAL_203)};
  assign _EVAL_157 = $signed(_EVAL_323) & $signed(-33'sh2000);
  assign _EVAL_195 = $signed(_EVAL_157);
  assign _EVAL_364 = $signed(_EVAL_195) == $signed(33'sh0);
  assign _EVAL_154 = _EVAL_14 ^ 32'h80000000;
  assign _EVAL_322 = {1'b0,$signed(_EVAL_154)};
  assign _EVAL_113 = $signed(_EVAL_322) & $signed(-33'sh20000);
  assign _EVAL_112 = $signed(_EVAL_113);
  assign _EVAL_352 = $signed(_EVAL_112) == $signed(33'sh0);
  assign _EVAL_270 = _EVAL_364 | _EVAL_352;
  assign _EVAL_303 = _EVAL_8 == 3'h6;
  assign _EVAL_186 = _EVAL_18 <= 4'h6;
  assign _EVAL_274 = _EVAL_186 & _EVAL_352;
  assign _EVAL_174 = _EVAL_14 ^ 32'hc000000;
  assign _EVAL_360 = {1'b0,$signed(_EVAL_174)};
  assign _EVAL_35 = $signed(_EVAL_360) & $signed(-33'sh4000000);
  assign _EVAL_337 = $signed(_EVAL_35);
  assign _EVAL_155 = $signed(_EVAL_337) == $signed(33'sh0);
  assign _EVAL_356 = _EVAL_104 | _EVAL_155;
  assign _EVAL_310 = _EVAL_14 ^ 32'h2000000;
  assign _EVAL_199 = {1'b0,$signed(_EVAL_310)};
  assign _EVAL_142 = $signed(_EVAL_199) & $signed(-33'sh10000);
  assign _EVAL_50 = $signed(_EVAL_142);
  assign _EVAL_44 = $signed(_EVAL_50) == $signed(33'sh0);
  assign _EVAL_162 = _EVAL_356 | _EVAL_44;
  assign _EVAL_219 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_19 = $signed(_EVAL_219) & $signed(-33'sh5000);
  assign _EVAL_137 = $signed(_EVAL_19);
  assign _EVAL_296 = $signed(_EVAL_137) == $signed(33'sh0);
  assign _EVAL_144 = _EVAL_88 == 1'h0;
  assign _EVAL_286 = _EVAL_288 == 1'h0;
  assign _EVAL_99 = _EVAL_144 & _EVAL_286;
  assign _EVAL_290 = _EVAL_109 & _EVAL_99;
  assign _EVAL_268 = 23'hff << _EVAL_18;
  assign _EVAL_27 = _EVAL_268[7:0];
  assign _EVAL_193 = ~ _EVAL_27;
  assign _EVAL_30 = _EVAL_8 == _EVAL_63;
  assign _EVAL_167 = _EVAL_30 | _EVAL_4;
  assign _EVAL_121 = _EVAL_167 == 1'h0;
  assign _EVAL_211 = _EVAL_172 | _EVAL_4;
  assign _EVAL_51 = _EVAL_3 == _EVAL_247;
  assign _EVAL_345 = _EVAL_51 | _EVAL_4;
  assign _EVAL_70 = _EVAL_168 | _EVAL_275;
  assign _EVAL_180 = _EVAL_16 >= 4'h2;
  assign _EVAL_114 = _EVAL_180 | _EVAL_4;
  assign _EVAL_77 = _EVAL_198 == 6'h0;
  assign _EVAL_169 = _EVAL_14 ^ 32'h20000000;
  assign _EVAL_289 = {1'b0,$signed(_EVAL_169)};
  assign _EVAL_207 = _EVAL_18 >= 4'h2;
  assign _EVAL_161 = _EVAL_206[1];
  assign _EVAL_69 = _EVAL_161 & _EVAL_88;
  assign _EVAL_228 = _EVAL_207 | _EVAL_69;
  assign _EVAL_217 = _EVAL_228 | _EVAL_282;
  assign _EVAL_129 = _EVAL_88 & _EVAL_286;
  assign _EVAL_145 = _EVAL_109 & _EVAL_129;
  assign _EVAL_353 = _EVAL_228 | _EVAL_145;
  assign _EVAL_341 = _EVAL_161 & _EVAL_144;
  assign _EVAL_238 = _EVAL_207 | _EVAL_341;
  assign _EVAL_115 = _EVAL_144 & _EVAL_288;
  assign _EVAL_262 = _EVAL_109 & _EVAL_115;
  assign _EVAL_55 = _EVAL_238 | _EVAL_262;
  assign _EVAL_300 = _EVAL_238 | _EVAL_290;
  assign _EVAL_150 = {_EVAL_217,_EVAL_353,_EVAL_55,_EVAL_300};
  assign _EVAL_215 = ~ _EVAL_150;
  assign _EVAL_358 = _EVAL_5 & _EVAL_215;
  assign _EVAL_20 = _EVAL_358 == 4'h0;
  assign _EVAL_266 = _EVAL_1[0];
  assign _EVAL_194 = ~ _EVAL_230;
  assign _EVAL_36 = _EVAL_194[7:2];
  assign _EVAL_237 = _EVAL_117 - 6'h1;
  assign _EVAL_54 = $signed(_EVAL_289) & $signed(-33'sh2000);
  assign _EVAL_118 = _EVAL_5 == _EVAL_150;
  assign _EVAL_362 = _EVAL <= 3'h4;
  assign _EVAL_185 = {{24'd0}, _EVAL_193};
  assign _EVAL_342 = _EVAL_14 & _EVAL_185;
  assign _EVAL_245 = _EVAL_342 == 32'h0;
  assign _EVAL_183 = _EVAL_245 | _EVAL_4;
  assign _EVAL_61 = _EVAL_183 == 1'h0;
  assign _EVAL_234 = _EVAL_87 == 6'h0;
  assign _EVAL_196 = _EVAL_3[5:3];
  assign _EVAL_349 = _EVAL_8 == 3'h7;
  assign _EVAL_317 = _EVAL_10 & _EVAL_349;
  assign _EVAL_212 = _EVAL_234 == 1'h0;
  assign _EVAL_170 = _EVAL_18 <= 4'h2;
  assign _EVAL_205 = _EVAL_168 != 33'h0;
  assign _EVAL_138 = _EVAL_6 == 6'h20;
  assign _EVAL_128 = _EVAL_39 == 3'h0;
  assign _EVAL_239 = _EVAL_138 | _EVAL_128;
  assign _EVAL_82 = _EVAL_239 | _EVAL_52;
  assign _EVAL_253 = _EVAL_39 == 3'h2;
  assign _EVAL_256 = _EVAL_82 | _EVAL_253;
  assign _EVAL_255 = _EVAL_39 == 3'h3;
  assign _EVAL_214 = _EVAL_256 | _EVAL_255;
  assign _EVAL_178 = _EVAL_214 | _EVAL_4;
  assign _EVAL_81 = _EVAL_178 == 1'h0;
  assign _EVAL_101 = _EVAL_162 | _EVAL_296;
  assign _EVAL_226 = _EVAL_101 | _EVAL_278;
  assign _EVAL_120 = _EVAL_14 ^ 32'h1900000;
  assign _EVAL_359 = {1'b0,$signed(_EVAL_120)};
  assign _EVAL_123 = $signed(_EVAL_359) & $signed(-33'sh2000);
  assign _EVAL_85 = $signed(_EVAL_123);
  assign _EVAL_285 = $signed(_EVAL_85) == $signed(33'sh0);
  assign _EVAL_328 = _EVAL_226 | _EVAL_285;
  assign _EVAL_130 = $signed(_EVAL_54);
  assign _EVAL_309 = $signed(_EVAL_130) == $signed(33'sh0);
  assign _EVAL_302 = _EVAL_328 | _EVAL_309;
  assign _EVAL_287 = _EVAL_170 & _EVAL_302;
  assign _EVAL_339 = _EVAL_287 | _EVAL_4;
  assign _EVAL_141 = _EVAL_339 == 1'h0;
  assign _EVAL_311 = _EVAL_1 == 3'h0;
  assign _EVAL_315 = _EVAL_87 - 6'h1;
  assign _EVAL_66 = _EVAL_4 == 1'h0;
  assign _EVAL_84 = _EVAL_192 | _EVAL_4;
  assign _EVAL_240 = _EVAL_84 == 1'h0;
  assign _EVAL_89 = ~ _EVAL_135;
  assign _EVAL_361 = _EVAL_70 & _EVAL_89;
  assign _EVAL_301 = _EVAL_198 - 6'h1;
  assign _EVAL_218 = _EVAL_2 == 1'h0;
  assign _EVAL_60 = _EVAL_218 | _EVAL_4;
  assign _EVAL_241 = _EVAL_60 == 1'h0;
  assign _EVAL_62 = _EVAL_8 == 3'h5;
  assign _EVAL_106 = _EVAL_18 == _EVAL_32;
  assign _EVAL_223 = _EVAL_7 == 1'h0;
  assign _EVAL_74 = _EVAL_223 | _EVAL_4;
  assign _EVAL_131 = _EVAL_9 == _EVAL_64;
  assign _EVAL_73 = _EVAL_297 | _EVAL_4;
  assign _EVAL_49 = _EVAL_73 == 1'h0;
  assign _EVAL_79 = _EVAL_218 | _EVAL_7;
  assign _EVAL_126 = _EVAL_79 | _EVAL_4;
  assign _EVAL_134 = _EVAL_126 == 1'h0;
  assign _EVAL_324 = _EVAL_205 == 1'h0;
  assign _EVAL_67 = plusarg_reader_out == 32'h0;
  assign _EVAL_221 = _EVAL_324 | _EVAL_67;
  assign _EVAL_25 = _EVAL_221 | _EVAL_90;
  assign _EVAL_281 = _EVAL_25 | _EVAL_4;
  assign _EVAL_97 = _EVAL_196 == 3'h0;
  assign _EVAL_184 = _EVAL_320 | _EVAL_97;
  assign _EVAL_140 = _EVAL_207 | _EVAL_4;
  assign _EVAL_246 = _EVAL_140 == 1'h0;
  assign _EVAL_100 = _EVAL_1 == 3'h1;
  assign _EVAL_136 = _EVAL_263[0];
  assign _EVAL_313 = _EVAL_136 | _EVAL_4;
  assign _EVAL_108 = _EVAL_193[7:2];
  assign _EVAL_271 = _EVAL_156 - 6'h1;
  assign _EVAL_244 = _EVAL_332 + 32'h1;
  assign _EVAL_95 = _EVAL_270 | _EVAL_155;
  assign _EVAL_94 = _EVAL_95 | _EVAL_44;
  assign _EVAL_102 = _EVAL_94 | _EVAL_296;
  assign _EVAL_153 = _EVAL != 3'h0;
  assign _EVAL_116 = _EVAL_196 == 3'h2;
  assign _EVAL_347 = _EVAL_164 | _EVAL_105;
  assign _EVAL_351 = _EVAL_106 | _EVAL_4;
  assign _EVAL_250 = _EVAL_351 == 1'h0;
  assign _EVAL_326 = _EVAL_165 | _EVAL_4;
  assign _EVAL_151 = _EVAL_326 == 1'h0;
  assign _EVAL_235 = _EVAL_12 != 2'h2;
  assign _EVAL_125 = _EVAL_17 & _EVAL_212;
  assign _EVAL_312 = _EVAL_235 | _EVAL_4;
  assign _EVAL_321 = _EVAL_312 == 1'h0;
  assign _EVAL_163 = _EVAL_102 | _EVAL_278;
  assign _EVAL_57 = _EVAL_163 | _EVAL_285;
  assign _EVAL_355 = _EVAL_57 | _EVAL_309;
  assign _EVAL_53 = _EVAL_186 & _EVAL_355;
  assign _EVAL_148 = _EVAL_53 | _EVAL_297;
  assign _EVAL_233 = _EVAL <= 3'h2;
  assign _EVAL_92 = _EVAL_17 & _EVAL_311;
  assign _EVAL_298 = _EVAL_281 == 1'h0;
  assign _EVAL_231 = _EVAL_8 == 3'h1;
  assign _EVAL_291 = _EVAL_211 == 1'h0;
  assign _EVAL_22 = _EVAL_12 <= 2'h2;
  assign _EVAL_48 = _EVAL_22 | _EVAL_4;
  assign _EVAL_330 = _EVAL_48 == 1'h0;
  assign _EVAL_248 = _EVAL_196 == 3'h1;
  assign _EVAL_179 = _EVAL_184 | _EVAL_248;
  assign _EVAL_143 = _EVAL_179 | _EVAL_116;
  assign _EVAL_146 = _EVAL_196 == 3'h3;
  assign _EVAL_242 = _EVAL_143 | _EVAL_146;
  assign _EVAL_293 = _EVAL_1 <= 3'h6;
  assign _EVAL_80 = _EVAL_6 == _EVAL_110;
  assign _EVAL_34 = _EVAL_77 == 1'h0;
  assign _EVAL_133 = _EVAL_10 & _EVAL_34;
  assign _EVAL_160 = _EVAL_362 | _EVAL_4;
  assign _EVAL_251 = _EVAL_160 == 1'h0;
  assign _EVAL_292 = _EVAL_8 == 3'h0;
  assign _EVAL_171 = _EVAL_10 & _EVAL_292;
  assign _EVAL_249 = _EVAL_0 == 1'h0;
  assign _EVAL_216 = _EVAL_249 | _EVAL_4;
  assign _EVAL_124 = _EVAL_118 | _EVAL_4;
  assign _EVAL_45 = _EVAL_124 == 1'h0;
  assign _EVAL_269 = _EVAL_20 | _EVAL_4;
  assign _EVAL_284 = ~ _EVAL_5;
  assign _EVAL_236 = _EVAL_284 == 4'h0;
  assign _EVAL_191 = _EVAL_236 | _EVAL_4;
  assign _EVAL_225 = _EVAL_293 | _EVAL_4;
  assign _EVAL_175 = _EVAL_225 == 1'h0;
  assign _EVAL_264 = _EVAL_8 == 3'h2;
  assign _EVAL_176 = _EVAL_10 & _EVAL_264;
  assign _EVAL_210 = _EVAL_14 == _EVAL_189;
  assign _EVAL_202 = _EVAL_210 | _EVAL_4;
  assign _EVAL_232 = _EVAL_202 == 1'h0;
  assign _EVAL_21 = _EVAL == _EVAL_119;
  assign _EVAL_68 = _EVAL_21 | _EVAL_4;
  assign _EVAL_56 = _EVAL_68 == 1'h0;
  assign _EVAL_83 = _EVAL_338 | _EVAL_4;
  assign _EVAL_272 = _EVAL_83 == 1'h0;
  assign _EVAL_209 = _EVAL_313 == 1'h0;
  assign _EVAL_122 = _EVAL_105 & _EVAL_234;
  assign _EVAL_26 = _EVAL_233 | _EVAL_4;
  assign _EVAL_58 = _EVAL_26 == 1'h0;
  assign _EVAL_29 = _EVAL_17 & _EVAL_331;
  assign _EVAL_305 = _EVAL_274 | _EVAL_4;
  assign _EVAL_333 = _EVAL_8 == 3'h4;
  assign _EVAL_265 = _EVAL_10 & _EVAL_333;
  assign _EVAL_38 = _EVAL_148 | _EVAL_4;
  assign _EVAL_354 = _EVAL_305 == 1'h0;
  assign _EVAL_258 = _EVAL_1 == _EVAL_107;
  assign _EVAL_24 = _EVAL_258 | _EVAL_4;
  assign _EVAL_28 = _EVAL_24 == 1'h0;
  assign _EVAL_98 = _EVAL_10 & _EVAL_303;
  assign _EVAL_224 = _EVAL_80 | _EVAL_4;
  assign _EVAL_33 = _EVAL_224 == 1'h0;
  assign _EVAL_47 = _EVAL_131 | _EVAL_4;
  assign _EVAL_257 = _EVAL_47 == 1'h0;
  assign _EVAL_72 = _EVAL_74 == 1'h0;
  assign _EVAL_273 = _EVAL_38 == 1'h0;
  assign _EVAL_304 = _EVAL_340 == 1'h0;
  assign _EVAL_188 = _EVAL_345 == 1'h0;
  assign _EVAL_308 = _EVAL_1 == 3'h5;
  assign _EVAL_295 = _EVAL_17 & _EVAL_308;
  assign _EVAL_252 = _EVAL_242 | _EVAL_4;
  assign _EVAL_91 = _EVAL_153 | _EVAL_4;
  assign _EVAL_346 = _EVAL_91 == 1'h0;
  assign _EVAL_42 = _EVAL_252 == 1'h0;
  assign _EVAL_96 = _EVAL_10 & _EVAL_46;
  assign _EVAL_319 = _EVAL_10 & _EVAL_231;
  assign _EVAL_227 = _EVAL_164 & _EVAL_77;
  assign _EVAL_182 = _EVAL_17 & _EVAL_100;
  assign _EVAL_127 = _EVAL_114 == 1'h0;
  assign _EVAL_283 = _EVAL_269 == 1'h0;
  assign _EVAL_75 = _EVAL_216 == 1'h0;
  assign _EVAL_147 = _EVAL_10 & _EVAL_62;
  assign _EVAL_152 = _EVAL_191 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_63 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_71 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_87 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_107 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_110 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_117 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_119 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_156 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _EVAL_168 = _RAND_10[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_189 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_198 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_200 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_222 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_247 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_332 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_11) begin
    if (_EVAL_227) begin
      _EVAL_32 <= _EVAL_18;
    end
    if (_EVAL_227) begin
      _EVAL_63 <= _EVAL_8;
    end
    if (_EVAL_122) begin
      _EVAL_64 <= _EVAL_9;
    end
    if (_EVAL_122) begin
      _EVAL_71 <= _EVAL_12;
    end
    if (_EVAL_4) begin
      _EVAL_87 <= 6'h0;
    end else begin
      if (_EVAL_105) begin
        if (_EVAL_234) begin
          if (_EVAL_266) begin
            _EVAL_87 <= _EVAL_36;
          end else begin
            _EVAL_87 <= 6'h0;
          end
        end else begin
          _EVAL_87 <= _EVAL_315;
        end
      end
    end
    if (_EVAL_122) begin
      _EVAL_107 <= _EVAL_1;
    end
    if (_EVAL_227) begin
      _EVAL_110 <= _EVAL_6;
    end
    if (_EVAL_4) begin
      _EVAL_117 <= 6'h0;
    end else begin
      if (_EVAL_105) begin
        if (_EVAL_65) begin
          if (_EVAL_266) begin
            _EVAL_117 <= _EVAL_36;
          end else begin
            _EVAL_117 <= 6'h0;
          end
        end else begin
          _EVAL_117 <= _EVAL_237;
        end
      end
    end
    if (_EVAL_227) begin
      _EVAL_119 <= _EVAL;
    end
    if (_EVAL_4) begin
      _EVAL_156 <= 6'h0;
    end else begin
      if (_EVAL_164) begin
        if (_EVAL_329) begin
          if (_EVAL_294) begin
            _EVAL_156 <= _EVAL_108;
          end else begin
            _EVAL_156 <= 6'h0;
          end
        end else begin
          _EVAL_156 <= _EVAL_271;
        end
      end
    end
    if (_EVAL_4) begin
      _EVAL_168 <= 33'h0;
    end else begin
      _EVAL_168 <= _EVAL_361;
    end
    if (_EVAL_227) begin
      _EVAL_189 <= _EVAL_14;
    end
    if (_EVAL_4) begin
      _EVAL_198 <= 6'h0;
    end else begin
      if (_EVAL_164) begin
        if (_EVAL_77) begin
          if (_EVAL_294) begin
            _EVAL_198 <= _EVAL_108;
          end else begin
            _EVAL_198 <= 6'h0;
          end
        end else begin
          _EVAL_198 <= _EVAL_301;
        end
      end
    end
    if (_EVAL_122) begin
      _EVAL_200 <= _EVAL_2;
    end
    if (_EVAL_122) begin
      _EVAL_222 <= _EVAL_16;
    end
    if (_EVAL_122) begin
      _EVAL_247 <= _EVAL_3;
    end
    if (_EVAL_4) begin
      _EVAL_332 <= 32'h0;
    end else begin
      if (_EVAL_347) begin
        _EVAL_332 <= 32'h0;
      end else begin
        _EVAL_332 <= _EVAL_244;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74ada32f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c37c27da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ddafa7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ef55a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96141eeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a85c81d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc3bb35d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bd4e5b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dffa9f26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aed79e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37ccef7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aee5314)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8929bfb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96c05be4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(896500ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50d128eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(850b7615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fd9a69d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c66d7360)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cb78638)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(386ccb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bb88fe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a4bc1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3d0b98f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a17b892a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9293334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7855d6ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(556c1488)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4809dbad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef419a2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(433b80ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cfe0101)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903784b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2ce5e37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65f85db6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07600b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9afee218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa142f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(800939f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d949250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8878fc7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8c00f05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47da62f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5d07ae0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53e36b76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(714da2a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5018c17b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa407584)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20a4198c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e4410d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1661818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87d30bd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b89425b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8af3a31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86a7bb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd37fa80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_346) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55712ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_346) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c78862b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(659fc996)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e869a49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bae9399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(572889ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(901579ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a2d9f15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f88f9526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc2e3e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92002278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7f49664)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eba50382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc6a9946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69dd4b2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e0c50f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d393506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d1ae095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f112d54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(200a1ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c7f7c2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76265ae1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81816ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bda47819)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3755c9a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cc582db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d4a2fc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3477427d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(123ed147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b44f040a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f45dbe1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3599ed4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
