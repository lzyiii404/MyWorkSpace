//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_3_assert(
  input  [3:0]  _EVAL,
  input  [31:0] _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input  [7:0]  _EVAL_8,
  input  [1:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  input  [1:0]  _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input  [3:0]  _EVAL_27,
  input  [2:0]  _EVAL_28,
  input         _EVAL_29,
  input  [2:0]  _EVAL_30,
  input  [3:0]  _EVAL_31,
  input         _EVAL_32
);
  wire [31:0] plusarg_reader_out;
  reg [4:0] _EVAL_37;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_168;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_201;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_203;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_235;
  reg [31:0] _RAND_4;
  reg [31:0] _EVAL_278;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_283;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_297;
  reg [31:0] _RAND_7;
  reg [4:0] _EVAL_316;
  reg [31:0] _RAND_8;
  reg [4:0] _EVAL_323;
  reg [31:0] _RAND_9;
  reg  _EVAL_351;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_360;
  reg [31:0] _RAND_11;
  reg [1:0] _EVAL_369;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_406;
  reg [31:0] _RAND_13;
  reg  _EVAL_407;
  reg [31:0] _RAND_14;
  reg [4:0] _EVAL_413;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_435;
  reg [31:0] _RAND_16;
  reg [4:0] _EVAL_442;
  reg [31:0] _RAND_17;
  reg [2:0] _EVAL_463;
  reg [31:0] _RAND_18;
  reg [3:0] _EVAL_464;
  reg [31:0] _RAND_19;
  reg [1:0] _EVAL_470;
  reg [31:0] _RAND_20;
  reg [2:0] _EVAL_474;
  reg [31:0] _RAND_21;
  reg [3:0] _EVAL_518;
  reg [31:0] _RAND_22;
  reg [2:0] _EVAL_557;
  reg [31:0] _RAND_23;
  reg [31:0] _EVAL_587;
  reg [31:0] _RAND_24;
  reg [31:0] _EVAL_605;
  reg [31:0] _RAND_25;
  reg [8:0] _EVAL_607;
  reg [31:0] _RAND_26;
  reg [3:0] _EVAL_628;
  reg [31:0] _RAND_27;
  wire [22:0] _EVAL_277;
  wire [31:0] _EVAL_332;
  wire [32:0] _EVAL_560;
  wire  _EVAL_59;
  wire  _EVAL_103;
  wire  _EVAL_525;
  wire  _EVAL_222;
  wire  _EVAL_329;
  wire  _EVAL_467;
  wire  _EVAL_217;
  wire  _EVAL_231;
  wire  _EVAL_595;
  wire [31:0] _EVAL_99;
  wire [32:0] _EVAL_322;
  wire [7:0] _EVAL_649;
  wire [7:0] _EVAL_394;
  wire [31:0] _EVAL_366;
  wire [31:0] _EVAL_264;
  wire  _EVAL_465;
  wire [31:0] _EVAL_335;
  wire [32:0] _EVAL_571;
  wire [32:0] _EVAL_519;
  wire [32:0] _EVAL_206;
  wire  _EVAL_111;
  wire [31:0] _EVAL_199;
  wire [32:0] _EVAL_656;
  wire [32:0] _EVAL_81;
  wire [32:0] _EVAL_128;
  wire  _EVAL_378;
  wire  _EVAL_270;
  wire [31:0] _EVAL_505;
  wire [32:0] _EVAL_559;
  wire [32:0] _EVAL_399;
  wire [32:0] _EVAL_334;
  wire  _EVAL_526;
  wire  _EVAL_379;
  wire  _EVAL_125;
  wire  _EVAL_487;
  wire  _EVAL_429;
  wire  _EVAL_589;
  wire  _EVAL_196;
  wire [22:0] _EVAL_408;
  wire [7:0] _EVAL_362;
  wire [1:0] _EVAL_263;
  wire [3:0] _EVAL_48;
  wire [2:0] _EVAL_621;
  wire [2:0] _EVAL_552;
  wire  _EVAL_570;
  wire  _EVAL_483;
  wire  _EVAL_363;
  wire  _EVAL_299;
  wire  _EVAL_82;
  wire  _EVAL_172;
  wire  _EVAL_148;
  wire  _EVAL_84;
  wire  _EVAL_476;
  wire  _EVAL_94;
  wire  _EVAL_73;
  wire  _EVAL_181;
  wire  _EVAL_508;
  wire  _EVAL_427;
  wire  _EVAL_305;
  wire  _EVAL_170;
  wire  _EVAL_496;
  wire  _EVAL_356;
  wire  _EVAL_510;
  wire  _EVAL_156;
  wire  _EVAL_255;
  wire [1:0] _EVAL_162;
  wire [1:0] _EVAL_236;
  wire [1:0] _EVAL_38;
  wire [1:0] _EVAL_669;
  wire  _EVAL_313;
  wire  _EVAL_419;
  wire [22:0] _EVAL_665;
  wire [7:0] _EVAL_53;
  wire [7:0] _EVAL_60;
  wire [4:0] _EVAL_578;
  wire [31:0] _EVAL_614;
  wire [32:0] _EVAL_618;
  wire [32:0] _EVAL_490;
  wire [32:0] _EVAL_401;
  wire  _EVAL_566;
  wire [31:0] _EVAL_319;
  wire [32:0] _EVAL_545;
  wire [32:0] _EVAL_136;
  wire [32:0] _EVAL_285;
  wire  _EVAL_232;
  wire  _EVAL_527;
  wire  _EVAL_484;
  wire  _EVAL_411;
  wire  _EVAL_253;
  wire  _EVAL_558;
  wire  _EVAL_542;
  wire  _EVAL_532;
  wire  _EVAL_287;
  wire [31:0] _EVAL_633;
  wire  _EVAL_503;
  wire  _EVAL_348;
  wire  _EVAL_108;
  wire  _EVAL_388;
  wire  _EVAL_548;
  wire  _EVAL_593;
  wire [31:0] _EVAL_439;
  wire [32:0] _EVAL_398;
  wire [32:0] _EVAL_135;
  wire [32:0] _EVAL_339;
  wire  _EVAL_134;
  wire [32:0] _EVAL_652;
  wire [32:0] _EVAL_610;
  wire  _EVAL_141;
  wire  _EVAL_132;
  wire [2:0] _EVAL_397;
  wire  _EVAL_296;
  wire  _EVAL_190;
  wire  _EVAL_543;
  wire  _EVAL_211;
  wire  _EVAL_89;
  wire  _EVAL_480;
  wire  _EVAL_343;
  wire  _EVAL_420;
  wire [7:0] _EVAL_572;
  wire [31:0] _EVAL_567;
  wire [31:0] _EVAL_314;
  wire [31:0] _EVAL_233;
  wire [31:0] _EVAL_35;
  wire  _EVAL_195;
  wire  _EVAL_205;
  wire  _EVAL_609;
  wire [31:0] _EVAL_506;
  wire [32:0] _EVAL_522;
  wire [32:0] _EVAL_352;
  wire  _EVAL_223;
  wire  _EVAL_51;
  wire  _EVAL_565;
  wire  _EVAL_70;
  wire  _EVAL_198;
  wire  _EVAL_240;
  wire  _EVAL_171;
  wire  _EVAL_377;
  wire  _EVAL_44;
  wire  _EVAL_336;
  wire  _EVAL_473;
  wire  _EVAL_234;
  wire  _EVAL_410;
  wire [32:0] _EVAL_662;
  wire  _EVAL_432;
  wire [31:0] _EVAL_42;
  wire [32:0] _EVAL_449;
  wire [32:0] _EVAL_426;
  wire  _EVAL_185;
  wire  _EVAL_486;
  wire [31:0] _EVAL_550;
  wire [32:0] _EVAL_177;
  wire [32:0] _EVAL_122;
  wire [32:0] _EVAL_668;
  wire  _EVAL_197;
  wire  _EVAL_462;
  wire  _EVAL_39;
  wire [31:0] _EVAL_380;
  wire [31:0] _EVAL_644;
  wire  _EVAL_159;
  wire  _EVAL_337;
  wire [32:0] _EVAL_133;
  wire [32:0] _EVAL_311;
  wire [32:0] _EVAL_274;
  wire [31:0] _EVAL_553;
  wire [32:0] _EVAL_100;
  wire  _EVAL_327;
  wire  _EVAL_276;
  wire  _EVAL_370;
  wire  _EVAL_445;
  wire [32:0] _EVAL_175;
  wire [32:0] _EVAL_229;
  wire [32:0] _EVAL_512;
  wire  _EVAL_166;
  wire  _EVAL_555;
  wire  _EVAL_528;
  wire  _EVAL_586;
  wire  _EVAL_200;
  wire  _EVAL_646;
  wire  _EVAL_228;
  wire [31:0] _EVAL_523;
  wire  _EVAL_326;
  wire [31:0] _EVAL_124;
  wire [32:0] _EVAL_541;
  wire [32:0] _EVAL_630;
  wire [32:0] _EVAL_386;
  wire  _EVAL_530;
  wire  _EVAL_387;
  wire [32:0] _EVAL_423;
  wire [32:0] _EVAL_180;
  wire [32:0] _EVAL_126;
  wire  _EVAL_357;
  wire  _EVAL_91;
  wire [32:0] _EVAL_214;
  wire [32:0] _EVAL_241;
  wire  _EVAL_491;
  wire  _EVAL_74;
  wire [31:0] _EVAL_41;
  wire [32:0] _EVAL_658;
  wire [32:0] _EVAL_105;
  wire [32:0] _EVAL_664;
  wire  _EVAL_342;
  wire  _EVAL_282;
  wire  _EVAL_49;
  wire  _EVAL_215;
  wire  _EVAL_433;
  wire  _EVAL_267;
  wire  _EVAL_626;
  wire  _EVAL_616;
  wire  _EVAL_295;
  wire  _EVAL_489;
  wire  _EVAL_153;
  wire  _EVAL_189;
  wire  _EVAL_385;
  wire  _EVAL_341;
  wire  _EVAL_376;
  wire  _EVAL_361;
  wire  _EVAL_301;
  wire  _EVAL_581;
  wire  _EVAL_67;
  wire  _EVAL_303;
  wire  _EVAL_194;
  wire  _EVAL_118;
  wire  _EVAL_627;
  wire  _EVAL_183;
  wire  _EVAL_62;
  wire  _EVAL_450;
  wire  _EVAL_271;
  wire  _EVAL_288;
  wire  _EVAL_86;
  wire  _EVAL_591;
  wire  _EVAL_637;
  wire  _EVAL_594;
  wire  _EVAL_247;
  wire  _EVAL_576;
  wire  _EVAL_538;
  wire  _EVAL_279;
  wire  _EVAL_254;
  wire  _EVAL_140;
  wire  _EVAL_210;
  wire  _EVAL_309;
  wire  _EVAL_373;
  wire  _EVAL_539;
  wire  _EVAL_258;
  wire  _EVAL_611;
  wire [7:0] _EVAL_226;
  wire [7:0] _EVAL_421;
  wire [7:0] _EVAL_142;
  wire  _EVAL_624;
  wire  _EVAL_515;
  wire  _EVAL_497;
  wire [7:0] _EVAL_573;
  wire  _EVAL_599;
  wire  _EVAL_615;
  wire  _EVAL_83;
  wire [4:0] _EVAL_425;
  wire  _EVAL_43;
  wire [31:0] _EVAL_350;
  wire [32:0] _EVAL_384;
  wire [32:0] _EVAL_116;
  wire [32:0] _EVAL_75;
  wire  _EVAL_209;
  wire  _EVAL_482;
  wire  _EVAL_479;
  wire  _EVAL_536;
  wire  _EVAL_227;
  wire  _EVAL_405;
  wire [32:0] _EVAL_239;
  wire [32:0] _EVAL_321;
  wire  _EVAL_120;
  wire [31:0] _EVAL_109;
  wire [32:0] _EVAL_601;
  wire  _EVAL_268;
  wire  _EVAL_102;
  wire  _EVAL_475;
  wire  _EVAL_556;
  wire  _EVAL_441;
  wire  _EVAL_174;
  wire  _EVAL_242;
  wire  _EVAL_547;
  wire  _EVAL_155;
  wire  _EVAL_96;
  wire  _EVAL_218;
  wire [31:0] _EVAL_72;
  wire [32:0] _EVAL_391;
  wire [32:0] _EVAL_382;
  wire [31:0] _EVAL_485;
  wire  _EVAL_353;
  wire  _EVAL_306;
  wire [32:0] _EVAL_597;
  wire [32:0] _EVAL_551;
  wire [32:0] _EVAL_293;
  wire  _EVAL_381;
  wire  _EVAL_638;
  wire  _EVAL_534;
  wire  _EVAL_88;
  wire [32:0] _EVAL_265;
  wire [32:0] _EVAL_390;
  wire [32:0] _EVAL_643;
  wire  _EVAL_76;
  wire  _EVAL_670;
  wire  _EVAL_667;
  wire  _EVAL_202;
  wire  _EVAL_225;
  wire  _EVAL_113;
  wire [15:0] _EVAL_651;
  wire [15:0] _EVAL_79;
  wire  _EVAL_540;
  wire  _EVAL_106;
  wire  _EVAL_354;
  wire  _EVAL_367;
  wire  _EVAL_167;
  wire [31:0] _EVAL_535;
  wire [32:0] _EVAL_448;
  wire [32:0] _EVAL_659;
  wire [4:0] _EVAL_207;
  wire  _EVAL_564;
  wire [31:0] _EVAL_68;
  wire [32:0] _EVAL_143;
  wire [1:0] _EVAL_359;
  wire [1:0] _EVAL_246;
  wire [1:0] _EVAL_191;
  wire [2:0] _EVAL_291;
  wire  _EVAL_434;
  wire [32:0] _EVAL_531;
  wire  _EVAL_502;
  wire  _EVAL_61;
  wire [32:0] _EVAL_36;
  wire  _EVAL_575;
  wire  _EVAL_606;
  wire [32:0] _EVAL_346;
  wire [32:0] _EVAL_308;
  wire [32:0] _EVAL_582;
  wire  _EVAL_163;
  wire  _EVAL_262;
  wire [31:0] _EVAL_290;
  wire [32:0] _EVAL_368;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_647;
  wire  _EVAL_65;
  wire  _EVAL_590;
  wire [32:0] _EVAL_468;
  wire [32:0] _EVAL_330;
  wire [32:0] _EVAL_119;
  wire  _EVAL_220;
  wire  _EVAL_46;
  wire [32:0] _EVAL_145;
  wire [32:0] _EVAL_230;
  wire  _EVAL_642;
  wire  _EVAL_412;
  wire  _EVAL_409;
  wire  _EVAL_603;
  wire [32:0] _EVAL_213;
  wire [32:0] _EVAL_121;
  wire [32:0] _EVAL_161;
  wire  _EVAL_454;
  wire  _EVAL_598;
  wire  _EVAL_157;
  wire [1:0] _EVAL_516;
  wire  _EVAL_57;
  wire  _EVAL_78;
  wire  _EVAL_192;
  wire  _EVAL_623;
  wire [1:0] _EVAL_47;
  wire  _EVAL_272;
  wire  _EVAL_493;
  wire  _EVAL_164;
  wire  _EVAL_273;
  wire  _EVAL_55;
  wire  _EVAL_107;
  wire  _EVAL_238;
  wire  _EVAL_114;
  wire  _EVAL_193;
  wire  _EVAL_251;
  wire  _EVAL_160;
  wire  _EVAL_619;
  wire [2:0] _EVAL_40;
  wire  _EVAL_440;
  wire  _EVAL_69;
  wire  _EVAL_592;
  wire  _EVAL_666;
  wire [15:0] _EVAL_501;
  wire  _EVAL_110;
  wire  _EVAL_537;
  wire  _EVAL_495;
  wire  _EVAL_585;
  wire  _EVAL_507;
  wire  _EVAL_396;
  wire  _EVAL_349;
  wire  _EVAL_645;
  wire  _EVAL_469;
  wire [4:0] _EVAL_472;
  wire [4:0] _EVAL_184;
  wire  _EVAL_579;
  wire  _EVAL_455;
  wire  _EVAL_95;
  wire  _EVAL_517;
  wire  _EVAL_150;
  wire  _EVAL_612;
  wire  _EVAL_613;
  wire  _EVAL_212;
  wire  _EVAL_554;
  wire [8:0] _EVAL_631;
  wire [8:0] _EVAL_204;
  wire  _EVAL_443;
  wire  _EVAL_625;
  wire [15:0] _EVAL_54;
  wire [8:0] _EVAL_66;
  wire [8:0] _EVAL_90;
  wire [8:0] _EVAL_580;
  wire  _EVAL_50;
  wire  _EVAL_452;
  wire  _EVAL_338;
  wire  _EVAL_252;
  wire  _EVAL_149;
  wire  _EVAL_617;
  wire  _EVAL_431;
  wire  _EVAL_604;
  wire  _EVAL_477;
  wire  _EVAL_488;
  wire  _EVAL_498;
  wire  _EVAL_648;
  wire  _EVAL_257;
  wire [8:0] _EVAL_393;
  wire  _EVAL_56;
  wire  _EVAL_492;
  wire  _EVAL_588;
  wire  _EVAL_459;
  wire  _EVAL_176;
  wire  _EVAL_151;
  wire  _EVAL_101;
  wire  _EVAL_112;
  wire  _EVAL_269;
  wire  _EVAL_216;
  wire  _EVAL_152;
  wire  _EVAL_655;
  wire  _EVAL_569;
  wire  _EVAL_178;
  wire  _EVAL_453;
  wire  _EVAL_248;
  wire  _EVAL_456;
  wire  _EVAL_131;
  wire  _EVAL_173;
  wire  _EVAL_358;
  wire  _EVAL_158;
  wire  _EVAL_138;
  wire  _EVAL_529;
  wire  _EVAL_620;
  wire  _EVAL_584;
  wire  _EVAL_544;
  wire  _EVAL_186;
  wire [32:0] _EVAL_402;
  wire [32:0] _EVAL_347;
  wire [32:0] _EVAL_165;
  wire  _EVAL_460;
  wire  _EVAL_123;
  wire [8:0] _EVAL_115;
  wire  _EVAL_400;
  wire  _EVAL_444;
  wire [1:0] _EVAL_446;
  wire  _EVAL_414;
  wire  _EVAL_511;
  wire  _EVAL_392;
  wire  _EVAL_436;
  wire  _EVAL_438;
  wire  _EVAL_608;
  wire  _EVAL_451;
  wire  _EVAL_117;
  wire  _EVAL_104;
  wire  _EVAL_404;
  wire  _EVAL_641;
  wire  _EVAL_640;
  wire  _EVAL_312;
  wire [31:0] _EVAL_514;
  wire  _EVAL_499;
  wire  _EVAL_513;
  wire  _EVAL_345;
  wire  _EVAL_494;
  wire  _EVAL_259;
  wire  _EVAL_395;
  wire  _EVAL_275;
  wire  _EVAL_34;
  wire  _EVAL_344;
  wire  _EVAL_635;
  wire [4:0] _EVAL_324;
  wire [4:0] _EVAL_208;
  wire  _EVAL_546;
  wire  _EVAL_415;
  wire  _EVAL_154;
  wire  _EVAL_521;
  wire  _EVAL_661;
  wire  _EVAL_98;
  wire  _EVAL_144;
  wire [8:0] _EVAL_256;
  wire  _EVAL_261;
  wire  _EVAL_221;
  wire  _EVAL_622;
  wire  _EVAL_328;
  wire  _EVAL_634;
  wire [4:0] _EVAL_219;
  wire  _EVAL_654;
  wire  _EVAL_561;
  wire  _EVAL_509;
  wire  _EVAL_602;
  wire  _EVAL_80;
  wire [32:0] _EVAL_280;
  wire [32:0] _EVAL_562;
  wire  _EVAL_93;
  wire  _EVAL_524;
  wire  _EVAL_307;
  wire  _EVAL_187;
  wire  _EVAL_310;
  wire  _EVAL_403;
  wire  _EVAL_430;
  wire [32:0] _EVAL_389;
  wire  _EVAL_245;
  wire  _EVAL_416;
  wire  _EVAL_600;
  wire [4:0] _EVAL_372;
  wire  _EVAL_281;
  wire  _EVAL_315;
  wire  _EVAL_224;
  wire  _EVAL_653;
  wire  _EVAL_182;
  wire  _EVAL_563;
  wire  _EVAL_533;
  wire  _EVAL_300;
  wire  _EVAL_63;
  wire  _EVAL_146;
  wire  _EVAL_466;
  wire  _EVAL_169;
  wire  _EVAL_478;
  wire  _EVAL_318;
  wire  _EVAL_294;
  wire  _EVAL_333;
  wire  _EVAL_457;
  wire  _EVAL_249;
  wire  _EVAL_77;
  wire  _EVAL_85;
  wire  _EVAL_355;
  wire  _EVAL_424;
  wire  _EVAL_596;
  wire  _EVAL_657;
  wire  _EVAL_374;
  wire  _EVAL_292;
  wire  _EVAL_520;
  wire  _EVAL_481;
  wire  _EVAL_129;
  wire  _EVAL_650;
  wire  _EVAL_660;
  wire  _EVAL_260;
  wire  _EVAL_639;
  wire  _EVAL_137;
  wire  _EVAL_284;
  wire  _EVAL_364;
  wire  _EVAL_500;
  wire  _EVAL_371;
  wire  _EVAL_340;
  wire  _EVAL_549;
  wire  _EVAL_325;
  wire  _EVAL_317;
  wire  _EVAL_365;
  wire  _EVAL_179;
  wire  _EVAL_629;
  wire  _EVAL_320;
  wire  _EVAL_127;
  wire  _EVAL_266;
  wire  _EVAL_243;
  wire  _EVAL_97;
  wire  _EVAL_577;
  wire  _EVAL_139;
  wire [4:0] _EVAL_583;
  wire  _EVAL_302;
  wire  _EVAL_87;
  wire  _EVAL_71;
  wire  _EVAL_447;
  wire  _EVAL_632;
  wire  _EVAL_45;
  wire  _EVAL_250;
  wire  _EVAL_422;
  wire  _EVAL_298;
  wire  _EVAL_188;
  wire  _EVAL_331;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_277 = 23'hff << _EVAL_15;
  assign _EVAL_332 = _EVAL_14 ^ 32'h20000000;
  assign _EVAL_560 = {1'b0,$signed(_EVAL_332)};
  assign _EVAL_59 = _EVAL_607 != 9'h0;
  assign _EVAL_103 = _EVAL_59 == 1'h0;
  assign _EVAL_525 = plusarg_reader_out == 32'h0;
  assign _EVAL_222 = _EVAL_103 | _EVAL_525;
  assign _EVAL_329 = _EVAL_235 < plusarg_reader_out;
  assign _EVAL_467 = _EVAL_222 | _EVAL_329;
  assign _EVAL_217 = _EVAL_16 & _EVAL_29;
  assign _EVAL_231 = _EVAL_17 & _EVAL_10;
  assign _EVAL_595 = _EVAL_217 | _EVAL_231;
  assign _EVAL_99 = _EVAL_0 ^ 32'h80000000;
  assign _EVAL_322 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_649 = _EVAL_277[7:0];
  assign _EVAL_394 = ~ _EVAL_649;
  assign _EVAL_366 = {{24'd0}, _EVAL_394};
  assign _EVAL_264 = _EVAL_0 & _EVAL_366;
  assign _EVAL_465 = _EVAL_264 == 32'h0;
  assign _EVAL_335 = _EVAL_14 ^ 32'h40000000;
  assign _EVAL_571 = {1'b0,$signed(_EVAL_335)};
  assign _EVAL_519 = $signed(_EVAL_571) & $signed(-33'sh2000);
  assign _EVAL_206 = $signed(_EVAL_519);
  assign _EVAL_111 = $signed(_EVAL_206) == $signed(33'sh0);
  assign _EVAL_199 = _EVAL_14 ^ 32'h80000000;
  assign _EVAL_656 = {1'b0,$signed(_EVAL_199)};
  assign _EVAL_81 = $signed(_EVAL_656) & $signed(-33'sh20000);
  assign _EVAL_128 = $signed(_EVAL_81);
  assign _EVAL_378 = $signed(_EVAL_128) == $signed(33'sh0);
  assign _EVAL_270 = _EVAL_111 | _EVAL_378;
  assign _EVAL_505 = _EVAL_14 ^ 32'h3000;
  assign _EVAL_559 = {1'b0,$signed(_EVAL_505)};
  assign _EVAL_399 = $signed(_EVAL_559) & $signed(-33'sh1000);
  assign _EVAL_334 = $signed(_EVAL_399);
  assign _EVAL_526 = $signed(_EVAL_334) == $signed(33'sh0);
  assign _EVAL_379 = _EVAL_270 | _EVAL_526;
  assign _EVAL_125 = _EVAL_9 <= 2'h2;
  assign _EVAL_487 = _EVAL_125 | _EVAL_32;
  assign _EVAL_429 = _EVAL_1 == 3'h5;
  assign _EVAL_589 = _EVAL_3 == 4'h8;
  assign _EVAL_196 = _EVAL_15 == _EVAL_628;
  assign _EVAL_408 = 23'hff << _EVAL_31;
  assign _EVAL_362 = _EVAL_408[7:0];
  assign _EVAL_263 = _EVAL_15[1:0];
  assign _EVAL_48 = 4'h1 << _EVAL_263;
  assign _EVAL_621 = _EVAL_48[2:0];
  assign _EVAL_552 = _EVAL_621 | 3'h1;
  assign _EVAL_570 = _EVAL_552[0];
  assign _EVAL_483 = _EVAL_0[2];
  assign _EVAL_363 = _EVAL_0[1];
  assign _EVAL_299 = _EVAL_363 == 1'h0;
  assign _EVAL_82 = _EVAL_483 & _EVAL_299;
  assign _EVAL_172 = _EVAL_0[0];
  assign _EVAL_148 = _EVAL_172 == 1'h0;
  assign _EVAL_84 = _EVAL_82 & _EVAL_148;
  assign _EVAL_476 = _EVAL_570 & _EVAL_84;
  assign _EVAL_94 = _EVAL_3 == _EVAL_360;
  assign _EVAL_73 = _EVAL_94 | _EVAL_32;
  assign _EVAL_181 = _EVAL_23 == 1'h0;
  assign _EVAL_508 = _EVAL_0 == _EVAL_587;
  assign _EVAL_427 = _EVAL_18 == 4'h0;
  assign _EVAL_305 = _EVAL_413 == 5'h0;
  assign _EVAL_170 = _EVAL_231 & _EVAL_305;
  assign _EVAL_496 = _EVAL_11[2];
  assign _EVAL_356 = _EVAL_11[1];
  assign _EVAL_510 = _EVAL_356 == 1'h0;
  assign _EVAL_156 = _EVAL_496 & _EVAL_510;
  assign _EVAL_255 = _EVAL_170 & _EVAL_156;
  assign _EVAL_162 = 2'h1 << _EVAL_24;
  assign _EVAL_236 = _EVAL_255 ? _EVAL_162 : 2'h0;
  assign _EVAL_38 = _EVAL_236 | _EVAL_470;
  assign _EVAL_669 = _EVAL_38 >> _EVAL_25;
  assign _EVAL_313 = _EVAL_669[0];
  assign _EVAL_419 = _EVAL_313 | _EVAL_32;
  assign _EVAL_665 = 23'hff << _EVAL;
  assign _EVAL_53 = _EVAL_665[7:0];
  assign _EVAL_60 = ~ _EVAL_53;
  assign _EVAL_578 = _EVAL_60[7:3];
  assign _EVAL_614 = _EVAL_7 ^ 32'h80000000;
  assign _EVAL_618 = {1'b0,$signed(_EVAL_614)};
  assign _EVAL_490 = $signed(_EVAL_618) & $signed(-33'sh20000);
  assign _EVAL_401 = $signed(_EVAL_490);
  assign _EVAL_566 = $signed(_EVAL_401) == $signed(33'sh0);
  assign _EVAL_319 = _EVAL_0 ^ 32'h20000000;
  assign _EVAL_545 = {1'b0,$signed(_EVAL_319)};
  assign _EVAL_136 = $signed(_EVAL_545) & $signed(-33'sh2000);
  assign _EVAL_285 = $signed(_EVAL_136);
  assign _EVAL_232 = $signed(_EVAL_285) == $signed(33'sh0);
  assign _EVAL_527 = _EVAL_1 == 3'h1;
  assign _EVAL_484 = _EVAL_406 == 5'h0;
  assign _EVAL_411 = _EVAL_30 == _EVAL_283;
  assign _EVAL_253 = _EVAL_411 | _EVAL_32;
  assign _EVAL_558 = _EVAL_28 == 3'h6;
  assign _EVAL_542 = _EVAL_6 & _EVAL_558;
  assign _EVAL_532 = _EVAL_323 == 5'h0;
  assign _EVAL_287 = _EVAL_532 == 1'h0;
  assign _EVAL_633 = _EVAL_14 ^ 32'h2000000;
  assign _EVAL_503 = _EVAL_1 == 3'h0;
  assign _EVAL_348 = _EVAL_28 == 3'h0;
  assign _EVAL_108 = _EVAL_6 & _EVAL_348;
  assign _EVAL_388 = _EVAL_37 == 5'h0;
  assign _EVAL_548 = _EVAL_388 == 1'h0;
  assign _EVAL_593 = _EVAL_27 == _EVAL_464;
  assign _EVAL_439 = _EVAL_0 ^ 32'h40000000;
  assign _EVAL_398 = {1'b0,$signed(_EVAL_439)};
  assign _EVAL_135 = $signed(_EVAL_398) & $signed(-33'sh2000);
  assign _EVAL_339 = $signed(_EVAL_135);
  assign _EVAL_134 = $signed(_EVAL_339) == $signed(33'sh0);
  assign _EVAL_652 = $signed(_EVAL_322) & $signed(-33'sh20000);
  assign _EVAL_610 = $signed(_EVAL_652);
  assign _EVAL_141 = $signed(_EVAL_610) == $signed(33'sh0);
  assign _EVAL_132 = _EVAL_134 | _EVAL_141;
  assign _EVAL_397 = _EVAL_18[2:0];
  assign _EVAL_296 = 3'h1 <= _EVAL_397;
  assign _EVAL_190 = _EVAL_19 != 3'h0;
  assign _EVAL_543 = _EVAL_190 | _EVAL_32;
  assign _EVAL_211 = _EVAL_3 == 4'h0;
  assign _EVAL_89 = 4'h6 == _EVAL_15;
  assign _EVAL_480 = _EVAL_211 ? _EVAL_89 : 1'h0;
  assign _EVAL_343 = _EVAL_480 | _EVAL_32;
  assign _EVAL_420 = _EVAL_343 == 1'h0;
  assign _EVAL_572 = ~ _EVAL_362;
  assign _EVAL_567 = {{24'd0}, _EVAL_572};
  assign _EVAL_314 = _EVAL_14 & _EVAL_567;
  assign _EVAL_233 = _EVAL_14 ^ 32'hc000000;
  assign _EVAL_35 = _EVAL_7 & 32'h3f;
  assign _EVAL_195 = _EVAL_35 == 32'h0;
  assign _EVAL_205 = _EVAL_195 | _EVAL_32;
  assign _EVAL_609 = _EVAL_205 == 1'h0;
  assign _EVAL_506 = _EVAL_7 ^ 32'h4000;
  assign _EVAL_522 = {1'b0,$signed(_EVAL_506)};
  assign _EVAL_352 = $signed(_EVAL_522) & $signed(-33'sh1000);
  assign _EVAL_223 = _EVAL_18 == 4'h8;
  assign _EVAL_51 = _EVAL_223 | _EVAL_427;
  assign _EVAL_565 = _EVAL_18[3:3];
  assign _EVAL_70 = _EVAL_565 == 1'h0;
  assign _EVAL_198 = _EVAL_70 & _EVAL_296;
  assign _EVAL_240 = _EVAL_51 | _EVAL_198;
  assign _EVAL_171 = _EVAL_240 | _EVAL_32;
  assign _EVAL_377 = _EVAL_1[2];
  assign _EVAL_44 = _EVAL_543 == 1'h0;
  assign _EVAL_336 = _EVAL_73 == 1'h0;
  assign _EVAL_473 = _EVAL_15 <= 4'h6;
  assign _EVAL_234 = _EVAL_473 & _EVAL_141;
  assign _EVAL_410 = _EVAL_28 == 3'h2;
  assign _EVAL_662 = $signed(_EVAL_352);
  assign _EVAL_432 = $signed(_EVAL_662) == $signed(33'sh0);
  assign _EVAL_42 = _EVAL_7 ^ 32'h40000000;
  assign _EVAL_449 = {1'b0,$signed(_EVAL_42)};
  assign _EVAL_426 = $signed(_EVAL_449) & $signed(-33'sh2000);
  assign _EVAL_185 = _EVAL_24 == _EVAL_351;
  assign _EVAL_486 = _EVAL_185 | _EVAL_32;
  assign _EVAL_550 = _EVAL_0 ^ 32'hc000000;
  assign _EVAL_177 = {1'b0,$signed(_EVAL_550)};
  assign _EVAL_122 = $signed(_EVAL_177) & $signed(-33'sh4000000);
  assign _EVAL_668 = $signed(_EVAL_122);
  assign _EVAL_197 = $signed(_EVAL_668) == $signed(33'sh0);
  assign _EVAL_462 = _EVAL_14 == _EVAL_278;
  assign _EVAL_39 = _EVAL_462 | _EVAL_32;
  assign _EVAL_380 = _EVAL_7 ^ 32'h20000000;
  assign _EVAL_644 = _EVAL_0 ^ 32'h3000;
  assign _EVAL_159 = _EVAL_26 == 1'h0;
  assign _EVAL_337 = _EVAL_159 | _EVAL_4;
  assign _EVAL_133 = {1'b0,$signed(_EVAL_633)};
  assign _EVAL_311 = $signed(_EVAL_133) & $signed(-33'sh10000);
  assign _EVAL_274 = $signed(_EVAL_311);
  assign _EVAL_553 = _EVAL_0 ^ 32'h1800000;
  assign _EVAL_100 = {1'b0,$signed(_EVAL_553)};
  assign _EVAL_327 = _EVAL_31 <= 4'h6;
  assign _EVAL_276 = _EVAL_327 & _EVAL_378;
  assign _EVAL_370 = _EVAL_276 | _EVAL_32;
  assign _EVAL_445 = _EVAL_370 == 1'h0;
  assign _EVAL_175 = {1'b0,$signed(_EVAL_644)};
  assign _EVAL_229 = $signed(_EVAL_175) & $signed(-33'sh1000);
  assign _EVAL_512 = $signed(_EVAL_229);
  assign _EVAL_166 = $signed(_EVAL_512) == $signed(33'sh0);
  assign _EVAL_555 = _EVAL_166 | _EVAL_197;
  assign _EVAL_528 = _EVAL_314 == 32'h0;
  assign _EVAL_586 = _EVAL_231 & _EVAL_388;
  assign _EVAL_200 = _EVAL_483 == 1'h0;
  assign _EVAL_646 = _EVAL_200 & _EVAL_363;
  assign _EVAL_228 = _EVAL_39 == 1'h0;
  assign _EVAL_523 = _EVAL_7 ^ 32'hc000000;
  assign _EVAL_326 = _EVAL_132 | _EVAL_197;
  assign _EVAL_124 = _EVAL_0 ^ 32'h2000000;
  assign _EVAL_541 = {1'b0,$signed(_EVAL_124)};
  assign _EVAL_630 = $signed(_EVAL_541) & $signed(-33'sh10000);
  assign _EVAL_386 = $signed(_EVAL_630);
  assign _EVAL_530 = $signed(_EVAL_386) == $signed(33'sh0);
  assign _EVAL_387 = _EVAL_326 | _EVAL_530;
  assign _EVAL_423 = {1'b0,$signed(_EVAL_0)};
  assign _EVAL_180 = $signed(_EVAL_423) & $signed(-33'sh5000);
  assign _EVAL_126 = $signed(_EVAL_180);
  assign _EVAL_357 = $signed(_EVAL_126) == $signed(33'sh0);
  assign _EVAL_91 = _EVAL_387 | _EVAL_357;
  assign _EVAL_214 = $signed(_EVAL_100) & $signed(-33'sh8000);
  assign _EVAL_241 = $signed(_EVAL_214);
  assign _EVAL_491 = $signed(_EVAL_241) == $signed(33'sh0);
  assign _EVAL_74 = _EVAL_91 | _EVAL_491;
  assign _EVAL_41 = _EVAL_0 ^ 32'h1900000;
  assign _EVAL_658 = {1'b0,$signed(_EVAL_41)};
  assign _EVAL_105 = $signed(_EVAL_658) & $signed(-33'sh2000);
  assign _EVAL_664 = $signed(_EVAL_105);
  assign _EVAL_342 = $signed(_EVAL_664) == $signed(33'sh0);
  assign _EVAL_282 = _EVAL_74 | _EVAL_342;
  assign _EVAL_49 = _EVAL_28 == 3'h5;
  assign _EVAL_215 = _EVAL_6 & _EVAL_49;
  assign _EVAL_433 = _EVAL_15 <= 4'h8;
  assign _EVAL_267 = _EVAL_15 >= 4'h3;
  assign _EVAL_626 = _EVAL_552[2];
  assign _EVAL_616 = _EVAL_626 & _EVAL_483;
  assign _EVAL_295 = _EVAL_267 | _EVAL_616;
  assign _EVAL_489 = _EVAL_552[1];
  assign _EVAL_153 = _EVAL_483 & _EVAL_363;
  assign _EVAL_189 = _EVAL_489 & _EVAL_153;
  assign _EVAL_385 = _EVAL_295 | _EVAL_189;
  assign _EVAL_341 = _EVAL_153 & _EVAL_172;
  assign _EVAL_376 = _EVAL_570 & _EVAL_341;
  assign _EVAL_361 = _EVAL_385 | _EVAL_376;
  assign _EVAL_301 = _EVAL_153 & _EVAL_148;
  assign _EVAL_581 = _EVAL_570 & _EVAL_301;
  assign _EVAL_67 = _EVAL_385 | _EVAL_581;
  assign _EVAL_303 = _EVAL_489 & _EVAL_82;
  assign _EVAL_194 = _EVAL_295 | _EVAL_303;
  assign _EVAL_118 = _EVAL_82 & _EVAL_172;
  assign _EVAL_627 = _EVAL_570 & _EVAL_118;
  assign _EVAL_183 = _EVAL_194 | _EVAL_627;
  assign _EVAL_62 = _EVAL_194 | _EVAL_476;
  assign _EVAL_450 = _EVAL_626 & _EVAL_200;
  assign _EVAL_271 = _EVAL_267 | _EVAL_450;
  assign _EVAL_288 = _EVAL_489 & _EVAL_646;
  assign _EVAL_86 = _EVAL_271 | _EVAL_288;
  assign _EVAL_591 = _EVAL_646 & _EVAL_172;
  assign _EVAL_637 = _EVAL_570 & _EVAL_591;
  assign _EVAL_594 = _EVAL_86 | _EVAL_637;
  assign _EVAL_247 = _EVAL_646 & _EVAL_148;
  assign _EVAL_576 = _EVAL_570 & _EVAL_247;
  assign _EVAL_538 = _EVAL_86 | _EVAL_576;
  assign _EVAL_279 = _EVAL_200 & _EVAL_299;
  assign _EVAL_254 = _EVAL_489 & _EVAL_279;
  assign _EVAL_140 = _EVAL_271 | _EVAL_254;
  assign _EVAL_210 = _EVAL_279 & _EVAL_172;
  assign _EVAL_309 = _EVAL_570 & _EVAL_210;
  assign _EVAL_373 = _EVAL_140 | _EVAL_309;
  assign _EVAL_539 = _EVAL_279 & _EVAL_148;
  assign _EVAL_258 = _EVAL_570 & _EVAL_539;
  assign _EVAL_611 = _EVAL_140 | _EVAL_258;
  assign _EVAL_226 = {_EVAL_361,_EVAL_67,_EVAL_183,_EVAL_62,_EVAL_594,_EVAL_538,_EVAL_373,_EVAL_611};
  assign _EVAL_421 = ~ _EVAL_226;
  assign _EVAL_142 = _EVAL_8 & _EVAL_421;
  assign _EVAL_624 = _EVAL_142 == 8'h0;
  assign _EVAL_515 = _EVAL_624 | _EVAL_32;
  assign _EVAL_497 = _EVAL_515 == 1'h0;
  assign _EVAL_573 = ~ _EVAL_8;
  assign _EVAL_599 = _EVAL_573 == 8'h0;
  assign _EVAL_615 = _EVAL_599 | _EVAL_32;
  assign _EVAL_83 = _EVAL_377 == 1'h0;
  assign _EVAL_425 = _EVAL_406 - 5'h1;
  assign _EVAL_43 = _EVAL_181 | _EVAL_32;
  assign _EVAL_350 = _EVAL_7 ^ 32'h1900000;
  assign _EVAL_384 = {1'b0,$signed(_EVAL_350)};
  assign _EVAL_116 = $signed(_EVAL_384) & $signed(-33'sh2000);
  assign _EVAL_75 = $signed(_EVAL_116);
  assign _EVAL_209 = $signed(_EVAL_75) == $signed(33'sh0);
  assign _EVAL_482 = _EVAL_11 == _EVAL_474;
  assign _EVAL_479 = _EVAL_482 | _EVAL_32;
  assign _EVAL_536 = _EVAL_479 == 1'h0;
  assign _EVAL_227 = _EVAL >= 4'h3;
  assign _EVAL_405 = _EVAL_555 | _EVAL_530;
  assign _EVAL_239 = $signed(_EVAL_560) & $signed(-33'sh2000);
  assign _EVAL_321 = $signed(_EVAL_239);
  assign _EVAL_120 = $signed(_EVAL_321) == $signed(33'sh0);
  assign _EVAL_109 = _EVAL_7 ^ 32'h1800000;
  assign _EVAL_601 = {1'b0,$signed(_EVAL_109)};
  assign _EVAL_268 = _EVAL_15 <= 4'h2;
  assign _EVAL_102 = _EVAL_405 | _EVAL_357;
  assign _EVAL_475 = _EVAL_102 | _EVAL_491;
  assign _EVAL_556 = _EVAL_475 | _EVAL_342;
  assign _EVAL_441 = _EVAL_556 | _EVAL_232;
  assign _EVAL_174 = _EVAL_268 & _EVAL_441;
  assign _EVAL_242 = _EVAL_174 | _EVAL_32;
  assign _EVAL_547 = _EVAL_242 == 1'h0;
  assign _EVAL_155 = _EVAL_201 == 5'h0;
  assign _EVAL_96 = _EVAL_155 == 1'h0;
  assign _EVAL_218 = _EVAL_2 & _EVAL_96;
  assign _EVAL_72 = _EVAL_7 ^ 32'h3000;
  assign _EVAL_391 = {1'b0,$signed(_EVAL_72)};
  assign _EVAL_382 = $signed(_EVAL_391) & $signed(-33'sh1000);
  assign _EVAL_485 = _EVAL_14 ^ 32'h1800000;
  assign _EVAL_353 = _EVAL_11 <= 3'h6;
  assign _EVAL_306 = _EVAL_353 | _EVAL_32;
  assign _EVAL_597 = {1'b0,$signed(_EVAL_233)};
  assign _EVAL_551 = $signed(_EVAL_597) & $signed(-33'sh4000000);
  assign _EVAL_293 = $signed(_EVAL_551);
  assign _EVAL_381 = $signed(_EVAL_293) == $signed(33'sh0);
  assign _EVAL_638 = _EVAL_379 | _EVAL_381;
  assign _EVAL_534 = $signed(_EVAL_274) == $signed(33'sh0);
  assign _EVAL_88 = _EVAL_638 | _EVAL_534;
  assign _EVAL_265 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_390 = $signed(_EVAL_265) & $signed(-33'sh1000);
  assign _EVAL_643 = $signed(_EVAL_390);
  assign _EVAL_76 = $signed(_EVAL_643) == $signed(33'sh0);
  assign _EVAL_670 = _EVAL_88 | _EVAL_76;
  assign _EVAL_667 = _EVAL_28 == 3'h4;
  assign _EVAL_202 = _EVAL_11 == 3'h6;
  assign _EVAL_225 = _EVAL_316 == 5'h0;
  assign _EVAL_113 = _EVAL_217 & _EVAL_225;
  assign _EVAL_651 = 16'h1 << _EVAL_3;
  assign _EVAL_79 = _EVAL_113 ? _EVAL_651 : 16'h0;
  assign _EVAL_540 = _EVAL_231 & _EVAL_484;
  assign _EVAL_106 = _EVAL_26 == _EVAL_407;
  assign _EVAL_354 = _EVAL_106 | _EVAL_32;
  assign _EVAL_367 = _EVAL_1 == _EVAL_168;
  assign _EVAL_167 = _EVAL_367 | _EVAL_32;
  assign _EVAL_535 = _EVAL_14 ^ 32'h4000;
  assign _EVAL_448 = {1'b0,$signed(_EVAL_535)};
  assign _EVAL_659 = $signed(_EVAL_448) & $signed(-33'sh1000);
  assign _EVAL_207 = _EVAL_201 - 5'h1;
  assign _EVAL_564 = _EVAL_589 | _EVAL_211;
  assign _EVAL_68 = _EVAL_14 ^ 32'h1900000;
  assign _EVAL_143 = {1'b0,$signed(_EVAL_68)};
  assign _EVAL_359 = _EVAL_470 | _EVAL_236;
  assign _EVAL_246 = 2'h1 << _EVAL_25;
  assign _EVAL_191 = _EVAL_22 ? _EVAL_246 : 2'h0;
  assign _EVAL_291 = _EVAL_3[2:0];
  assign _EVAL_434 = 3'h1 <= _EVAL_291;
  assign _EVAL_531 = $signed(_EVAL_426);
  assign _EVAL_502 = $signed(_EVAL_531) == $signed(33'sh0);
  assign _EVAL_61 = _EVAL_502 | _EVAL_566;
  assign _EVAL_36 = $signed(_EVAL_382);
  assign _EVAL_575 = $signed(_EVAL_36) == $signed(33'sh0);
  assign _EVAL_606 = _EVAL_61 | _EVAL_575;
  assign _EVAL_346 = {1'b0,$signed(_EVAL_523)};
  assign _EVAL_308 = $signed(_EVAL_346) & $signed(-33'sh4000000);
  assign _EVAL_582 = $signed(_EVAL_308);
  assign _EVAL_163 = $signed(_EVAL_582) == $signed(33'sh0);
  assign _EVAL_262 = _EVAL_606 | _EVAL_163;
  assign _EVAL_290 = _EVAL_7 ^ 32'h2000000;
  assign _EVAL_368 = {1'b0,$signed(_EVAL_290)};
  assign _EVAL_130 = $signed(_EVAL_368) & $signed(-33'sh10000);
  assign _EVAL_647 = $signed(_EVAL_130);
  assign _EVAL_65 = $signed(_EVAL_647) == $signed(33'sh0);
  assign _EVAL_590 = _EVAL_262 | _EVAL_65;
  assign _EVAL_468 = {1'b0,$signed(_EVAL_7)};
  assign _EVAL_330 = $signed(_EVAL_468) & $signed(-33'sh1000);
  assign _EVAL_119 = $signed(_EVAL_330);
  assign _EVAL_220 = $signed(_EVAL_119) == $signed(33'sh0);
  assign _EVAL_46 = _EVAL_590 | _EVAL_220;
  assign _EVAL_145 = $signed(_EVAL_601) & $signed(-33'sh8000);
  assign _EVAL_230 = $signed(_EVAL_145);
  assign _EVAL_642 = $signed(_EVAL_230) == $signed(33'sh0);
  assign _EVAL_412 = _EVAL_46 | _EVAL_642;
  assign _EVAL_409 = _EVAL_412 | _EVAL_209;
  assign _EVAL_603 = _EVAL_409 | _EVAL_432;
  assign _EVAL_213 = {1'b0,$signed(_EVAL_380)};
  assign _EVAL_121 = $signed(_EVAL_213) & $signed(-33'sh2000);
  assign _EVAL_161 = $signed(_EVAL_121);
  assign _EVAL_454 = $signed(_EVAL_161) == $signed(33'sh0);
  assign _EVAL_598 = _EVAL_603 | _EVAL_454;
  assign _EVAL_157 = _EVAL_598 | _EVAL_32;
  assign _EVAL_516 = _EVAL_470 >> _EVAL_24;
  assign _EVAL_57 = _EVAL_516[0];
  assign _EVAL_78 = _EVAL_57 == 1'h0;
  assign _EVAL_192 = _EVAL_78 | _EVAL_32;
  assign _EVAL_623 = _EVAL_192 == 1'h0;
  assign _EVAL_47 = ~ _EVAL_191;
  assign _EVAL_272 = _EVAL_354 == 1'h0;
  assign _EVAL_493 = _EVAL_8 == _EVAL_226;
  assign _EVAL_164 = _EVAL_493 | _EVAL_32;
  assign _EVAL_273 = _EVAL_164 == 1'h0;
  assign _EVAL_55 = _EVAL_28 == _EVAL_557;
  assign _EVAL_107 = _EVAL_55 | _EVAL_32;
  assign _EVAL_238 = _EVAL_31 >= 4'h3;
  assign _EVAL_114 = _EVAL_238 | _EVAL_32;
  assign _EVAL_193 = _EVAL_9 != 2'h2;
  assign _EVAL_251 = _EVAL_193 | _EVAL_32;
  assign _EVAL_160 = _EVAL_282 | _EVAL_232;
  assign _EVAL_619 = _EVAL_11[0];
  assign _EVAL_40 = _EVAL_27[2:0];
  assign _EVAL_440 = 3'h1 <= _EVAL_40;
  assign _EVAL_69 = _EVAL_528 | _EVAL_32;
  assign _EVAL_592 = _EVAL_69 == 1'h0;
  assign _EVAL_666 = _EVAL_487 == 1'h0;
  assign _EVAL_501 = 16'h1 << _EVAL_27;
  assign _EVAL_110 = _EVAL_19 <= 3'h2;
  assign _EVAL_537 = _EVAL_110 | _EVAL_32;
  assign _EVAL_495 = _EVAL_537 == 1'h0;
  assign _EVAL_585 = _EVAL_3[3:3];
  assign _EVAL_507 = _EVAL_585 == 1'h0;
  assign _EVAL_396 = _EVAL_507 & _EVAL_434;
  assign _EVAL_349 = _EVAL_107 == 1'h0;
  assign _EVAL_645 = _EVAL_11 == 3'h1;
  assign _EVAL_469 = _EVAL_442 == 5'h0;
  assign _EVAL_472 = _EVAL_394[7:3];
  assign _EVAL_184 = _EVAL_442 - 5'h1;
  assign _EVAL_579 = _EVAL_20 <= 2'h2;
  assign _EVAL_455 = _EVAL_579 | _EVAL_32;
  assign _EVAL_95 = _EVAL_455 == 1'h0;
  assign _EVAL_517 = _EVAL_28 == 3'h1;
  assign _EVAL_150 = _EVAL_6 & _EVAL_517;
  assign _EVAL_612 = _EVAL_465 | _EVAL_32;
  assign _EVAL_613 = _EVAL_612 == 1'h0;
  assign _EVAL_212 = _EVAL_9 == _EVAL_369;
  assign _EVAL_554 = _EVAL_212 | _EVAL_32;
  assign _EVAL_631 = _EVAL_79[8:0];
  assign _EVAL_204 = _EVAL_607 | _EVAL_631;
  assign _EVAL_443 = _EVAL_202 == 1'h0;
  assign _EVAL_625 = _EVAL_540 & _EVAL_443;
  assign _EVAL_54 = _EVAL_625 ? _EVAL_501 : 16'h0;
  assign _EVAL_66 = _EVAL_54[8:0];
  assign _EVAL_90 = ~ _EVAL_66;
  assign _EVAL_580 = _EVAL_204 & _EVAL_90;
  assign _EVAL_50 = _EVAL_11 == 3'h0;
  assign _EVAL_452 = _EVAL_10 & _EVAL_50;
  assign _EVAL_338 = _EVAL_6 & _EVAL_410;
  assign _EVAL_252 = _EVAL_253 == 1'h0;
  assign _EVAL_149 = _EVAL_27 == 4'h8;
  assign _EVAL_617 = _EVAL_30 <= 3'h2;
  assign _EVAL_431 = _EVAL_617 | _EVAL_32;
  assign _EVAL_604 = _EVAL_431 == 1'h0;
  assign _EVAL_477 = _EVAL_508 | _EVAL_32;
  assign _EVAL_488 = _EVAL_157 == 1'h0;
  assign _EVAL_498 = _EVAL_227 | _EVAL_32;
  assign _EVAL_648 = _EVAL_498 == 1'h0;
  assign _EVAL_257 = _EVAL_11 == 3'h4;
  assign _EVAL_393 = _EVAL_631 | _EVAL_607;
  assign _EVAL_56 = _EVAL_19 == 3'h0;
  assign _EVAL_492 = _EVAL_56 | _EVAL_32;
  assign _EVAL_588 = _EVAL_492 == 1'h0;
  assign _EVAL_459 = _EVAL_4 == 1'h0;
  assign _EVAL_176 = _EVAL_30 == 3'h0;
  assign _EVAL_151 = _EVAL_433 & _EVAL_166;
  assign _EVAL_101 = _EVAL_151 | _EVAL_32;
  assign _EVAL_112 = _EVAL_30 <= 3'h5;
  assign _EVAL_269 = _EVAL_112 | _EVAL_32;
  assign _EVAL_216 = _EVAL_18 == _EVAL_435;
  assign _EVAL_152 = _EVAL_216 | _EVAL_32;
  assign _EVAL_655 = _EVAL_152 == 1'h0;
  assign _EVAL_569 = _EVAL_11 == 3'h2;
  assign _EVAL_178 = _EVAL_10 & _EVAL_569;
  assign _EVAL_453 = _EVAL_267 | _EVAL_32;
  assign _EVAL_248 = _EVAL_5 == 1'h0;
  assign _EVAL_456 = _EVAL_248 | _EVAL_32;
  assign _EVAL_131 = _EVAL_564 | _EVAL_396;
  assign _EVAL_173 = _EVAL_131 | _EVAL_32;
  assign _EVAL_358 = _EVAL_631 != 9'h0;
  assign _EVAL_158 = _EVAL_358 == 1'h0;
  assign _EVAL_138 = _EVAL_12 & _EVAL_2;
  assign _EVAL_529 = _EVAL_234 | _EVAL_32;
  assign _EVAL_620 = _EVAL_529 == 1'h0;
  assign _EVAL_584 = _EVAL_10 & _EVAL_202;
  assign _EVAL_544 = _EVAL_6 & _EVAL_287;
  assign _EVAL_186 = _EVAL_453 == 1'h0;
  assign _EVAL_402 = {1'b0,$signed(_EVAL_485)};
  assign _EVAL_347 = $signed(_EVAL_402) & $signed(-33'sh8000);
  assign _EVAL_165 = $signed(_EVAL_347);
  assign _EVAL_460 = $signed(_EVAL_165) == $signed(33'sh0);
  assign _EVAL_123 = _EVAL_593 | _EVAL_32;
  assign _EVAL_115 = _EVAL_607 >> _EVAL_3;
  assign _EVAL_400 = _EVAL_115[0];
  assign _EVAL_444 = _EVAL_631 != _EVAL_66;
  assign _EVAL_446 = _EVAL_359 & _EVAL_47;
  assign _EVAL_414 = _EVAL_473 & _EVAL_160;
  assign _EVAL_511 = _EVAL_414 | _EVAL_151;
  assign _EVAL_392 = _EVAL_511 | _EVAL_32;
  assign _EVAL_436 = _EVAL_20 == _EVAL_203;
  assign _EVAL_438 = _EVAL_436 | _EVAL_32;
  assign _EVAL_608 = _EVAL_477 == 1'h0;
  assign _EVAL_451 = _EVAL_1 == 3'h6;
  assign _EVAL_117 = _EVAL_29 & _EVAL_451;
  assign _EVAL_104 = 4'h6 == _EVAL_31;
  assign _EVAL_404 = _EVAL_427 ? _EVAL_104 : 1'h0;
  assign _EVAL_641 = _EVAL_404 | _EVAL_32;
  assign _EVAL_640 = _EVAL_641 == 1'h0;
  assign _EVAL_312 = _EVAL_171 == 1'h0;
  assign _EVAL_514 = _EVAL_235 + 32'h1;
  assign _EVAL_499 = _EVAL_1 == 3'h7;
  assign _EVAL_513 = _EVAL_28 == 3'h7;
  assign _EVAL_345 = _EVAL_6 & _EVAL_513;
  assign _EVAL_494 = _EVAL_7 == _EVAL_605;
  assign _EVAL_259 = _EVAL_27 == 4'h0;
  assign _EVAL_395 = _EVAL_149 | _EVAL_259;
  assign _EVAL_275 = _EVAL_27[3:3];
  assign _EVAL_34 = _EVAL_275 == 1'h0;
  assign _EVAL_344 = _EVAL_34 & _EVAL_440;
  assign _EVAL_635 = _EVAL_395 | _EVAL_344;
  assign _EVAL_324 = _EVAL_37 - 5'h1;
  assign _EVAL_208 = _EVAL_413 - 5'h1;
  assign _EVAL_546 = _EVAL_138 & _EVAL_155;
  assign _EVAL_415 = _EVAL_196 | _EVAL_32;
  assign _EVAL_154 = _EVAL_415 == 1'h0;
  assign _EVAL_521 = _EVAL_176 | _EVAL_32;
  assign _EVAL_661 = _EVAL_521 == 1'h0;
  assign _EVAL_98 = _EVAL_337 | _EVAL_32;
  assign _EVAL_144 = _EVAL_98 == 1'h0;
  assign _EVAL_256 = _EVAL_393 >> _EVAL_27;
  assign _EVAL_261 = _EVAL_256[0];
  assign _EVAL_221 = _EVAL_261 | _EVAL_32;
  assign _EVAL_622 = _EVAL_221 == 1'h0;
  assign _EVAL_328 = _EVAL_1 == 3'h4;
  assign _EVAL_634 = _EVAL_28[0];
  assign _EVAL_219 = _EVAL_572[7:3];
  assign _EVAL_654 = _EVAL_1 == 3'h3;
  assign _EVAL_561 = _EVAL_10 & _EVAL_548;
  assign _EVAL_509 = _EVAL_635 | _EVAL_32;
  assign _EVAL_602 = _EVAL_670 | _EVAL_460;
  assign _EVAL_80 = _EVAL_494 | _EVAL_32;
  assign _EVAL_280 = $signed(_EVAL_143) & $signed(-33'sh2000);
  assign _EVAL_562 = $signed(_EVAL_280);
  assign _EVAL_93 = $signed(_EVAL_562) == $signed(33'sh0);
  assign _EVAL_524 = _EVAL_602 | _EVAL_93;
  assign _EVAL_307 = _EVAL_21 & _EVAL_6;
  assign _EVAL_187 = _EVAL_31 == _EVAL_297;
  assign _EVAL_310 = _EVAL_187 | _EVAL_32;
  assign _EVAL_403 = _EVAL_310 == 1'h0;
  assign _EVAL_430 = _EVAL_392 == 1'h0;
  assign _EVAL_389 = $signed(_EVAL_659);
  assign _EVAL_245 = $signed(_EVAL_389) == $signed(33'sh0);
  assign _EVAL_416 = _EVAL_524 | _EVAL_245;
  assign _EVAL_600 = _EVAL_416 | _EVAL_120;
  assign _EVAL_372 = _EVAL_316 - 5'h1;
  assign _EVAL_281 = _EVAL_467 | _EVAL_32;
  assign _EVAL_315 = _EVAL_400 == 1'h0;
  assign _EVAL_224 = _EVAL_315 | _EVAL_32;
  assign _EVAL_653 = _EVAL_469 == 1'h0;
  assign _EVAL_182 = _EVAL_217 & _EVAL_469;
  assign _EVAL_563 = _EVAL_19 == _EVAL_463;
  assign _EVAL_533 = _EVAL_9 == 2'h0;
  assign _EVAL_300 = _EVAL_19 <= 3'h3;
  assign _EVAL_63 = _EVAL_300 | _EVAL_32;
  assign _EVAL_146 = _EVAL_29 & _EVAL_527;
  assign _EVAL_466 = _EVAL_444 | _EVAL_158;
  assign _EVAL_169 = _EVAL_466 | _EVAL_32;
  assign _EVAL_478 = _EVAL_554 == 1'h0;
  assign _EVAL_318 = _EVAL_173 == 1'h0;
  assign _EVAL_294 = _EVAL_19 <= 3'h4;
  assign _EVAL_333 = _EVAL_600 | _EVAL_32;
  assign _EVAL_457 = _EVAL_333 == 1'h0;
  assign _EVAL_249 = _EVAL_456 == 1'h0;
  assign _EVAL_77 = _EVAL_281 == 1'h0;
  assign _EVAL_85 = _EVAL_169 == 1'h0;
  assign _EVAL_355 = _EVAL_509 == 1'h0;
  assign _EVAL_424 = _EVAL_533 | _EVAL_32;
  assign _EVAL_596 = _EVAL_424 == 1'h0;
  assign _EVAL_657 = _EVAL_306 == 1'h0;
  assign _EVAL_374 = _EVAL_29 & _EVAL_429;
  assign _EVAL_292 = _EVAL_159 | _EVAL_32;
  assign _EVAL_520 = _EVAL_292 == 1'h0;
  assign _EVAL_481 = _EVAL_251 == 1'h0;
  assign _EVAL_129 = _EVAL_114 == 1'h0;
  assign _EVAL_650 = _EVAL_459 | _EVAL_32;
  assign _EVAL_660 = _EVAL_650 == 1'h0;
  assign _EVAL_260 = _EVAL_438 == 1'h0;
  assign _EVAL_639 = _EVAL_6 & _EVAL_667;
  assign _EVAL_137 = _EVAL_1 == 3'h2;
  assign _EVAL_284 = _EVAL_563 | _EVAL_32;
  assign _EVAL_364 = _EVAL_284 == 1'h0;
  assign _EVAL_500 = _EVAL_101 == 1'h0;
  assign _EVAL_371 = _EVAL_615 == 1'h0;
  assign _EVAL_340 = _EVAL_11 == 3'h5;
  assign _EVAL_549 = _EVAL_10 & _EVAL_340;
  assign _EVAL_325 = _EVAL_294 | _EVAL_32;
  assign _EVAL_317 = _EVAL_10 & _EVAL_257;
  assign _EVAL_365 = _EVAL_29 & _EVAL_499;
  assign _EVAL_179 = _EVAL == _EVAL_518;
  assign _EVAL_629 = _EVAL_486 == 1'h0;
  assign _EVAL_320 = _EVAL_167 == 1'h0;
  assign _EVAL_127 = _EVAL_307 & _EVAL_532;
  assign _EVAL_266 = _EVAL_179 | _EVAL_32;
  assign _EVAL_243 = _EVAL_266 == 1'h0;
  assign _EVAL_97 = _EVAL_29 & _EVAL_328;
  assign _EVAL_577 = _EVAL_10 & _EVAL_645;
  assign _EVAL_139 = _EVAL_29 & _EVAL_653;
  assign _EVAL_583 = _EVAL_323 - 5'h1;
  assign _EVAL_302 = _EVAL_419 == 1'h0;
  assign _EVAL_87 = _EVAL_80 == 1'h0;
  assign _EVAL_71 = _EVAL_325 == 1'h0;
  assign _EVAL_447 = _EVAL_63 == 1'h0;
  assign _EVAL_632 = _EVAL_123 == 1'h0;
  assign _EVAL_45 = _EVAL_269 == 1'h0;
  assign _EVAL_250 = _EVAL_29 & _EVAL_654;
  assign _EVAL_422 = _EVAL_29 & _EVAL_503;
  assign _EVAL_298 = _EVAL_43 == 1'h0;
  assign _EVAL_188 = _EVAL_224 == 1'h0;
  assign _EVAL_331 = _EVAL_29 & _EVAL_137;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_37 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_168 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_201 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_203 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_235 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_278 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_283 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_297 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_316 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_323 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_351 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_360 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_369 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_406 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_407 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_413 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_435 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_442 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_463 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_464 = _RAND_19[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_470 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_474 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_518 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_557 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_587 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_605 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_607 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_628 = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_13) begin
    if (_EVAL_32) begin
      _EVAL_37 <= 5'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_388) begin
          if (_EVAL_619) begin
            _EVAL_37 <= _EVAL_578;
          end else begin
            _EVAL_37 <= 5'h0;
          end
        end else begin
          _EVAL_37 <= _EVAL_324;
        end
      end
    end
    if (_EVAL_182) begin
      _EVAL_168 <= _EVAL_1;
    end
    if (_EVAL_32) begin
      _EVAL_201 <= 5'h0;
    end else begin
      if (_EVAL_138) begin
        if (_EVAL_155) begin
          _EVAL_201 <= 5'h0;
        end else begin
          _EVAL_201 <= _EVAL_207;
        end
      end
    end
    if (_EVAL_546) begin
      _EVAL_203 <= _EVAL_20;
    end
    if (_EVAL_32) begin
      _EVAL_235 <= 32'h0;
    end else begin
      if (_EVAL_595) begin
        _EVAL_235 <= 32'h0;
      end else begin
        _EVAL_235 <= _EVAL_514;
      end
    end
    if (_EVAL_127) begin
      _EVAL_278 <= _EVAL_14;
    end
    if (_EVAL_127) begin
      _EVAL_283 <= _EVAL_30;
    end
    if (_EVAL_127) begin
      _EVAL_297 <= _EVAL_31;
    end
    if (_EVAL_32) begin
      _EVAL_316 <= 5'h0;
    end else begin
      if (_EVAL_217) begin
        if (_EVAL_225) begin
          if (_EVAL_83) begin
            _EVAL_316 <= _EVAL_472;
          end else begin
            _EVAL_316 <= 5'h0;
          end
        end else begin
          _EVAL_316 <= _EVAL_372;
        end
      end
    end
    if (_EVAL_32) begin
      _EVAL_323 <= 5'h0;
    end else begin
      if (_EVAL_307) begin
        if (_EVAL_532) begin
          if (_EVAL_634) begin
            _EVAL_323 <= _EVAL_219;
          end else begin
            _EVAL_323 <= 5'h0;
          end
        end else begin
          _EVAL_323 <= _EVAL_583;
        end
      end
    end
    if (_EVAL_586) begin
      _EVAL_351 <= _EVAL_24;
    end
    if (_EVAL_182) begin
      _EVAL_360 <= _EVAL_3;
    end
    if (_EVAL_586) begin
      _EVAL_369 <= _EVAL_9;
    end
    if (_EVAL_32) begin
      _EVAL_406 <= 5'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_484) begin
          if (_EVAL_619) begin
            _EVAL_406 <= _EVAL_578;
          end else begin
            _EVAL_406 <= 5'h0;
          end
        end else begin
          _EVAL_406 <= _EVAL_425;
        end
      end
    end
    if (_EVAL_586) begin
      _EVAL_407 <= _EVAL_26;
    end
    if (_EVAL_32) begin
      _EVAL_413 <= 5'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_305) begin
          if (_EVAL_619) begin
            _EVAL_413 <= _EVAL_578;
          end else begin
            _EVAL_413 <= 5'h0;
          end
        end else begin
          _EVAL_413 <= _EVAL_208;
        end
      end
    end
    if (_EVAL_127) begin
      _EVAL_435 <= _EVAL_18;
    end
    if (_EVAL_32) begin
      _EVAL_442 <= 5'h0;
    end else begin
      if (_EVAL_217) begin
        if (_EVAL_469) begin
          if (_EVAL_83) begin
            _EVAL_442 <= _EVAL_472;
          end else begin
            _EVAL_442 <= 5'h0;
          end
        end else begin
          _EVAL_442 <= _EVAL_184;
        end
      end
    end
    if (_EVAL_182) begin
      _EVAL_463 <= _EVAL_19;
    end
    if (_EVAL_586) begin
      _EVAL_464 <= _EVAL_27;
    end
    if (_EVAL_32) begin
      _EVAL_470 <= 2'h0;
    end else begin
      _EVAL_470 <= _EVAL_446;
    end
    if (_EVAL_586) begin
      _EVAL_474 <= _EVAL_11;
    end
    if (_EVAL_586) begin
      _EVAL_518 <= _EVAL;
    end
    if (_EVAL_127) begin
      _EVAL_557 <= _EVAL_28;
    end
    if (_EVAL_182) begin
      _EVAL_587 <= _EVAL_0;
    end
    if (_EVAL_546) begin
      _EVAL_605 <= _EVAL_7;
    end
    if (_EVAL_32) begin
      _EVAL_607 <= 9'h0;
    end else begin
      _EVAL_607 <= _EVAL_580;
    end
    if (_EVAL_182) begin
      _EVAL_628 <= _EVAL_15;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_660) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07709a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74f6c6db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a78a0371)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bee9e888)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_403) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5faa636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_481) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bcf1293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_661) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79d60916)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6026c1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_481) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e8828f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_620) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41816eae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(193f5604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dc85f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_660) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5303c13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d651fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b10069b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_655) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(318f0f06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e139a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_629) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29e6f0d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_596) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_609) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_660) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5366c7c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_481) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_497) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_596) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f17260e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_547) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54b1f283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d741591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_661) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_430) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_596) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f79d51e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b154c9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_596) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca25a84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8a63c9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6514abd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dd2dd8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_648) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b18defb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_608) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da9d20d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_666) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4bca6e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_320) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6af1682a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_536) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9fc6024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_655) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ff9add)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e60c077)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2640c93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_336) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e42e854d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_648) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9062184a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(330dd068)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_336) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_445) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d821994a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ddfb83d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e29064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(533b38c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5038b5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d2009bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9039e6e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_488) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_625 & _EVAL_622) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ee41bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_445) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_661) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beb89e39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f0cd124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_620) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50861b1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_478) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5d63e7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e3ca7b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_420) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af86018)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_420) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(926e7cef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9f72d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_481) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(680a82c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_588) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cc5fbe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_495) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_588) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2562ae46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fdff968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8971637c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f09f371)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_497) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1697b0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8c47bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_640) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dae5588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_430) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b76a9529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9677efdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edf0a3cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e0fa88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_640) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_371) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d031d3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_495) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e899e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_661) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b953d64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bbd16b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_520) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(320a1b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_445) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_447) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_320) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_488) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0019ce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf525092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_623) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_547) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80716266)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_661) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0298b7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_596) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b8a02f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_420) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_596) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(897f1ded)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_349) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1918b8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea8e9a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_660) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d26e1c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_478) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43c9da5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_623) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d410849c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_588) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e6366d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec7e481e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_666) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f70e26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27bfea60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_625 & _EVAL_622) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_430) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f118fa15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_588) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b666d14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_495) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e5f3f01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_371) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba6623c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_640) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c368c3ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_648) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_447) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1ba89d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a456deba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fce64991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_547) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_648) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ead679)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c24a7c0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_620) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(280bb58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93ceef1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_349) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd559709)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_657) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81a2c49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(867d1b09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(552480c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e89ce957)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c8b3b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2337c61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e6d2257)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31e27270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d5c73d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_536) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c36ce2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_403) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_661) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cba465d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_588) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c20c3c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_445) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17697d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_547) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_371) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380b9f6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f550495a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_608) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b92c16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_648) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(772edca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_596) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_520) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(814162a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a935eae5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_430) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d3142d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_596) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_640) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_500) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e906ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_648) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_500) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30d300e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_588) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c14686f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_420) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd09bc2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_495) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7d56945)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34441912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e183671a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2e908c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c98e128e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_620) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_592) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8532fc03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_609) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a2319b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_592) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7244ebae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_629) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_430) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_613) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6f4884b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_430) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d33498c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(155af4e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_371) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b64be954)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_657) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28630975)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
