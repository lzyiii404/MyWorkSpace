//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_134_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [25:0] _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [6:0]  _EVAL_13,
  input  [6:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_18;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_45;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_72;
  reg [31:0] _RAND_2;
  reg [72:0] _EVAL_112;
  reg [95:0] _RAND_3;
  reg [2:0] _EVAL_153;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_156;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_197;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_212;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_213;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_215;
  reg [31:0] _RAND_9;
  reg [6:0] _EVAL_222;
  reg [31:0] _RAND_10;
  reg [6:0] _EVAL_226;
  reg [31:0] _RAND_11;
  reg [25:0] _EVAL_250;
  reg [31:0] _RAND_12;
  reg [3:0] _EVAL_262;
  reg [31:0] _RAND_13;
  wire  _EVAL_155;
  wire  _EVAL_259;
  wire  _EVAL_141;
  wire  _EVAL_267;
  wire  _EVAL_118;
  wire  _EVAL_192;
  wire  _EVAL_264;
  wire  _EVAL_60;
  wire [3:0] _EVAL_274;
  wire  _EVAL_201;
  wire [1:0] _EVAL_126;
  wire [1:0] _EVAL_16;
  wire  _EVAL_19;
  wire  _EVAL_239;
  wire  _EVAL_122;
  wire  _EVAL_158;
  wire [3:0] _EVAL_268;
  wire  _EVAL_91;
  wire  _EVAL_234;
  wire [3:0] _EVAL_70;
  wire  _EVAL_20;
  wire  _EVAL_140;
  wire  _EVAL_245;
  wire  _EVAL_49;
  wire  _EVAL_261;
  wire  _EVAL_177;
  wire [3:0] _EVAL_196;
  wire  _EVAL_58;
  wire [2:0] _EVAL_164;
  wire  _EVAL_179;
  wire  _EVAL_251;
  wire  _EVAL_223;
  wire  _EVAL_199;
  wire  _EVAL_195;
  wire  _EVAL_38;
  wire  _EVAL_131;
  wire  _EVAL_152;
  wire  _EVAL_186;
  wire  _EVAL_260;
  wire  _EVAL_54;
  wire  _EVAL_257;
  wire  _EVAL_147;
  wire  _EVAL_92;
  wire  _EVAL_28;
  wire  _EVAL_182;
  wire  _EVAL_129;
  wire  _EVAL_144;
  wire  _EVAL_79;
  wire [127:0] _EVAL_178;
  wire [127:0] _EVAL_273;
  wire [72:0] _EVAL_145;
  wire [72:0] _EVAL_138;
  wire [72:0] _EVAL_214;
  wire  _EVAL_76;
  wire  _EVAL_66;
  wire  _EVAL_189;
  wire [12:0] _EVAL_105;
  wire [31:0] _EVAL_256;
  wire  _EVAL_143;
  wire  _EVAL_89;
  wire  _EVAL_163;
  wire  _EVAL_123;
  wire  _EVAL_31;
  wire  _EVAL_26;
  wire  _EVAL_104;
  wire  _EVAL_90;
  wire  _EVAL_77;
  wire  _EVAL_24;
  wire  _EVAL_94;
  wire  _EVAL_108;
  wire  _EVAL_208;
  wire  _EVAL_229;
  wire  _EVAL_73;
  wire  _EVAL_50;
  wire  _EVAL_40;
  wire  _EVAL_210;
  wire [2:0] _EVAL_238;
  wire  _EVAL_148;
  wire  _EVAL_278;
  wire [5:0] _EVAL_282;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_67;
  wire  _EVAL_252;
  wire  _EVAL_151;
  wire [12:0] _EVAL_249;
  wire [5:0] _EVAL_279;
  wire [5:0] _EVAL_146;
  wire [3:0] _EVAL_231;
  wire  _EVAL_246;
  wire  _EVAL_181;
  wire  _EVAL_188;
  wire  _EVAL_42;
  wire  _EVAL_27;
  wire  _EVAL_217;
  wire  _EVAL_87;
  wire  _EVAL_132;
  wire  _EVAL_110;
  wire  _EVAL_220;
  wire  _EVAL_206;
  wire  _EVAL_63;
  wire  _EVAL_173;
  wire  _EVAL_106;
  wire  _EVAL_183;
  wire  _EVAL_198;
  wire  _EVAL_254;
  wire  _EVAL_221;
  wire  _EVAL_228;
  wire  _EVAL_81;
  wire  _EVAL_205;
  wire  _EVAL_175;
  wire  _EVAL_17;
  wire [127:0] _EVAL_133;
  wire [127:0] _EVAL_265;
  wire [72:0] _EVAL_275;
  wire [72:0] _EVAL_136;
  wire  _EVAL_244;
  wire  _EVAL_117;
  wire [3:0] _EVAL_51;
  wire  _EVAL_237;
  wire  _EVAL_53;
  wire  _EVAL_211;
  wire  _EVAL_241;
  wire  _EVAL_95;
  wire  _EVAL_193;
  wire  _EVAL_232;
  wire  _EVAL_224;
  wire  _EVAL_52;
  wire  _EVAL_47;
  wire  _EVAL_167;
  wire  _EVAL_22;
  wire  _EVAL_266;
  wire  _EVAL_187;
  wire  _EVAL_41;
  wire  _EVAL_124;
  wire  _EVAL_101;
  wire  _EVAL_154;
  wire  _EVAL_82;
  wire  _EVAL_15;
  wire  _EVAL_21;
  wire  _EVAL_174;
  wire [3:0] _EVAL_64;
  wire  _EVAL_281;
  wire  _EVAL_37;
  wire [25:0] _EVAL_99;
  wire [26:0] _EVAL_243;
  wire [26:0] _EVAL_159;
  wire [26:0] _EVAL_277;
  wire  _EVAL_227;
  wire  _EVAL_34;
  wire  _EVAL_65;
  wire  _EVAL_236;
  wire  _EVAL_130;
  wire  _EVAL_253;
  wire  _EVAL_242;
  wire  _EVAL_48;
  wire  _EVAL_71;
  wire  _EVAL_46;
  wire  _EVAL_233;
  wire  _EVAL_98;
  wire [5:0] _EVAL_113;
  wire  _EVAL_230;
  wire  _EVAL_209;
  wire  _EVAL_202;
  wire  _EVAL_235;
  wire  _EVAL_184;
  wire  _EVAL_134;
  wire  _EVAL_30;
  wire [3:0] _EVAL_125;
  wire [3:0] _EVAL_119;
  wire  _EVAL_190;
  wire  _EVAL_35;
  wire [3:0] _EVAL_57;
  wire [72:0] _EVAL_172;
  wire  _EVAL_137;
  wire  _EVAL_165;
  wire  _EVAL_102;
  wire  _EVAL_255;
  wire  _EVAL_218;
  wire  _EVAL_116;
  wire  _EVAL_109;
  wire [25:0] _EVAL_160;
  wire [25:0] _EVAL_62;
  wire  _EVAL_150;
  wire  _EVAL_142;
  wire [3:0] _EVAL_162;
  wire [3:0] _EVAL_139;
  wire  _EVAL_135;
  wire  _EVAL_127;
  wire  _EVAL_29;
  wire  _EVAL_93;
  wire  _EVAL_200;
  wire  _EVAL_59;
  wire  _EVAL_225;
  wire  _EVAL_107;
  wire  _EVAL_43;
  wire  _EVAL_86;
  wire  _EVAL_161;
  wire  _EVAL_114;
  wire  _EVAL_276;
  wire  _EVAL_55;
  wire  _EVAL_84;
  wire  _EVAL_120;
  wire  _EVAL_269;
  wire  _EVAL_111;
  wire  _EVAL_194;
  wire  _EVAL_169;
  wire  _EVAL_23;
  wire  _EVAL_216;
  wire  _EVAL_240;
  wire  _EVAL_149;
  wire  _EVAL_36;
  wire  _EVAL_263;
  wire  _EVAL_248;
  wire  _EVAL_168;
  wire  _EVAL_280;
  wire  _EVAL_170;
  wire  _EVAL_25;
  wire  _EVAL_157;
  wire  _EVAL_258;
  wire [72:0] _EVAL_61;
  wire [72:0] _EVAL_128;
  wire  _EVAL_272;
  wire  _EVAL_83;
  wire  _EVAL_68;
  wire  _EVAL_96;
  wire  _EVAL_33;
  wire  _EVAL_185;
  wire  _EVAL_85;
  wire  _EVAL_191;
  wire  _EVAL_121;
  wire  _EVAL_69;
  wire  _EVAL_80;
  wire  _EVAL_219;
  wire  _EVAL_166;
  wire  _EVAL_207;
  wire  _EVAL_56;
  wire  _EVAL_39;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_155 = _EVAL_0 >= 3'h2;
  assign _EVAL_259 = _EVAL_155 | _EVAL_3;
  assign _EVAL_141 = _EVAL_259 == 1'h0;
  assign _EVAL_267 = _EVAL_13 == _EVAL_222;
  assign _EVAL_118 = _EVAL_267 | _EVAL_3;
  assign _EVAL_192 = _EVAL_7 == 3'h0;
  assign _EVAL_264 = _EVAL_192 | _EVAL_3;
  assign _EVAL_60 = _EVAL_264 == 1'h0;
  assign _EVAL_274 = _EVAL_262 - 4'h1;
  assign _EVAL_201 = _EVAL_2[0];
  assign _EVAL_126 = 2'h1 << _EVAL_201;
  assign _EVAL_16 = _EVAL_126 | 2'h1;
  assign _EVAL_19 = _EVAL_16[1];
  assign _EVAL_239 = _EVAL_10[1];
  assign _EVAL_122 = _EVAL_239 == 1'h0;
  assign _EVAL_158 = _EVAL_19 & _EVAL_122;
  assign _EVAL_268 = _EVAL_13[6:3];
  assign _EVAL_91 = _EVAL_268 == 4'h2;
  assign _EVAL_234 = _EVAL_5 == 3'h6;
  assign _EVAL_70 = ~ _EVAL_12;
  assign _EVAL_20 = _EVAL_70 == 4'h0;
  assign _EVAL_140 = _EVAL_20 | _EVAL_3;
  assign _EVAL_245 = _EVAL_140 == 1'h0;
  assign _EVAL_49 = _EVAL_14 == 7'h48;
  assign _EVAL_261 = _EVAL_14 == 7'h40;
  assign _EVAL_177 = _EVAL_49 | _EVAL_261;
  assign _EVAL_196 = _EVAL_14[6:3];
  assign _EVAL_58 = _EVAL_196 == 4'h8;
  assign _EVAL_164 = _EVAL_14[2:0];
  assign _EVAL_179 = 3'h1 <= _EVAL_164;
  assign _EVAL_251 = _EVAL_58 & _EVAL_179;
  assign _EVAL_223 = _EVAL_177 | _EVAL_251;
  assign _EVAL_199 = _EVAL_14 == 7'h20;
  assign _EVAL_195 = _EVAL_223 | _EVAL_199;
  assign _EVAL_38 = _EVAL_196 == 4'h0;
  assign _EVAL_131 = _EVAL_195 | _EVAL_38;
  assign _EVAL_152 = _EVAL_196 == 4'h1;
  assign _EVAL_186 = _EVAL_131 | _EVAL_152;
  assign _EVAL_260 = _EVAL_196 == 4'h2;
  assign _EVAL_54 = _EVAL_186 | _EVAL_260;
  assign _EVAL_257 = _EVAL_196 == 4'h3;
  assign _EVAL_147 = _EVAL_54 | _EVAL_257;
  assign _EVAL_92 = _EVAL_7 != 3'h0;
  assign _EVAL_28 = _EVAL_92 | _EVAL_3;
  assign _EVAL_182 = _EVAL_28 == 1'h0;
  assign _EVAL_129 = _EVAL_6 & _EVAL_11;
  assign _EVAL_144 = _EVAL_18 == 4'h0;
  assign _EVAL_79 = _EVAL_129 & _EVAL_144;
  assign _EVAL_178 = 128'h1 << _EVAL_14;
  assign _EVAL_273 = _EVAL_79 ? _EVAL_178 : 128'h0;
  assign _EVAL_145 = _EVAL_273[72:0];
  assign _EVAL_138 = _EVAL_145 | _EVAL_112;
  assign _EVAL_214 = _EVAL_138 >> _EVAL_13;
  assign _EVAL_76 = _EVAL_72 == 4'h0;
  assign _EVAL_66 = _EVAL_7 <= 3'h2;
  assign _EVAL_189 = _EVAL_234 == 1'h0;
  assign _EVAL_105 = 13'h3f << _EVAL_2;
  assign _EVAL_256 = _EVAL_45 + 32'h1;
  assign _EVAL_143 = _EVAL_0 == _EVAL_215;
  assign _EVAL_89 = _EVAL_143 | _EVAL_3;
  assign _EVAL_163 = _EVAL_89 == 1'h0;
  assign _EVAL_123 = _EVAL_1 == 3'h2;
  assign _EVAL_31 = _EVAL_16[0];
  assign _EVAL_26 = _EVAL_10[0];
  assign _EVAL_104 = _EVAL_239 & _EVAL_26;
  assign _EVAL_90 = _EVAL_31 & _EVAL_104;
  assign _EVAL_77 = _EVAL_13 == 7'h20;
  assign _EVAL_24 = _EVAL_5 == 3'h2;
  assign _EVAL_94 = _EVAL_7 <= 3'h4;
  assign _EVAL_108 = _EVAL_156 == 4'h0;
  assign _EVAL_208 = _EVAL_108 == 1'h0;
  assign _EVAL_229 = _EVAL & _EVAL_208;
  assign _EVAL_73 = 3'h6 == _EVAL_2;
  assign _EVAL_50 = _EVAL_261 ? _EVAL_73 : 1'h0;
  assign _EVAL_40 = _EVAL_2 >= 3'h2;
  assign _EVAL_210 = _EVAL_268 == 4'h8;
  assign _EVAL_238 = _EVAL_13[2:0];
  assign _EVAL_148 = 3'h1 <= _EVAL_238;
  assign _EVAL_278 = _EVAL_210 & _EVAL_148;
  assign _EVAL_282 = _EVAL_105[5:0];
  assign _EVAL_74 = _EVAL_7 == _EVAL_212;
  assign _EVAL_75 = _EVAL_74 | _EVAL_3;
  assign _EVAL_67 = _EVAL_75 == 1'h0;
  assign _EVAL_252 = _EVAL_13 == 7'h40;
  assign _EVAL_151 = _EVAL_9 == 1'h0;
  assign _EVAL_249 = 13'h3f << _EVAL_0;
  assign _EVAL_279 = _EVAL_249[5:0];
  assign _EVAL_146 = ~ _EVAL_279;
  assign _EVAL_231 = _EVAL_146[5:2];
  assign _EVAL_246 = _EVAL_1 == 3'h5;
  assign _EVAL_181 = _EVAL_13 == 7'h48;
  assign _EVAL_188 = _EVAL_181 | _EVAL_252;
  assign _EVAL_42 = _EVAL_188 | _EVAL_278;
  assign _EVAL_27 = _EVAL_42 | _EVAL_77;
  assign _EVAL_217 = _EVAL_268 == 4'h0;
  assign _EVAL_87 = _EVAL_27 | _EVAL_217;
  assign _EVAL_132 = _EVAL_268 == 4'h1;
  assign _EVAL_110 = _EVAL_87 | _EVAL_132;
  assign _EVAL_220 = _EVAL_110 | _EVAL_91;
  assign _EVAL_206 = _EVAL_268 == 4'h3;
  assign _EVAL_63 = _EVAL_220 | _EVAL_206;
  assign _EVAL_173 = _EVAL_63 | _EVAL_3;
  assign _EVAL_106 = _EVAL_173 == 1'h0;
  assign _EVAL_183 = _EVAL_1 == 3'h6;
  assign _EVAL_198 = _EVAL_50 | _EVAL_3;
  assign _EVAL_254 = _EVAL_5 == _EVAL_197;
  assign _EVAL_221 = _EVAL_254 | _EVAL_3;
  assign _EVAL_228 = _EVAL_221 == 1'h0;
  assign _EVAL_81 = _EVAL_1 == 3'h1;
  assign _EVAL_205 = _EVAL_8 & _EVAL;
  assign _EVAL_175 = _EVAL_205 & _EVAL_76;
  assign _EVAL_17 = _EVAL_175 & _EVAL_189;
  assign _EVAL_133 = 128'h1 << _EVAL_13;
  assign _EVAL_265 = _EVAL_17 ? _EVAL_133 : 128'h0;
  assign _EVAL_275 = _EVAL_265[72:0];
  assign _EVAL_136 = ~ _EVAL_275;
  assign _EVAL_244 = _EVAL_2 == _EVAL_153;
  assign _EVAL_117 = _EVAL_5[0];
  assign _EVAL_51 = _EVAL_72 - 4'h1;
  assign _EVAL_237 = _EVAL_112 != 73'h0;
  assign _EVAL_53 = _EVAL_237 == 1'h0;
  assign _EVAL_211 = plusarg_reader_out == 32'h0;
  assign _EVAL_241 = _EVAL_53 | _EVAL_211;
  assign _EVAL_95 = _EVAL_45 < plusarg_reader_out;
  assign _EVAL_193 = _EVAL_241 | _EVAL_95;
  assign _EVAL_232 = _EVAL_19 & _EVAL_239;
  assign _EVAL_224 = _EVAL_193 | _EVAL_3;
  assign _EVAL_52 = _EVAL_224 == 1'h0;
  assign _EVAL_47 = _EVAL_40 | _EVAL_232;
  assign _EVAL_167 = _EVAL_47 | _EVAL_90;
  assign _EVAL_22 = _EVAL_26 == 1'h0;
  assign _EVAL_266 = _EVAL_239 & _EVAL_22;
  assign _EVAL_187 = _EVAL_31 & _EVAL_266;
  assign _EVAL_41 = _EVAL_47 | _EVAL_187;
  assign _EVAL_124 = _EVAL_40 | _EVAL_158;
  assign _EVAL_101 = _EVAL_122 & _EVAL_26;
  assign _EVAL_154 = _EVAL_31 & _EVAL_101;
  assign _EVAL_82 = _EVAL_124 | _EVAL_154;
  assign _EVAL_15 = _EVAL_122 & _EVAL_22;
  assign _EVAL_21 = _EVAL_31 & _EVAL_15;
  assign _EVAL_174 = _EVAL_124 | _EVAL_21;
  assign _EVAL_64 = {_EVAL_167,_EVAL_41,_EVAL_82,_EVAL_174};
  assign _EVAL_281 = _EVAL_12 == _EVAL_64;
  assign _EVAL_37 = _EVAL_2 <= 3'h6;
  assign _EVAL_99 = _EVAL_10 ^ 26'h2000000;
  assign _EVAL_243 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_159 = $signed(_EVAL_243) & $signed(-27'sh10000);
  assign _EVAL_277 = $signed(_EVAL_159);
  assign _EVAL_227 = $signed(_EVAL_277) == $signed(27'sh0);
  assign _EVAL_34 = _EVAL_37 & _EVAL_227;
  assign _EVAL_65 = _EVAL_34 | _EVAL_3;
  assign _EVAL_236 = _EVAL_65 == 1'h0;
  assign _EVAL_130 = _EVAL_1 == 3'h7;
  assign _EVAL_253 = _EVAL_1 == 3'h4;
  assign _EVAL_242 = _EVAL_5 == 3'h1;
  assign _EVAL_48 = _EVAL & _EVAL_242;
  assign _EVAL_71 = _EVAL_5 <= 3'h6;
  assign _EVAL_46 = _EVAL_71 | _EVAL_3;
  assign _EVAL_233 = _EVAL_46 == 1'h0;
  assign _EVAL_98 = _EVAL_151 | _EVAL_3;
  assign _EVAL_113 = ~ _EVAL_282;
  assign _EVAL_230 = _EVAL_198 == 1'h0;
  assign _EVAL_209 = _EVAL & _EVAL_234;
  assign _EVAL_202 = _EVAL_129 | _EVAL_205;
  assign _EVAL_235 = _EVAL & _EVAL_24;
  assign _EVAL_184 = _EVAL_94 | _EVAL_3;
  assign _EVAL_134 = _EVAL_1[2];
  assign _EVAL_30 = _EVAL_134 == 1'h0;
  assign _EVAL_125 = _EVAL_113[5:2];
  assign _EVAL_119 = _EVAL_18 - 4'h1;
  assign _EVAL_190 = _EVAL_184 == 1'h0;
  assign _EVAL_35 = _EVAL_3 == 1'h0;
  assign _EVAL_57 = _EVAL_156 - 4'h1;
  assign _EVAL_172 = _EVAL_112 >> _EVAL_14;
  assign _EVAL_137 = _EVAL_262 == 4'h0;
  assign _EVAL_165 = _EVAL_129 & _EVAL_137;
  assign _EVAL_102 = _EVAL_5 == 3'h0;
  assign _EVAL_255 = _EVAL & _EVAL_102;
  assign _EVAL_218 = _EVAL_214[0];
  assign _EVAL_116 = _EVAL_281 | _EVAL_3;
  assign _EVAL_109 = _EVAL_116 == 1'h0;
  assign _EVAL_160 = {{20'd0}, _EVAL_113};
  assign _EVAL_62 = _EVAL_10 & _EVAL_160;
  assign _EVAL_150 = _EVAL_62 == 26'h0;
  assign _EVAL_142 = _EVAL_150 | _EVAL_3;
  assign _EVAL_162 = ~ _EVAL_64;
  assign _EVAL_139 = _EVAL_12 & _EVAL_162;
  assign _EVAL_135 = _EVAL_137 == 1'h0;
  assign _EVAL_127 = _EVAL_11 & _EVAL_135;
  assign _EVAL_29 = _EVAL_11 & _EVAL_246;
  assign _EVAL_93 = _EVAL_14 == _EVAL_226;
  assign _EVAL_200 = _EVAL_1 == 3'h0;
  assign _EVAL_59 = _EVAL_11 & _EVAL_200;
  assign _EVAL_225 = _EVAL_11 & _EVAL_183;
  assign _EVAL_107 = _EVAL_139 == 4'h0;
  assign _EVAL_43 = _EVAL_107 | _EVAL_3;
  assign _EVAL_86 = _EVAL_172[0];
  assign _EVAL_161 = _EVAL_66 | _EVAL_3;
  assign _EVAL_114 = _EVAL_10 == _EVAL_250;
  assign _EVAL_276 = _EVAL_7 <= 3'h3;
  assign _EVAL_55 = _EVAL_161 == 1'h0;
  assign _EVAL_84 = _EVAL_5 == 3'h4;
  assign _EVAL_120 = _EVAL_40 | _EVAL_3;
  assign _EVAL_269 = _EVAL_142 == 1'h0;
  assign _EVAL_111 = _EVAL_86 == 1'h0;
  assign _EVAL_194 = _EVAL_111 | _EVAL_3;
  assign _EVAL_169 = _EVAL_276 | _EVAL_3;
  assign _EVAL_23 = _EVAL_194 == 1'h0;
  assign _EVAL_216 = _EVAL_120 == 1'h0;
  assign _EVAL_240 = _EVAL_114 | _EVAL_3;
  assign _EVAL_149 = _EVAL_240 == 1'h0;
  assign _EVAL_36 = _EVAL_147 | _EVAL_3;
  assign _EVAL_263 = _EVAL_11 & _EVAL_130;
  assign _EVAL_248 = _EVAL_93 | _EVAL_3;
  assign _EVAL_168 = _EVAL_248 == 1'h0;
  assign _EVAL_280 = _EVAL_36 == 1'h0;
  assign _EVAL_170 = _EVAL_118 == 1'h0;
  assign _EVAL_25 = _EVAL_1 == 3'h3;
  assign _EVAL_157 = _EVAL_1 == _EVAL_213;
  assign _EVAL_258 = _EVAL_205 & _EVAL_108;
  assign _EVAL_61 = _EVAL_112 | _EVAL_145;
  assign _EVAL_128 = _EVAL_61 & _EVAL_136;
  assign _EVAL_272 = _EVAL_11 & _EVAL_123;
  assign _EVAL_83 = _EVAL_169 == 1'h0;
  assign _EVAL_68 = _EVAL_218 | _EVAL_3;
  assign _EVAL_96 = _EVAL_68 == 1'h0;
  assign _EVAL_33 = _EVAL_43 == 1'h0;
  assign _EVAL_185 = _EVAL_98 == 1'h0;
  assign _EVAL_85 = _EVAL_244 | _EVAL_3;
  assign _EVAL_191 = _EVAL_85 == 1'h0;
  assign _EVAL_121 = _EVAL_157 | _EVAL_3;
  assign _EVAL_69 = _EVAL_121 == 1'h0;
  assign _EVAL_80 = _EVAL_5 == 3'h5;
  assign _EVAL_219 = _EVAL_11 & _EVAL_25;
  assign _EVAL_166 = _EVAL & _EVAL_84;
  assign _EVAL_207 = _EVAL_11 & _EVAL_253;
  assign _EVAL_56 = _EVAL & _EVAL_80;
  assign _EVAL_39 = _EVAL_11 & _EVAL_81;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_18 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_45 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_72 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  _EVAL_112 = _RAND_3[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_153 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_156 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_197 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_212 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_213 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_215 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_222 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_226 = _RAND_11[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_250 = _RAND_12[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_262 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_3) begin
      _EVAL_18 <= 4'h0;
    end else begin
      if (_EVAL_129) begin
        if (_EVAL_144) begin
          if (_EVAL_30) begin
            _EVAL_18 <= _EVAL_125;
          end else begin
            _EVAL_18 <= 4'h0;
          end
        end else begin
          _EVAL_18 <= _EVAL_119;
        end
      end
    end
    if (_EVAL_3) begin
      _EVAL_45 <= 32'h0;
    end else begin
      if (_EVAL_202) begin
        _EVAL_45 <= 32'h0;
      end else begin
        _EVAL_45 <= _EVAL_256;
      end
    end
    if (_EVAL_3) begin
      _EVAL_72 <= 4'h0;
    end else begin
      if (_EVAL_205) begin
        if (_EVAL_76) begin
          if (_EVAL_117) begin
            _EVAL_72 <= _EVAL_231;
          end else begin
            _EVAL_72 <= 4'h0;
          end
        end else begin
          _EVAL_72 <= _EVAL_51;
        end
      end
    end
    if (_EVAL_3) begin
      _EVAL_112 <= 73'h0;
    end else begin
      _EVAL_112 <= _EVAL_128;
    end
    if (_EVAL_165) begin
      _EVAL_153 <= _EVAL_2;
    end
    if (_EVAL_3) begin
      _EVAL_156 <= 4'h0;
    end else begin
      if (_EVAL_205) begin
        if (_EVAL_108) begin
          if (_EVAL_117) begin
            _EVAL_156 <= _EVAL_231;
          end else begin
            _EVAL_156 <= 4'h0;
          end
        end else begin
          _EVAL_156 <= _EVAL_57;
        end
      end
    end
    if (_EVAL_258) begin
      _EVAL_197 <= _EVAL_5;
    end
    if (_EVAL_165) begin
      _EVAL_212 <= _EVAL_7;
    end
    if (_EVAL_165) begin
      _EVAL_213 <= _EVAL_1;
    end
    if (_EVAL_258) begin
      _EVAL_215 <= _EVAL_0;
    end
    if (_EVAL_258) begin
      _EVAL_222 <= _EVAL_13;
    end
    if (_EVAL_165) begin
      _EVAL_226 <= _EVAL_14;
    end
    if (_EVAL_165) begin
      _EVAL_250 <= _EVAL_10;
    end
    if (_EVAL_3) begin
      _EVAL_262 <= 4'h0;
    end else begin
      if (_EVAL_129) begin
        if (_EVAL_137) begin
          if (_EVAL_30) begin
            _EVAL_262 <= _EVAL_125;
          end else begin
            _EVAL_262 <= 4'h0;
          end
        end else begin
          _EVAL_262 <= _EVAL_274;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48cadb78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1dca7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daa2611a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c87e887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84b6535b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72c9fd57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b2c46b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d456cecb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5773f769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aa4f6de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b99217ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6c4337f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eab4ea1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f29d434)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc78c402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ddc981f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc011b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a6a99c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(750fda10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(116cc29a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0e7055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3779ed6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd9dbfae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d17ce97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18cf13a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14df7a30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9e2e26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c326347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc3c8216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3160d7ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef184c5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3a65f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25255f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7935dc35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(538d1f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea6a619c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(683d725c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c6b6d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db98b04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d2ad7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(deee5e90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81be8d03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76d5faeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58e3b918)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e1e110)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f147c180)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b62a51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f0900d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1256d84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32129a5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b4ea8f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1af1cada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44b76b8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4b1fe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f0c7a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c2b1c8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae36b963)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(159f3672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ddbb342)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e78bf84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58244ae9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d47e59ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d528aee4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdfd81f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee5213f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bd7cc7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82907d53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da31c85f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d70d53c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(216459b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f14dd19c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
