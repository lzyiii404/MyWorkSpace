//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_179(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  output [3:0]  _EVAL_3,
  output [1:0]  _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  output [3:0]  _EVAL_9,
  input  [6:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  output        _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output [29:0] _EVAL_17,
  input         _EVAL_18,
  output [2:0]  _EVAL_19,
  input  [3:0]  _EVAL_20,
  output [6:0]  _EVAL_21,
  output        _EVAL_22,
  input  [3:0]  _EVAL_23,
  output        _EVAL_24,
  input  [6:0]  _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  output [31:0] _EVAL_28,
  input  [31:0] _EVAL_29,
  output [6:0]  _EVAL_30,
  input  [29:0] _EVAL_31,
  output [31:0] _EVAL_32,
  output        _EVAL_33,
  output [3:0]  _EVAL_34,
  input  [2:0]  _EVAL_35,
  input         _EVAL_36,
  output [2:0]  _EVAL_37,
  output [2:0]  _EVAL_38,
  input         _EVAL_39,
  output        _EVAL_40
);
  assign _EVAL_28 = _EVAL_29;
  assign _EVAL_34 = _EVAL_23;
  assign _EVAL_3 = _EVAL_7;
  assign _EVAL_22 = _EVAL_0;
  assign _EVAL_33 = _EVAL_14;
  assign _EVAL_21 = _EVAL_10;
  assign _EVAL_32 = _EVAL_13;
  assign _EVAL_37 = _EVAL;
  assign _EVAL_12 = _EVAL_8;
  assign _EVAL_38 = _EVAL_11;
  assign _EVAL_16 = _EVAL_1;
  assign _EVAL_26 = _EVAL_39;
  assign _EVAL_4 = _EVAL_2;
  assign _EVAL_9 = _EVAL_20;
  assign _EVAL_5 = _EVAL_18;
  assign _EVAL_40 = _EVAL_36;
  assign _EVAL_24 = _EVAL_6;
  assign _EVAL_30 = _EVAL_25;
  assign _EVAL_19 = _EVAL_35;
  assign _EVAL_17 = _EVAL_31;
endmodule
