//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_17(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  output [2:0]  _EVAL_1,
  input  [63:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output [63:0] _EVAL_5,
  output [1:0]  _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [31:0] _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output [1:0]  _EVAL_14,
  output [1:0]  _EVAL_15,
  output [1:0]  _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [63:0] _EVAL_20,
  output [31:0] _EVAL_21,
  input  [2:0]  _EVAL_22,
  input  [3:0]  _EVAL_23,
  input  [3:0]  _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  output [63:0] _EVAL_27,
  input  [1:0]  _EVAL_28,
  input  [1:0]  _EVAL_29,
  input  [1:0]  _EVAL_30,
  input         _EVAL_31,
  output [2:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input  [3:0]  _EVAL_34,
  input  [2:0]  _EVAL_35,
  input  [2:0]  _EVAL_36,
  output        _EVAL_37,
  input         _EVAL_38,
  output [1:0]  _EVAL_39,
  output [3:0]  _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  input  [1:0]  _EVAL_43,
  input  [1:0]  _EVAL_44,
  output [3:0]  _EVAL_45,
  output        _EVAL_46,
  input  [7:0]  _EVAL_47,
  input  [3:0]  _EVAL_48,
  output [3:0]  _EVAL_49,
  output [63:0] _EVAL_50,
  output [1:0]  _EVAL_51,
  input  [2:0]  _EVAL_52,
  input  [3:0]  _EVAL_53,
  input         _EVAL_54,
  input  [3:0]  _EVAL_55,
  output [3:0]  _EVAL_56,
  input  [2:0]  _EVAL_57,
  input  [3:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  output        _EVAL_60,
  output        _EVAL_61,
  input         _EVAL_62,
  input  [3:0]  _EVAL_63,
  input  [2:0]  _EVAL_64,
  output [31:0] _EVAL_65,
  input         _EVAL_66,
  output        _EVAL_67,
  output [2:0]  _EVAL_68,
  input  [1:0]  _EVAL_69,
  output        _EVAL_70,
  input  [3:0]  _EVAL_71,
  input  [31:0] _EVAL_72,
  output        _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  output [1:0]  _EVAL_77,
  input  [2:0]  _EVAL_78,
  output        _EVAL_79,
  output [3:0]  _EVAL_80,
  output        _EVAL_81,
  input         _EVAL_82,
  output [7:0]  _EVAL_83,
  output [31:0] _EVAL_84,
  input  [31:0] _EVAL_85,
  input  [3:0]  _EVAL_86,
  input  [1:0]  _EVAL_87,
  input  [63:0] _EVAL_88,
  output        _EVAL_89,
  output [31:0] _EVAL_90,
  input  [63:0] _EVAL_91,
  output [3:0]  _EVAL_92,
  input         _EVAL_93,
  output [1:0]  _EVAL_94,
  output [3:0]  _EVAL_95,
  output [63:0] _EVAL_96,
  input  [7:0]  _EVAL_97,
  input  [31:0] _EVAL_98,
  output [1:0]  _EVAL_99,
  input         _EVAL_100,
  output [2:0]  _EVAL_101,
  input  [63:0] _EVAL_102,
  output        _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  output        _EVAL_106,
  output        _EVAL_107
);
  wire [2:0] RationalCrossingSink_1__EVAL;
  wire [3:0] RationalCrossingSink_1__EVAL_0;
  wire [2:0] RationalCrossingSink_1__EVAL_1;
  wire [2:0] RationalCrossingSink_1__EVAL_2;
  wire  RationalCrossingSink_1__EVAL_3;
  wire  RationalCrossingSink_1__EVAL_4;
  wire  RationalCrossingSink_1__EVAL_5;
  wire [3:0] RationalCrossingSink_1__EVAL_6;
  wire  RationalCrossingSink_1__EVAL_7;
  wire [3:0] RationalCrossingSink_1__EVAL_8;
  wire [1:0] RationalCrossingSink_1__EVAL_9;
  wire [63:0] RationalCrossingSink_1__EVAL_10;
  wire [3:0] RationalCrossingSink_1__EVAL_11;
  wire [31:0] RationalCrossingSink_1__EVAL_12;
  wire  RationalCrossingSink_1__EVAL_13;
  wire [31:0] RationalCrossingSink_1__EVAL_14;
  wire  RationalCrossingSink_1__EVAL_15;
  wire  RationalCrossingSink_1__EVAL_16;
  wire [1:0] RationalCrossingSink_1__EVAL_17;
  wire  RationalCrossingSink_1__EVAL_18;
  wire [31:0] RationalCrossingSink_1__EVAL_19;
  wire [2:0] RationalCrossingSink_1__EVAL_20;
  wire [3:0] RationalCrossingSink_1__EVAL_21;
  wire [2:0] RationalCrossingSink_1__EVAL_22;
  wire [2:0] RationalCrossingSink_1__EVAL_23;
  wire [63:0] RationalCrossingSink_1__EVAL_24;
  wire  RationalCrossingSink_1__EVAL_25;
  wire [3:0] RationalCrossingSink_1__EVAL_26;
  wire [63:0] RationalCrossingSink_1__EVAL_27;
  wire  RationalCrossingSink_2__EVAL;
  wire  RationalCrossingSink_2__EVAL_0;
  wire  RationalCrossingSink_2__EVAL_1;
  wire  RationalCrossingSink_2__EVAL_2;
  wire  RationalCrossingSink_2__EVAL_3;
  wire  RationalCrossingSink_2__EVAL_4;
  wire  RationalCrossingSink_2__EVAL_5;
  wire  RationalCrossingSink_2__EVAL_6;
  wire [1:0] RationalCrossingSink_2__EVAL_7;
  wire [1:0] RationalCrossingSink_2__EVAL_8;
  wire  RationalCrossingSource__EVAL;
  wire  RationalCrossingSource__EVAL_0;
  wire  RationalCrossingSource__EVAL_1;
  wire [2:0] RationalCrossingSource__EVAL_2;
  wire [2:0] RationalCrossingSource__EVAL_3;
  wire  RationalCrossingSource__EVAL_4;
  wire  RationalCrossingSource__EVAL_5;
  wire  RationalCrossingSource__EVAL_6;
  wire  RationalCrossingSource__EVAL_7;
  wire  RationalCrossingSource__EVAL_8;
  wire  RationalCrossingSource__EVAL_9;
  wire [3:0] RationalCrossingSource__EVAL_10;
  wire  RationalCrossingSource__EVAL_11;
  wire [63:0] RationalCrossingSource__EVAL_12;
  wire  RationalCrossingSource__EVAL_13;
  wire  RationalCrossingSource__EVAL_14;
  wire [1:0] RationalCrossingSource__EVAL_15;
  wire  RationalCrossingSource__EVAL_16;
  wire [1:0] RationalCrossingSource__EVAL_17;
  wire  RationalCrossingSource__EVAL_18;
  wire [1:0] RationalCrossingSource__EVAL_19;
  wire [3:0] RationalCrossingSource__EVAL_20;
  wire [3:0] RationalCrossingSource__EVAL_21;
  wire [3:0] RationalCrossingSource__EVAL_22;
  wire  RationalCrossingSource__EVAL_23;
  wire [63:0] RationalCrossingSource__EVAL_24;
  wire [1:0] RationalCrossingSource__EVAL_25;
  wire [3:0] RationalCrossingSource__EVAL_26;
  wire [3:0] RationalCrossingSource__EVAL_27;
  wire [1:0] RationalCrossingSource__EVAL_28;
  wire [2:0] RationalCrossingSource__EVAL_29;
  wire [63:0] RationalCrossingSource__EVAL_30;
  wire  RationalCrossingSource_1__EVAL;
  wire [1:0] RationalCrossingSource_1__EVAL_0;
  wire  RationalCrossingSource_1__EVAL_1;
  wire  RationalCrossingSource_1__EVAL_2;
  wire  RationalCrossingSource_1__EVAL_3;
  wire [31:0] RationalCrossingSource_1__EVAL_4;
  wire  RationalCrossingSource_1__EVAL_5;
  wire [1:0] RationalCrossingSource_1__EVAL_6;
  wire [1:0] RationalCrossingSource_1__EVAL_7;
  wire [1:0] RationalCrossingSource_1__EVAL_8;
  wire [1:0] RationalCrossingSource_1__EVAL_9;
  wire [31:0] RationalCrossingSource_1__EVAL_10;
  wire  RationalCrossingSource_1__EVAL_11;
  wire [31:0] RationalCrossingSource_1__EVAL_12;
  wire [2:0] RationalCrossingSink__EVAL;
  wire [7:0] RationalCrossingSink__EVAL_0;
  wire  RationalCrossingSink__EVAL_1;
  wire  RationalCrossingSink__EVAL_2;
  wire [3:0] RationalCrossingSink__EVAL_3;
  wire [2:0] RationalCrossingSink__EVAL_4;
  wire [3:0] RationalCrossingSink__EVAL_5;
  wire [31:0] RationalCrossingSink__EVAL_6;
  wire  RationalCrossingSink__EVAL_7;
  wire [1:0] RationalCrossingSink__EVAL_8;
  wire [63:0] RationalCrossingSink__EVAL_9;
  wire  RationalCrossingSink__EVAL_10;
  wire [1:0] RationalCrossingSink__EVAL_11;
  wire [3:0] RationalCrossingSink__EVAL_12;
  wire [2:0] RationalCrossingSink__EVAL_13;
  wire [31:0] RationalCrossingSink__EVAL_14;
  wire [3:0] RationalCrossingSink__EVAL_15;
  wire [3:0] RationalCrossingSink__EVAL_16;
  wire [63:0] RationalCrossingSink__EVAL_17;
  wire [2:0] RationalCrossingSink__EVAL_18;
  wire [3:0] RationalCrossingSink__EVAL_19;
  wire  RationalCrossingSink__EVAL_20;
  wire [31:0] RationalCrossingSink__EVAL_21;
  wire [63:0] RationalCrossingSink__EVAL_22;
  wire  RationalCrossingSink__EVAL_23;
  wire [7:0] RationalCrossingSink__EVAL_24;
  wire [2:0] RationalCrossingSink__EVAL_25;
  wire [7:0] RationalCrossingSink__EVAL_26;
  wire [2:0] RationalCrossingSink__EVAL_27;
  wire  RationalCrossingSink__EVAL_28;
  wire  RationalCrossingSink__EVAL_29;
  wire  RationalCrossingSink__EVAL_30;
  SiFive__EVAL_14 RationalCrossingSink_1 (
    ._EVAL(RationalCrossingSink_1__EVAL),
    ._EVAL_0(RationalCrossingSink_1__EVAL_0),
    ._EVAL_1(RationalCrossingSink_1__EVAL_1),
    ._EVAL_2(RationalCrossingSink_1__EVAL_2),
    ._EVAL_3(RationalCrossingSink_1__EVAL_3),
    ._EVAL_4(RationalCrossingSink_1__EVAL_4),
    ._EVAL_5(RationalCrossingSink_1__EVAL_5),
    ._EVAL_6(RationalCrossingSink_1__EVAL_6),
    ._EVAL_7(RationalCrossingSink_1__EVAL_7),
    ._EVAL_8(RationalCrossingSink_1__EVAL_8),
    ._EVAL_9(RationalCrossingSink_1__EVAL_9),
    ._EVAL_10(RationalCrossingSink_1__EVAL_10),
    ._EVAL_11(RationalCrossingSink_1__EVAL_11),
    ._EVAL_12(RationalCrossingSink_1__EVAL_12),
    ._EVAL_13(RationalCrossingSink_1__EVAL_13),
    ._EVAL_14(RationalCrossingSink_1__EVAL_14),
    ._EVAL_15(RationalCrossingSink_1__EVAL_15),
    ._EVAL_16(RationalCrossingSink_1__EVAL_16),
    ._EVAL_17(RationalCrossingSink_1__EVAL_17),
    ._EVAL_18(RationalCrossingSink_1__EVAL_18),
    ._EVAL_19(RationalCrossingSink_1__EVAL_19),
    ._EVAL_20(RationalCrossingSink_1__EVAL_20),
    ._EVAL_21(RationalCrossingSink_1__EVAL_21),
    ._EVAL_22(RationalCrossingSink_1__EVAL_22),
    ._EVAL_23(RationalCrossingSink_1__EVAL_23),
    ._EVAL_24(RationalCrossingSink_1__EVAL_24),
    ._EVAL_25(RationalCrossingSink_1__EVAL_25),
    ._EVAL_26(RationalCrossingSink_1__EVAL_26),
    ._EVAL_27(RationalCrossingSink_1__EVAL_27)
  );
  SiFive__EVAL_16 RationalCrossingSink_2 (
    ._EVAL(RationalCrossingSink_2__EVAL),
    ._EVAL_0(RationalCrossingSink_2__EVAL_0),
    ._EVAL_1(RationalCrossingSink_2__EVAL_1),
    ._EVAL_2(RationalCrossingSink_2__EVAL_2),
    ._EVAL_3(RationalCrossingSink_2__EVAL_3),
    ._EVAL_4(RationalCrossingSink_2__EVAL_4),
    ._EVAL_5(RationalCrossingSink_2__EVAL_5),
    ._EVAL_6(RationalCrossingSink_2__EVAL_6),
    ._EVAL_7(RationalCrossingSink_2__EVAL_7),
    ._EVAL_8(RationalCrossingSink_2__EVAL_8)
  );
  SiFive__EVAL_10 RationalCrossingSource (
    ._EVAL(RationalCrossingSource__EVAL),
    ._EVAL_0(RationalCrossingSource__EVAL_0),
    ._EVAL_1(RationalCrossingSource__EVAL_1),
    ._EVAL_2(RationalCrossingSource__EVAL_2),
    ._EVAL_3(RationalCrossingSource__EVAL_3),
    ._EVAL_4(RationalCrossingSource__EVAL_4),
    ._EVAL_5(RationalCrossingSource__EVAL_5),
    ._EVAL_6(RationalCrossingSource__EVAL_6),
    ._EVAL_7(RationalCrossingSource__EVAL_7),
    ._EVAL_8(RationalCrossingSource__EVAL_8),
    ._EVAL_9(RationalCrossingSource__EVAL_9),
    ._EVAL_10(RationalCrossingSource__EVAL_10),
    ._EVAL_11(RationalCrossingSource__EVAL_11),
    ._EVAL_12(RationalCrossingSource__EVAL_12),
    ._EVAL_13(RationalCrossingSource__EVAL_13),
    ._EVAL_14(RationalCrossingSource__EVAL_14),
    ._EVAL_15(RationalCrossingSource__EVAL_15),
    ._EVAL_16(RationalCrossingSource__EVAL_16),
    ._EVAL_17(RationalCrossingSource__EVAL_17),
    ._EVAL_18(RationalCrossingSource__EVAL_18),
    ._EVAL_19(RationalCrossingSource__EVAL_19),
    ._EVAL_20(RationalCrossingSource__EVAL_20),
    ._EVAL_21(RationalCrossingSource__EVAL_21),
    ._EVAL_22(RationalCrossingSource__EVAL_22),
    ._EVAL_23(RationalCrossingSource__EVAL_23),
    ._EVAL_24(RationalCrossingSource__EVAL_24),
    ._EVAL_25(RationalCrossingSource__EVAL_25),
    ._EVAL_26(RationalCrossingSource__EVAL_26),
    ._EVAL_27(RationalCrossingSource__EVAL_27),
    ._EVAL_28(RationalCrossingSource__EVAL_28),
    ._EVAL_29(RationalCrossingSource__EVAL_29),
    ._EVAL_30(RationalCrossingSource__EVAL_30)
  );
  SiFive__EVAL_12 RationalCrossingSource_1 (
    ._EVAL(RationalCrossingSource_1__EVAL),
    ._EVAL_0(RationalCrossingSource_1__EVAL_0),
    ._EVAL_1(RationalCrossingSource_1__EVAL_1),
    ._EVAL_2(RationalCrossingSource_1__EVAL_2),
    ._EVAL_3(RationalCrossingSource_1__EVAL_3),
    ._EVAL_4(RationalCrossingSource_1__EVAL_4),
    ._EVAL_5(RationalCrossingSource_1__EVAL_5),
    ._EVAL_6(RationalCrossingSource_1__EVAL_6),
    ._EVAL_7(RationalCrossingSource_1__EVAL_7),
    ._EVAL_8(RationalCrossingSource_1__EVAL_8),
    ._EVAL_9(RationalCrossingSource_1__EVAL_9),
    ._EVAL_10(RationalCrossingSource_1__EVAL_10),
    ._EVAL_11(RationalCrossingSource_1__EVAL_11),
    ._EVAL_12(RationalCrossingSource_1__EVAL_12)
  );
  SiFive__EVAL_8 RationalCrossingSink (
    ._EVAL(RationalCrossingSink__EVAL),
    ._EVAL_0(RationalCrossingSink__EVAL_0),
    ._EVAL_1(RationalCrossingSink__EVAL_1),
    ._EVAL_2(RationalCrossingSink__EVAL_2),
    ._EVAL_3(RationalCrossingSink__EVAL_3),
    ._EVAL_4(RationalCrossingSink__EVAL_4),
    ._EVAL_5(RationalCrossingSink__EVAL_5),
    ._EVAL_6(RationalCrossingSink__EVAL_6),
    ._EVAL_7(RationalCrossingSink__EVAL_7),
    ._EVAL_8(RationalCrossingSink__EVAL_8),
    ._EVAL_9(RationalCrossingSink__EVAL_9),
    ._EVAL_10(RationalCrossingSink__EVAL_10),
    ._EVAL_11(RationalCrossingSink__EVAL_11),
    ._EVAL_12(RationalCrossingSink__EVAL_12),
    ._EVAL_13(RationalCrossingSink__EVAL_13),
    ._EVAL_14(RationalCrossingSink__EVAL_14),
    ._EVAL_15(RationalCrossingSink__EVAL_15),
    ._EVAL_16(RationalCrossingSink__EVAL_16),
    ._EVAL_17(RationalCrossingSink__EVAL_17),
    ._EVAL_18(RationalCrossingSink__EVAL_18),
    ._EVAL_19(RationalCrossingSink__EVAL_19),
    ._EVAL_20(RationalCrossingSink__EVAL_20),
    ._EVAL_21(RationalCrossingSink__EVAL_21),
    ._EVAL_22(RationalCrossingSink__EVAL_22),
    ._EVAL_23(RationalCrossingSink__EVAL_23),
    ._EVAL_24(RationalCrossingSink__EVAL_24),
    ._EVAL_25(RationalCrossingSink__EVAL_25),
    ._EVAL_26(RationalCrossingSink__EVAL_26),
    ._EVAL_27(RationalCrossingSink__EVAL_27),
    ._EVAL_28(RationalCrossingSink__EVAL_28),
    ._EVAL_29(RationalCrossingSink__EVAL_29),
    ._EVAL_30(RationalCrossingSink__EVAL_30)
  );
  assign RationalCrossingSink_1__EVAL_26 = _EVAL_63;
  assign RationalCrossingSink_1__EVAL_7 = _EVAL_17;
  assign _EVAL_73 = RationalCrossingSource__EVAL_9;
  assign _EVAL_5 = RationalCrossingSource__EVAL_12;
  assign RationalCrossingSink__EVAL_16 = _EVAL_71;
  assign RationalCrossingSink_1__EVAL_12 = _EVAL_33;
  assign RationalCrossingSource_1__EVAL_5 = _EVAL_31;
  assign RationalCrossingSource__EVAL_26 = _EVAL_58;
  assign _EVAL_107 = RationalCrossingSink_2__EVAL_3;
  assign _EVAL_14 = RationalCrossingSource__EVAL_25;
  assign RationalCrossingSink__EVAL_25 = _EVAL_78;
  assign RationalCrossingSink__EVAL_19 = _EVAL_23;
  assign _EVAL_18 = RationalCrossingSource__EVAL_14;
  assign _EVAL_89 = RationalCrossingSource__EVAL_23;
  assign RationalCrossingSink_2__EVAL_5 = _EVAL_66;
  assign RationalCrossingSource__EVAL_13 = _EVAL_75;
  assign RationalCrossingSink_1__EVAL_15 = _EVAL_104;
  assign _EVAL_77 = RationalCrossingSink_2__EVAL_7;
  assign RationalCrossingSink_1__EVAL_10 = _EVAL_91;
  assign _EVAL_103 = RationalCrossingSink__EVAL_20;
  assign RationalCrossingSource__EVAL_11 = _EVAL_100;
  assign RationalCrossingSource__EVAL_21 = _EVAL_55;
  assign _EVAL_21 = RationalCrossingSink_1__EVAL_19;
  assign RationalCrossingSink_1__EVAL_20 = _EVAL_36;
  assign _EVAL_56 = RationalCrossingSource__EVAL_22;
  assign RationalCrossingSource__EVAL_19 = _EVAL_29;
  assign RationalCrossingSink__EVAL_22 = _EVAL_20;
  assign RationalCrossingSource__EVAL_1 = _EVAL_105;
  assign _EVAL_92 = RationalCrossingSource__EVAL_20;
  assign _EVAL_16 = RationalCrossingSource_1__EVAL_7;
  assign RationalCrossingSink__EVAL_3 = _EVAL_24;
  assign _EVAL_94 = RationalCrossingSource__EVAL_28;
  assign RationalCrossingSink_2__EVAL_0 = _EVAL_74;
  assign RationalCrossingSource__EVAL_0 = _EVAL_82;
  assign RationalCrossingSink__EVAL_21 = _EVAL_72;
  assign _EVAL_6 = RationalCrossingSink__EVAL_11;
  assign _EVAL_106 = RationalCrossingSink_2__EVAL_6;
  assign _EVAL_1 = RationalCrossingSink__EVAL_13;
  assign RationalCrossingSink_1__EVAL_5 = _EVAL_3;
  assign _EVAL_8 = RationalCrossingSink_1__EVAL_13;
  assign _EVAL_60 = RationalCrossingSource__EVAL_7;
  assign RationalCrossingSink_2__EVAL_2 = _EVAL_4;
  assign RationalCrossingSink__EVAL_27 = _EVAL_35;
  assign RationalCrossingSink_1__EVAL_25 = _EVAL_31;
  assign RationalCrossingSink__EVAL_10 = _EVAL_31;
  assign _EVAL_49 = RationalCrossingSink__EVAL_5;
  assign RationalCrossingSource_1__EVAL_10 = _EVAL_98;
  assign _EVAL_84 = RationalCrossingSource_1__EVAL_12;
  assign RationalCrossingSink__EVAL_7 = _EVAL_76;
  assign _EVAL_80 = RationalCrossingSink_1__EVAL_11;
  assign RationalCrossingSink_1__EVAL_27 = _EVAL_88;
  assign RationalCrossingSink__EVAL_30 = _EVAL_93;
  assign RationalCrossingSource__EVAL_17 = _EVAL_44;
  assign _EVAL_90 = RationalCrossingSink__EVAL_14;
  assign RationalCrossingSink__EVAL = _EVAL_64;
  assign _EVAL_50 = RationalCrossingSink_1__EVAL_24;
  assign _EVAL_46 = RationalCrossingSource_1__EVAL_11;
  assign RationalCrossingSink_1__EVAL_16 = _EVAL_26;
  assign RationalCrossingSink_1__EVAL_22 = _EVAL_25;
  assign _EVAL_65 = RationalCrossingSource_1__EVAL_4;
  assign RationalCrossingSink__EVAL_24 = _EVAL_47;
  assign _EVAL_7 = RationalCrossingSource__EVAL_8;
  assign RationalCrossingSource_1__EVAL_2 = _EVAL_66;
  assign _EVAL_51 = RationalCrossingSource__EVAL_15;
  assign _EVAL_0 = RationalCrossingSink_1__EVAL;
  assign _EVAL_32 = RationalCrossingSink__EVAL_18;
  assign _EVAL_39 = RationalCrossingSource_1__EVAL_0;
  assign RationalCrossingSink__EVAL_28 = _EVAL_66;
  assign RationalCrossingSource__EVAL_16 = _EVAL_31;
  assign _EVAL_79 = RationalCrossingSource_1__EVAL_1;
  assign _EVAL_27 = RationalCrossingSink__EVAL_9;
  assign _EVAL_67 = RationalCrossingSource__EVAL;
  assign RationalCrossingSink_1__EVAL_21 = _EVAL_86;
  assign _EVAL_45 = RationalCrossingSource__EVAL_10;
  assign _EVAL_83 = RationalCrossingSink__EVAL_26;
  assign RationalCrossingSource__EVAL_5 = _EVAL_66;
  assign RationalCrossingSink__EVAL_17 = _EVAL_102;
  assign _EVAL_41 = RationalCrossingSource__EVAL_6;
  assign _EVAL_81 = RationalCrossingSink_1__EVAL_4;
  assign RationalCrossingSink_1__EVAL_14 = _EVAL_85;
  assign _EVAL_99 = RationalCrossingSource_1__EVAL_8;
  assign _EVAL_61 = RationalCrossingSource__EVAL_18;
  assign _EVAL_15 = RationalCrossingSink_1__EVAL_9;
  assign RationalCrossingSink__EVAL_29 = _EVAL_12;
  assign _EVAL_96 = RationalCrossingSource__EVAL_24;
  assign _EVAL_59 = RationalCrossingSink_1__EVAL_8;
  assign RationalCrossingSink_2__EVAL_1 = _EVAL_31;
  assign _EVAL_40 = RationalCrossingSource__EVAL_27;
  assign RationalCrossingSink_1__EVAL_3 = _EVAL_66;
  assign _EVAL_95 = RationalCrossingSink__EVAL_15;
  assign _EVAL_42 = RationalCrossingSink_2__EVAL;
  assign RationalCrossingSink_2__EVAL_4 = _EVAL_19;
  assign RationalCrossingSource_1__EVAL = _EVAL;
  assign RationalCrossingSource__EVAL_4 = _EVAL_62;
  assign RationalCrossingSource__EVAL_30 = _EVAL_2;
  assign RationalCrossingSink_1__EVAL_0 = _EVAL_53;
  assign RationalCrossingSource__EVAL_29 = _EVAL_10;
  assign RationalCrossingSink__EVAL_6 = _EVAL_11;
  assign RationalCrossingSource_1__EVAL_9 = _EVAL_43;
  assign _EVAL_68 = RationalCrossingSource__EVAL_3;
  assign RationalCrossingSink__EVAL_4 = _EVAL_22;
  assign RationalCrossingSink_1__EVAL_6 = _EVAL_34;
  assign RationalCrossingSink_2__EVAL_8 = _EVAL_69;
  assign RationalCrossingSource_1__EVAL_3 = _EVAL_38;
  assign RationalCrossingSink_1__EVAL_1 = _EVAL_52;
  assign RationalCrossingSink_1__EVAL_17 = _EVAL_87;
  assign RationalCrossingSource_1__EVAL_6 = _EVAL_28;
  assign _EVAL_9 = RationalCrossingSink_1__EVAL_2;
  assign _EVAL_101 = RationalCrossingSource__EVAL_2;
  assign _EVAL_37 = RationalCrossingSink__EVAL_23;
  assign RationalCrossingSink__EVAL_8 = _EVAL_30;
  assign RationalCrossingSink__EVAL_2 = _EVAL_54;
  assign _EVAL_13 = RationalCrossingSink__EVAL_1;
  assign _EVAL_70 = RationalCrossingSink_1__EVAL_18;
  assign RationalCrossingSink__EVAL_12 = _EVAL_48;
  assign RationalCrossingSink__EVAL_0 = _EVAL_97;
  assign RationalCrossingSink_1__EVAL_23 = _EVAL_57;
endmodule
