//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_112_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_9,
  input         _EVAL_11,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  input  [29:0] _EVAL_16,
  input  [6:0]  _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [3:0]  _EVAL_31,
  input  [6:0]  _EVAL_34,
  input         _EVAL_39,
  input  [3:0]  _EVAL_40,
  input         _EVAL_43,
  input         _EVAL_90,
  input         _EVAL_99,
  input         _EVAL_141,
  input         _EVAL_170,
  input         _EVAL_173,
  input         _EVAL_204,
  input         _EVAL_212,
  input         _EVAL_219,
  input         _EVAL_273,
  input         _EVAL_293,
  input         _EVAL_296,
  input         _EVAL_344,
  input         _EVAL_357,
  input         _EVAL_358,
  input         _EVAL_370,
  input         _EVAL_401,
  input         _EVAL_410,
  input         _EVAL_413,
  input         _EVAL_476,
  input         _EVAL_490,
  input         _EVAL_491,
  input         _EVAL_501,
  input         _EVAL_511,
  input         _EVAL_556,
  input         _EVAL_598,
  input         _EVAL_603,
  input         _EVAL_623,
  input         _EVAL_630,
  input         _EVAL_634,
  input         _EVAL_640,
  input         _EVAL_97,
  input         _EVAL_557,
  input         _EVAL_266,
  input         _EVAL_562,
  input         _EVAL_589
);
  wire [2:0] TLMonitor__EVAL;
  wire [6:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire [3:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire [3:0] TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire [3:0] TLMonitor__EVAL_8;
  wire [2:0] TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire  TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [6:0] TLMonitor__EVAL_14;
  wire [1:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire [2:0] TLMonitor__EVAL_17;
  wire [29:0] TLMonitor__EVAL_18;
  reg  _EVAL_47;
  reg [31:0] _RAND_0;
  reg  _EVAL_67;
  reg [31:0] _RAND_1;
  reg  _EVAL_78;
  reg [31:0] _RAND_2;
  reg  _EVAL_98;
  reg [31:0] _RAND_3;
  reg  _EVAL_108;
  reg [31:0] _RAND_4;
  reg  _EVAL_119;
  reg [31:0] _RAND_5;
  reg  _EVAL_128;
  reg [31:0] _RAND_6;
  reg  _EVAL_203;
  reg [31:0] _RAND_7;
  reg  _EVAL_205;
  reg [31:0] _RAND_8;
  reg  _EVAL_224;
  reg [31:0] _RAND_9;
  reg  _EVAL_252;
  reg [31:0] _RAND_10;
  reg  _EVAL_269;
  reg [31:0] _RAND_11;
  reg  _EVAL_271;
  reg [31:0] _RAND_12;
  reg  _EVAL_279;
  reg [31:0] _RAND_13;
  reg  _EVAL_289;
  reg [31:0] _RAND_14;
  reg  _EVAL_315;
  reg [31:0] _RAND_15;
  reg  _EVAL_340;
  reg [31:0] _RAND_16;
  reg  _EVAL_351;
  reg [31:0] _RAND_17;
  reg  _EVAL_377;
  reg [31:0] _RAND_18;
  reg  _EVAL_382;
  reg [31:0] _RAND_19;
  reg  _EVAL_390;
  reg [31:0] _RAND_20;
  reg  _EVAL_432;
  reg [31:0] _RAND_21;
  reg  _EVAL_437;
  reg [31:0] _RAND_22;
  reg  _EVAL_448;
  reg [31:0] _RAND_23;
  reg  _EVAL_466;
  reg [31:0] _RAND_24;
  reg  _EVAL_471;
  reg [31:0] _RAND_25;
  reg  _EVAL_484;
  reg [31:0] _RAND_26;
  reg  _EVAL_517;
  reg [31:0] _RAND_27;
  reg  _EVAL_555;
  reg [31:0] _RAND_28;
  reg  _EVAL_559;
  reg [31:0] _RAND_29;
  reg  _EVAL_564;
  reg [31:0] _RAND_30;
  reg  _EVAL_594;
  reg [31:0] _RAND_31;
  reg [72:0] _EVAL_608;
  reg [95:0] _RAND_32;
  reg  _EVAL_627;
  reg [31:0] _RAND_33;
  reg  _EVAL_633;
  reg [31:0] _RAND_34;
  wire  _EVAL_117;
  wire  _EVAL_573;
  wire  _EVAL_280;
  wire  _EVAL_609;
  wire  _EVAL_50;
  wire  _EVAL_209;
  wire  _EVAL_425;
  wire  _EVAL_328;
  wire  _EVAL_475;
  wire  _EVAL_583;
  wire  _EVAL_77;
  wire  _EVAL_427;
  wire  _EVAL_621;
  wire  _EVAL_622;
  wire  _EVAL_576;
  wire  _EVAL_318;
  wire  _EVAL_365;
  wire  _EVAL_247;
  wire  _EVAL_136;
  wire  _EVAL_659;
  wire  _EVAL_597;
  wire  _EVAL_60;
  wire  _EVAL_214;
  wire  _EVAL_95;
  wire  _EVAL_592;
  wire  _EVAL_193;
  wire  _EVAL_498;
  wire  _EVAL_254;
  wire  _EVAL_121;
  wire  _EVAL_488;
  wire  _EVAL_560;
  wire  _EVAL_506;
  wire  _EVAL_435;
  wire  _EVAL_540;
  wire  _EVAL_309;
  wire  _EVAL_185;
  wire  _EVAL_657;
  wire  _EVAL_147;
  wire  _EVAL_364;
  wire  _EVAL_165;
  wire  _EVAL_155;
  wire  _EVAL_157;
  wire  _EVAL_620;
  wire  _EVAL_584;
  wire  _EVAL_639;
  wire  _EVAL_325;
  wire  _EVAL_213;
  wire  _EVAL_600;
  wire [127:0] _EVAL_248;
  wire [127:0] _EVAL_563;
  wire [72:0] _EVAL_406;
  wire  _EVAL_643;
  wire  _EVAL_459;
  wire  _EVAL_581;
  wire  _EVAL_468;
  wire  _EVAL_274;
  wire  _EVAL_69;
  wire  _EVAL_316;
  wire  _EVAL_94;
  wire  _EVAL_126;
  wire [127:0] _EVAL_587;
  wire [127:0] _EVAL_101;
  wire [72:0] _EVAL_195;
  wire  _EVAL_450;
  wire  _EVAL_551;
  wire  _EVAL_225;
  wire  _EVAL_72;
  wire  _EVAL_159;
  wire  _EVAL_384;
  wire  _EVAL_470;
  wire  _EVAL_172;
  wire  _EVAL_138;
  wire  _EVAL_652;
  wire  _EVAL_526;
  wire  _EVAL_402;
  wire [72:0] _EVAL_423;
  wire  _EVAL_412;
  wire  _EVAL_123;
  SiFive__EVAL_111_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18)
  );
  assign _EVAL_117 = _EVAL_97 | _EVAL_634;
  assign _EVAL_573 = _EVAL_117 | _EVAL_141;
  assign _EVAL_280 = _EVAL_573 | _EVAL_598;
  assign _EVAL_609 = _EVAL_280 | _EVAL_293;
  assign _EVAL_50 = _EVAL_609 | _EVAL_170;
  assign _EVAL_209 = _EVAL_50 | _EVAL_603;
  assign _EVAL_425 = _EVAL_209 | _EVAL_410;
  assign _EVAL_328 = _EVAL_425 | _EVAL_173;
  assign _EVAL_475 = _EVAL_328 | _EVAL_556;
  assign _EVAL_583 = _EVAL_475 | _EVAL_99;
  assign _EVAL_77 = _EVAL_583 | _EVAL_296;
  assign _EVAL_427 = _EVAL_77 | _EVAL_490;
  assign _EVAL_621 = _EVAL_427 | _EVAL_511;
  assign _EVAL_622 = _EVAL_621 | _EVAL_623;
  assign _EVAL_576 = _EVAL_622 | _EVAL_204;
  assign _EVAL_318 = _EVAL_576 | _EVAL_90;
  assign _EVAL_365 = _EVAL_318 | _EVAL_219;
  assign _EVAL_247 = _EVAL_365 | _EVAL_413;
  assign _EVAL_136 = _EVAL_247 | _EVAL_640;
  assign _EVAL_659 = _EVAL_136 | _EVAL_357;
  assign _EVAL_597 = _EVAL_659 | _EVAL_212;
  assign _EVAL_60 = _EVAL_597 | _EVAL_491;
  assign _EVAL_214 = _EVAL_60 | _EVAL_358;
  assign _EVAL_95 = _EVAL_214 | _EVAL_401;
  assign _EVAL_592 = _EVAL_95 | _EVAL_279;
  assign _EVAL_193 = _EVAL_592 | _EVAL_67;
  assign _EVAL_498 = _EVAL_193 | _EVAL_437;
  assign _EVAL_254 = _EVAL_498 | _EVAL_269;
  assign _EVAL_121 = _EVAL_254 | _EVAL_564;
  assign _EVAL_488 = _EVAL_121 | _EVAL_377;
  assign _EVAL_560 = _EVAL_488 | _EVAL_466;
  assign _EVAL_506 = _EVAL_560 | _EVAL_432;
  assign _EVAL_435 = _EVAL_506 | _EVAL_224;
  assign _EVAL_540 = _EVAL_435 | _EVAL_594;
  assign _EVAL_309 = _EVAL_540 | _EVAL_555;
  assign _EVAL_185 = _EVAL_309 | _EVAL_252;
  assign _EVAL_657 = _EVAL_185 | _EVAL_382;
  assign _EVAL_147 = _EVAL_657 | _EVAL_484;
  assign _EVAL_364 = _EVAL_147 | _EVAL_448;
  assign _EVAL_165 = _EVAL_364 | _EVAL_627;
  assign _EVAL_155 = _EVAL_165 | _EVAL_271;
  assign _EVAL_157 = _EVAL_155 | _EVAL_340;
  assign _EVAL_620 = _EVAL_157 | _EVAL_289;
  assign _EVAL_584 = _EVAL_620 | _EVAL_315;
  assign _EVAL_639 = _EVAL_584 | _EVAL_390;
  assign _EVAL_325 = _EVAL_639 | _EVAL_47;
  assign _EVAL_213 = _EVAL_325 | _EVAL_559;
  assign _EVAL_600 = _EVAL_213 | _EVAL_205;
  assign _EVAL_248 = 128'h1 << _EVAL_34;
  assign _EVAL_563 = _EVAL_562 ? _EVAL_248 : 128'h0;
  assign _EVAL_406 = _EVAL_563[72:0];
  assign _EVAL_643 = _EVAL_600 | _EVAL_351;
  assign _EVAL_459 = _EVAL_643 | _EVAL_633;
  assign _EVAL_581 = _EVAL_459 | _EVAL_203;
  assign _EVAL_468 = _EVAL_581 | _EVAL_517;
  assign _EVAL_274 = _EVAL_468 | _EVAL_108;
  assign _EVAL_69 = _EVAL_274 | _EVAL_78;
  assign _EVAL_316 = _EVAL_69 | _EVAL_128;
  assign _EVAL_94 = _EVAL_316 | _EVAL_98;
  assign _EVAL_126 = _EVAL_94 | _EVAL_119;
  assign _EVAL_587 = 128'h1 << _EVAL_21;
  assign _EVAL_101 = _EVAL_589 ? _EVAL_587 : 128'h0;
  assign _EVAL_195 = _EVAL_101[72:0];
  assign _EVAL_450 = _EVAL_195 > 73'h0;
  assign _EVAL_551 = _EVAL_11 == 1'h0;
  assign _EVAL_225 = _EVAL_126 | _EVAL_370;
  assign _EVAL_72 = _EVAL_225 | _EVAL_501;
  assign _EVAL_159 = _EVAL_608 == 73'h1ffffffffffffffffff;
  assign _EVAL_384 = _EVAL_406 > 73'h0;
  assign _EVAL_470 = _EVAL_72 | _EVAL_630;
  assign _EVAL_172 = _EVAL_470 | _EVAL_344;
  assign _EVAL_138 = _EVAL_172 | _EVAL_476;
  assign _EVAL_652 = _EVAL_138 | _EVAL_43;
  assign _EVAL_526 = _EVAL_652 | _EVAL_273;
  assign _EVAL_402 = _EVAL_9 & _EVAL_557;
  assign _EVAL_423 = _EVAL_608 | _EVAL_406;
  assign _EVAL_412 = _EVAL_526 | _EVAL_471;
  assign _EVAL_123 = _EVAL_412 == 1'h0;
  assign TLMonitor__EVAL_2 = _EVAL_14;
  assign TLMonitor__EVAL_17 = _EVAL_2;
  assign TLMonitor__EVAL_4 = _EVAL_3;
  assign TLMonitor__EVAL_8 = _EVAL_31;
  assign TLMonitor__EVAL_12 = _EVAL_11;
  assign TLMonitor__EVAL_6 = _EVAL_40;
  assign TLMonitor__EVAL_0 = _EVAL_21;
  assign TLMonitor__EVAL_5 = _EVAL_24 & _EVAL_266;
  assign TLMonitor__EVAL = _EVAL_22;
  assign TLMonitor__EVAL_1 = _EVAL_23;
  assign TLMonitor__EVAL_16 = _EVAL_9;
  assign TLMonitor__EVAL_11 = _EVAL_1;
  assign TLMonitor__EVAL_15 = _EVAL_15;
  assign TLMonitor__EVAL_10 = _EVAL_5;
  assign TLMonitor__EVAL_18 = _EVAL_16;
  assign TLMonitor__EVAL_13 = _EVAL_4;
  assign TLMonitor__EVAL_3 = _EVAL_0;
  assign TLMonitor__EVAL_7 = _EVAL_39;
  assign TLMonitor__EVAL_9 = _EVAL;
  assign TLMonitor__EVAL_14 = _EVAL_34;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_47 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_67 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_78 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_98 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_108 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_119 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_128 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_203 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_205 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_224 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_252 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_269 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_271 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_279 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_289 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_315 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_340 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_351 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_377 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_382 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_390 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_432 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_437 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_448 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_466 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_471 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_484 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_517 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_555 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_559 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_564 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_594 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {3{`RANDOM}};
  _EVAL_608 = _RAND_32[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_627 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_633 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_11) begin
      _EVAL_47 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h35 == _EVAL_21) begin
          _EVAL_47 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h35 == _EVAL_34) begin
              _EVAL_47 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h35 == _EVAL_34) begin
            _EVAL_47 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_67 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h21 == _EVAL_21) begin
          _EVAL_67 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h21 == _EVAL_34) begin
              _EVAL_67 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h21 == _EVAL_34) begin
            _EVAL_67 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_78 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3d == _EVAL_21) begin
          _EVAL_78 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3d == _EVAL_34) begin
              _EVAL_78 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3d == _EVAL_34) begin
            _EVAL_78 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_98 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3f == _EVAL_21) begin
          _EVAL_98 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3f == _EVAL_34) begin
              _EVAL_98 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3f == _EVAL_34) begin
            _EVAL_98 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_108 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3c == _EVAL_21) begin
          _EVAL_108 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3c == _EVAL_34) begin
              _EVAL_108 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3c == _EVAL_34) begin
            _EVAL_108 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_119 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h40 == _EVAL_21) begin
          _EVAL_119 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h40 == _EVAL_34) begin
              _EVAL_119 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h40 == _EVAL_34) begin
            _EVAL_119 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_128 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3e == _EVAL_21) begin
          _EVAL_128 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3e == _EVAL_34) begin
              _EVAL_128 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3e == _EVAL_34) begin
            _EVAL_128 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_203 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3a == _EVAL_21) begin
          _EVAL_203 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3a == _EVAL_34) begin
              _EVAL_203 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3a == _EVAL_34) begin
            _EVAL_203 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_205 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h37 == _EVAL_21) begin
          _EVAL_205 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h37 == _EVAL_34) begin
              _EVAL_205 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h37 == _EVAL_34) begin
            _EVAL_205 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_224 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h28 == _EVAL_21) begin
          _EVAL_224 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h28 == _EVAL_34) begin
              _EVAL_224 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h28 == _EVAL_34) begin
            _EVAL_224 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_252 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2b == _EVAL_21) begin
          _EVAL_252 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2b == _EVAL_34) begin
              _EVAL_252 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2b == _EVAL_34) begin
            _EVAL_252 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_269 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h23 == _EVAL_21) begin
          _EVAL_269 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h23 == _EVAL_34) begin
              _EVAL_269 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h23 == _EVAL_34) begin
            _EVAL_269 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_271 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h30 == _EVAL_21) begin
          _EVAL_271 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h30 == _EVAL_34) begin
              _EVAL_271 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h30 == _EVAL_34) begin
            _EVAL_271 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_279 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h20 == _EVAL_21) begin
          _EVAL_279 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h20 == _EVAL_34) begin
              _EVAL_279 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h20 == _EVAL_34) begin
            _EVAL_279 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_289 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h32 == _EVAL_21) begin
          _EVAL_289 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h32 == _EVAL_34) begin
              _EVAL_289 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h32 == _EVAL_34) begin
            _EVAL_289 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_315 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h33 == _EVAL_21) begin
          _EVAL_315 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h33 == _EVAL_34) begin
              _EVAL_315 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h33 == _EVAL_34) begin
            _EVAL_315 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_340 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h31 == _EVAL_21) begin
          _EVAL_340 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h31 == _EVAL_34) begin
              _EVAL_340 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h31 == _EVAL_34) begin
            _EVAL_340 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_351 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h38 == _EVAL_21) begin
          _EVAL_351 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h38 == _EVAL_34) begin
              _EVAL_351 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h38 == _EVAL_34) begin
            _EVAL_351 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_377 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h25 == _EVAL_21) begin
          _EVAL_377 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h25 == _EVAL_34) begin
              _EVAL_377 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h25 == _EVAL_34) begin
            _EVAL_377 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_382 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2c == _EVAL_21) begin
          _EVAL_382 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2c == _EVAL_34) begin
              _EVAL_382 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2c == _EVAL_34) begin
            _EVAL_382 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_390 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h34 == _EVAL_21) begin
          _EVAL_390 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h34 == _EVAL_34) begin
              _EVAL_390 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h34 == _EVAL_34) begin
            _EVAL_390 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_432 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h27 == _EVAL_21) begin
          _EVAL_432 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h27 == _EVAL_34) begin
              _EVAL_432 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h27 == _EVAL_34) begin
            _EVAL_432 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_437 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h22 == _EVAL_21) begin
          _EVAL_437 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h22 == _EVAL_34) begin
              _EVAL_437 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h22 == _EVAL_34) begin
            _EVAL_437 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_448 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2e == _EVAL_21) begin
          _EVAL_448 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2e == _EVAL_34) begin
              _EVAL_448 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2e == _EVAL_34) begin
            _EVAL_448 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_466 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h26 == _EVAL_21) begin
          _EVAL_466 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h26 == _EVAL_34) begin
              _EVAL_466 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h26 == _EVAL_34) begin
            _EVAL_466 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_471 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h48 == _EVAL_21) begin
          _EVAL_471 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h48 == _EVAL_34) begin
              _EVAL_471 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h48 == _EVAL_34) begin
            _EVAL_471 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_484 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2d == _EVAL_21) begin
          _EVAL_484 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2d == _EVAL_34) begin
              _EVAL_484 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2d == _EVAL_34) begin
            _EVAL_484 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_517 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3b == _EVAL_21) begin
          _EVAL_517 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3b == _EVAL_34) begin
              _EVAL_517 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3b == _EVAL_34) begin
            _EVAL_517 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_555 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2a == _EVAL_21) begin
          _EVAL_555 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2a == _EVAL_34) begin
              _EVAL_555 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2a == _EVAL_34) begin
            _EVAL_555 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_559 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h36 == _EVAL_21) begin
          _EVAL_559 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h36 == _EVAL_34) begin
              _EVAL_559 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h36 == _EVAL_34) begin
            _EVAL_559 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_564 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h24 == _EVAL_21) begin
          _EVAL_564 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h24 == _EVAL_34) begin
              _EVAL_564 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h24 == _EVAL_34) begin
            _EVAL_564 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_594 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h29 == _EVAL_21) begin
          _EVAL_594 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h29 == _EVAL_34) begin
              _EVAL_594 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h29 == _EVAL_34) begin
            _EVAL_594 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_608 <= 73'h0;
    end else begin
      _EVAL_608 <= _EVAL_423;
    end
    if (_EVAL_11) begin
      _EVAL_627 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2f == _EVAL_21) begin
          _EVAL_627 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2f == _EVAL_34) begin
              _EVAL_627 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2f == _EVAL_34) begin
            _EVAL_627 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_633 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h39 == _EVAL_21) begin
          _EVAL_633 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h39 == _EVAL_34) begin
              _EVAL_633 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h39 == _EVAL_34) begin
            _EVAL_633 <= 1'h1;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_551) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf26c64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_450 & _EVAL_551) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(687f9502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_551) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e982a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_402 & _EVAL_551) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cee430f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_551) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b98e21ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
