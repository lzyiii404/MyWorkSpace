//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module CoreIPSubsystemAllPortRAMTestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  system_clock;
  wire  system_reset;
  wire  system_debug_psd_test_mode;
  wire  system_debug_psd_test_mode_reset;
  wire  system_debug_systemjtag_jtag_TCK;
  wire  system_debug_systemjtag_jtag_TMS;
  wire  system_debug_systemjtag_jtag_TDI;
  wire  system_debug_systemjtag_jtag_TDO_data;
  wire  system_debug_systemjtag_jtag_TDO_driven;
  wire  system_debug_systemjtag_reset;
  wire [10:0] system_debug_systemjtag_mfr_id;
  wire  system_debug_ndreset;
  wire  system_debug_dmactive;
  wire  system_core_clock_0;
  wire [31:0] system_reset_vector_0;
  wire  system_rtc_toggle;
  wire [126:0] system_global_interrupts;
  wire  system_mem_port_axi4_0_aw_ready;
  wire  system_mem_port_axi4_0_aw_valid;
  wire [3:0] system_mem_port_axi4_0_aw_bits_id;
  wire [31:0] system_mem_port_axi4_0_aw_bits_addr;
  wire [7:0] system_mem_port_axi4_0_aw_bits_len;
  wire [2:0] system_mem_port_axi4_0_aw_bits_size;
  wire [1:0] system_mem_port_axi4_0_aw_bits_burst;
  wire  system_mem_port_axi4_0_aw_bits_lock;
  wire [3:0] system_mem_port_axi4_0_aw_bits_cache;
  wire [2:0] system_mem_port_axi4_0_aw_bits_prot;
  wire [3:0] system_mem_port_axi4_0_aw_bits_qos;
  wire  system_mem_port_axi4_0_w_ready;
  wire  system_mem_port_axi4_0_w_valid;
  wire [63:0] system_mem_port_axi4_0_w_bits_data;
  wire [7:0] system_mem_port_axi4_0_w_bits_strb;
  wire  system_mem_port_axi4_0_w_bits_last;
  wire  system_mem_port_axi4_0_w_bits_corrupt;
  wire  system_mem_port_axi4_0_b_ready;
  wire  system_mem_port_axi4_0_b_valid;
  wire [3:0] system_mem_port_axi4_0_b_bits_id;
  wire [1:0] system_mem_port_axi4_0_b_bits_resp;
  wire  system_mem_port_axi4_0_ar_ready;
  wire  system_mem_port_axi4_0_ar_valid;
  wire [3:0] system_mem_port_axi4_0_ar_bits_id;
  wire [31:0] system_mem_port_axi4_0_ar_bits_addr;
  wire [7:0] system_mem_port_axi4_0_ar_bits_len;
  wire [2:0] system_mem_port_axi4_0_ar_bits_size;
  wire [1:0] system_mem_port_axi4_0_ar_bits_burst;
  wire  system_mem_port_axi4_0_ar_bits_lock;
  wire [3:0] system_mem_port_axi4_0_ar_bits_cache;
  wire [2:0] system_mem_port_axi4_0_ar_bits_prot;
  wire [3:0] system_mem_port_axi4_0_ar_bits_qos;
  wire  system_mem_port_axi4_0_r_ready;
  wire  system_mem_port_axi4_0_r_valid;
  wire [3:0] system_mem_port_axi4_0_r_bits_id;
  wire [63:0] system_mem_port_axi4_0_r_bits_data;
  wire [1:0] system_mem_port_axi4_0_r_bits_resp;
  wire  system_mem_port_axi4_0_r_bits_last;
  wire  system_sys_port_axi4_0_aw_ready;
  wire  system_sys_port_axi4_0_aw_valid;
  wire [3:0] system_sys_port_axi4_0_aw_bits_id;
  wire [30:0] system_sys_port_axi4_0_aw_bits_addr;
  wire [7:0] system_sys_port_axi4_0_aw_bits_len;
  wire [2:0] system_sys_port_axi4_0_aw_bits_size;
  wire [1:0] system_sys_port_axi4_0_aw_bits_burst;
  wire  system_sys_port_axi4_0_aw_bits_lock;
  wire [3:0] system_sys_port_axi4_0_aw_bits_cache;
  wire [2:0] system_sys_port_axi4_0_aw_bits_prot;
  wire [3:0] system_sys_port_axi4_0_aw_bits_qos;
  wire  system_sys_port_axi4_0_w_ready;
  wire  system_sys_port_axi4_0_w_valid;
  wire [31:0] system_sys_port_axi4_0_w_bits_data;
  wire [3:0] system_sys_port_axi4_0_w_bits_strb;
  wire  system_sys_port_axi4_0_w_bits_last;
  wire  system_sys_port_axi4_0_b_ready;
  wire  system_sys_port_axi4_0_b_valid;
  wire [3:0] system_sys_port_axi4_0_b_bits_id;
  wire [1:0] system_sys_port_axi4_0_b_bits_resp;
  wire  system_sys_port_axi4_0_ar_ready;
  wire  system_sys_port_axi4_0_ar_valid;
  wire [3:0] system_sys_port_axi4_0_ar_bits_id;
  wire [30:0] system_sys_port_axi4_0_ar_bits_addr;
  wire [7:0] system_sys_port_axi4_0_ar_bits_len;
  wire [2:0] system_sys_port_axi4_0_ar_bits_size;
  wire [1:0] system_sys_port_axi4_0_ar_bits_burst;
  wire  system_sys_port_axi4_0_ar_bits_lock;
  wire [3:0] system_sys_port_axi4_0_ar_bits_cache;
  wire [2:0] system_sys_port_axi4_0_ar_bits_prot;
  wire [3:0] system_sys_port_axi4_0_ar_bits_qos;
  wire  system_sys_port_axi4_0_r_ready;
  wire  system_sys_port_axi4_0_r_valid;
  wire [3:0] system_sys_port_axi4_0_r_bits_id;
  wire [31:0] system_sys_port_axi4_0_r_bits_data;
  wire [1:0] system_sys_port_axi4_0_r_bits_resp;
  wire  system_sys_port_axi4_0_r_bits_last;
  wire  system_periph_port_axi4_0_aw_ready;
  wire  system_periph_port_axi4_0_aw_valid;
  wire  system_periph_port_axi4_0_aw_bits_id;
  wire [29:0] system_periph_port_axi4_0_aw_bits_addr;
  wire [7:0] system_periph_port_axi4_0_aw_bits_len;
  wire [2:0] system_periph_port_axi4_0_aw_bits_size;
  wire [1:0] system_periph_port_axi4_0_aw_bits_burst;
  wire  system_periph_port_axi4_0_aw_bits_lock;
  wire [3:0] system_periph_port_axi4_0_aw_bits_cache;
  wire [2:0] system_periph_port_axi4_0_aw_bits_prot;
  wire [3:0] system_periph_port_axi4_0_aw_bits_qos;
  wire  system_periph_port_axi4_0_w_ready;
  wire  system_periph_port_axi4_0_w_valid;
  wire [31:0] system_periph_port_axi4_0_w_bits_data;
  wire [3:0] system_periph_port_axi4_0_w_bits_strb;
  wire  system_periph_port_axi4_0_w_bits_last;
  wire  system_periph_port_axi4_0_b_ready;
  wire  system_periph_port_axi4_0_b_valid;
  wire  system_periph_port_axi4_0_b_bits_id;
  wire [1:0] system_periph_port_axi4_0_b_bits_resp;
  wire  system_periph_port_axi4_0_ar_ready;
  wire  system_periph_port_axi4_0_ar_valid;
  wire  system_periph_port_axi4_0_ar_bits_id;
  wire [29:0] system_periph_port_axi4_0_ar_bits_addr;
  wire [7:0] system_periph_port_axi4_0_ar_bits_len;
  wire [2:0] system_periph_port_axi4_0_ar_bits_size;
  wire [1:0] system_periph_port_axi4_0_ar_bits_burst;
  wire  system_periph_port_axi4_0_ar_bits_lock;
  wire [3:0] system_periph_port_axi4_0_ar_bits_cache;
  wire [2:0] system_periph_port_axi4_0_ar_bits_prot;
  wire [3:0] system_periph_port_axi4_0_ar_bits_qos;
  wire  system_periph_port_axi4_0_r_ready;
  wire  system_periph_port_axi4_0_r_valid;
  wire  system_periph_port_axi4_0_r_bits_id;
  wire [31:0] system_periph_port_axi4_0_r_bits_data;
  wire [1:0] system_periph_port_axi4_0_r_bits_resp;
  wire  system_periph_port_axi4_0_r_bits_last;
  wire  system_front_port_axi4_0_aw_ready;
  wire  system_front_port_axi4_0_aw_valid;
  wire [7:0] system_front_port_axi4_0_aw_bits_id;
  wire [31:0] system_front_port_axi4_0_aw_bits_addr;
  wire [7:0] system_front_port_axi4_0_aw_bits_len;
  wire [2:0] system_front_port_axi4_0_aw_bits_size;
  wire [1:0] system_front_port_axi4_0_aw_bits_burst;
  wire  system_front_port_axi4_0_aw_bits_lock;
  wire [3:0] system_front_port_axi4_0_aw_bits_cache;
  wire [2:0] system_front_port_axi4_0_aw_bits_prot;
  wire [3:0] system_front_port_axi4_0_aw_bits_qos;
  wire  system_front_port_axi4_0_w_ready;
  wire  system_front_port_axi4_0_w_valid;
  wire [31:0] system_front_port_axi4_0_w_bits_data;
  wire [3:0] system_front_port_axi4_0_w_bits_strb;
  wire  system_front_port_axi4_0_w_bits_last;
  wire  system_front_port_axi4_0_b_ready;
  wire  system_front_port_axi4_0_b_valid;
  wire [7:0] system_front_port_axi4_0_b_bits_id;
  wire [1:0] system_front_port_axi4_0_b_bits_resp;
  wire  system_front_port_axi4_0_ar_ready;
  wire  system_front_port_axi4_0_ar_valid;
  wire [7:0] system_front_port_axi4_0_ar_bits_id;
  wire [31:0] system_front_port_axi4_0_ar_bits_addr;
  wire [7:0] system_front_port_axi4_0_ar_bits_len;
  wire [2:0] system_front_port_axi4_0_ar_bits_size;
  wire [1:0] system_front_port_axi4_0_ar_bits_burst;
  wire  system_front_port_axi4_0_ar_bits_lock;
  wire [3:0] system_front_port_axi4_0_ar_bits_cache;
  wire [2:0] system_front_port_axi4_0_ar_bits_prot;
  wire [3:0] system_front_port_axi4_0_ar_bits_qos;
  wire  system_front_port_axi4_0_r_ready;
  wire  system_front_port_axi4_0_r_valid;
  wire [7:0] system_front_port_axi4_0_r_bits_id;
  wire [31:0] system_front_port_axi4_0_r_bits_data;
  wire [1:0] system_front_port_axi4_0_r_bits_resp;
  wire  system_front_port_axi4_0_r_bits_last;
  wire  func_clock_clock;
  wire  func_clock_io_clock_out;
  wire  ClockSkew_clkin;
  wire  ClockSkew_clkout;
  wire  Pow2ClockDivider_clock;
  wire  Pow2ClockDivider_io_clock_out;
  wire  dpiClockGate_clock_in;
  wire  dpiClockGate_clock_out;
  wire  c_core_reset_driver_clock;
  wire  DataTap_5__1_clock;
  wire  DataTap_5__1_reset;
  wire [31:0] DataTap_5__1_hartid;
  wire [31:0] DataTap_5__1_timer;
  wire  DataTap_5__1_valid;
  wire [31:0] DataTap_5__1_pc;
  wire [4:0] DataTap_5__1_wrdst;
  wire [31:0] DataTap_5__1_wrdata;
  wire  DataTap_5__1_wren;
  wire [4:0] DataTap_5__1_rd0src;
  wire [31:0] DataTap_5__1_rd0val;
  wire [4:0] DataTap_5__1_rd1src;
  wire [31:0] DataTap_5__1_rd1val;
  wire [31:0] DataTap_5__1_inst;
  wire  DataTap_5__0_clock;
  wire  DataTap_5__0_reset;
  wire [31:0] DataTap_5__0_hartid;
  wire [31:0] DataTap_5__0_timer;
  wire  DataTap_5__0_valid;
  wire [31:0] DataTap_5__0_pc;
  wire [4:0] DataTap_5__0_wrdst;
  wire [31:0] DataTap_5__0_wrdata;
  wire  DataTap_5__0_wren;
  wire [4:0] DataTap_5__0_rd0src;
  wire [31:0] DataTap_5__0_rd0val;
  wire [4:0] DataTap_5__0_rd1src;
  wire [31:0] DataTap_5__0_rd1val;
  wire [31:0] DataTap_5__0_inst;
  wire  testRAM_clock;
  wire  testRAM_reset;
  wire  testRAM_io_axi4_0_aw_ready;
  wire  testRAM_io_axi4_0_aw_valid;
  wire  testRAM_io_axi4_0_aw_bits_id;
  wire [29:0] testRAM_io_axi4_0_aw_bits_addr;
  wire [7:0] testRAM_io_axi4_0_aw_bits_len;
  wire [2:0] testRAM_io_axi4_0_aw_bits_size;
  wire [1:0] testRAM_io_axi4_0_aw_bits_burst;
  wire  testRAM_io_axi4_0_aw_bits_lock;
  wire [3:0] testRAM_io_axi4_0_aw_bits_cache;
  wire [2:0] testRAM_io_axi4_0_aw_bits_prot;
  wire [3:0] testRAM_io_axi4_0_aw_bits_qos;
  wire  testRAM_io_axi4_0_w_ready;
  wire  testRAM_io_axi4_0_w_valid;
  wire [31:0] testRAM_io_axi4_0_w_bits_data;
  wire [3:0] testRAM_io_axi4_0_w_bits_strb;
  wire  testRAM_io_axi4_0_w_bits_last;
  wire  testRAM_io_axi4_0_b_ready;
  wire  testRAM_io_axi4_0_b_valid;
  wire  testRAM_io_axi4_0_b_bits_id;
  wire [1:0] testRAM_io_axi4_0_b_bits_resp;
  wire  testRAM_io_axi4_0_ar_ready;
  wire  testRAM_io_axi4_0_ar_valid;
  wire  testRAM_io_axi4_0_ar_bits_id;
  wire [29:0] testRAM_io_axi4_0_ar_bits_addr;
  wire [7:0] testRAM_io_axi4_0_ar_bits_len;
  wire [2:0] testRAM_io_axi4_0_ar_bits_size;
  wire [1:0] testRAM_io_axi4_0_ar_bits_burst;
  wire  testRAM_io_axi4_0_ar_bits_lock;
  wire [3:0] testRAM_io_axi4_0_ar_bits_cache;
  wire [2:0] testRAM_io_axi4_0_ar_bits_prot;
  wire [3:0] testRAM_io_axi4_0_ar_bits_qos;
  wire  testRAM_io_axi4_0_r_ready;
  wire  testRAM_io_axi4_0_r_valid;
  wire  testRAM_io_axi4_0_r_bits_id;
  wire [31:0] testRAM_io_axi4_0_r_bits_data;
  wire [1:0] testRAM_io_axi4_0_r_bits_resp;
  wire  testRAM_io_axi4_0_r_bits_last;
  wire  testRAM_1_clock;
  wire  testRAM_1_reset;
  wire  testRAM_1_io_axi4_0_aw_ready;
  wire  testRAM_1_io_axi4_0_aw_valid;
  wire [3:0] testRAM_1_io_axi4_0_aw_bits_id;
  wire [30:0] testRAM_1_io_axi4_0_aw_bits_addr;
  wire [7:0] testRAM_1_io_axi4_0_aw_bits_len;
  wire [2:0] testRAM_1_io_axi4_0_aw_bits_size;
  wire [1:0] testRAM_1_io_axi4_0_aw_bits_burst;
  wire  testRAM_1_io_axi4_0_aw_bits_lock;
  wire [3:0] testRAM_1_io_axi4_0_aw_bits_cache;
  wire [2:0] testRAM_1_io_axi4_0_aw_bits_prot;
  wire [3:0] testRAM_1_io_axi4_0_aw_bits_qos;
  wire  testRAM_1_io_axi4_0_w_ready;
  wire  testRAM_1_io_axi4_0_w_valid;
  wire [31:0] testRAM_1_io_axi4_0_w_bits_data;
  wire [3:0] testRAM_1_io_axi4_0_w_bits_strb;
  wire  testRAM_1_io_axi4_0_w_bits_last;
  wire  testRAM_1_io_axi4_0_b_ready;
  wire  testRAM_1_io_axi4_0_b_valid;
  wire [3:0] testRAM_1_io_axi4_0_b_bits_id;
  wire [1:0] testRAM_1_io_axi4_0_b_bits_resp;
  wire  testRAM_1_io_axi4_0_ar_ready;
  wire  testRAM_1_io_axi4_0_ar_valid;
  wire [3:0] testRAM_1_io_axi4_0_ar_bits_id;
  wire [30:0] testRAM_1_io_axi4_0_ar_bits_addr;
  wire [7:0] testRAM_1_io_axi4_0_ar_bits_len;
  wire [2:0] testRAM_1_io_axi4_0_ar_bits_size;
  wire [1:0] testRAM_1_io_axi4_0_ar_bits_burst;
  wire  testRAM_1_io_axi4_0_ar_bits_lock;
  wire [3:0] testRAM_1_io_axi4_0_ar_bits_cache;
  wire [2:0] testRAM_1_io_axi4_0_ar_bits_prot;
  wire [3:0] testRAM_1_io_axi4_0_ar_bits_qos;
  wire  testRAM_1_io_axi4_0_r_ready;
  wire  testRAM_1_io_axi4_0_r_valid;
  wire [3:0] testRAM_1_io_axi4_0_r_bits_id;
  wire [31:0] testRAM_1_io_axi4_0_r_bits_data;
  wire [1:0] testRAM_1_io_axi4_0_r_bits_resp;
  wire  testRAM_1_io_axi4_0_r_bits_last;
  wire  testRAM_2_clock;
  wire  testRAM_2_reset;
  wire  testRAM_2_io_axi4_0_aw_ready;
  wire  testRAM_2_io_axi4_0_aw_valid;
  wire [3:0] testRAM_2_io_axi4_0_aw_bits_id;
  wire [31:0] testRAM_2_io_axi4_0_aw_bits_addr;
  wire [7:0] testRAM_2_io_axi4_0_aw_bits_len;
  wire [2:0] testRAM_2_io_axi4_0_aw_bits_size;
  wire [1:0] testRAM_2_io_axi4_0_aw_bits_burst;
  wire  testRAM_2_io_axi4_0_aw_bits_lock;
  wire [3:0] testRAM_2_io_axi4_0_aw_bits_cache;
  wire [2:0] testRAM_2_io_axi4_0_aw_bits_prot;
  wire [3:0] testRAM_2_io_axi4_0_aw_bits_qos;
  wire  testRAM_2_io_axi4_0_w_ready;
  wire  testRAM_2_io_axi4_0_w_valid;
  wire [63:0] testRAM_2_io_axi4_0_w_bits_data;
  wire [7:0] testRAM_2_io_axi4_0_w_bits_strb;
  wire  testRAM_2_io_axi4_0_w_bits_last;
  wire  testRAM_2_io_axi4_0_b_ready;
  wire  testRAM_2_io_axi4_0_b_valid;
  wire [3:0] testRAM_2_io_axi4_0_b_bits_id;
  wire [1:0] testRAM_2_io_axi4_0_b_bits_resp;
  wire  testRAM_2_io_axi4_0_ar_ready;
  wire  testRAM_2_io_axi4_0_ar_valid;
  wire [3:0] testRAM_2_io_axi4_0_ar_bits_id;
  wire [31:0] testRAM_2_io_axi4_0_ar_bits_addr;
  wire [7:0] testRAM_2_io_axi4_0_ar_bits_len;
  wire [2:0] testRAM_2_io_axi4_0_ar_bits_size;
  wire [1:0] testRAM_2_io_axi4_0_ar_bits_burst;
  wire  testRAM_2_io_axi4_0_ar_bits_lock;
  wire [3:0] testRAM_2_io_axi4_0_ar_bits_cache;
  wire [2:0] testRAM_2_io_axi4_0_ar_bits_prot;
  wire [3:0] testRAM_2_io_axi4_0_ar_bits_qos;
  wire  testRAM_2_io_axi4_0_r_ready;
  wire  testRAM_2_io_axi4_0_r_valid;
  wire [3:0] testRAM_2_io_axi4_0_r_bits_id;
  wire [63:0] testRAM_2_io_axi4_0_r_bits_data;
  wire [1:0] testRAM_2_io_axi4_0_r_bits_resp;
  wire  testRAM_2_io_axi4_0_r_bits_last;
  wire  DPIJTAGDriver_clock;
  wire  DPIJTAGDriver_reset;
  wire  DPIJTAGDriver_jtag_TRSTn;
  wire  DPIJTAGDriver_jtag_TCK;
  wire  DPIJTAGDriver_jtag_TMS;
  wire  DPIJTAGDriver_jtag_TDI;
  wire  DPIJTAGDriver_jtag_TDO_data;
  wire  DPIJTAGDriver_jtag_TDO_driven;
  wire  system_reset_driver_clock;
  wire  system_reset_driver_out;
  wire [31:0] plusarg_reader_out;
  wire  CountAndDriver_clock;
  wire  CountAndDriver_reset;
  wire  CountAndDriver_io_default_value;
  wire [15:0] CountAndDriver_io_count;
  wire  CountAndDriver_io_driven_value;
  wire  core_reset_driver_clock;
  wire  core_monitor_m_0_clock;
  wire  core_monitor_m_0_reset;
  wire [31:0] core_monitor_m_0_hartid;
  wire [31:0] core_monitor_m_0_timer;
  wire  core_monitor_m_0_valid;
  wire [31:0] core_monitor_m_0_pc;
  wire [4:0] core_monitor_m_0_wrdst;
  wire [31:0] core_monitor_m_0_wrdata;
  wire  core_monitor_m_0_wren;
  wire [4:0] core_monitor_m_0_rd0src;
  wire [31:0] core_monitor_m_0_rd0val;
  wire [4:0] core_monitor_m_0_rd1src;
  wire [31:0] core_monitor_m_0_rd1val;
  wire [31:0] core_monitor_m_0_inst;
  wire  core_monitor_m_1_clock;
  wire  core_monitor_m_1_reset;
  wire [31:0] core_monitor_m_1_hartid;
  wire [31:0] core_monitor_m_1_timer;
  wire  core_monitor_m_1_valid;
  wire [31:0] core_monitor_m_1_pc;
  wire [4:0] core_monitor_m_1_wrdst;
  wire [31:0] core_monitor_m_1_wrdata;
  wire  core_monitor_m_1_wren;
  wire [4:0] core_monitor_m_1_rd0src;
  wire [31:0] core_monitor_m_1_rd0val;
  wire [4:0] core_monitor_m_1_rd1src;
  wire [31:0] core_monitor_m_1_rd1val;
  wire [31:0] core_monitor_m_1_inst;
  wire [31:0] plusarg_reader_1_out;
  wire  InterruptsDriver_clock;
  wire  InterruptsDriver_reset;
  wire  dpitbh_clock;
  wire  dpitbh_reset;
  wire [31:0] plusarg_reader_2_out;
  reg [4:0] _T;
  reg [31:0] _RAND_0;
  reg  _T_1;
  reg [31:0] _RAND_1;
  wire [4:0] _T_3;
  wire  _T_4;
  wire  _T_5;
  wire  _T_14;
  wire  ndm_reset;
  wire  _T_28;
  wire [31:0] _T_30;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_39;
  wire  _T_43;
  reg [6:0] value_1;
  reg [31:0] _RAND_2;
  wire  _T_45;
  wire [6:0] _T_47;
  wire [31:0] _T_44;
  wire  _T_48;
  wire  _T_49;
  wire  _T_51;
  wire  _T_179;
  reg [6:0] value_2;
  reg [31:0] _RAND_3;
  wire  _T_180;
  wire [6:0] _T_182;
  wire [127:0] _T_184;
  wire  _T_185;
  reg [15:0] _T_186;
  reg [31:0] _RAND_4;
  wire  _T_187;
  wire  _T_188;
  wire  _T_189;
  wire  _T_190;
  wire  _T_191;
  wire  _T_192;
  wire  _T_193;
  wire  _T_194;
  wire [14:0] _T_195;
  wire [15:0] _T_196;
  reg [15:0] _T_198;
  reg [31:0] _RAND_5;
  wire  _T_199;
  wire  _T_200;
  wire  _T_201;
  wire  _T_202;
  wire  _T_203;
  wire  _T_204;
  wire  _T_205;
  wire  _T_206;
  wire [14:0] _T_207;
  wire [15:0] _T_208;
  reg [15:0] _T_210;
  reg [31:0] _RAND_6;
  wire  _T_211;
  wire  _T_212;
  wire  _T_213;
  wire  _T_214;
  wire  _T_215;
  wire  _T_216;
  wire  _T_217;
  wire  _T_218;
  wire [14:0] _T_219;
  wire [15:0] _T_220;
  reg [15:0] _T_222;
  reg [31:0] _RAND_7;
  wire  _T_223;
  wire  _T_224;
  wire  _T_225;
  wire  _T_226;
  wire  _T_227;
  wire  _T_228;
  wire  _T_229;
  wire  _T_230;
  wire [14:0] _T_231;
  wire [15:0] _T_232;
  reg [15:0] _T_234;
  reg [31:0] _RAND_8;
  wire  _T_235;
  wire  _T_236;
  wire  _T_237;
  wire  _T_238;
  wire  _T_239;
  wire  _T_240;
  wire  _T_241;
  wire  _T_242;
  wire [14:0] _T_243;
  wire [15:0] _T_244;
  reg [15:0] _T_246;
  reg [31:0] _RAND_9;
  wire  _T_247;
  wire  _T_248;
  wire  _T_249;
  wire  _T_250;
  wire  _T_251;
  wire  _T_252;
  wire  _T_253;
  wire  _T_254;
  wire [14:0] _T_255;
  wire [15:0] _T_256;
  reg [15:0] _T_258;
  reg [31:0] _RAND_10;
  wire  _T_259;
  wire  _T_260;
  wire  _T_261;
  wire  _T_262;
  wire  _T_263;
  wire  _T_264;
  wire  _T_265;
  wire  _T_266;
  wire [14:0] _T_267;
  wire [15:0] _T_268;
  reg [15:0] _T_270;
  reg [31:0] _RAND_11;
  wire  _T_271;
  wire  _T_272;
  wire  _T_273;
  wire  _T_274;
  wire  _T_275;
  wire  _T_276;
  wire  _T_277;
  wire  _T_278;
  wire [14:0] _T_279;
  wire [15:0] _T_280;
  reg [15:0] _T_282;
  reg [31:0] _RAND_12;
  wire  _T_283;
  wire  _T_284;
  wire  _T_285;
  wire  _T_286;
  wire  _T_287;
  wire  _T_288;
  wire  _T_289;
  wire  _T_290;
  wire [14:0] _T_291;
  wire [15:0] _T_292;
  reg [15:0] _T_294;
  reg [31:0] _RAND_13;
  wire  _T_295;
  wire  _T_296;
  wire  _T_297;
  wire  _T_298;
  wire  _T_299;
  wire  _T_300;
  wire  _T_301;
  wire  _T_302;
  wire [14:0] _T_303;
  wire [15:0] _T_304;
  reg [15:0] _T_306;
  reg [31:0] _RAND_14;
  wire  _T_307;
  wire  _T_308;
  wire  _T_309;
  wire  _T_310;
  wire  _T_311;
  wire  _T_312;
  wire  _T_313;
  wire  _T_314;
  wire [14:0] _T_315;
  wire [15:0] _T_316;
  reg [15:0] _T_318;
  reg [31:0] _RAND_15;
  wire  _T_319;
  wire  _T_320;
  wire  _T_321;
  wire  _T_322;
  wire  _T_323;
  wire  _T_324;
  wire  _T_325;
  wire  _T_326;
  wire [14:0] _T_327;
  wire [15:0] _T_328;
  reg [15:0] _T_330;
  reg [31:0] _RAND_16;
  wire  _T_331;
  wire  _T_332;
  wire  _T_333;
  wire  _T_334;
  wire  _T_335;
  wire  _T_336;
  wire  _T_337;
  wire  _T_338;
  wire [14:0] _T_339;
  wire [15:0] _T_340;
  reg [15:0] _T_342;
  reg [31:0] _RAND_17;
  wire  _T_343;
  wire  _T_344;
  wire  _T_345;
  wire  _T_346;
  wire  _T_347;
  wire  _T_348;
  wire  _T_349;
  wire  _T_350;
  wire [14:0] _T_351;
  wire [15:0] _T_352;
  reg [15:0] _T_354;
  reg [31:0] _RAND_18;
  wire  _T_355;
  wire  _T_356;
  wire  _T_357;
  wire  _T_358;
  wire  _T_359;
  wire  _T_360;
  wire  _T_361;
  wire  _T_362;
  wire [14:0] _T_363;
  wire [15:0] _T_364;
  reg [15:0] _T_366;
  reg [31:0] _RAND_19;
  wire  _T_367;
  wire  _T_368;
  wire  _T_369;
  wire  _T_370;
  wire  _T_371;
  wire  _T_372;
  wire  _T_373;
  wire  _T_374;
  wire [14:0] _T_375;
  wire [15:0] _T_376;
  reg [15:0] _T_378;
  reg [31:0] _RAND_20;
  wire  _T_379;
  wire  _T_380;
  wire  _T_381;
  wire  _T_382;
  wire  _T_383;
  wire  _T_384;
  wire  _T_385;
  wire  _T_386;
  wire [14:0] _T_387;
  wire [15:0] _T_388;
  reg [15:0] _T_390;
  reg [31:0] _RAND_21;
  wire  _T_391;
  wire  _T_392;
  wire  _T_393;
  wire  _T_394;
  wire  _T_395;
  wire  _T_396;
  wire  _T_397;
  wire  _T_398;
  wire [14:0] _T_399;
  wire [15:0] _T_400;
  reg [15:0] _T_402;
  reg [31:0] _RAND_22;
  wire  _T_403;
  wire  _T_404;
  wire  _T_405;
  wire  _T_406;
  wire  _T_407;
  wire  _T_408;
  wire  _T_409;
  wire  _T_410;
  wire [14:0] _T_411;
  wire [15:0] _T_412;
  reg [15:0] _T_414;
  reg [31:0] _RAND_23;
  wire  _T_415;
  wire  _T_416;
  wire  _T_417;
  wire  _T_418;
  wire  _T_419;
  wire  _T_420;
  wire  _T_421;
  wire  _T_422;
  wire [14:0] _T_423;
  wire [15:0] _T_424;
  reg [15:0] _T_426;
  reg [31:0] _RAND_24;
  wire  _T_427;
  wire  _T_428;
  wire  _T_429;
  wire  _T_430;
  wire  _T_431;
  wire  _T_432;
  wire  _T_433;
  wire  _T_434;
  wire [14:0] _T_435;
  wire [15:0] _T_436;
  reg [15:0] _T_438;
  reg [31:0] _RAND_25;
  wire  _T_439;
  wire  _T_440;
  wire  _T_441;
  wire  _T_442;
  wire  _T_443;
  wire  _T_444;
  wire  _T_445;
  wire  _T_446;
  wire [14:0] _T_447;
  wire [15:0] _T_448;
  reg [15:0] _T_450;
  reg [31:0] _RAND_26;
  wire  _T_451;
  wire  _T_452;
  wire  _T_453;
  wire  _T_454;
  wire  _T_455;
  wire  _T_456;
  wire  _T_457;
  wire  _T_458;
  wire [14:0] _T_459;
  wire [15:0] _T_460;
  reg [15:0] _T_462;
  reg [31:0] _RAND_27;
  wire  _T_463;
  wire  _T_464;
  wire  _T_465;
  wire  _T_466;
  wire  _T_467;
  wire  _T_468;
  wire  _T_469;
  wire  _T_470;
  wire [14:0] _T_471;
  wire [15:0] _T_472;
  reg [15:0] _T_474;
  reg [31:0] _RAND_28;
  wire  _T_475;
  wire  _T_476;
  wire  _T_477;
  wire  _T_478;
  wire  _T_479;
  wire  _T_480;
  wire  _T_481;
  wire  _T_482;
  wire [14:0] _T_483;
  wire [15:0] _T_484;
  reg [15:0] _T_486;
  reg [31:0] _RAND_29;
  wire  _T_487;
  wire  _T_488;
  wire  _T_489;
  wire  _T_490;
  wire  _T_491;
  wire  _T_492;
  wire  _T_493;
  wire  _T_494;
  wire [14:0] _T_495;
  wire [15:0] _T_496;
  reg [15:0] _T_498;
  reg [31:0] _RAND_30;
  wire  _T_499;
  wire  _T_500;
  wire  _T_501;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_506;
  wire [14:0] _T_507;
  wire [15:0] _T_508;
  reg [15:0] _T_510;
  reg [31:0] _RAND_31;
  wire  _T_511;
  wire  _T_512;
  wire  _T_513;
  wire  _T_514;
  wire  _T_515;
  wire  _T_516;
  wire  _T_517;
  wire  _T_518;
  wire [14:0] _T_519;
  wire [15:0] _T_520;
  reg [15:0] _T_522;
  reg [31:0] _RAND_32;
  wire  _T_523;
  wire  _T_524;
  wire  _T_525;
  wire  _T_526;
  wire  _T_527;
  wire  _T_528;
  wire  _T_529;
  wire  _T_530;
  wire [14:0] _T_531;
  wire [15:0] _T_532;
  reg [15:0] _T_534;
  reg [31:0] _RAND_33;
  wire  _T_535;
  wire  _T_536;
  wire  _T_537;
  wire  _T_538;
  wire  _T_539;
  wire  _T_540;
  wire  _T_541;
  wire  _T_542;
  wire [14:0] _T_543;
  wire [15:0] _T_544;
  reg [15:0] _T_546;
  reg [31:0] _RAND_34;
  wire  _T_547;
  wire  _T_548;
  wire  _T_549;
  wire  _T_550;
  wire  _T_551;
  wire  _T_552;
  wire  _T_553;
  wire  _T_554;
  wire [14:0] _T_555;
  wire [15:0] _T_556;
  reg [15:0] _T_558;
  reg [31:0] _RAND_35;
  wire  _T_559;
  wire  _T_560;
  wire  _T_561;
  wire  _T_562;
  wire  _T_563;
  wire  _T_564;
  wire  _T_565;
  wire  _T_566;
  wire [14:0] _T_567;
  wire [15:0] _T_568;
  reg [15:0] _T_570;
  reg [31:0] _RAND_36;
  wire  _T_571;
  wire  _T_572;
  wire  _T_573;
  wire  _T_574;
  wire  _T_575;
  wire  _T_576;
  wire  _T_577;
  wire  _T_578;
  wire [14:0] _T_579;
  wire [15:0] _T_580;
  reg [15:0] _T_582;
  reg [31:0] _RAND_37;
  wire  _T_583;
  wire  _T_584;
  wire  _T_585;
  wire  _T_586;
  wire  _T_587;
  wire  _T_588;
  wire  _T_589;
  wire  _T_590;
  wire [14:0] _T_591;
  wire [15:0] _T_592;
  reg [15:0] _T_594;
  reg [31:0] _RAND_38;
  wire  _T_595;
  wire  _T_596;
  wire  _T_597;
  wire  _T_598;
  wire  _T_599;
  wire  _T_600;
  wire  _T_601;
  wire  _T_602;
  wire [14:0] _T_603;
  wire [15:0] _T_604;
  reg [15:0] _T_606;
  reg [31:0] _RAND_39;
  wire  _T_607;
  wire  _T_608;
  wire  _T_609;
  wire  _T_610;
  wire  _T_611;
  wire  _T_612;
  wire  _T_613;
  wire  _T_614;
  wire [14:0] _T_615;
  wire [15:0] _T_616;
  reg [15:0] _T_618;
  reg [31:0] _RAND_40;
  wire  _T_619;
  wire  _T_620;
  wire  _T_621;
  wire  _T_622;
  wire  _T_623;
  wire  _T_624;
  wire  _T_625;
  wire  _T_626;
  wire [14:0] _T_627;
  wire [15:0] _T_628;
  reg [15:0] _T_630;
  reg [31:0] _RAND_41;
  wire  _T_631;
  wire  _T_632;
  wire  _T_633;
  wire  _T_634;
  wire  _T_635;
  wire  _T_636;
  wire  _T_637;
  wire  _T_638;
  wire [14:0] _T_639;
  wire [15:0] _T_640;
  reg [15:0] _T_642;
  reg [31:0] _RAND_42;
  wire  _T_643;
  wire  _T_644;
  wire  _T_645;
  wire  _T_646;
  wire  _T_647;
  wire  _T_648;
  wire  _T_649;
  wire  _T_650;
  wire [14:0] _T_651;
  wire [15:0] _T_652;
  reg [15:0] _T_654;
  reg [31:0] _RAND_43;
  wire  _T_655;
  wire  _T_656;
  wire  _T_657;
  wire  _T_658;
  wire  _T_659;
  wire  _T_660;
  wire  _T_661;
  wire  _T_662;
  wire [14:0] _T_663;
  wire [15:0] _T_664;
  reg [15:0] _T_666;
  reg [31:0] _RAND_44;
  wire  _T_667;
  wire  _T_668;
  wire  _T_669;
  wire  _T_670;
  wire  _T_671;
  wire  _T_672;
  wire  _T_673;
  wire  _T_674;
  wire [14:0] _T_675;
  wire [15:0] _T_676;
  reg [15:0] _T_678;
  reg [31:0] _RAND_45;
  wire  _T_679;
  wire  _T_680;
  wire  _T_681;
  wire  _T_682;
  wire  _T_683;
  wire  _T_684;
  wire  _T_685;
  wire  _T_686;
  wire [14:0] _T_687;
  wire [15:0] _T_688;
  reg [15:0] _T_690;
  reg [31:0] _RAND_46;
  wire  _T_691;
  wire  _T_692;
  wire  _T_693;
  wire  _T_694;
  wire  _T_695;
  wire  _T_696;
  wire  _T_697;
  wire  _T_698;
  wire [14:0] _T_699;
  wire [15:0] _T_700;
  reg [15:0] _T_702;
  reg [31:0] _RAND_47;
  wire  _T_703;
  wire  _T_704;
  wire  _T_705;
  wire  _T_706;
  wire  _T_707;
  wire  _T_708;
  wire  _T_709;
  wire  _T_710;
  wire [14:0] _T_711;
  wire [15:0] _T_712;
  reg [15:0] _T_714;
  reg [31:0] _RAND_48;
  wire  _T_715;
  wire  _T_716;
  wire  _T_717;
  wire  _T_718;
  wire  _T_719;
  wire  _T_720;
  wire  _T_721;
  wire  _T_722;
  wire [14:0] _T_723;
  wire [15:0] _T_724;
  reg [15:0] _T_726;
  reg [31:0] _RAND_49;
  wire  _T_727;
  wire  _T_728;
  wire  _T_729;
  wire  _T_730;
  wire  _T_731;
  wire  _T_732;
  wire  _T_733;
  wire  _T_734;
  wire [14:0] _T_735;
  wire [15:0] _T_736;
  reg [15:0] _T_738;
  reg [31:0] _RAND_50;
  wire  _T_739;
  wire  _T_740;
  wire  _T_741;
  wire  _T_742;
  wire  _T_743;
  wire  _T_744;
  wire  _T_745;
  wire  _T_746;
  wire [14:0] _T_747;
  wire [15:0] _T_748;
  reg [15:0] _T_750;
  reg [31:0] _RAND_51;
  wire  _T_751;
  wire  _T_752;
  wire  _T_753;
  wire  _T_754;
  wire  _T_755;
  wire  _T_756;
  wire  _T_757;
  wire  _T_758;
  wire [14:0] _T_759;
  wire [15:0] _T_760;
  reg [15:0] _T_762;
  reg [31:0] _RAND_52;
  wire  _T_763;
  wire  _T_764;
  wire  _T_765;
  wire  _T_766;
  wire  _T_767;
  wire  _T_768;
  wire  _T_769;
  wire  _T_770;
  wire [14:0] _T_771;
  wire [15:0] _T_772;
  reg [15:0] _T_774;
  reg [31:0] _RAND_53;
  wire  _T_775;
  wire  _T_776;
  wire  _T_777;
  wire  _T_778;
  wire  _T_779;
  wire  _T_780;
  wire  _T_781;
  wire  _T_782;
  wire [14:0] _T_783;
  wire [15:0] _T_784;
  reg [15:0] _T_786;
  reg [31:0] _RAND_54;
  wire  _T_787;
  wire  _T_788;
  wire  _T_789;
  wire  _T_790;
  wire  _T_791;
  wire  _T_792;
  wire  _T_793;
  wire  _T_794;
  wire [14:0] _T_795;
  wire [15:0] _T_796;
  reg [15:0] _T_798;
  reg [31:0] _RAND_55;
  wire  _T_799;
  wire  _T_800;
  wire  _T_801;
  wire  _T_802;
  wire  _T_803;
  wire  _T_804;
  wire  _T_805;
  wire  _T_806;
  wire [14:0] _T_807;
  wire [15:0] _T_808;
  reg [15:0] _T_810;
  reg [31:0] _RAND_56;
  wire  _T_811;
  wire  _T_812;
  wire  _T_813;
  wire  _T_814;
  wire  _T_815;
  wire  _T_816;
  wire  _T_817;
  wire  _T_818;
  wire [14:0] _T_819;
  wire [15:0] _T_820;
  reg [15:0] _T_822;
  reg [31:0] _RAND_57;
  wire  _T_823;
  wire  _T_824;
  wire  _T_825;
  wire  _T_826;
  wire  _T_827;
  wire  _T_828;
  wire  _T_829;
  wire  _T_830;
  wire [14:0] _T_831;
  wire [15:0] _T_832;
  reg [15:0] _T_834;
  reg [31:0] _RAND_58;
  wire  _T_835;
  wire  _T_836;
  wire  _T_837;
  wire  _T_838;
  wire  _T_839;
  wire  _T_840;
  wire  _T_841;
  wire  _T_842;
  wire [14:0] _T_843;
  wire [15:0] _T_844;
  reg [15:0] _T_846;
  reg [31:0] _RAND_59;
  wire  _T_847;
  wire  _T_848;
  wire  _T_849;
  wire  _T_850;
  wire  _T_851;
  wire  _T_852;
  wire  _T_853;
  wire  _T_854;
  wire [14:0] _T_855;
  wire [15:0] _T_856;
  reg [15:0] _T_858;
  reg [31:0] _RAND_60;
  wire  _T_859;
  wire  _T_860;
  wire  _T_861;
  wire  _T_862;
  wire  _T_863;
  wire  _T_864;
  wire  _T_865;
  wire  _T_866;
  wire [14:0] _T_867;
  wire [15:0] _T_868;
  reg [15:0] _T_870;
  reg [31:0] _RAND_61;
  wire  _T_871;
  wire  _T_872;
  wire  _T_873;
  wire  _T_874;
  wire  _T_875;
  wire  _T_876;
  wire  _T_877;
  wire  _T_878;
  wire [14:0] _T_879;
  wire [15:0] _T_880;
  reg [15:0] _T_882;
  reg [31:0] _RAND_62;
  wire  _T_883;
  wire  _T_884;
  wire  _T_885;
  wire  _T_886;
  wire  _T_887;
  wire  _T_888;
  wire  _T_889;
  wire  _T_890;
  wire [14:0] _T_891;
  wire [15:0] _T_892;
  reg [15:0] _T_894;
  reg [31:0] _RAND_63;
  wire  _T_895;
  wire  _T_896;
  wire  _T_897;
  wire  _T_898;
  wire  _T_899;
  wire  _T_900;
  wire  _T_901;
  wire  _T_902;
  wire [14:0] _T_903;
  wire [15:0] _T_904;
  reg [15:0] _T_906;
  reg [31:0] _RAND_64;
  wire  _T_907;
  wire  _T_908;
  wire  _T_909;
  wire  _T_910;
  wire  _T_911;
  wire  _T_912;
  wire  _T_913;
  wire  _T_914;
  wire [14:0] _T_915;
  wire [15:0] _T_916;
  reg [15:0] _T_918;
  reg [31:0] _RAND_65;
  wire  _T_919;
  wire  _T_920;
  wire  _T_921;
  wire  _T_922;
  wire  _T_923;
  wire  _T_924;
  wire  _T_925;
  wire  _T_926;
  wire [14:0] _T_927;
  wire [15:0] _T_928;
  reg [15:0] _T_930;
  reg [31:0] _RAND_66;
  wire  _T_931;
  wire  _T_932;
  wire  _T_933;
  wire  _T_934;
  wire  _T_935;
  wire  _T_936;
  wire  _T_937;
  wire  _T_938;
  wire [14:0] _T_939;
  wire [15:0] _T_940;
  reg [15:0] _T_942;
  reg [31:0] _RAND_67;
  wire  _T_943;
  wire  _T_944;
  wire  _T_945;
  wire  _T_946;
  wire  _T_947;
  wire  _T_948;
  wire  _T_949;
  wire  _T_950;
  wire [14:0] _T_951;
  wire [15:0] _T_952;
  reg [15:0] _T_954;
  reg [31:0] _RAND_68;
  wire  _T_955;
  wire  _T_956;
  wire  _T_957;
  wire  _T_958;
  wire  _T_959;
  wire  _T_960;
  wire  _T_961;
  wire  _T_962;
  wire [14:0] _T_963;
  wire [15:0] _T_964;
  reg [15:0] _T_966;
  reg [31:0] _RAND_69;
  wire  _T_967;
  wire  _T_968;
  wire  _T_969;
  wire  _T_970;
  wire  _T_971;
  wire  _T_972;
  wire  _T_973;
  wire  _T_974;
  wire [14:0] _T_975;
  wire [15:0] _T_976;
  reg [15:0] _T_978;
  reg [31:0] _RAND_70;
  wire  _T_979;
  wire  _T_980;
  wire  _T_981;
  wire  _T_982;
  wire  _T_983;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire [14:0] _T_987;
  wire [15:0] _T_988;
  reg [15:0] _T_990;
  reg [31:0] _RAND_71;
  wire  _T_991;
  wire  _T_992;
  wire  _T_993;
  wire  _T_994;
  wire  _T_995;
  wire  _T_996;
  wire  _T_997;
  wire  _T_998;
  wire [14:0] _T_999;
  wire [15:0] _T_1000;
  reg [15:0] _T_1002;
  reg [31:0] _RAND_72;
  wire  _T_1003;
  wire  _T_1004;
  wire  _T_1005;
  wire  _T_1006;
  wire  _T_1007;
  wire  _T_1008;
  wire  _T_1009;
  wire  _T_1010;
  wire [14:0] _T_1011;
  wire [15:0] _T_1012;
  reg [15:0] _T_1014;
  reg [31:0] _RAND_73;
  wire  _T_1015;
  wire  _T_1016;
  wire  _T_1017;
  wire  _T_1018;
  wire  _T_1019;
  wire  _T_1020;
  wire  _T_1021;
  wire  _T_1022;
  wire [14:0] _T_1023;
  wire [15:0] _T_1024;
  reg [15:0] _T_1026;
  reg [31:0] _RAND_74;
  wire  _T_1027;
  wire  _T_1028;
  wire  _T_1029;
  wire  _T_1030;
  wire  _T_1031;
  wire  _T_1032;
  wire  _T_1033;
  wire  _T_1034;
  wire [14:0] _T_1035;
  wire [15:0] _T_1036;
  reg [15:0] _T_1038;
  reg [31:0] _RAND_75;
  wire  _T_1039;
  wire  _T_1040;
  wire  _T_1041;
  wire  _T_1042;
  wire  _T_1043;
  wire  _T_1044;
  wire  _T_1045;
  wire  _T_1046;
  wire [14:0] _T_1047;
  wire [15:0] _T_1048;
  reg [15:0] _T_1050;
  reg [31:0] _RAND_76;
  wire  _T_1051;
  wire  _T_1052;
  wire  _T_1053;
  wire  _T_1054;
  wire  _T_1055;
  wire  _T_1056;
  wire  _T_1057;
  wire  _T_1058;
  wire [14:0] _T_1059;
  wire [15:0] _T_1060;
  reg [15:0] _T_1062;
  reg [31:0] _RAND_77;
  wire  _T_1063;
  wire  _T_1064;
  wire  _T_1065;
  wire  _T_1066;
  wire  _T_1067;
  wire  _T_1068;
  wire  _T_1069;
  wire  _T_1070;
  wire [14:0] _T_1071;
  wire [15:0] _T_1072;
  reg [15:0] _T_1074;
  reg [31:0] _RAND_78;
  wire  _T_1075;
  wire  _T_1076;
  wire  _T_1077;
  wire  _T_1078;
  wire  _T_1079;
  wire  _T_1080;
  wire  _T_1081;
  wire  _T_1082;
  wire [14:0] _T_1083;
  wire [15:0] _T_1084;
  reg [15:0] _T_1086;
  reg [31:0] _RAND_79;
  wire  _T_1087;
  wire  _T_1088;
  wire  _T_1089;
  wire  _T_1090;
  wire  _T_1091;
  wire  _T_1092;
  wire  _T_1093;
  wire  _T_1094;
  wire [14:0] _T_1095;
  wire [15:0] _T_1096;
  reg [15:0] _T_1098;
  reg [31:0] _RAND_80;
  wire  _T_1099;
  wire  _T_1100;
  wire  _T_1101;
  wire  _T_1102;
  wire  _T_1103;
  wire  _T_1104;
  wire  _T_1105;
  wire  _T_1106;
  wire [14:0] _T_1107;
  wire [15:0] _T_1108;
  reg [15:0] _T_1110;
  reg [31:0] _RAND_81;
  wire  _T_1111;
  wire  _T_1112;
  wire  _T_1113;
  wire  _T_1114;
  wire  _T_1115;
  wire  _T_1116;
  wire  _T_1117;
  wire  _T_1118;
  wire [14:0] _T_1119;
  wire [15:0] _T_1120;
  reg [15:0] _T_1122;
  reg [31:0] _RAND_82;
  wire  _T_1123;
  wire  _T_1124;
  wire  _T_1125;
  wire  _T_1126;
  wire  _T_1127;
  wire  _T_1128;
  wire  _T_1129;
  wire  _T_1130;
  wire [14:0] _T_1131;
  wire [15:0] _T_1132;
  reg [15:0] _T_1134;
  reg [31:0] _RAND_83;
  wire  _T_1135;
  wire  _T_1136;
  wire  _T_1137;
  wire  _T_1138;
  wire  _T_1139;
  wire  _T_1140;
  wire  _T_1141;
  wire  _T_1142;
  wire [14:0] _T_1143;
  wire [15:0] _T_1144;
  reg [15:0] _T_1146;
  reg [31:0] _RAND_84;
  wire  _T_1147;
  wire  _T_1148;
  wire  _T_1149;
  wire  _T_1150;
  wire  _T_1151;
  wire  _T_1152;
  wire  _T_1153;
  wire  _T_1154;
  wire [14:0] _T_1155;
  wire [15:0] _T_1156;
  reg [15:0] _T_1158;
  reg [31:0] _RAND_85;
  wire  _T_1159;
  wire  _T_1160;
  wire  _T_1161;
  wire  _T_1162;
  wire  _T_1163;
  wire  _T_1164;
  wire  _T_1165;
  wire  _T_1166;
  wire [14:0] _T_1167;
  wire [15:0] _T_1168;
  reg [15:0] _T_1170;
  reg [31:0] _RAND_86;
  wire  _T_1171;
  wire  _T_1172;
  wire  _T_1173;
  wire  _T_1174;
  wire  _T_1175;
  wire  _T_1176;
  wire  _T_1177;
  wire  _T_1178;
  wire [14:0] _T_1179;
  wire [15:0] _T_1180;
  reg [15:0] _T_1182;
  reg [31:0] _RAND_87;
  wire  _T_1183;
  wire  _T_1184;
  wire  _T_1185;
  wire  _T_1186;
  wire  _T_1187;
  wire  _T_1188;
  wire  _T_1189;
  wire  _T_1190;
  wire [14:0] _T_1191;
  wire [15:0] _T_1192;
  reg [15:0] _T_1194;
  reg [31:0] _RAND_88;
  wire  _T_1195;
  wire  _T_1196;
  wire  _T_1197;
  wire  _T_1198;
  wire  _T_1199;
  wire  _T_1200;
  wire  _T_1201;
  wire  _T_1202;
  wire [14:0] _T_1203;
  wire [15:0] _T_1204;
  reg [15:0] _T_1206;
  reg [31:0] _RAND_89;
  wire  _T_1207;
  wire  _T_1208;
  wire  _T_1209;
  wire  _T_1210;
  wire  _T_1211;
  wire  _T_1212;
  wire  _T_1213;
  wire  _T_1214;
  wire [14:0] _T_1215;
  wire [15:0] _T_1216;
  reg [15:0] _T_1218;
  reg [31:0] _RAND_90;
  wire  _T_1219;
  wire  _T_1220;
  wire  _T_1221;
  wire  _T_1222;
  wire  _T_1223;
  wire  _T_1224;
  wire  _T_1225;
  wire  _T_1226;
  wire [14:0] _T_1227;
  wire [15:0] _T_1228;
  reg [15:0] _T_1230;
  reg [31:0] _RAND_91;
  wire  _T_1231;
  wire  _T_1232;
  wire  _T_1233;
  wire  _T_1234;
  wire  _T_1235;
  wire  _T_1236;
  wire  _T_1237;
  wire  _T_1238;
  wire [14:0] _T_1239;
  wire [15:0] _T_1240;
  reg [15:0] _T_1242;
  reg [31:0] _RAND_92;
  wire  _T_1243;
  wire  _T_1244;
  wire  _T_1245;
  wire  _T_1246;
  wire  _T_1247;
  wire  _T_1248;
  wire  _T_1249;
  wire  _T_1250;
  wire [14:0] _T_1251;
  wire [15:0] _T_1252;
  reg [15:0] _T_1254;
  reg [31:0] _RAND_93;
  wire  _T_1255;
  wire  _T_1256;
  wire  _T_1257;
  wire  _T_1258;
  wire  _T_1259;
  wire  _T_1260;
  wire  _T_1261;
  wire  _T_1262;
  wire [14:0] _T_1263;
  wire [15:0] _T_1264;
  reg [15:0] _T_1266;
  reg [31:0] _RAND_94;
  wire  _T_1267;
  wire  _T_1268;
  wire  _T_1269;
  wire  _T_1270;
  wire  _T_1271;
  wire  _T_1272;
  wire  _T_1273;
  wire  _T_1274;
  wire [14:0] _T_1275;
  wire [15:0] _T_1276;
  reg [15:0] _T_1278;
  reg [31:0] _RAND_95;
  wire  _T_1279;
  wire  _T_1280;
  wire  _T_1281;
  wire  _T_1282;
  wire  _T_1283;
  wire  _T_1284;
  wire  _T_1285;
  wire  _T_1286;
  wire [14:0] _T_1287;
  wire [15:0] _T_1288;
  reg [15:0] _T_1290;
  reg [31:0] _RAND_96;
  wire  _T_1291;
  wire  _T_1292;
  wire  _T_1293;
  wire  _T_1294;
  wire  _T_1295;
  wire  _T_1296;
  wire  _T_1297;
  wire  _T_1298;
  wire [14:0] _T_1299;
  wire [15:0] _T_1300;
  reg [15:0] _T_1302;
  reg [31:0] _RAND_97;
  wire  _T_1303;
  wire  _T_1304;
  wire  _T_1305;
  wire  _T_1306;
  wire  _T_1307;
  wire  _T_1308;
  wire  _T_1309;
  wire  _T_1310;
  wire [14:0] _T_1311;
  wire [15:0] _T_1312;
  reg [15:0] _T_1314;
  reg [31:0] _RAND_98;
  wire  _T_1315;
  wire  _T_1316;
  wire  _T_1317;
  wire  _T_1318;
  wire  _T_1319;
  wire  _T_1320;
  wire  _T_1321;
  wire  _T_1322;
  wire [14:0] _T_1323;
  wire [15:0] _T_1324;
  reg [15:0] _T_1326;
  reg [31:0] _RAND_99;
  wire  _T_1327;
  wire  _T_1328;
  wire  _T_1329;
  wire  _T_1330;
  wire  _T_1331;
  wire  _T_1332;
  wire  _T_1333;
  wire  _T_1334;
  wire [14:0] _T_1335;
  wire [15:0] _T_1336;
  reg [15:0] _T_1338;
  reg [31:0] _RAND_100;
  wire  _T_1339;
  wire  _T_1340;
  wire  _T_1341;
  wire  _T_1342;
  wire  _T_1343;
  wire  _T_1344;
  wire  _T_1345;
  wire  _T_1346;
  wire [14:0] _T_1347;
  wire [15:0] _T_1348;
  reg [15:0] _T_1350;
  reg [31:0] _RAND_101;
  wire  _T_1351;
  wire  _T_1352;
  wire  _T_1353;
  wire  _T_1354;
  wire  _T_1355;
  wire  _T_1356;
  wire  _T_1357;
  wire  _T_1358;
  wire [14:0] _T_1359;
  wire [15:0] _T_1360;
  reg [15:0] _T_1362;
  reg [31:0] _RAND_102;
  wire  _T_1363;
  wire  _T_1364;
  wire  _T_1365;
  wire  _T_1366;
  wire  _T_1367;
  wire  _T_1368;
  wire  _T_1369;
  wire  _T_1370;
  wire [14:0] _T_1371;
  wire [15:0] _T_1372;
  reg [15:0] _T_1374;
  reg [31:0] _RAND_103;
  wire  _T_1375;
  wire  _T_1376;
  wire  _T_1377;
  wire  _T_1378;
  wire  _T_1379;
  wire  _T_1380;
  wire  _T_1381;
  wire  _T_1382;
  wire [14:0] _T_1383;
  wire [15:0] _T_1384;
  reg [15:0] _T_1386;
  reg [31:0] _RAND_104;
  wire  _T_1387;
  wire  _T_1388;
  wire  _T_1389;
  wire  _T_1390;
  wire  _T_1391;
  wire  _T_1392;
  wire  _T_1393;
  wire  _T_1394;
  wire [14:0] _T_1395;
  wire [15:0] _T_1396;
  reg [15:0] _T_1398;
  reg [31:0] _RAND_105;
  wire  _T_1399;
  wire  _T_1400;
  wire  _T_1401;
  wire  _T_1402;
  wire  _T_1403;
  wire  _T_1404;
  wire  _T_1405;
  wire  _T_1406;
  wire [14:0] _T_1407;
  wire [15:0] _T_1408;
  reg [15:0] _T_1410;
  reg [31:0] _RAND_106;
  wire  _T_1411;
  wire  _T_1412;
  wire  _T_1413;
  wire  _T_1414;
  wire  _T_1415;
  wire  _T_1416;
  wire  _T_1417;
  wire  _T_1418;
  wire [14:0] _T_1419;
  wire [15:0] _T_1420;
  reg [15:0] _T_1422;
  reg [31:0] _RAND_107;
  wire  _T_1423;
  wire  _T_1424;
  wire  _T_1425;
  wire  _T_1426;
  wire  _T_1427;
  wire  _T_1428;
  wire  _T_1429;
  wire  _T_1430;
  wire [14:0] _T_1431;
  wire [15:0] _T_1432;
  reg [15:0] _T_1434;
  reg [31:0] _RAND_108;
  wire  _T_1435;
  wire  _T_1436;
  wire  _T_1437;
  wire  _T_1438;
  wire  _T_1439;
  wire  _T_1440;
  wire  _T_1441;
  wire  _T_1442;
  wire [14:0] _T_1443;
  wire [15:0] _T_1444;
  reg [15:0] _T_1446;
  reg [31:0] _RAND_109;
  wire  _T_1447;
  wire  _T_1448;
  wire  _T_1449;
  wire  _T_1450;
  wire  _T_1451;
  wire  _T_1452;
  wire  _T_1453;
  wire  _T_1454;
  wire [14:0] _T_1455;
  wire [15:0] _T_1456;
  reg [15:0] _T_1458;
  reg [31:0] _RAND_110;
  wire  _T_1459;
  wire  _T_1460;
  wire  _T_1461;
  wire  _T_1462;
  wire  _T_1463;
  wire  _T_1464;
  wire  _T_1465;
  wire  _T_1466;
  wire [14:0] _T_1467;
  wire [15:0] _T_1468;
  reg [15:0] _T_1470;
  reg [31:0] _RAND_111;
  wire  _T_1471;
  wire  _T_1472;
  wire  _T_1473;
  wire  _T_1474;
  wire  _T_1475;
  wire  _T_1476;
  wire  _T_1477;
  wire  _T_1478;
  wire [14:0] _T_1479;
  wire [15:0] _T_1480;
  reg [15:0] _T_1482;
  reg [31:0] _RAND_112;
  wire  _T_1483;
  wire  _T_1484;
  wire  _T_1485;
  wire  _T_1486;
  wire  _T_1487;
  wire  _T_1488;
  wire  _T_1489;
  wire  _T_1490;
  wire [14:0] _T_1491;
  wire [15:0] _T_1492;
  reg [15:0] _T_1494;
  reg [31:0] _RAND_113;
  wire  _T_1495;
  wire  _T_1496;
  wire  _T_1497;
  wire  _T_1498;
  wire  _T_1499;
  wire  _T_1500;
  wire  _T_1501;
  wire  _T_1502;
  wire [14:0] _T_1503;
  wire [15:0] _T_1504;
  reg [15:0] _T_1506;
  reg [31:0] _RAND_114;
  wire  _T_1507;
  wire  _T_1508;
  wire  _T_1509;
  wire  _T_1510;
  wire  _T_1511;
  wire  _T_1512;
  wire  _T_1513;
  wire  _T_1514;
  wire [14:0] _T_1515;
  wire [15:0] _T_1516;
  reg [15:0] _T_1518;
  reg [31:0] _RAND_115;
  wire  _T_1519;
  wire  _T_1520;
  wire  _T_1521;
  wire  _T_1522;
  wire  _T_1523;
  wire  _T_1524;
  wire  _T_1525;
  wire  _T_1526;
  wire [14:0] _T_1527;
  wire [15:0] _T_1528;
  reg [15:0] _T_1530;
  reg [31:0] _RAND_116;
  wire  _T_1531;
  wire  _T_1532;
  wire  _T_1533;
  wire  _T_1534;
  wire  _T_1535;
  wire  _T_1536;
  wire  _T_1537;
  wire  _T_1538;
  wire [14:0] _T_1539;
  wire [15:0] _T_1540;
  reg [15:0] _T_1542;
  reg [31:0] _RAND_117;
  wire  _T_1543;
  wire  _T_1544;
  wire  _T_1545;
  wire  _T_1546;
  wire  _T_1547;
  wire  _T_1548;
  wire  _T_1549;
  wire  _T_1550;
  wire [14:0] _T_1551;
  wire [15:0] _T_1552;
  reg [15:0] _T_1554;
  reg [31:0] _RAND_118;
  wire  _T_1555;
  wire  _T_1556;
  wire  _T_1557;
  wire  _T_1558;
  wire  _T_1559;
  wire  _T_1560;
  wire  _T_1561;
  wire  _T_1562;
  wire [14:0] _T_1563;
  wire [15:0] _T_1564;
  reg [15:0] _T_1566;
  reg [31:0] _RAND_119;
  wire  _T_1567;
  wire  _T_1568;
  wire  _T_1569;
  wire  _T_1570;
  wire  _T_1571;
  wire  _T_1572;
  wire  _T_1573;
  wire  _T_1574;
  wire [14:0] _T_1575;
  wire [15:0] _T_1576;
  reg [15:0] _T_1578;
  reg [31:0] _RAND_120;
  wire  _T_1579;
  wire  _T_1580;
  wire  _T_1581;
  wire  _T_1582;
  wire  _T_1583;
  wire  _T_1584;
  wire  _T_1585;
  wire  _T_1586;
  wire [14:0] _T_1587;
  wire [15:0] _T_1588;
  reg [15:0] _T_1590;
  reg [31:0] _RAND_121;
  wire  _T_1591;
  wire  _T_1592;
  wire  _T_1593;
  wire  _T_1594;
  wire  _T_1595;
  wire  _T_1596;
  wire  _T_1597;
  wire  _T_1598;
  wire [14:0] _T_1599;
  wire [15:0] _T_1600;
  reg [15:0] _T_1602;
  reg [31:0] _RAND_122;
  wire  _T_1603;
  wire  _T_1604;
  wire  _T_1605;
  wire  _T_1606;
  wire  _T_1607;
  wire  _T_1608;
  wire  _T_1609;
  wire  _T_1610;
  wire [14:0] _T_1611;
  wire [15:0] _T_1612;
  reg [15:0] _T_1614;
  reg [31:0] _RAND_123;
  wire  _T_1615;
  wire  _T_1616;
  wire  _T_1617;
  wire  _T_1618;
  wire  _T_1619;
  wire  _T_1620;
  wire  _T_1621;
  wire  _T_1622;
  wire [14:0] _T_1623;
  wire [15:0] _T_1624;
  reg [15:0] _T_1626;
  reg [31:0] _RAND_124;
  wire  _T_1627;
  wire  _T_1628;
  wire  _T_1629;
  wire  _T_1630;
  wire  _T_1631;
  wire  _T_1632;
  wire  _T_1633;
  wire  _T_1634;
  wire [14:0] _T_1635;
  wire [15:0] _T_1636;
  reg [15:0] _T_1638;
  reg [31:0] _RAND_125;
  wire  _T_1639;
  wire  _T_1640;
  wire  _T_1641;
  wire  _T_1642;
  wire  _T_1643;
  wire  _T_1644;
  wire  _T_1645;
  wire  _T_1646;
  wire [14:0] _T_1647;
  wire [15:0] _T_1648;
  reg [15:0] _T_1650;
  reg [31:0] _RAND_126;
  wire  _T_1651;
  wire  _T_1652;
  wire  _T_1653;
  wire  _T_1654;
  wire  _T_1655;
  wire  _T_1656;
  wire  _T_1657;
  wire  _T_1658;
  wire [14:0] _T_1659;
  wire [15:0] _T_1660;
  reg [15:0] _T_1662;
  reg [31:0] _RAND_127;
  wire  _T_1663;
  wire  _T_1664;
  wire  _T_1665;
  wire  _T_1666;
  wire  _T_1667;
  wire  _T_1668;
  wire  _T_1669;
  wire  _T_1670;
  wire [14:0] _T_1671;
  wire [15:0] _T_1672;
  reg [15:0] _T_1674;
  reg [31:0] _RAND_128;
  wire  _T_1675;
  wire  _T_1676;
  wire  _T_1677;
  wire  _T_1678;
  wire  _T_1679;
  wire  _T_1680;
  wire  _T_1681;
  wire  _T_1682;
  wire [14:0] _T_1683;
  wire [15:0] _T_1684;
  reg [15:0] _T_1686;
  reg [31:0] _RAND_129;
  wire  _T_1687;
  wire  _T_1688;
  wire  _T_1689;
  wire  _T_1690;
  wire  _T_1691;
  wire  _T_1692;
  wire  _T_1693;
  wire  _T_1694;
  wire [14:0] _T_1695;
  wire [15:0] _T_1696;
  reg [15:0] _T_1698;
  reg [31:0] _RAND_130;
  wire  _T_1699;
  wire  _T_1700;
  wire  _T_1701;
  wire  _T_1702;
  wire  _T_1703;
  wire  _T_1704;
  wire  _T_1705;
  wire  _T_1706;
  wire [14:0] _T_1707;
  wire [15:0] _T_1708;
  reg [15:0] _T_1712;
  reg [31:0] _RAND_131;
  wire  _T_1713;
  wire  _T_1714;
  wire  _T_1715;
  wire  _T_1716;
  wire  _T_1717;
  wire  _T_1718;
  wire  _T_1719;
  wire  _T_1720;
  wire [14:0] _T_1721;
  wire [15:0] _T_1722;
  reg [15:0] _T_1724;
  reg [31:0] _RAND_132;
  wire  _T_1725;
  wire  _T_1726;
  wire  _T_1727;
  wire  _T_1728;
  wire  _T_1729;
  wire  _T_1730;
  wire  _T_1731;
  wire  _T_1732;
  wire [14:0] _T_1733;
  wire [15:0] _T_1734;
  reg [15:0] _T_1736;
  reg [31:0] _RAND_133;
  wire  _T_1737;
  wire  _T_1738;
  wire  _T_1739;
  wire  _T_1740;
  wire  _T_1741;
  wire  _T_1742;
  wire  _T_1743;
  wire  _T_1744;
  wire [14:0] _T_1745;
  wire [15:0] _T_1746;
  reg [15:0] _T_1748;
  reg [31:0] _RAND_134;
  wire  _T_1749;
  wire  _T_1750;
  wire  _T_1751;
  wire  _T_1752;
  wire  _T_1753;
  wire  _T_1754;
  wire  _T_1755;
  wire  _T_1756;
  wire [14:0] _T_1757;
  wire [15:0] _T_1758;
  reg [15:0] _T_1760;
  reg [31:0] _RAND_135;
  wire  _T_1761;
  wire  _T_1762;
  wire  _T_1763;
  wire  _T_1764;
  wire  _T_1765;
  wire  _T_1766;
  wire  _T_1767;
  wire  _T_1768;
  wire [14:0] _T_1769;
  wire [15:0] _T_1770;
  reg [15:0] _T_1772;
  reg [31:0] _RAND_136;
  wire  _T_1773;
  wire  _T_1774;
  wire  _T_1775;
  wire  _T_1776;
  wire  _T_1777;
  wire  _T_1778;
  wire  _T_1779;
  wire  _T_1780;
  wire [14:0] _T_1781;
  wire [15:0] _T_1782;
  reg [15:0] _T_1784;
  reg [31:0] _RAND_137;
  wire  _T_1785;
  wire  _T_1786;
  wire  _T_1787;
  wire  _T_1788;
  wire  _T_1789;
  wire  _T_1790;
  wire  _T_1791;
  wire  _T_1792;
  wire [14:0] _T_1793;
  wire [15:0] _T_1794;
  reg [15:0] _T_1796;
  reg [31:0] _RAND_138;
  wire  _T_1797;
  wire  _T_1798;
  wire  _T_1799;
  wire  _T_1800;
  wire  _T_1801;
  wire  _T_1802;
  wire  _T_1803;
  wire  _T_1804;
  wire [14:0] _T_1805;
  wire [15:0] _T_1806;
  reg [15:0] _T_1808;
  reg [31:0] _RAND_139;
  wire  _T_1809;
  wire  _T_1810;
  wire  _T_1811;
  wire  _T_1812;
  wire  _T_1813;
  wire  _T_1814;
  wire  _T_1815;
  wire  _T_1816;
  wire [14:0] _T_1817;
  wire [15:0] _T_1818;
  reg [15:0] _T_1820;
  reg [31:0] _RAND_140;
  wire  _T_1821;
  wire  _T_1822;
  wire  _T_1823;
  wire  _T_1824;
  wire  _T_1825;
  wire  _T_1826;
  wire  _T_1827;
  wire  _T_1828;
  wire [14:0] _T_1829;
  wire [15:0] _T_1830;
  reg [15:0] _T_1832;
  reg [31:0] _RAND_141;
  wire  _T_1833;
  wire  _T_1834;
  wire  _T_1835;
  wire  _T_1836;
  wire  _T_1837;
  wire  _T_1838;
  wire  _T_1839;
  wire  _T_1840;
  wire [14:0] _T_1841;
  wire [15:0] _T_1842;
  reg [15:0] _T_1844;
  reg [31:0] _RAND_142;
  wire  _T_1845;
  wire  _T_1846;
  wire  _T_1847;
  wire  _T_1848;
  wire  _T_1849;
  wire  _T_1850;
  wire  _T_1851;
  wire  _T_1852;
  wire [14:0] _T_1853;
  wire [15:0] _T_1854;
  reg [15:0] _T_1856;
  reg [31:0] _RAND_143;
  wire  _T_1857;
  wire  _T_1858;
  wire  _T_1859;
  wire  _T_1860;
  wire  _T_1861;
  wire  _T_1862;
  wire  _T_1863;
  wire  _T_1864;
  wire [14:0] _T_1865;
  wire [15:0] _T_1866;
  reg [15:0] _T_1868;
  reg [31:0] _RAND_144;
  wire  _T_1869;
  wire  _T_1870;
  wire  _T_1871;
  wire  _T_1872;
  wire  _T_1873;
  wire  _T_1874;
  wire  _T_1875;
  wire  _T_1876;
  wire [14:0] _T_1877;
  wire [15:0] _T_1878;
  reg [15:0] _T_1880;
  reg [31:0] _RAND_145;
  wire  _T_1881;
  wire  _T_1882;
  wire  _T_1883;
  wire  _T_1884;
  wire  _T_1885;
  wire  _T_1886;
  wire  _T_1887;
  wire  _T_1888;
  wire [14:0] _T_1889;
  wire [15:0] _T_1890;
  reg [15:0] _T_1892;
  reg [31:0] _RAND_146;
  wire  _T_1893;
  wire  _T_1894;
  wire  _T_1895;
  wire  _T_1896;
  wire  _T_1897;
  wire  _T_1898;
  wire  _T_1899;
  wire  _T_1900;
  wire [14:0] _T_1901;
  wire [15:0] _T_1902;
  reg [15:0] _T_1904;
  reg [31:0] _RAND_147;
  wire  _T_1905;
  wire  _T_1906;
  wire  _T_1907;
  wire  _T_1908;
  wire  _T_1909;
  wire  _T_1910;
  wire  _T_1911;
  wire  _T_1912;
  wire [14:0] _T_1913;
  wire [15:0] _T_1914;
  reg [15:0] _T_1916;
  reg [31:0] _RAND_148;
  wire  _T_1917;
  wire  _T_1918;
  wire  _T_1919;
  wire  _T_1920;
  wire  _T_1921;
  wire  _T_1922;
  wire  _T_1923;
  wire  _T_1924;
  wire [14:0] _T_1925;
  wire [15:0] _T_1926;
  reg [15:0] _T_1928;
  reg [31:0] _RAND_149;
  wire  _T_1929;
  wire  _T_1930;
  wire  _T_1931;
  wire  _T_1932;
  wire  _T_1933;
  wire  _T_1934;
  wire  _T_1935;
  wire  _T_1936;
  wire [14:0] _T_1937;
  wire [15:0] _T_1938;
  reg [15:0] _T_1940;
  reg [31:0] _RAND_150;
  wire  _T_1941;
  wire  _T_1942;
  wire  _T_1943;
  wire  _T_1944;
  wire  _T_1945;
  wire  _T_1946;
  wire  _T_1947;
  wire  _T_1948;
  wire [14:0] _T_1949;
  wire [15:0] _T_1950;
  reg [15:0] _T_1952;
  reg [31:0] _RAND_151;
  wire  _T_1953;
  wire  _T_1954;
  wire  _T_1955;
  wire  _T_1956;
  wire  _T_1957;
  wire  _T_1958;
  wire  _T_1959;
  wire  _T_1960;
  wire [14:0] _T_1961;
  wire [15:0] _T_1962;
  reg [15:0] _T_1964;
  reg [31:0] _RAND_152;
  wire  _T_1965;
  wire  _T_1966;
  wire  _T_1967;
  wire  _T_1968;
  wire  _T_1969;
  wire  _T_1970;
  wire  _T_1971;
  wire  _T_1972;
  wire [14:0] _T_1973;
  wire [15:0] _T_1974;
  reg [15:0] _T_1976;
  reg [31:0] _RAND_153;
  wire  _T_1977;
  wire  _T_1978;
  wire  _T_1979;
  wire  _T_1980;
  wire  _T_1981;
  wire  _T_1982;
  wire  _T_1983;
  wire  _T_1984;
  wire [14:0] _T_1985;
  wire [15:0] _T_1986;
  reg [15:0] _T_1988;
  reg [31:0] _RAND_154;
  wire  _T_1989;
  wire  _T_1990;
  wire  _T_1991;
  wire  _T_1992;
  wire  _T_1993;
  wire  _T_1994;
  wire  _T_1995;
  wire  _T_1996;
  wire [14:0] _T_1997;
  wire [15:0] _T_1998;
  reg [15:0] _T_2000;
  reg [31:0] _RAND_155;
  wire  _T_2001;
  wire  _T_2002;
  wire  _T_2003;
  wire  _T_2004;
  wire  _T_2005;
  wire  _T_2006;
  wire  _T_2007;
  wire  _T_2008;
  wire [14:0] _T_2009;
  wire [15:0] _T_2010;
  reg [15:0] _T_2012;
  reg [31:0] _RAND_156;
  wire  _T_2013;
  wire  _T_2014;
  wire  _T_2015;
  wire  _T_2016;
  wire  _T_2017;
  wire  _T_2018;
  wire  _T_2019;
  wire  _T_2020;
  wire [14:0] _T_2021;
  wire [15:0] _T_2022;
  reg [15:0] _T_2024;
  reg [31:0] _RAND_157;
  wire  _T_2025;
  wire  _T_2026;
  wire  _T_2027;
  wire  _T_2028;
  wire  _T_2029;
  wire  _T_2030;
  wire  _T_2031;
  wire  _T_2032;
  wire [14:0] _T_2033;
  wire [15:0] _T_2034;
  reg [15:0] _T_2036;
  reg [31:0] _RAND_158;
  wire  _T_2037;
  wire  _T_2038;
  wire  _T_2039;
  wire  _T_2040;
  wire  _T_2041;
  wire  _T_2042;
  wire  _T_2043;
  wire  _T_2044;
  wire [14:0] _T_2045;
  wire [15:0] _T_2046;
  reg [15:0] _T_2048;
  reg [31:0] _RAND_159;
  wire  _T_2049;
  wire  _T_2050;
  wire  _T_2051;
  wire  _T_2052;
  wire  _T_2053;
  wire  _T_2054;
  wire  _T_2055;
  wire  _T_2056;
  wire [14:0] _T_2057;
  wire [15:0] _T_2058;
  reg [15:0] _T_2060;
  reg [31:0] _RAND_160;
  wire  _T_2061;
  wire  _T_2062;
  wire  _T_2063;
  wire  _T_2064;
  wire  _T_2065;
  wire  _T_2066;
  wire  _T_2067;
  wire  _T_2068;
  wire [14:0] _T_2069;
  wire [15:0] _T_2070;
  reg [15:0] _T_2072;
  reg [31:0] _RAND_161;
  wire  _T_2073;
  wire  _T_2074;
  wire  _T_2075;
  wire  _T_2076;
  wire  _T_2077;
  wire  _T_2078;
  wire  _T_2079;
  wire  _T_2080;
  wire [14:0] _T_2081;
  wire [15:0] _T_2082;
  reg [15:0] _T_2084;
  reg [31:0] _RAND_162;
  wire  _T_2085;
  wire  _T_2086;
  wire  _T_2087;
  wire  _T_2088;
  wire  _T_2089;
  wire  _T_2090;
  wire  _T_2091;
  wire  _T_2092;
  wire [14:0] _T_2093;
  wire [15:0] _T_2094;
  reg [15:0] _T_2096;
  reg [31:0] _RAND_163;
  wire  _T_2097;
  wire  _T_2098;
  wire  _T_2099;
  wire  _T_2100;
  wire  _T_2101;
  wire  _T_2102;
  wire  _T_2103;
  wire  _T_2104;
  wire [14:0] _T_2105;
  wire [15:0] _T_2106;
  reg [15:0] _T_2108;
  reg [31:0] _RAND_164;
  wire  _T_2109;
  wire  _T_2110;
  wire  _T_2111;
  wire  _T_2112;
  wire  _T_2113;
  wire  _T_2114;
  wire  _T_2115;
  wire  _T_2116;
  wire [14:0] _T_2117;
  wire [15:0] _T_2118;
  reg [15:0] _T_2120;
  reg [31:0] _RAND_165;
  wire  _T_2121;
  wire  _T_2122;
  wire  _T_2123;
  wire  _T_2124;
  wire  _T_2125;
  wire  _T_2126;
  wire  _T_2127;
  wire  _T_2128;
  wire [14:0] _T_2129;
  wire [15:0] _T_2130;
  reg [15:0] _T_2132;
  reg [31:0] _RAND_166;
  wire  _T_2133;
  wire  _T_2134;
  wire  _T_2135;
  wire  _T_2136;
  wire  _T_2137;
  wire  _T_2138;
  wire  _T_2139;
  wire  _T_2140;
  wire [14:0] _T_2141;
  wire [15:0] _T_2142;
  reg [15:0] _T_2144;
  reg [31:0] _RAND_167;
  wire  _T_2145;
  wire  _T_2146;
  wire  _T_2147;
  wire  _T_2148;
  wire  _T_2149;
  wire  _T_2150;
  wire  _T_2151;
  wire  _T_2152;
  wire [14:0] _T_2153;
  wire [15:0] _T_2154;
  reg [15:0] _T_2156;
  reg [31:0] _RAND_168;
  wire  _T_2157;
  wire  _T_2158;
  wire  _T_2159;
  wire  _T_2160;
  wire  _T_2161;
  wire  _T_2162;
  wire  _T_2163;
  wire  _T_2164;
  wire [14:0] _T_2165;
  wire [15:0] _T_2166;
  reg [15:0] _T_2168;
  reg [31:0] _RAND_169;
  wire  _T_2169;
  wire  _T_2170;
  wire  _T_2171;
  wire  _T_2172;
  wire  _T_2173;
  wire  _T_2174;
  wire  _T_2175;
  wire  _T_2176;
  wire [14:0] _T_2177;
  wire [15:0] _T_2178;
  reg [15:0] _T_2180;
  reg [31:0] _RAND_170;
  wire  _T_2181;
  wire  _T_2182;
  wire  _T_2183;
  wire  _T_2184;
  wire  _T_2185;
  wire  _T_2186;
  wire  _T_2187;
  wire  _T_2188;
  wire [14:0] _T_2189;
  wire [15:0] _T_2190;
  reg [15:0] _T_2192;
  reg [31:0] _RAND_171;
  wire  _T_2193;
  wire  _T_2194;
  wire  _T_2195;
  wire  _T_2196;
  wire  _T_2197;
  wire  _T_2198;
  wire  _T_2199;
  wire  _T_2200;
  wire [14:0] _T_2201;
  wire [15:0] _T_2202;
  reg [15:0] _T_2204;
  reg [31:0] _RAND_172;
  wire  _T_2205;
  wire  _T_2206;
  wire  _T_2207;
  wire  _T_2208;
  wire  _T_2209;
  wire  _T_2210;
  wire  _T_2211;
  wire  _T_2212;
  wire [14:0] _T_2213;
  wire [15:0] _T_2214;
  reg [15:0] _T_2216;
  reg [31:0] _RAND_173;
  wire  _T_2217;
  wire  _T_2218;
  wire  _T_2219;
  wire  _T_2220;
  wire  _T_2221;
  wire  _T_2222;
  wire  _T_2223;
  wire  _T_2224;
  wire [14:0] _T_2225;
  wire [15:0] _T_2226;
  reg [15:0] _T_2228;
  reg [31:0] _RAND_174;
  wire  _T_2229;
  wire  _T_2230;
  wire  _T_2231;
  wire  _T_2232;
  wire  _T_2233;
  wire  _T_2234;
  wire  _T_2235;
  wire  _T_2236;
  wire [14:0] _T_2237;
  wire [15:0] _T_2238;
  reg [15:0] _T_2240;
  reg [31:0] _RAND_175;
  wire  _T_2241;
  wire  _T_2242;
  wire  _T_2243;
  wire  _T_2244;
  wire  _T_2245;
  wire  _T_2246;
  wire  _T_2247;
  wire  _T_2248;
  wire [14:0] _T_2249;
  wire [15:0] _T_2250;
  reg [15:0] _T_2252;
  reg [31:0] _RAND_176;
  wire  _T_2253;
  wire  _T_2254;
  wire  _T_2255;
  wire  _T_2256;
  wire  _T_2257;
  wire  _T_2258;
  wire  _T_2259;
  wire  _T_2260;
  wire [14:0] _T_2261;
  wire [15:0] _T_2262;
  reg [15:0] _T_2264;
  reg [31:0] _RAND_177;
  wire  _T_2265;
  wire  _T_2266;
  wire  _T_2267;
  wire  _T_2268;
  wire  _T_2269;
  wire  _T_2270;
  wire  _T_2271;
  wire  _T_2272;
  wire [14:0] _T_2273;
  wire [15:0] _T_2274;
  reg [15:0] _T_2276;
  reg [31:0] _RAND_178;
  wire  _T_2277;
  wire  _T_2278;
  wire  _T_2279;
  wire  _T_2280;
  wire  _T_2281;
  wire  _T_2282;
  wire  _T_2283;
  wire  _T_2284;
  wire [14:0] _T_2285;
  wire [15:0] _T_2286;
  reg [15:0] _T_2288;
  reg [31:0] _RAND_179;
  wire  _T_2289;
  wire  _T_2290;
  wire  _T_2291;
  wire  _T_2292;
  wire  _T_2293;
  wire  _T_2294;
  wire  _T_2295;
  wire  _T_2296;
  wire [14:0] _T_2297;
  wire [15:0] _T_2298;
  reg [15:0] _T_2300;
  reg [31:0] _RAND_180;
  wire  _T_2301;
  wire  _T_2302;
  wire  _T_2303;
  wire  _T_2304;
  wire  _T_2305;
  wire  _T_2306;
  wire  _T_2307;
  wire  _T_2308;
  wire [14:0] _T_2309;
  wire [15:0] _T_2310;
  reg [15:0] _T_2312;
  reg [31:0] _RAND_181;
  wire  _T_2313;
  wire  _T_2314;
  wire  _T_2315;
  wire  _T_2316;
  wire  _T_2317;
  wire  _T_2318;
  wire  _T_2319;
  wire  _T_2320;
  wire [14:0] _T_2321;
  wire [15:0] _T_2322;
  reg [15:0] _T_2324;
  reg [31:0] _RAND_182;
  wire  _T_2325;
  wire  _T_2326;
  wire  _T_2327;
  wire  _T_2328;
  wire  _T_2329;
  wire  _T_2330;
  wire  _T_2331;
  wire  _T_2332;
  wire [14:0] _T_2333;
  wire [15:0] _T_2334;
  reg [15:0] _T_2336;
  reg [31:0] _RAND_183;
  wire  _T_2337;
  wire  _T_2338;
  wire  _T_2339;
  wire  _T_2340;
  wire  _T_2341;
  wire  _T_2342;
  wire  _T_2343;
  wire  _T_2344;
  wire [14:0] _T_2345;
  wire [15:0] _T_2346;
  reg [15:0] _T_2348;
  reg [31:0] _RAND_184;
  wire  _T_2349;
  wire  _T_2350;
  wire  _T_2351;
  wire  _T_2352;
  wire  _T_2353;
  wire  _T_2354;
  wire  _T_2355;
  wire  _T_2356;
  wire [14:0] _T_2357;
  wire [15:0] _T_2358;
  reg [15:0] _T_2360;
  reg [31:0] _RAND_185;
  wire  _T_2361;
  wire  _T_2362;
  wire  _T_2363;
  wire  _T_2364;
  wire  _T_2365;
  wire  _T_2366;
  wire  _T_2367;
  wire  _T_2368;
  wire [14:0] _T_2369;
  wire [15:0] _T_2370;
  reg [15:0] _T_2372;
  reg [31:0] _RAND_186;
  wire  _T_2373;
  wire  _T_2374;
  wire  _T_2375;
  wire  _T_2376;
  wire  _T_2377;
  wire  _T_2378;
  wire  _T_2379;
  wire  _T_2380;
  wire [14:0] _T_2381;
  wire [15:0] _T_2382;
  reg [15:0] _T_2384;
  reg [31:0] _RAND_187;
  wire  _T_2385;
  wire  _T_2386;
  wire  _T_2387;
  wire  _T_2388;
  wire  _T_2389;
  wire  _T_2390;
  wire  _T_2391;
  wire  _T_2392;
  wire [14:0] _T_2393;
  wire [15:0] _T_2394;
  reg [15:0] _T_2396;
  reg [31:0] _RAND_188;
  wire  _T_2397;
  wire  _T_2398;
  wire  _T_2399;
  wire  _T_2400;
  wire  _T_2401;
  wire  _T_2402;
  wire  _T_2403;
  wire  _T_2404;
  wire [14:0] _T_2405;
  wire [15:0] _T_2406;
  reg [15:0] _T_2408;
  reg [31:0] _RAND_189;
  wire  _T_2409;
  wire  _T_2410;
  wire  _T_2411;
  wire  _T_2412;
  wire  _T_2413;
  wire  _T_2414;
  wire  _T_2415;
  wire  _T_2416;
  wire [14:0] _T_2417;
  wire [15:0] _T_2418;
  reg [15:0] _T_2420;
  reg [31:0] _RAND_190;
  wire  _T_2421;
  wire  _T_2422;
  wire  _T_2423;
  wire  _T_2424;
  wire  _T_2425;
  wire  _T_2426;
  wire  _T_2427;
  wire  _T_2428;
  wire [14:0] _T_2429;
  wire [15:0] _T_2430;
  reg [15:0] _T_2432;
  reg [31:0] _RAND_191;
  wire  _T_2433;
  wire  _T_2434;
  wire  _T_2435;
  wire  _T_2436;
  wire  _T_2437;
  wire  _T_2438;
  wire  _T_2439;
  wire  _T_2440;
  wire [14:0] _T_2441;
  wire [15:0] _T_2442;
  reg [15:0] _T_2444;
  reg [31:0] _RAND_192;
  wire  _T_2445;
  wire  _T_2446;
  wire  _T_2447;
  wire  _T_2448;
  wire  _T_2449;
  wire  _T_2450;
  wire  _T_2451;
  wire  _T_2452;
  wire [14:0] _T_2453;
  wire [15:0] _T_2454;
  reg [15:0] _T_2456;
  reg [31:0] _RAND_193;
  wire  _T_2457;
  wire  _T_2458;
  wire  _T_2459;
  wire  _T_2460;
  wire  _T_2461;
  wire  _T_2462;
  wire  _T_2463;
  wire  _T_2464;
  wire [14:0] _T_2465;
  wire [15:0] _T_2466;
  reg [15:0] _T_2468;
  reg [31:0] _RAND_194;
  wire  _T_2469;
  wire  _T_2470;
  wire  _T_2471;
  wire  _T_2472;
  wire  _T_2473;
  wire  _T_2474;
  wire  _T_2475;
  wire  _T_2476;
  wire [14:0] _T_2477;
  wire [15:0] _T_2478;
  reg [15:0] _T_2480;
  reg [31:0] _RAND_195;
  wire  _T_2481;
  wire  _T_2482;
  wire  _T_2483;
  wire  _T_2484;
  wire  _T_2485;
  wire  _T_2486;
  wire  _T_2487;
  wire  _T_2488;
  wire [14:0] _T_2489;
  wire [15:0] _T_2490;
  reg [15:0] _T_2492;
  reg [31:0] _RAND_196;
  wire  _T_2493;
  wire  _T_2494;
  wire  _T_2495;
  wire  _T_2496;
  wire  _T_2497;
  wire  _T_2498;
  wire  _T_2499;
  wire  _T_2500;
  wire [14:0] _T_2501;
  wire [15:0] _T_2502;
  reg [15:0] _T_2504;
  reg [31:0] _RAND_197;
  wire  _T_2505;
  wire  _T_2506;
  wire  _T_2507;
  wire  _T_2508;
  wire  _T_2509;
  wire  _T_2510;
  wire  _T_2511;
  wire  _T_2512;
  wire [14:0] _T_2513;
  wire [15:0] _T_2514;
  reg [15:0] _T_2516;
  reg [31:0] _RAND_198;
  wire  _T_2517;
  wire  _T_2518;
  wire  _T_2519;
  wire  _T_2520;
  wire  _T_2521;
  wire  _T_2522;
  wire  _T_2523;
  wire  _T_2524;
  wire [14:0] _T_2525;
  wire [15:0] _T_2526;
  reg [15:0] _T_2528;
  reg [31:0] _RAND_199;
  wire  _T_2529;
  wire  _T_2530;
  wire  _T_2531;
  wire  _T_2532;
  wire  _T_2533;
  wire  _T_2534;
  wire  _T_2535;
  wire  _T_2536;
  wire [14:0] _T_2537;
  wire [15:0] _T_2538;
  reg [15:0] _T_2540;
  reg [31:0] _RAND_200;
  wire  _T_2541;
  wire  _T_2542;
  wire  _T_2543;
  wire  _T_2544;
  wire  _T_2545;
  wire  _T_2546;
  wire  _T_2547;
  wire  _T_2548;
  wire [14:0] _T_2549;
  wire [15:0] _T_2550;
  reg [15:0] _T_2552;
  reg [31:0] _RAND_201;
  wire  _T_2553;
  wire  _T_2554;
  wire  _T_2555;
  wire  _T_2556;
  wire  _T_2557;
  wire  _T_2558;
  wire  _T_2559;
  wire  _T_2560;
  wire [14:0] _T_2561;
  wire [15:0] _T_2562;
  reg [15:0] _T_2564;
  reg [31:0] _RAND_202;
  wire  _T_2565;
  wire  _T_2566;
  wire  _T_2567;
  wire  _T_2568;
  wire  _T_2569;
  wire  _T_2570;
  wire  _T_2571;
  wire  _T_2572;
  wire [14:0] _T_2573;
  wire [15:0] _T_2574;
  reg [15:0] _T_2576;
  reg [31:0] _RAND_203;
  wire  _T_2577;
  wire  _T_2578;
  wire  _T_2579;
  wire  _T_2580;
  wire  _T_2581;
  wire  _T_2582;
  wire  _T_2583;
  wire  _T_2584;
  wire [14:0] _T_2585;
  wire [15:0] _T_2586;
  reg [15:0] _T_2588;
  reg [31:0] _RAND_204;
  wire  _T_2589;
  wire  _T_2590;
  wire  _T_2591;
  wire  _T_2592;
  wire  _T_2593;
  wire  _T_2594;
  wire  _T_2595;
  wire  _T_2596;
  wire [14:0] _T_2597;
  wire [15:0] _T_2598;
  reg [15:0] _T_2600;
  reg [31:0] _RAND_205;
  wire  _T_2601;
  wire  _T_2602;
  wire  _T_2603;
  wire  _T_2604;
  wire  _T_2605;
  wire  _T_2606;
  wire  _T_2607;
  wire  _T_2608;
  wire [14:0] _T_2609;
  wire [15:0] _T_2610;
  reg [15:0] _T_2612;
  reg [31:0] _RAND_206;
  wire  _T_2613;
  wire  _T_2614;
  wire  _T_2615;
  wire  _T_2616;
  wire  _T_2617;
  wire  _T_2618;
  wire  _T_2619;
  wire  _T_2620;
  wire [14:0] _T_2621;
  wire [15:0] _T_2622;
  reg [15:0] _T_2624;
  reg [31:0] _RAND_207;
  wire  _T_2625;
  wire  _T_2626;
  wire  _T_2627;
  wire  _T_2628;
  wire  _T_2629;
  wire  _T_2630;
  wire  _T_2631;
  wire  _T_2632;
  wire [14:0] _T_2633;
  wire [15:0] _T_2634;
  reg [15:0] _T_2636;
  reg [31:0] _RAND_208;
  wire  _T_2637;
  wire  _T_2638;
  wire  _T_2639;
  wire  _T_2640;
  wire  _T_2641;
  wire  _T_2642;
  wire  _T_2643;
  wire  _T_2644;
  wire [14:0] _T_2645;
  wire [15:0] _T_2646;
  reg [15:0] _T_2648;
  reg [31:0] _RAND_209;
  wire  _T_2649;
  wire  _T_2650;
  wire  _T_2651;
  wire  _T_2652;
  wire  _T_2653;
  wire  _T_2654;
  wire  _T_2655;
  wire  _T_2656;
  wire [14:0] _T_2657;
  wire [15:0] _T_2658;
  reg [15:0] _T_2660;
  reg [31:0] _RAND_210;
  wire  _T_2661;
  wire  _T_2662;
  wire  _T_2663;
  wire  _T_2664;
  wire  _T_2665;
  wire  _T_2666;
  wire  _T_2667;
  wire  _T_2668;
  wire [14:0] _T_2669;
  wire [15:0] _T_2670;
  reg [15:0] _T_2672;
  reg [31:0] _RAND_211;
  wire  _T_2673;
  wire  _T_2674;
  wire  _T_2675;
  wire  _T_2676;
  wire  _T_2677;
  wire  _T_2678;
  wire  _T_2679;
  wire  _T_2680;
  wire [14:0] _T_2681;
  wire [15:0] _T_2682;
  reg [15:0] _T_2684;
  reg [31:0] _RAND_212;
  wire  _T_2685;
  wire  _T_2686;
  wire  _T_2687;
  wire  _T_2688;
  wire  _T_2689;
  wire  _T_2690;
  wire  _T_2691;
  wire  _T_2692;
  wire [14:0] _T_2693;
  wire [15:0] _T_2694;
  reg [15:0] _T_2696;
  reg [31:0] _RAND_213;
  wire  _T_2697;
  wire  _T_2698;
  wire  _T_2699;
  wire  _T_2700;
  wire  _T_2701;
  wire  _T_2702;
  wire  _T_2703;
  wire  _T_2704;
  wire [14:0] _T_2705;
  wire [15:0] _T_2706;
  reg [15:0] _T_2708;
  reg [31:0] _RAND_214;
  wire  _T_2709;
  wire  _T_2710;
  wire  _T_2711;
  wire  _T_2712;
  wire  _T_2713;
  wire  _T_2714;
  wire  _T_2715;
  wire  _T_2716;
  wire [14:0] _T_2717;
  wire [15:0] _T_2718;
  reg [15:0] _T_2720;
  reg [31:0] _RAND_215;
  wire  _T_2721;
  wire  _T_2722;
  wire  _T_2723;
  wire  _T_2724;
  wire  _T_2725;
  wire  _T_2726;
  wire  _T_2727;
  wire  _T_2728;
  wire [14:0] _T_2729;
  wire [15:0] _T_2730;
  reg [15:0] _T_2732;
  reg [31:0] _RAND_216;
  wire  _T_2733;
  wire  _T_2734;
  wire  _T_2735;
  wire  _T_2736;
  wire  _T_2737;
  wire  _T_2738;
  wire  _T_2739;
  wire  _T_2740;
  wire [14:0] _T_2741;
  wire [15:0] _T_2742;
  reg [15:0] _T_2744;
  reg [31:0] _RAND_217;
  wire  _T_2745;
  wire  _T_2746;
  wire  _T_2747;
  wire  _T_2748;
  wire  _T_2749;
  wire  _T_2750;
  wire  _T_2751;
  wire  _T_2752;
  wire [14:0] _T_2753;
  wire [15:0] _T_2754;
  reg [15:0] _T_2756;
  reg [31:0] _RAND_218;
  wire  _T_2757;
  wire  _T_2758;
  wire  _T_2759;
  wire  _T_2760;
  wire  _T_2761;
  wire  _T_2762;
  wire  _T_2763;
  wire  _T_2764;
  wire [14:0] _T_2765;
  wire [15:0] _T_2766;
  reg [15:0] _T_2768;
  reg [31:0] _RAND_219;
  wire  _T_2769;
  wire  _T_2770;
  wire  _T_2771;
  wire  _T_2772;
  wire  _T_2773;
  wire  _T_2774;
  wire  _T_2775;
  wire  _T_2776;
  wire [14:0] _T_2777;
  wire [15:0] _T_2778;
  reg [15:0] _T_2780;
  reg [31:0] _RAND_220;
  wire  _T_2781;
  wire  _T_2782;
  wire  _T_2783;
  wire  _T_2784;
  wire  _T_2785;
  wire  _T_2786;
  wire  _T_2787;
  wire  _T_2788;
  wire [14:0] _T_2789;
  wire [15:0] _T_2790;
  reg [15:0] _T_2792;
  reg [31:0] _RAND_221;
  wire  _T_2793;
  wire  _T_2794;
  wire  _T_2795;
  wire  _T_2796;
  wire  _T_2797;
  wire  _T_2798;
  wire  _T_2799;
  wire  _T_2800;
  wire [14:0] _T_2801;
  wire [15:0] _T_2802;
  reg [15:0] _T_2804;
  reg [31:0] _RAND_222;
  wire  _T_2805;
  wire  _T_2806;
  wire  _T_2807;
  wire  _T_2808;
  wire  _T_2809;
  wire  _T_2810;
  wire  _T_2811;
  wire  _T_2812;
  wire [14:0] _T_2813;
  wire [15:0] _T_2814;
  reg [15:0] _T_2816;
  reg [31:0] _RAND_223;
  wire  _T_2817;
  wire  _T_2818;
  wire  _T_2819;
  wire  _T_2820;
  wire  _T_2821;
  wire  _T_2822;
  wire  _T_2823;
  wire  _T_2824;
  wire [14:0] _T_2825;
  wire [15:0] _T_2826;
  reg [15:0] _T_2828;
  reg [31:0] _RAND_224;
  wire  _T_2829;
  wire  _T_2830;
  wire  _T_2831;
  wire  _T_2832;
  wire  _T_2833;
  wire  _T_2834;
  wire  _T_2835;
  wire  _T_2836;
  wire [14:0] _T_2837;
  wire [15:0] _T_2838;
  reg [15:0] _T_2840;
  reg [31:0] _RAND_225;
  wire  _T_2841;
  wire  _T_2842;
  wire  _T_2843;
  wire  _T_2844;
  wire  _T_2845;
  wire  _T_2846;
  wire  _T_2847;
  wire  _T_2848;
  wire [14:0] _T_2849;
  wire [15:0] _T_2850;
  reg [15:0] _T_2852;
  reg [31:0] _RAND_226;
  wire  _T_2853;
  wire  _T_2854;
  wire  _T_2855;
  wire  _T_2856;
  wire  _T_2857;
  wire  _T_2858;
  wire  _T_2859;
  wire  _T_2860;
  wire [14:0] _T_2861;
  wire [15:0] _T_2862;
  reg [15:0] _T_2864;
  reg [31:0] _RAND_227;
  wire  _T_2865;
  wire  _T_2866;
  wire  _T_2867;
  wire  _T_2868;
  wire  _T_2869;
  wire  _T_2870;
  wire  _T_2871;
  wire  _T_2872;
  wire [14:0] _T_2873;
  wire [15:0] _T_2874;
  reg [15:0] _T_2876;
  reg [31:0] _RAND_228;
  wire  _T_2877;
  wire  _T_2878;
  wire  _T_2879;
  wire  _T_2880;
  wire  _T_2881;
  wire  _T_2882;
  wire  _T_2883;
  wire  _T_2884;
  wire [14:0] _T_2885;
  wire [15:0] _T_2886;
  reg [15:0] _T_2888;
  reg [31:0] _RAND_229;
  wire  _T_2889;
  wire  _T_2890;
  wire  _T_2891;
  wire  _T_2892;
  wire  _T_2893;
  wire  _T_2894;
  wire  _T_2895;
  wire  _T_2896;
  wire [14:0] _T_2897;
  wire [15:0] _T_2898;
  reg [15:0] _T_2900;
  reg [31:0] _RAND_230;
  wire  _T_2901;
  wire  _T_2902;
  wire  _T_2903;
  wire  _T_2904;
  wire  _T_2905;
  wire  _T_2906;
  wire  _T_2907;
  wire  _T_2908;
  wire [14:0] _T_2909;
  wire [15:0] _T_2910;
  reg [15:0] _T_2912;
  reg [31:0] _RAND_231;
  wire  _T_2913;
  wire  _T_2914;
  wire  _T_2915;
  wire  _T_2916;
  wire  _T_2917;
  wire  _T_2918;
  wire  _T_2919;
  wire  _T_2920;
  wire [14:0] _T_2921;
  wire [15:0] _T_2922;
  reg [15:0] _T_2924;
  reg [31:0] _RAND_232;
  wire  _T_2925;
  wire  _T_2926;
  wire  _T_2927;
  wire  _T_2928;
  wire  _T_2929;
  wire  _T_2930;
  wire  _T_2931;
  wire  _T_2932;
  wire [14:0] _T_2933;
  wire [15:0] _T_2934;
  reg [15:0] _T_2936;
  reg [31:0] _RAND_233;
  wire  _T_2937;
  wire  _T_2938;
  wire  _T_2939;
  wire  _T_2940;
  wire  _T_2941;
  wire  _T_2942;
  wire  _T_2943;
  wire  _T_2944;
  wire [14:0] _T_2945;
  wire [15:0] _T_2946;
  reg [15:0] _T_2948;
  reg [31:0] _RAND_234;
  wire  _T_2949;
  wire  _T_2950;
  wire  _T_2951;
  wire  _T_2952;
  wire  _T_2953;
  wire  _T_2954;
  wire  _T_2955;
  wire  _T_2956;
  wire [14:0] _T_2957;
  wire [15:0] _T_2958;
  reg [15:0] _T_2960;
  reg [31:0] _RAND_235;
  wire  _T_2961;
  wire  _T_2962;
  wire  _T_2963;
  wire  _T_2964;
  wire  _T_2965;
  wire  _T_2966;
  wire  _T_2967;
  wire  _T_2968;
  wire [14:0] _T_2969;
  wire [15:0] _T_2970;
  reg [15:0] _T_2972;
  reg [31:0] _RAND_236;
  wire  _T_2973;
  wire  _T_2974;
  wire  _T_2975;
  wire  _T_2976;
  wire  _T_2977;
  wire  _T_2978;
  wire  _T_2979;
  wire  _T_2980;
  wire [14:0] _T_2981;
  wire [15:0] _T_2982;
  reg [15:0] _T_2984;
  reg [31:0] _RAND_237;
  wire  _T_2985;
  wire  _T_2986;
  wire  _T_2987;
  wire  _T_2988;
  wire  _T_2989;
  wire  _T_2990;
  wire  _T_2991;
  wire  _T_2992;
  wire [14:0] _T_2993;
  wire [15:0] _T_2994;
  reg [15:0] _T_2996;
  reg [31:0] _RAND_238;
  wire  _T_2997;
  wire  _T_2998;
  wire  _T_2999;
  wire  _T_3000;
  wire  _T_3001;
  wire  _T_3002;
  wire  _T_3003;
  wire  _T_3004;
  wire [14:0] _T_3005;
  wire [15:0] _T_3006;
  reg [15:0] _T_3008;
  reg [31:0] _RAND_239;
  wire  _T_3009;
  wire  _T_3010;
  wire  _T_3011;
  wire  _T_3012;
  wire  _T_3013;
  wire  _T_3014;
  wire  _T_3015;
  wire  _T_3016;
  wire [14:0] _T_3017;
  wire [15:0] _T_3018;
  reg [15:0] _T_3020;
  reg [31:0] _RAND_240;
  wire  _T_3021;
  wire  _T_3022;
  wire  _T_3023;
  wire  _T_3024;
  wire  _T_3025;
  wire  _T_3026;
  wire  _T_3027;
  wire  _T_3028;
  wire [14:0] _T_3029;
  wire [15:0] _T_3030;
  reg [15:0] _T_3032;
  reg [31:0] _RAND_241;
  wire  _T_3033;
  wire  _T_3034;
  wire  _T_3035;
  wire  _T_3036;
  wire  _T_3037;
  wire  _T_3038;
  wire  _T_3039;
  wire  _T_3040;
  wire [14:0] _T_3041;
  wire [15:0] _T_3042;
  reg [15:0] _T_3044;
  reg [31:0] _RAND_242;
  wire  _T_3045;
  wire  _T_3046;
  wire  _T_3047;
  wire  _T_3048;
  wire  _T_3049;
  wire  _T_3050;
  wire  _T_3051;
  wire  _T_3052;
  wire [14:0] _T_3053;
  wire [15:0] _T_3054;
  reg [15:0] _T_3056;
  reg [31:0] _RAND_243;
  wire  _T_3057;
  wire  _T_3058;
  wire  _T_3059;
  wire  _T_3060;
  wire  _T_3061;
  wire  _T_3062;
  wire  _T_3063;
  wire  _T_3064;
  wire [14:0] _T_3065;
  wire [15:0] _T_3066;
  reg [15:0] _T_3068;
  reg [31:0] _RAND_244;
  wire  _T_3069;
  wire  _T_3070;
  wire  _T_3071;
  wire  _T_3072;
  wire  _T_3073;
  wire  _T_3074;
  wire  _T_3075;
  wire  _T_3076;
  wire [14:0] _T_3077;
  wire [15:0] _T_3078;
  reg [15:0] _T_3080;
  reg [31:0] _RAND_245;
  wire  _T_3081;
  wire  _T_3082;
  wire  _T_3083;
  wire  _T_3084;
  wire  _T_3085;
  wire  _T_3086;
  wire  _T_3087;
  wire  _T_3088;
  wire [14:0] _T_3089;
  wire [15:0] _T_3090;
  reg [15:0] _T_3092;
  reg [31:0] _RAND_246;
  wire  _T_3093;
  wire  _T_3094;
  wire  _T_3095;
  wire  _T_3096;
  wire  _T_3097;
  wire  _T_3098;
  wire  _T_3099;
  wire  _T_3100;
  wire [14:0] _T_3101;
  wire [15:0] _T_3102;
  reg [15:0] _T_3104;
  reg [31:0] _RAND_247;
  wire  _T_3105;
  wire  _T_3106;
  wire  _T_3107;
  wire  _T_3108;
  wire  _T_3109;
  wire  _T_3110;
  wire  _T_3111;
  wire  _T_3112;
  wire [14:0] _T_3113;
  wire [15:0] _T_3114;
  reg [15:0] _T_3116;
  reg [31:0] _RAND_248;
  wire  _T_3117;
  wire  _T_3118;
  wire  _T_3119;
  wire  _T_3120;
  wire  _T_3121;
  wire  _T_3122;
  wire  _T_3123;
  wire  _T_3124;
  wire [14:0] _T_3125;
  wire [15:0] _T_3126;
  reg [15:0] _T_3128;
  reg [31:0] _RAND_249;
  wire  _T_3129;
  wire  _T_3130;
  wire  _T_3131;
  wire  _T_3132;
  wire  _T_3133;
  wire  _T_3134;
  wire  _T_3135;
  wire  _T_3136;
  wire [14:0] _T_3137;
  wire [15:0] _T_3138;
  reg [15:0] _T_3140;
  reg [31:0] _RAND_250;
  wire  _T_3141;
  wire  _T_3142;
  wire  _T_3143;
  wire  _T_3144;
  wire  _T_3145;
  wire  _T_3146;
  wire  _T_3147;
  wire  _T_3148;
  wire [14:0] _T_3149;
  wire [15:0] _T_3150;
  reg [15:0] _T_3152;
  reg [31:0] _RAND_251;
  wire  _T_3153;
  wire  _T_3154;
  wire  _T_3155;
  wire  _T_3156;
  wire  _T_3157;
  wire  _T_3158;
  wire  _T_3159;
  wire  _T_3160;
  wire [14:0] _T_3161;
  wire [15:0] _T_3162;
  reg [15:0] _T_3164;
  reg [31:0] _RAND_252;
  wire  _T_3165;
  wire  _T_3166;
  wire  _T_3167;
  wire  _T_3168;
  wire  _T_3169;
  wire  _T_3170;
  wire  _T_3171;
  wire  _T_3172;
  wire [14:0] _T_3173;
  wire [15:0] _T_3174;
  reg [15:0] _T_3176;
  reg [31:0] _RAND_253;
  wire  _T_3177;
  wire  _T_3178;
  wire  _T_3179;
  wire  _T_3180;
  wire  _T_3181;
  wire  _T_3182;
  wire  _T_3183;
  wire  _T_3184;
  wire [14:0] _T_3185;
  wire [15:0] _T_3186;
  reg [15:0] _T_3188;
  reg [31:0] _RAND_254;
  wire  _T_3189;
  wire  _T_3190;
  wire  _T_3191;
  wire  _T_3192;
  wire  _T_3193;
  wire  _T_3194;
  wire  _T_3195;
  wire  _T_3196;
  wire [14:0] _T_3197;
  wire [15:0] _T_3198;
  reg [15:0] _T_3200;
  reg [31:0] _RAND_255;
  wire  _T_3201;
  wire  _T_3202;
  wire  _T_3203;
  wire  _T_3204;
  wire  _T_3205;
  wire  _T_3206;
  wire  _T_3207;
  wire  _T_3208;
  wire [14:0] _T_3209;
  wire [15:0] _T_3210;
  reg [15:0] _T_3212;
  reg [31:0] _RAND_256;
  wire  _T_3213;
  wire  _T_3214;
  wire  _T_3215;
  wire  _T_3216;
  wire  _T_3217;
  wire  _T_3218;
  wire  _T_3219;
  wire  _T_3220;
  wire [14:0] _T_3221;
  wire [15:0] _T_3222;
  reg [15:0] _T_3224;
  reg [31:0] _RAND_257;
  wire  _T_3225;
  wire  _T_3226;
  wire  _T_3227;
  wire  _T_3228;
  wire  _T_3229;
  wire  _T_3230;
  wire  _T_3231;
  wire  _T_3232;
  wire [14:0] _T_3233;
  wire [15:0] _T_3234;
  wire [6:0] _T_3243;
  wire [14:0] _T_3251;
  wire [7:0] _T_3258;
  wire [30:0] _T_3267;
  wire [7:0] _T_3274;
  wire [15:0] _T_3282;
  wire [7:0] _T_3289;
  wire [31:0] _T_3298;
  wire [7:0] _T_3306;
  wire [15:0] _T_3314;
  wire [7:0] _T_3321;
  wire [31:0] _T_3330;
  wire [7:0] _T_3337;
  wire [15:0] _T_3345;
  wire [7:0] _T_3352;
  wire [31:0] _T_3361;
  wire [126:0] _T_3363;
  wire [126:0] _GEN_513;
  wire [127:0] _GEN_514;
  wire [127:0] _GEN_515;
  wire [127:0] _GEN_516;
  wire [127:0] _GEN_517;
  wire  _GEN_518;
  wire  _GEN_519;
  wire  _GEN_520;
  wire  _GEN_521;
  wire  _GEN_522;
  wire  _GEN_523;
  wire  _GEN_524;
  wire  _GEN_525;
  wire  _GEN_526;
  wire  _GEN_527;
  wire  _GEN_528;
  wire  _GEN_540;
  wire  _GEN_541;
  wire  _GEN_542;
  wire  _GEN_543;
  wire  _GEN_544;
  wire  _GEN_545;
  wire  _GEN_546;
  wire  _GEN_547;
  wire  _GEN_548;
  SiFive_CoreIPSubsystem system (
    .clock(system_clock),
    .reset(system_reset),
    .debug_psd_test_mode(system_debug_psd_test_mode),
    .debug_psd_test_mode_reset(system_debug_psd_test_mode_reset),
    .debug_systemjtag_jtag_TCK(system_debug_systemjtag_jtag_TCK),
    .debug_systemjtag_jtag_TMS(system_debug_systemjtag_jtag_TMS),
    .debug_systemjtag_jtag_TDI(system_debug_systemjtag_jtag_TDI),
    .debug_systemjtag_jtag_TDO_data(system_debug_systemjtag_jtag_TDO_data),
    .debug_systemjtag_jtag_TDO_driven(system_debug_systemjtag_jtag_TDO_driven),
    .debug_systemjtag_reset(system_debug_systemjtag_reset),
    .debug_systemjtag_mfr_id(system_debug_systemjtag_mfr_id),
    .debug_ndreset(system_debug_ndreset),
    .debug_dmactive(system_debug_dmactive),
    .core_clock_0(system_core_clock_0),
    .reset_vector_0(system_reset_vector_0),
    .rtc_toggle(system_rtc_toggle),
    .global_interrupts(system_global_interrupts),
    .mem_port_axi4_0_aw_ready(system_mem_port_axi4_0_aw_ready),
    .mem_port_axi4_0_aw_valid(system_mem_port_axi4_0_aw_valid),
    .mem_port_axi4_0_aw_bits_id(system_mem_port_axi4_0_aw_bits_id),
    .mem_port_axi4_0_aw_bits_addr(system_mem_port_axi4_0_aw_bits_addr),
    .mem_port_axi4_0_aw_bits_len(system_mem_port_axi4_0_aw_bits_len),
    .mem_port_axi4_0_aw_bits_size(system_mem_port_axi4_0_aw_bits_size),
    .mem_port_axi4_0_aw_bits_burst(system_mem_port_axi4_0_aw_bits_burst),
    .mem_port_axi4_0_aw_bits_lock(system_mem_port_axi4_0_aw_bits_lock),
    .mem_port_axi4_0_aw_bits_cache(system_mem_port_axi4_0_aw_bits_cache),
    .mem_port_axi4_0_aw_bits_prot(system_mem_port_axi4_0_aw_bits_prot),
    .mem_port_axi4_0_aw_bits_qos(system_mem_port_axi4_0_aw_bits_qos),
    .mem_port_axi4_0_w_ready(system_mem_port_axi4_0_w_ready),
    .mem_port_axi4_0_w_valid(system_mem_port_axi4_0_w_valid),
    .mem_port_axi4_0_w_bits_data(system_mem_port_axi4_0_w_bits_data),
    .mem_port_axi4_0_w_bits_strb(system_mem_port_axi4_0_w_bits_strb),
    .mem_port_axi4_0_w_bits_last(system_mem_port_axi4_0_w_bits_last),
    .mem_port_axi4_0_w_bits_corrupt(system_mem_port_axi4_0_w_bits_corrupt),
    .mem_port_axi4_0_b_ready(system_mem_port_axi4_0_b_ready),
    .mem_port_axi4_0_b_valid(system_mem_port_axi4_0_b_valid),
    .mem_port_axi4_0_b_bits_id(system_mem_port_axi4_0_b_bits_id),
    .mem_port_axi4_0_b_bits_resp(system_mem_port_axi4_0_b_bits_resp),
    .mem_port_axi4_0_ar_ready(system_mem_port_axi4_0_ar_ready),
    .mem_port_axi4_0_ar_valid(system_mem_port_axi4_0_ar_valid),
    .mem_port_axi4_0_ar_bits_id(system_mem_port_axi4_0_ar_bits_id),
    .mem_port_axi4_0_ar_bits_addr(system_mem_port_axi4_0_ar_bits_addr),
    .mem_port_axi4_0_ar_bits_len(system_mem_port_axi4_0_ar_bits_len),
    .mem_port_axi4_0_ar_bits_size(system_mem_port_axi4_0_ar_bits_size),
    .mem_port_axi4_0_ar_bits_burst(system_mem_port_axi4_0_ar_bits_burst),
    .mem_port_axi4_0_ar_bits_lock(system_mem_port_axi4_0_ar_bits_lock),
    .mem_port_axi4_0_ar_bits_cache(system_mem_port_axi4_0_ar_bits_cache),
    .mem_port_axi4_0_ar_bits_prot(system_mem_port_axi4_0_ar_bits_prot),
    .mem_port_axi4_0_ar_bits_qos(system_mem_port_axi4_0_ar_bits_qos),
    .mem_port_axi4_0_r_ready(system_mem_port_axi4_0_r_ready),
    .mem_port_axi4_0_r_valid(system_mem_port_axi4_0_r_valid),
    .mem_port_axi4_0_r_bits_id(system_mem_port_axi4_0_r_bits_id),
    .mem_port_axi4_0_r_bits_data(system_mem_port_axi4_0_r_bits_data),
    .mem_port_axi4_0_r_bits_resp(system_mem_port_axi4_0_r_bits_resp),
    .mem_port_axi4_0_r_bits_last(system_mem_port_axi4_0_r_bits_last),
    .sys_port_axi4_0_aw_ready(system_sys_port_axi4_0_aw_ready),
    .sys_port_axi4_0_aw_valid(system_sys_port_axi4_0_aw_valid),
    .sys_port_axi4_0_aw_bits_id(system_sys_port_axi4_0_aw_bits_id),
    .sys_port_axi4_0_aw_bits_addr(system_sys_port_axi4_0_aw_bits_addr),
    .sys_port_axi4_0_aw_bits_len(system_sys_port_axi4_0_aw_bits_len),
    .sys_port_axi4_0_aw_bits_size(system_sys_port_axi4_0_aw_bits_size),
    .sys_port_axi4_0_aw_bits_burst(system_sys_port_axi4_0_aw_bits_burst),
    .sys_port_axi4_0_aw_bits_lock(system_sys_port_axi4_0_aw_bits_lock),
    .sys_port_axi4_0_aw_bits_cache(system_sys_port_axi4_0_aw_bits_cache),
    .sys_port_axi4_0_aw_bits_prot(system_sys_port_axi4_0_aw_bits_prot),
    .sys_port_axi4_0_aw_bits_qos(system_sys_port_axi4_0_aw_bits_qos),
    .sys_port_axi4_0_w_ready(system_sys_port_axi4_0_w_ready),
    .sys_port_axi4_0_w_valid(system_sys_port_axi4_0_w_valid),
    .sys_port_axi4_0_w_bits_data(system_sys_port_axi4_0_w_bits_data),
    .sys_port_axi4_0_w_bits_strb(system_sys_port_axi4_0_w_bits_strb),
    .sys_port_axi4_0_w_bits_last(system_sys_port_axi4_0_w_bits_last),
    .sys_port_axi4_0_b_ready(system_sys_port_axi4_0_b_ready),
    .sys_port_axi4_0_b_valid(system_sys_port_axi4_0_b_valid),
    .sys_port_axi4_0_b_bits_id(system_sys_port_axi4_0_b_bits_id),
    .sys_port_axi4_0_b_bits_resp(system_sys_port_axi4_0_b_bits_resp),
    .sys_port_axi4_0_ar_ready(system_sys_port_axi4_0_ar_ready),
    .sys_port_axi4_0_ar_valid(system_sys_port_axi4_0_ar_valid),
    .sys_port_axi4_0_ar_bits_id(system_sys_port_axi4_0_ar_bits_id),
    .sys_port_axi4_0_ar_bits_addr(system_sys_port_axi4_0_ar_bits_addr),
    .sys_port_axi4_0_ar_bits_len(system_sys_port_axi4_0_ar_bits_len),
    .sys_port_axi4_0_ar_bits_size(system_sys_port_axi4_0_ar_bits_size),
    .sys_port_axi4_0_ar_bits_burst(system_sys_port_axi4_0_ar_bits_burst),
    .sys_port_axi4_0_ar_bits_lock(system_sys_port_axi4_0_ar_bits_lock),
    .sys_port_axi4_0_ar_bits_cache(system_sys_port_axi4_0_ar_bits_cache),
    .sys_port_axi4_0_ar_bits_prot(system_sys_port_axi4_0_ar_bits_prot),
    .sys_port_axi4_0_ar_bits_qos(system_sys_port_axi4_0_ar_bits_qos),
    .sys_port_axi4_0_r_ready(system_sys_port_axi4_0_r_ready),
    .sys_port_axi4_0_r_valid(system_sys_port_axi4_0_r_valid),
    .sys_port_axi4_0_r_bits_id(system_sys_port_axi4_0_r_bits_id),
    .sys_port_axi4_0_r_bits_data(system_sys_port_axi4_0_r_bits_data),
    .sys_port_axi4_0_r_bits_resp(system_sys_port_axi4_0_r_bits_resp),
    .sys_port_axi4_0_r_bits_last(system_sys_port_axi4_0_r_bits_last),
    .periph_port_axi4_0_aw_ready(system_periph_port_axi4_0_aw_ready),
    .periph_port_axi4_0_aw_valid(system_periph_port_axi4_0_aw_valid),
    .periph_port_axi4_0_aw_bits_id(system_periph_port_axi4_0_aw_bits_id),
    .periph_port_axi4_0_aw_bits_addr(system_periph_port_axi4_0_aw_bits_addr),
    .periph_port_axi4_0_aw_bits_len(system_periph_port_axi4_0_aw_bits_len),
    .periph_port_axi4_0_aw_bits_size(system_periph_port_axi4_0_aw_bits_size),
    .periph_port_axi4_0_aw_bits_burst(system_periph_port_axi4_0_aw_bits_burst),
    .periph_port_axi4_0_aw_bits_lock(system_periph_port_axi4_0_aw_bits_lock),
    .periph_port_axi4_0_aw_bits_cache(system_periph_port_axi4_0_aw_bits_cache),
    .periph_port_axi4_0_aw_bits_prot(system_periph_port_axi4_0_aw_bits_prot),
    .periph_port_axi4_0_aw_bits_qos(system_periph_port_axi4_0_aw_bits_qos),
    .periph_port_axi4_0_w_ready(system_periph_port_axi4_0_w_ready),
    .periph_port_axi4_0_w_valid(system_periph_port_axi4_0_w_valid),
    .periph_port_axi4_0_w_bits_data(system_periph_port_axi4_0_w_bits_data),
    .periph_port_axi4_0_w_bits_strb(system_periph_port_axi4_0_w_bits_strb),
    .periph_port_axi4_0_w_bits_last(system_periph_port_axi4_0_w_bits_last),
    .periph_port_axi4_0_b_ready(system_periph_port_axi4_0_b_ready),
    .periph_port_axi4_0_b_valid(system_periph_port_axi4_0_b_valid),
    .periph_port_axi4_0_b_bits_id(system_periph_port_axi4_0_b_bits_id),
    .periph_port_axi4_0_b_bits_resp(system_periph_port_axi4_0_b_bits_resp),
    .periph_port_axi4_0_ar_ready(system_periph_port_axi4_0_ar_ready),
    .periph_port_axi4_0_ar_valid(system_periph_port_axi4_0_ar_valid),
    .periph_port_axi4_0_ar_bits_id(system_periph_port_axi4_0_ar_bits_id),
    .periph_port_axi4_0_ar_bits_addr(system_periph_port_axi4_0_ar_bits_addr),
    .periph_port_axi4_0_ar_bits_len(system_periph_port_axi4_0_ar_bits_len),
    .periph_port_axi4_0_ar_bits_size(system_periph_port_axi4_0_ar_bits_size),
    .periph_port_axi4_0_ar_bits_burst(system_periph_port_axi4_0_ar_bits_burst),
    .periph_port_axi4_0_ar_bits_lock(system_periph_port_axi4_0_ar_bits_lock),
    .periph_port_axi4_0_ar_bits_cache(system_periph_port_axi4_0_ar_bits_cache),
    .periph_port_axi4_0_ar_bits_prot(system_periph_port_axi4_0_ar_bits_prot),
    .periph_port_axi4_0_ar_bits_qos(system_periph_port_axi4_0_ar_bits_qos),
    .periph_port_axi4_0_r_ready(system_periph_port_axi4_0_r_ready),
    .periph_port_axi4_0_r_valid(system_periph_port_axi4_0_r_valid),
    .periph_port_axi4_0_r_bits_id(system_periph_port_axi4_0_r_bits_id),
    .periph_port_axi4_0_r_bits_data(system_periph_port_axi4_0_r_bits_data),
    .periph_port_axi4_0_r_bits_resp(system_periph_port_axi4_0_r_bits_resp),
    .periph_port_axi4_0_r_bits_last(system_periph_port_axi4_0_r_bits_last),
    .front_port_axi4_0_aw_ready(system_front_port_axi4_0_aw_ready),
    .front_port_axi4_0_aw_valid(system_front_port_axi4_0_aw_valid),
    .front_port_axi4_0_aw_bits_id(system_front_port_axi4_0_aw_bits_id),
    .front_port_axi4_0_aw_bits_addr(system_front_port_axi4_0_aw_bits_addr),
    .front_port_axi4_0_aw_bits_len(system_front_port_axi4_0_aw_bits_len),
    .front_port_axi4_0_aw_bits_size(system_front_port_axi4_0_aw_bits_size),
    .front_port_axi4_0_aw_bits_burst(system_front_port_axi4_0_aw_bits_burst),
    .front_port_axi4_0_aw_bits_lock(system_front_port_axi4_0_aw_bits_lock),
    .front_port_axi4_0_aw_bits_cache(system_front_port_axi4_0_aw_bits_cache),
    .front_port_axi4_0_aw_bits_prot(system_front_port_axi4_0_aw_bits_prot),
    .front_port_axi4_0_aw_bits_qos(system_front_port_axi4_0_aw_bits_qos),
    .front_port_axi4_0_w_ready(system_front_port_axi4_0_w_ready),
    .front_port_axi4_0_w_valid(system_front_port_axi4_0_w_valid),
    .front_port_axi4_0_w_bits_data(system_front_port_axi4_0_w_bits_data),
    .front_port_axi4_0_w_bits_strb(system_front_port_axi4_0_w_bits_strb),
    .front_port_axi4_0_w_bits_last(system_front_port_axi4_0_w_bits_last),
    .front_port_axi4_0_b_ready(system_front_port_axi4_0_b_ready),
    .front_port_axi4_0_b_valid(system_front_port_axi4_0_b_valid),
    .front_port_axi4_0_b_bits_id(system_front_port_axi4_0_b_bits_id),
    .front_port_axi4_0_b_bits_resp(system_front_port_axi4_0_b_bits_resp),
    .front_port_axi4_0_ar_ready(system_front_port_axi4_0_ar_ready),
    .front_port_axi4_0_ar_valid(system_front_port_axi4_0_ar_valid),
    .front_port_axi4_0_ar_bits_id(system_front_port_axi4_0_ar_bits_id),
    .front_port_axi4_0_ar_bits_addr(system_front_port_axi4_0_ar_bits_addr),
    .front_port_axi4_0_ar_bits_len(system_front_port_axi4_0_ar_bits_len),
    .front_port_axi4_0_ar_bits_size(system_front_port_axi4_0_ar_bits_size),
    .front_port_axi4_0_ar_bits_burst(system_front_port_axi4_0_ar_bits_burst),
    .front_port_axi4_0_ar_bits_lock(system_front_port_axi4_0_ar_bits_lock),
    .front_port_axi4_0_ar_bits_cache(system_front_port_axi4_0_ar_bits_cache),
    .front_port_axi4_0_ar_bits_prot(system_front_port_axi4_0_ar_bits_prot),
    .front_port_axi4_0_ar_bits_qos(system_front_port_axi4_0_ar_bits_qos),
    .front_port_axi4_0_r_ready(system_front_port_axi4_0_r_ready),
    .front_port_axi4_0_r_valid(system_front_port_axi4_0_r_valid),
    .front_port_axi4_0_r_bits_id(system_front_port_axi4_0_r_bits_id),
    .front_port_axi4_0_r_bits_data(system_front_port_axi4_0_r_bits_data),
    .front_port_axi4_0_r_bits_resp(system_front_port_axi4_0_r_bits_resp),
    .front_port_axi4_0_r_bits_last(system_front_port_axi4_0_r_bits_last)
  );
  Pow2ClockDivider func_clock (
    .clock(func_clock_clock),
    .io_clock_out(func_clock_io_clock_out)
  );
  ClockSkew #(.DELAY_RTL(0.0), .DELAY_GL(0.0)) ClockSkew (
    .clkin(ClockSkew_clkin),
    .clkout(ClockSkew_clkout)
  );
  Pow2ClockDivider_1 Pow2ClockDivider (
    .clock(Pow2ClockDivider_clock),
    .io_clock_out(Pow2ClockDivider_io_clock_out)
  );
  system_clock_en dpiClockGate (
    .clock_in(dpiClockGate_clock_in),
    .clock_out(dpiClockGate_clock_out)
  );
  c_core_reset_driver c_core_reset_driver (
    .clock(c_core_reset_driver_clock)
  );
  DataTap_5 DataTap_5 (
    ._1_clock(DataTap_5__1_clock),
    ._1_reset(DataTap_5__1_reset),
    ._1_hartid(DataTap_5__1_hartid),
    ._1_timer(DataTap_5__1_timer),
    ._1_valid(DataTap_5__1_valid),
    ._1_pc(DataTap_5__1_pc),
    ._1_wrdst(DataTap_5__1_wrdst),
    ._1_wrdata(DataTap_5__1_wrdata),
    ._1_wren(DataTap_5__1_wren),
    ._1_rd0src(DataTap_5__1_rd0src),
    ._1_rd0val(DataTap_5__1_rd0val),
    ._1_rd1src(DataTap_5__1_rd1src),
    ._1_rd1val(DataTap_5__1_rd1val),
    ._1_inst(DataTap_5__1_inst),
    ._0_clock(DataTap_5__0_clock),
    ._0_reset(DataTap_5__0_reset),
    ._0_hartid(DataTap_5__0_hartid),
    ._0_timer(DataTap_5__0_timer),
    ._0_valid(DataTap_5__0_valid),
    ._0_pc(DataTap_5__0_pc),
    ._0_wrdst(DataTap_5__0_wrdst),
    ._0_wrdata(DataTap_5__0_wrdata),
    ._0_wren(DataTap_5__0_wren),
    ._0_rd0src(DataTap_5__0_rd0src),
    ._0_rd0val(DataTap_5__0_rd0val),
    ._0_rd1src(DataTap_5__0_rd1src),
    ._0_rd1val(DataTap_5__0_rd1val),
    ._0_inst(DataTap_5__0_inst)
  );
  AXI4PortRAMSlave testRAM (
    .clock(testRAM_clock),
    .reset(testRAM_reset),
    .io_axi4_0_aw_ready(testRAM_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(testRAM_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(testRAM_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(testRAM_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(testRAM_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(testRAM_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(testRAM_io_axi4_0_aw_bits_burst),
    .io_axi4_0_aw_bits_lock(testRAM_io_axi4_0_aw_bits_lock),
    .io_axi4_0_aw_bits_cache(testRAM_io_axi4_0_aw_bits_cache),
    .io_axi4_0_aw_bits_prot(testRAM_io_axi4_0_aw_bits_prot),
    .io_axi4_0_aw_bits_qos(testRAM_io_axi4_0_aw_bits_qos),
    .io_axi4_0_w_ready(testRAM_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(testRAM_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(testRAM_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(testRAM_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(testRAM_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(testRAM_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(testRAM_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(testRAM_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(testRAM_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(testRAM_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(testRAM_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(testRAM_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(testRAM_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(testRAM_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(testRAM_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(testRAM_io_axi4_0_ar_bits_burst),
    .io_axi4_0_ar_bits_lock(testRAM_io_axi4_0_ar_bits_lock),
    .io_axi4_0_ar_bits_cache(testRAM_io_axi4_0_ar_bits_cache),
    .io_axi4_0_ar_bits_prot(testRAM_io_axi4_0_ar_bits_prot),
    .io_axi4_0_ar_bits_qos(testRAM_io_axi4_0_ar_bits_qos),
    .io_axi4_0_r_ready(testRAM_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(testRAM_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(testRAM_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(testRAM_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(testRAM_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(testRAM_io_axi4_0_r_bits_last)
  );
  AXI4PortRAMSlave_1 testRAM_1 (
    .clock(testRAM_1_clock),
    .reset(testRAM_1_reset),
    .io_axi4_0_aw_ready(testRAM_1_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(testRAM_1_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(testRAM_1_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(testRAM_1_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(testRAM_1_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(testRAM_1_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(testRAM_1_io_axi4_0_aw_bits_burst),
    .io_axi4_0_aw_bits_lock(testRAM_1_io_axi4_0_aw_bits_lock),
    .io_axi4_0_aw_bits_cache(testRAM_1_io_axi4_0_aw_bits_cache),
    .io_axi4_0_aw_bits_prot(testRAM_1_io_axi4_0_aw_bits_prot),
    .io_axi4_0_aw_bits_qos(testRAM_1_io_axi4_0_aw_bits_qos),
    .io_axi4_0_w_ready(testRAM_1_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(testRAM_1_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(testRAM_1_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(testRAM_1_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(testRAM_1_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(testRAM_1_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(testRAM_1_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(testRAM_1_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(testRAM_1_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(testRAM_1_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(testRAM_1_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(testRAM_1_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(testRAM_1_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(testRAM_1_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(testRAM_1_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(testRAM_1_io_axi4_0_ar_bits_burst),
    .io_axi4_0_ar_bits_lock(testRAM_1_io_axi4_0_ar_bits_lock),
    .io_axi4_0_ar_bits_cache(testRAM_1_io_axi4_0_ar_bits_cache),
    .io_axi4_0_ar_bits_prot(testRAM_1_io_axi4_0_ar_bits_prot),
    .io_axi4_0_ar_bits_qos(testRAM_1_io_axi4_0_ar_bits_qos),
    .io_axi4_0_r_ready(testRAM_1_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(testRAM_1_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(testRAM_1_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(testRAM_1_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(testRAM_1_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(testRAM_1_io_axi4_0_r_bits_last)
  );
  AXI4PortRAMSlave_2 testRAM_2 (
    .clock(testRAM_2_clock),
    .reset(testRAM_2_reset),
    .io_axi4_0_aw_ready(testRAM_2_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(testRAM_2_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(testRAM_2_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(testRAM_2_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(testRAM_2_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(testRAM_2_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(testRAM_2_io_axi4_0_aw_bits_burst),
    .io_axi4_0_aw_bits_lock(testRAM_2_io_axi4_0_aw_bits_lock),
    .io_axi4_0_aw_bits_cache(testRAM_2_io_axi4_0_aw_bits_cache),
    .io_axi4_0_aw_bits_prot(testRAM_2_io_axi4_0_aw_bits_prot),
    .io_axi4_0_aw_bits_qos(testRAM_2_io_axi4_0_aw_bits_qos),
    .io_axi4_0_w_ready(testRAM_2_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(testRAM_2_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(testRAM_2_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(testRAM_2_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(testRAM_2_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(testRAM_2_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(testRAM_2_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(testRAM_2_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(testRAM_2_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(testRAM_2_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(testRAM_2_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(testRAM_2_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(testRAM_2_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(testRAM_2_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(testRAM_2_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(testRAM_2_io_axi4_0_ar_bits_burst),
    .io_axi4_0_ar_bits_lock(testRAM_2_io_axi4_0_ar_bits_lock),
    .io_axi4_0_ar_bits_cache(testRAM_2_io_axi4_0_ar_bits_cache),
    .io_axi4_0_ar_bits_prot(testRAM_2_io_axi4_0_ar_bits_prot),
    .io_axi4_0_ar_bits_qos(testRAM_2_io_axi4_0_ar_bits_qos),
    .io_axi4_0_r_ready(testRAM_2_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(testRAM_2_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(testRAM_2_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(testRAM_2_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(testRAM_2_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(testRAM_2_io_axi4_0_r_bits_last)
  );
  DPIJTAGDriver DPIJTAGDriver (
    .clock(DPIJTAGDriver_clock),
    .reset(DPIJTAGDriver_reset),
    .jtag_TRSTn(DPIJTAGDriver_jtag_TRSTn),
    .jtag_TCK(DPIJTAGDriver_jtag_TCK),
    .jtag_TMS(DPIJTAGDriver_jtag_TMS),
    .jtag_TDI(DPIJTAGDriver_jtag_TDI),
    .jtag_TDO_data(DPIJTAGDriver_jtag_TDO_data),
    .jtag_TDO_driven(DPIJTAGDriver_jtag_TDO_driven)
  );
  system_reset_driver system_reset_driver (
    .clock(system_reset_driver_clock),
    .out(system_reset_driver_out)
  );
  plusarg_reader #(.FORMAT("system_reset_delay=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  CountAndDriver CountAndDriver (
    .clock(CountAndDriver_clock),
    .reset(CountAndDriver_reset),
    .io_default_value(CountAndDriver_io_default_value),
    .io_count(CountAndDriver_io_count),
    .io_driven_value(CountAndDriver_io_driven_value)
  );
  core_reset_driver core_reset_driver (
    .clock(core_reset_driver_clock)
  );
  core_monitor core_monitor (
    .m_0_clock(core_monitor_m_0_clock),
    .m_0_reset(core_monitor_m_0_reset),
    .m_0_hartid(core_monitor_m_0_hartid),
    .m_0_timer(core_monitor_m_0_timer),
    .m_0_valid(core_monitor_m_0_valid),
    .m_0_pc(core_monitor_m_0_pc),
    .m_0_wrdst(core_monitor_m_0_wrdst),
    .m_0_wrdata(core_monitor_m_0_wrdata),
    .m_0_wren(core_monitor_m_0_wren),
    .m_0_rd0src(core_monitor_m_0_rd0src),
    .m_0_rd0val(core_monitor_m_0_rd0val),
    .m_0_rd1src(core_monitor_m_0_rd1src),
    .m_0_rd1val(core_monitor_m_0_rd1val),
    .m_0_inst(core_monitor_m_0_inst),
    .m_1_clock(core_monitor_m_1_clock),
    .m_1_reset(core_monitor_m_1_reset),
    .m_1_hartid(core_monitor_m_1_hartid),
    .m_1_timer(core_monitor_m_1_timer),
    .m_1_valid(core_monitor_m_1_valid),
    .m_1_pc(core_monitor_m_1_pc),
    .m_1_wrdst(core_monitor_m_1_wrdst),
    .m_1_wrdata(core_monitor_m_1_wrdata),
    .m_1_wren(core_monitor_m_1_wren),
    .m_1_rd0src(core_monitor_m_1_rd0src),
    .m_1_rd0val(core_monitor_m_1_rd0val),
    .m_1_rd1src(core_monitor_m_1_rd1src),
    .m_1_rd1val(core_monitor_m_1_rd1val),
    .m_1_inst(core_monitor_m_1_inst)
  );
  plusarg_reader #(.FORMAT("drive_local_interrupt_type=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 (
    .out(plusarg_reader_1_out)
  );
  InterruptsDriver InterruptsDriver (
    .clock(InterruptsDriver_clock),
    .reset(InterruptsDriver_reset)
  );
  DPITestbenchHooks dpitbh (
    .clock(dpitbh_clock),
    .reset(dpitbh_reset)
  );
  plusarg_reader #(.FORMAT("drive_global_interrupt_type=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_2 (
    .out(plusarg_reader_2_out)
  );
  assign _T_3 = _T + 5'h1;
  assign _T_4 = _T == 5'h0;
  assign _T_5 = ~ _T_1;
  assign _T_14 = system_debug_ndreset;
  assign ndm_reset = reset | _T_14;
  assign _T_28 = system_reset_driver_out;
  assign _T_30 = plusarg_reader_1_out;
  assign _T_34 = _T_30 == 32'h0;
  assign _T_35 = _T_30 == 32'h1;
  assign _T_36 = _T_30 == 32'h2;
  assign _T_37 = _T_30 == 32'h3;
  assign _T_38 = _T_30 == 32'h4;
  assign _T_39 = _T_30 == 32'h5;
  assign _T_43 = reset == 1'h0;
  assign _T_45 = value_1 == 7'h63;
  assign _T_47 = value_1 + 7'h1;
  assign _T_44 = plusarg_reader_2_out;
  assign _T_48 = _T_44 == 32'h0;
  assign _T_49 = _T_44 == 32'h1;
  assign _T_51 = _T_44 == 32'h2;
  assign _T_179 = _T_44 == 32'h3;
  assign _T_180 = value_2 == 7'h7e;
  assign _T_182 = value_2 + 7'h1;
  assign _T_184 = 128'h1 << value_2;
  assign _T_185 = _T_44 == 32'h4;
  assign _T_187 = _T_186 == 16'h0;
  assign _T_188 = _T_186[0];
  assign _T_189 = _T_186[2];
  assign _T_190 = _T_188 ^ _T_189;
  assign _T_191 = _T_186[3];
  assign _T_192 = _T_190 ^ _T_191;
  assign _T_193 = _T_186[5];
  assign _T_194 = _T_192 ^ _T_193;
  assign _T_195 = _T_186[15:1];
  assign _T_196 = {_T_194,_T_195};
  assign _T_199 = _T_198 == 16'h0;
  assign _T_200 = _T_198[0];
  assign _T_201 = _T_198[2];
  assign _T_202 = _T_200 ^ _T_201;
  assign _T_203 = _T_198[3];
  assign _T_204 = _T_202 ^ _T_203;
  assign _T_205 = _T_198[5];
  assign _T_206 = _T_204 ^ _T_205;
  assign _T_207 = _T_198[15:1];
  assign _T_208 = {_T_206,_T_207};
  assign _T_211 = _T_210 == 16'h0;
  assign _T_212 = _T_210[0];
  assign _T_213 = _T_210[2];
  assign _T_214 = _T_212 ^ _T_213;
  assign _T_215 = _T_210[3];
  assign _T_216 = _T_214 ^ _T_215;
  assign _T_217 = _T_210[5];
  assign _T_218 = _T_216 ^ _T_217;
  assign _T_219 = _T_210[15:1];
  assign _T_220 = {_T_218,_T_219};
  assign _T_223 = _T_222 == 16'h0;
  assign _T_224 = _T_222[0];
  assign _T_225 = _T_222[2];
  assign _T_226 = _T_224 ^ _T_225;
  assign _T_227 = _T_222[3];
  assign _T_228 = _T_226 ^ _T_227;
  assign _T_229 = _T_222[5];
  assign _T_230 = _T_228 ^ _T_229;
  assign _T_231 = _T_222[15:1];
  assign _T_232 = {_T_230,_T_231};
  assign _T_235 = _T_234 == 16'h0;
  assign _T_236 = _T_234[0];
  assign _T_237 = _T_234[2];
  assign _T_238 = _T_236 ^ _T_237;
  assign _T_239 = _T_234[3];
  assign _T_240 = _T_238 ^ _T_239;
  assign _T_241 = _T_234[5];
  assign _T_242 = _T_240 ^ _T_241;
  assign _T_243 = _T_234[15:1];
  assign _T_244 = {_T_242,_T_243};
  assign _T_247 = _T_246 == 16'h0;
  assign _T_248 = _T_246[0];
  assign _T_249 = _T_246[2];
  assign _T_250 = _T_248 ^ _T_249;
  assign _T_251 = _T_246[3];
  assign _T_252 = _T_250 ^ _T_251;
  assign _T_253 = _T_246[5];
  assign _T_254 = _T_252 ^ _T_253;
  assign _T_255 = _T_246[15:1];
  assign _T_256 = {_T_254,_T_255};
  assign _T_259 = _T_258 == 16'h0;
  assign _T_260 = _T_258[0];
  assign _T_261 = _T_258[2];
  assign _T_262 = _T_260 ^ _T_261;
  assign _T_263 = _T_258[3];
  assign _T_264 = _T_262 ^ _T_263;
  assign _T_265 = _T_258[5];
  assign _T_266 = _T_264 ^ _T_265;
  assign _T_267 = _T_258[15:1];
  assign _T_268 = {_T_266,_T_267};
  assign _T_271 = _T_270 == 16'h0;
  assign _T_272 = _T_270[0];
  assign _T_273 = _T_270[2];
  assign _T_274 = _T_272 ^ _T_273;
  assign _T_275 = _T_270[3];
  assign _T_276 = _T_274 ^ _T_275;
  assign _T_277 = _T_270[5];
  assign _T_278 = _T_276 ^ _T_277;
  assign _T_279 = _T_270[15:1];
  assign _T_280 = {_T_278,_T_279};
  assign _T_283 = _T_282 == 16'h0;
  assign _T_284 = _T_282[0];
  assign _T_285 = _T_282[2];
  assign _T_286 = _T_284 ^ _T_285;
  assign _T_287 = _T_282[3];
  assign _T_288 = _T_286 ^ _T_287;
  assign _T_289 = _T_282[5];
  assign _T_290 = _T_288 ^ _T_289;
  assign _T_291 = _T_282[15:1];
  assign _T_292 = {_T_290,_T_291};
  assign _T_295 = _T_294 == 16'h0;
  assign _T_296 = _T_294[0];
  assign _T_297 = _T_294[2];
  assign _T_298 = _T_296 ^ _T_297;
  assign _T_299 = _T_294[3];
  assign _T_300 = _T_298 ^ _T_299;
  assign _T_301 = _T_294[5];
  assign _T_302 = _T_300 ^ _T_301;
  assign _T_303 = _T_294[15:1];
  assign _T_304 = {_T_302,_T_303};
  assign _T_307 = _T_306 == 16'h0;
  assign _T_308 = _T_306[0];
  assign _T_309 = _T_306[2];
  assign _T_310 = _T_308 ^ _T_309;
  assign _T_311 = _T_306[3];
  assign _T_312 = _T_310 ^ _T_311;
  assign _T_313 = _T_306[5];
  assign _T_314 = _T_312 ^ _T_313;
  assign _T_315 = _T_306[15:1];
  assign _T_316 = {_T_314,_T_315};
  assign _T_319 = _T_318 == 16'h0;
  assign _T_320 = _T_318[0];
  assign _T_321 = _T_318[2];
  assign _T_322 = _T_320 ^ _T_321;
  assign _T_323 = _T_318[3];
  assign _T_324 = _T_322 ^ _T_323;
  assign _T_325 = _T_318[5];
  assign _T_326 = _T_324 ^ _T_325;
  assign _T_327 = _T_318[15:1];
  assign _T_328 = {_T_326,_T_327};
  assign _T_331 = _T_330 == 16'h0;
  assign _T_332 = _T_330[0];
  assign _T_333 = _T_330[2];
  assign _T_334 = _T_332 ^ _T_333;
  assign _T_335 = _T_330[3];
  assign _T_336 = _T_334 ^ _T_335;
  assign _T_337 = _T_330[5];
  assign _T_338 = _T_336 ^ _T_337;
  assign _T_339 = _T_330[15:1];
  assign _T_340 = {_T_338,_T_339};
  assign _T_343 = _T_342 == 16'h0;
  assign _T_344 = _T_342[0];
  assign _T_345 = _T_342[2];
  assign _T_346 = _T_344 ^ _T_345;
  assign _T_347 = _T_342[3];
  assign _T_348 = _T_346 ^ _T_347;
  assign _T_349 = _T_342[5];
  assign _T_350 = _T_348 ^ _T_349;
  assign _T_351 = _T_342[15:1];
  assign _T_352 = {_T_350,_T_351};
  assign _T_355 = _T_354 == 16'h0;
  assign _T_356 = _T_354[0];
  assign _T_357 = _T_354[2];
  assign _T_358 = _T_356 ^ _T_357;
  assign _T_359 = _T_354[3];
  assign _T_360 = _T_358 ^ _T_359;
  assign _T_361 = _T_354[5];
  assign _T_362 = _T_360 ^ _T_361;
  assign _T_363 = _T_354[15:1];
  assign _T_364 = {_T_362,_T_363};
  assign _T_367 = _T_366 == 16'h0;
  assign _T_368 = _T_366[0];
  assign _T_369 = _T_366[2];
  assign _T_370 = _T_368 ^ _T_369;
  assign _T_371 = _T_366[3];
  assign _T_372 = _T_370 ^ _T_371;
  assign _T_373 = _T_366[5];
  assign _T_374 = _T_372 ^ _T_373;
  assign _T_375 = _T_366[15:1];
  assign _T_376 = {_T_374,_T_375};
  assign _T_379 = _T_378 == 16'h0;
  assign _T_380 = _T_378[0];
  assign _T_381 = _T_378[2];
  assign _T_382 = _T_380 ^ _T_381;
  assign _T_383 = _T_378[3];
  assign _T_384 = _T_382 ^ _T_383;
  assign _T_385 = _T_378[5];
  assign _T_386 = _T_384 ^ _T_385;
  assign _T_387 = _T_378[15:1];
  assign _T_388 = {_T_386,_T_387};
  assign _T_391 = _T_390 == 16'h0;
  assign _T_392 = _T_390[0];
  assign _T_393 = _T_390[2];
  assign _T_394 = _T_392 ^ _T_393;
  assign _T_395 = _T_390[3];
  assign _T_396 = _T_394 ^ _T_395;
  assign _T_397 = _T_390[5];
  assign _T_398 = _T_396 ^ _T_397;
  assign _T_399 = _T_390[15:1];
  assign _T_400 = {_T_398,_T_399};
  assign _T_403 = _T_402 == 16'h0;
  assign _T_404 = _T_402[0];
  assign _T_405 = _T_402[2];
  assign _T_406 = _T_404 ^ _T_405;
  assign _T_407 = _T_402[3];
  assign _T_408 = _T_406 ^ _T_407;
  assign _T_409 = _T_402[5];
  assign _T_410 = _T_408 ^ _T_409;
  assign _T_411 = _T_402[15:1];
  assign _T_412 = {_T_410,_T_411};
  assign _T_415 = _T_414 == 16'h0;
  assign _T_416 = _T_414[0];
  assign _T_417 = _T_414[2];
  assign _T_418 = _T_416 ^ _T_417;
  assign _T_419 = _T_414[3];
  assign _T_420 = _T_418 ^ _T_419;
  assign _T_421 = _T_414[5];
  assign _T_422 = _T_420 ^ _T_421;
  assign _T_423 = _T_414[15:1];
  assign _T_424 = {_T_422,_T_423};
  assign _T_427 = _T_426 == 16'h0;
  assign _T_428 = _T_426[0];
  assign _T_429 = _T_426[2];
  assign _T_430 = _T_428 ^ _T_429;
  assign _T_431 = _T_426[3];
  assign _T_432 = _T_430 ^ _T_431;
  assign _T_433 = _T_426[5];
  assign _T_434 = _T_432 ^ _T_433;
  assign _T_435 = _T_426[15:1];
  assign _T_436 = {_T_434,_T_435};
  assign _T_439 = _T_438 == 16'h0;
  assign _T_440 = _T_438[0];
  assign _T_441 = _T_438[2];
  assign _T_442 = _T_440 ^ _T_441;
  assign _T_443 = _T_438[3];
  assign _T_444 = _T_442 ^ _T_443;
  assign _T_445 = _T_438[5];
  assign _T_446 = _T_444 ^ _T_445;
  assign _T_447 = _T_438[15:1];
  assign _T_448 = {_T_446,_T_447};
  assign _T_451 = _T_450 == 16'h0;
  assign _T_452 = _T_450[0];
  assign _T_453 = _T_450[2];
  assign _T_454 = _T_452 ^ _T_453;
  assign _T_455 = _T_450[3];
  assign _T_456 = _T_454 ^ _T_455;
  assign _T_457 = _T_450[5];
  assign _T_458 = _T_456 ^ _T_457;
  assign _T_459 = _T_450[15:1];
  assign _T_460 = {_T_458,_T_459};
  assign _T_463 = _T_462 == 16'h0;
  assign _T_464 = _T_462[0];
  assign _T_465 = _T_462[2];
  assign _T_466 = _T_464 ^ _T_465;
  assign _T_467 = _T_462[3];
  assign _T_468 = _T_466 ^ _T_467;
  assign _T_469 = _T_462[5];
  assign _T_470 = _T_468 ^ _T_469;
  assign _T_471 = _T_462[15:1];
  assign _T_472 = {_T_470,_T_471};
  assign _T_475 = _T_474 == 16'h0;
  assign _T_476 = _T_474[0];
  assign _T_477 = _T_474[2];
  assign _T_478 = _T_476 ^ _T_477;
  assign _T_479 = _T_474[3];
  assign _T_480 = _T_478 ^ _T_479;
  assign _T_481 = _T_474[5];
  assign _T_482 = _T_480 ^ _T_481;
  assign _T_483 = _T_474[15:1];
  assign _T_484 = {_T_482,_T_483};
  assign _T_487 = _T_486 == 16'h0;
  assign _T_488 = _T_486[0];
  assign _T_489 = _T_486[2];
  assign _T_490 = _T_488 ^ _T_489;
  assign _T_491 = _T_486[3];
  assign _T_492 = _T_490 ^ _T_491;
  assign _T_493 = _T_486[5];
  assign _T_494 = _T_492 ^ _T_493;
  assign _T_495 = _T_486[15:1];
  assign _T_496 = {_T_494,_T_495};
  assign _T_499 = _T_498 == 16'h0;
  assign _T_500 = _T_498[0];
  assign _T_501 = _T_498[2];
  assign _T_502 = _T_500 ^ _T_501;
  assign _T_503 = _T_498[3];
  assign _T_504 = _T_502 ^ _T_503;
  assign _T_505 = _T_498[5];
  assign _T_506 = _T_504 ^ _T_505;
  assign _T_507 = _T_498[15:1];
  assign _T_508 = {_T_506,_T_507};
  assign _T_511 = _T_510 == 16'h0;
  assign _T_512 = _T_510[0];
  assign _T_513 = _T_510[2];
  assign _T_514 = _T_512 ^ _T_513;
  assign _T_515 = _T_510[3];
  assign _T_516 = _T_514 ^ _T_515;
  assign _T_517 = _T_510[5];
  assign _T_518 = _T_516 ^ _T_517;
  assign _T_519 = _T_510[15:1];
  assign _T_520 = {_T_518,_T_519};
  assign _T_523 = _T_522 == 16'h0;
  assign _T_524 = _T_522[0];
  assign _T_525 = _T_522[2];
  assign _T_526 = _T_524 ^ _T_525;
  assign _T_527 = _T_522[3];
  assign _T_528 = _T_526 ^ _T_527;
  assign _T_529 = _T_522[5];
  assign _T_530 = _T_528 ^ _T_529;
  assign _T_531 = _T_522[15:1];
  assign _T_532 = {_T_530,_T_531};
  assign _T_535 = _T_534 == 16'h0;
  assign _T_536 = _T_534[0];
  assign _T_537 = _T_534[2];
  assign _T_538 = _T_536 ^ _T_537;
  assign _T_539 = _T_534[3];
  assign _T_540 = _T_538 ^ _T_539;
  assign _T_541 = _T_534[5];
  assign _T_542 = _T_540 ^ _T_541;
  assign _T_543 = _T_534[15:1];
  assign _T_544 = {_T_542,_T_543};
  assign _T_547 = _T_546 == 16'h0;
  assign _T_548 = _T_546[0];
  assign _T_549 = _T_546[2];
  assign _T_550 = _T_548 ^ _T_549;
  assign _T_551 = _T_546[3];
  assign _T_552 = _T_550 ^ _T_551;
  assign _T_553 = _T_546[5];
  assign _T_554 = _T_552 ^ _T_553;
  assign _T_555 = _T_546[15:1];
  assign _T_556 = {_T_554,_T_555};
  assign _T_559 = _T_558 == 16'h0;
  assign _T_560 = _T_558[0];
  assign _T_561 = _T_558[2];
  assign _T_562 = _T_560 ^ _T_561;
  assign _T_563 = _T_558[3];
  assign _T_564 = _T_562 ^ _T_563;
  assign _T_565 = _T_558[5];
  assign _T_566 = _T_564 ^ _T_565;
  assign _T_567 = _T_558[15:1];
  assign _T_568 = {_T_566,_T_567};
  assign _T_571 = _T_570 == 16'h0;
  assign _T_572 = _T_570[0];
  assign _T_573 = _T_570[2];
  assign _T_574 = _T_572 ^ _T_573;
  assign _T_575 = _T_570[3];
  assign _T_576 = _T_574 ^ _T_575;
  assign _T_577 = _T_570[5];
  assign _T_578 = _T_576 ^ _T_577;
  assign _T_579 = _T_570[15:1];
  assign _T_580 = {_T_578,_T_579};
  assign _T_583 = _T_582 == 16'h0;
  assign _T_584 = _T_582[0];
  assign _T_585 = _T_582[2];
  assign _T_586 = _T_584 ^ _T_585;
  assign _T_587 = _T_582[3];
  assign _T_588 = _T_586 ^ _T_587;
  assign _T_589 = _T_582[5];
  assign _T_590 = _T_588 ^ _T_589;
  assign _T_591 = _T_582[15:1];
  assign _T_592 = {_T_590,_T_591};
  assign _T_595 = _T_594 == 16'h0;
  assign _T_596 = _T_594[0];
  assign _T_597 = _T_594[2];
  assign _T_598 = _T_596 ^ _T_597;
  assign _T_599 = _T_594[3];
  assign _T_600 = _T_598 ^ _T_599;
  assign _T_601 = _T_594[5];
  assign _T_602 = _T_600 ^ _T_601;
  assign _T_603 = _T_594[15:1];
  assign _T_604 = {_T_602,_T_603};
  assign _T_607 = _T_606 == 16'h0;
  assign _T_608 = _T_606[0];
  assign _T_609 = _T_606[2];
  assign _T_610 = _T_608 ^ _T_609;
  assign _T_611 = _T_606[3];
  assign _T_612 = _T_610 ^ _T_611;
  assign _T_613 = _T_606[5];
  assign _T_614 = _T_612 ^ _T_613;
  assign _T_615 = _T_606[15:1];
  assign _T_616 = {_T_614,_T_615};
  assign _T_619 = _T_618 == 16'h0;
  assign _T_620 = _T_618[0];
  assign _T_621 = _T_618[2];
  assign _T_622 = _T_620 ^ _T_621;
  assign _T_623 = _T_618[3];
  assign _T_624 = _T_622 ^ _T_623;
  assign _T_625 = _T_618[5];
  assign _T_626 = _T_624 ^ _T_625;
  assign _T_627 = _T_618[15:1];
  assign _T_628 = {_T_626,_T_627};
  assign _T_631 = _T_630 == 16'h0;
  assign _T_632 = _T_630[0];
  assign _T_633 = _T_630[2];
  assign _T_634 = _T_632 ^ _T_633;
  assign _T_635 = _T_630[3];
  assign _T_636 = _T_634 ^ _T_635;
  assign _T_637 = _T_630[5];
  assign _T_638 = _T_636 ^ _T_637;
  assign _T_639 = _T_630[15:1];
  assign _T_640 = {_T_638,_T_639};
  assign _T_643 = _T_642 == 16'h0;
  assign _T_644 = _T_642[0];
  assign _T_645 = _T_642[2];
  assign _T_646 = _T_644 ^ _T_645;
  assign _T_647 = _T_642[3];
  assign _T_648 = _T_646 ^ _T_647;
  assign _T_649 = _T_642[5];
  assign _T_650 = _T_648 ^ _T_649;
  assign _T_651 = _T_642[15:1];
  assign _T_652 = {_T_650,_T_651};
  assign _T_655 = _T_654 == 16'h0;
  assign _T_656 = _T_654[0];
  assign _T_657 = _T_654[2];
  assign _T_658 = _T_656 ^ _T_657;
  assign _T_659 = _T_654[3];
  assign _T_660 = _T_658 ^ _T_659;
  assign _T_661 = _T_654[5];
  assign _T_662 = _T_660 ^ _T_661;
  assign _T_663 = _T_654[15:1];
  assign _T_664 = {_T_662,_T_663};
  assign _T_667 = _T_666 == 16'h0;
  assign _T_668 = _T_666[0];
  assign _T_669 = _T_666[2];
  assign _T_670 = _T_668 ^ _T_669;
  assign _T_671 = _T_666[3];
  assign _T_672 = _T_670 ^ _T_671;
  assign _T_673 = _T_666[5];
  assign _T_674 = _T_672 ^ _T_673;
  assign _T_675 = _T_666[15:1];
  assign _T_676 = {_T_674,_T_675};
  assign _T_679 = _T_678 == 16'h0;
  assign _T_680 = _T_678[0];
  assign _T_681 = _T_678[2];
  assign _T_682 = _T_680 ^ _T_681;
  assign _T_683 = _T_678[3];
  assign _T_684 = _T_682 ^ _T_683;
  assign _T_685 = _T_678[5];
  assign _T_686 = _T_684 ^ _T_685;
  assign _T_687 = _T_678[15:1];
  assign _T_688 = {_T_686,_T_687};
  assign _T_691 = _T_690 == 16'h0;
  assign _T_692 = _T_690[0];
  assign _T_693 = _T_690[2];
  assign _T_694 = _T_692 ^ _T_693;
  assign _T_695 = _T_690[3];
  assign _T_696 = _T_694 ^ _T_695;
  assign _T_697 = _T_690[5];
  assign _T_698 = _T_696 ^ _T_697;
  assign _T_699 = _T_690[15:1];
  assign _T_700 = {_T_698,_T_699};
  assign _T_703 = _T_702 == 16'h0;
  assign _T_704 = _T_702[0];
  assign _T_705 = _T_702[2];
  assign _T_706 = _T_704 ^ _T_705;
  assign _T_707 = _T_702[3];
  assign _T_708 = _T_706 ^ _T_707;
  assign _T_709 = _T_702[5];
  assign _T_710 = _T_708 ^ _T_709;
  assign _T_711 = _T_702[15:1];
  assign _T_712 = {_T_710,_T_711};
  assign _T_715 = _T_714 == 16'h0;
  assign _T_716 = _T_714[0];
  assign _T_717 = _T_714[2];
  assign _T_718 = _T_716 ^ _T_717;
  assign _T_719 = _T_714[3];
  assign _T_720 = _T_718 ^ _T_719;
  assign _T_721 = _T_714[5];
  assign _T_722 = _T_720 ^ _T_721;
  assign _T_723 = _T_714[15:1];
  assign _T_724 = {_T_722,_T_723};
  assign _T_727 = _T_726 == 16'h0;
  assign _T_728 = _T_726[0];
  assign _T_729 = _T_726[2];
  assign _T_730 = _T_728 ^ _T_729;
  assign _T_731 = _T_726[3];
  assign _T_732 = _T_730 ^ _T_731;
  assign _T_733 = _T_726[5];
  assign _T_734 = _T_732 ^ _T_733;
  assign _T_735 = _T_726[15:1];
  assign _T_736 = {_T_734,_T_735};
  assign _T_739 = _T_738 == 16'h0;
  assign _T_740 = _T_738[0];
  assign _T_741 = _T_738[2];
  assign _T_742 = _T_740 ^ _T_741;
  assign _T_743 = _T_738[3];
  assign _T_744 = _T_742 ^ _T_743;
  assign _T_745 = _T_738[5];
  assign _T_746 = _T_744 ^ _T_745;
  assign _T_747 = _T_738[15:1];
  assign _T_748 = {_T_746,_T_747};
  assign _T_751 = _T_750 == 16'h0;
  assign _T_752 = _T_750[0];
  assign _T_753 = _T_750[2];
  assign _T_754 = _T_752 ^ _T_753;
  assign _T_755 = _T_750[3];
  assign _T_756 = _T_754 ^ _T_755;
  assign _T_757 = _T_750[5];
  assign _T_758 = _T_756 ^ _T_757;
  assign _T_759 = _T_750[15:1];
  assign _T_760 = {_T_758,_T_759};
  assign _T_763 = _T_762 == 16'h0;
  assign _T_764 = _T_762[0];
  assign _T_765 = _T_762[2];
  assign _T_766 = _T_764 ^ _T_765;
  assign _T_767 = _T_762[3];
  assign _T_768 = _T_766 ^ _T_767;
  assign _T_769 = _T_762[5];
  assign _T_770 = _T_768 ^ _T_769;
  assign _T_771 = _T_762[15:1];
  assign _T_772 = {_T_770,_T_771};
  assign _T_775 = _T_774 == 16'h0;
  assign _T_776 = _T_774[0];
  assign _T_777 = _T_774[2];
  assign _T_778 = _T_776 ^ _T_777;
  assign _T_779 = _T_774[3];
  assign _T_780 = _T_778 ^ _T_779;
  assign _T_781 = _T_774[5];
  assign _T_782 = _T_780 ^ _T_781;
  assign _T_783 = _T_774[15:1];
  assign _T_784 = {_T_782,_T_783};
  assign _T_787 = _T_786 == 16'h0;
  assign _T_788 = _T_786[0];
  assign _T_789 = _T_786[2];
  assign _T_790 = _T_788 ^ _T_789;
  assign _T_791 = _T_786[3];
  assign _T_792 = _T_790 ^ _T_791;
  assign _T_793 = _T_786[5];
  assign _T_794 = _T_792 ^ _T_793;
  assign _T_795 = _T_786[15:1];
  assign _T_796 = {_T_794,_T_795};
  assign _T_799 = _T_798 == 16'h0;
  assign _T_800 = _T_798[0];
  assign _T_801 = _T_798[2];
  assign _T_802 = _T_800 ^ _T_801;
  assign _T_803 = _T_798[3];
  assign _T_804 = _T_802 ^ _T_803;
  assign _T_805 = _T_798[5];
  assign _T_806 = _T_804 ^ _T_805;
  assign _T_807 = _T_798[15:1];
  assign _T_808 = {_T_806,_T_807};
  assign _T_811 = _T_810 == 16'h0;
  assign _T_812 = _T_810[0];
  assign _T_813 = _T_810[2];
  assign _T_814 = _T_812 ^ _T_813;
  assign _T_815 = _T_810[3];
  assign _T_816 = _T_814 ^ _T_815;
  assign _T_817 = _T_810[5];
  assign _T_818 = _T_816 ^ _T_817;
  assign _T_819 = _T_810[15:1];
  assign _T_820 = {_T_818,_T_819};
  assign _T_823 = _T_822 == 16'h0;
  assign _T_824 = _T_822[0];
  assign _T_825 = _T_822[2];
  assign _T_826 = _T_824 ^ _T_825;
  assign _T_827 = _T_822[3];
  assign _T_828 = _T_826 ^ _T_827;
  assign _T_829 = _T_822[5];
  assign _T_830 = _T_828 ^ _T_829;
  assign _T_831 = _T_822[15:1];
  assign _T_832 = {_T_830,_T_831};
  assign _T_835 = _T_834 == 16'h0;
  assign _T_836 = _T_834[0];
  assign _T_837 = _T_834[2];
  assign _T_838 = _T_836 ^ _T_837;
  assign _T_839 = _T_834[3];
  assign _T_840 = _T_838 ^ _T_839;
  assign _T_841 = _T_834[5];
  assign _T_842 = _T_840 ^ _T_841;
  assign _T_843 = _T_834[15:1];
  assign _T_844 = {_T_842,_T_843};
  assign _T_847 = _T_846 == 16'h0;
  assign _T_848 = _T_846[0];
  assign _T_849 = _T_846[2];
  assign _T_850 = _T_848 ^ _T_849;
  assign _T_851 = _T_846[3];
  assign _T_852 = _T_850 ^ _T_851;
  assign _T_853 = _T_846[5];
  assign _T_854 = _T_852 ^ _T_853;
  assign _T_855 = _T_846[15:1];
  assign _T_856 = {_T_854,_T_855};
  assign _T_859 = _T_858 == 16'h0;
  assign _T_860 = _T_858[0];
  assign _T_861 = _T_858[2];
  assign _T_862 = _T_860 ^ _T_861;
  assign _T_863 = _T_858[3];
  assign _T_864 = _T_862 ^ _T_863;
  assign _T_865 = _T_858[5];
  assign _T_866 = _T_864 ^ _T_865;
  assign _T_867 = _T_858[15:1];
  assign _T_868 = {_T_866,_T_867};
  assign _T_871 = _T_870 == 16'h0;
  assign _T_872 = _T_870[0];
  assign _T_873 = _T_870[2];
  assign _T_874 = _T_872 ^ _T_873;
  assign _T_875 = _T_870[3];
  assign _T_876 = _T_874 ^ _T_875;
  assign _T_877 = _T_870[5];
  assign _T_878 = _T_876 ^ _T_877;
  assign _T_879 = _T_870[15:1];
  assign _T_880 = {_T_878,_T_879};
  assign _T_883 = _T_882 == 16'h0;
  assign _T_884 = _T_882[0];
  assign _T_885 = _T_882[2];
  assign _T_886 = _T_884 ^ _T_885;
  assign _T_887 = _T_882[3];
  assign _T_888 = _T_886 ^ _T_887;
  assign _T_889 = _T_882[5];
  assign _T_890 = _T_888 ^ _T_889;
  assign _T_891 = _T_882[15:1];
  assign _T_892 = {_T_890,_T_891};
  assign _T_895 = _T_894 == 16'h0;
  assign _T_896 = _T_894[0];
  assign _T_897 = _T_894[2];
  assign _T_898 = _T_896 ^ _T_897;
  assign _T_899 = _T_894[3];
  assign _T_900 = _T_898 ^ _T_899;
  assign _T_901 = _T_894[5];
  assign _T_902 = _T_900 ^ _T_901;
  assign _T_903 = _T_894[15:1];
  assign _T_904 = {_T_902,_T_903};
  assign _T_907 = _T_906 == 16'h0;
  assign _T_908 = _T_906[0];
  assign _T_909 = _T_906[2];
  assign _T_910 = _T_908 ^ _T_909;
  assign _T_911 = _T_906[3];
  assign _T_912 = _T_910 ^ _T_911;
  assign _T_913 = _T_906[5];
  assign _T_914 = _T_912 ^ _T_913;
  assign _T_915 = _T_906[15:1];
  assign _T_916 = {_T_914,_T_915};
  assign _T_919 = _T_918 == 16'h0;
  assign _T_920 = _T_918[0];
  assign _T_921 = _T_918[2];
  assign _T_922 = _T_920 ^ _T_921;
  assign _T_923 = _T_918[3];
  assign _T_924 = _T_922 ^ _T_923;
  assign _T_925 = _T_918[5];
  assign _T_926 = _T_924 ^ _T_925;
  assign _T_927 = _T_918[15:1];
  assign _T_928 = {_T_926,_T_927};
  assign _T_931 = _T_930 == 16'h0;
  assign _T_932 = _T_930[0];
  assign _T_933 = _T_930[2];
  assign _T_934 = _T_932 ^ _T_933;
  assign _T_935 = _T_930[3];
  assign _T_936 = _T_934 ^ _T_935;
  assign _T_937 = _T_930[5];
  assign _T_938 = _T_936 ^ _T_937;
  assign _T_939 = _T_930[15:1];
  assign _T_940 = {_T_938,_T_939};
  assign _T_943 = _T_942 == 16'h0;
  assign _T_944 = _T_942[0];
  assign _T_945 = _T_942[2];
  assign _T_946 = _T_944 ^ _T_945;
  assign _T_947 = _T_942[3];
  assign _T_948 = _T_946 ^ _T_947;
  assign _T_949 = _T_942[5];
  assign _T_950 = _T_948 ^ _T_949;
  assign _T_951 = _T_942[15:1];
  assign _T_952 = {_T_950,_T_951};
  assign _T_955 = _T_954 == 16'h0;
  assign _T_956 = _T_954[0];
  assign _T_957 = _T_954[2];
  assign _T_958 = _T_956 ^ _T_957;
  assign _T_959 = _T_954[3];
  assign _T_960 = _T_958 ^ _T_959;
  assign _T_961 = _T_954[5];
  assign _T_962 = _T_960 ^ _T_961;
  assign _T_963 = _T_954[15:1];
  assign _T_964 = {_T_962,_T_963};
  assign _T_967 = _T_966 == 16'h0;
  assign _T_968 = _T_966[0];
  assign _T_969 = _T_966[2];
  assign _T_970 = _T_968 ^ _T_969;
  assign _T_971 = _T_966[3];
  assign _T_972 = _T_970 ^ _T_971;
  assign _T_973 = _T_966[5];
  assign _T_974 = _T_972 ^ _T_973;
  assign _T_975 = _T_966[15:1];
  assign _T_976 = {_T_974,_T_975};
  assign _T_979 = _T_978 == 16'h0;
  assign _T_980 = _T_978[0];
  assign _T_981 = _T_978[2];
  assign _T_982 = _T_980 ^ _T_981;
  assign _T_983 = _T_978[3];
  assign _T_984 = _T_982 ^ _T_983;
  assign _T_985 = _T_978[5];
  assign _T_986 = _T_984 ^ _T_985;
  assign _T_987 = _T_978[15:1];
  assign _T_988 = {_T_986,_T_987};
  assign _T_991 = _T_990 == 16'h0;
  assign _T_992 = _T_990[0];
  assign _T_993 = _T_990[2];
  assign _T_994 = _T_992 ^ _T_993;
  assign _T_995 = _T_990[3];
  assign _T_996 = _T_994 ^ _T_995;
  assign _T_997 = _T_990[5];
  assign _T_998 = _T_996 ^ _T_997;
  assign _T_999 = _T_990[15:1];
  assign _T_1000 = {_T_998,_T_999};
  assign _T_1003 = _T_1002 == 16'h0;
  assign _T_1004 = _T_1002[0];
  assign _T_1005 = _T_1002[2];
  assign _T_1006 = _T_1004 ^ _T_1005;
  assign _T_1007 = _T_1002[3];
  assign _T_1008 = _T_1006 ^ _T_1007;
  assign _T_1009 = _T_1002[5];
  assign _T_1010 = _T_1008 ^ _T_1009;
  assign _T_1011 = _T_1002[15:1];
  assign _T_1012 = {_T_1010,_T_1011};
  assign _T_1015 = _T_1014 == 16'h0;
  assign _T_1016 = _T_1014[0];
  assign _T_1017 = _T_1014[2];
  assign _T_1018 = _T_1016 ^ _T_1017;
  assign _T_1019 = _T_1014[3];
  assign _T_1020 = _T_1018 ^ _T_1019;
  assign _T_1021 = _T_1014[5];
  assign _T_1022 = _T_1020 ^ _T_1021;
  assign _T_1023 = _T_1014[15:1];
  assign _T_1024 = {_T_1022,_T_1023};
  assign _T_1027 = _T_1026 == 16'h0;
  assign _T_1028 = _T_1026[0];
  assign _T_1029 = _T_1026[2];
  assign _T_1030 = _T_1028 ^ _T_1029;
  assign _T_1031 = _T_1026[3];
  assign _T_1032 = _T_1030 ^ _T_1031;
  assign _T_1033 = _T_1026[5];
  assign _T_1034 = _T_1032 ^ _T_1033;
  assign _T_1035 = _T_1026[15:1];
  assign _T_1036 = {_T_1034,_T_1035};
  assign _T_1039 = _T_1038 == 16'h0;
  assign _T_1040 = _T_1038[0];
  assign _T_1041 = _T_1038[2];
  assign _T_1042 = _T_1040 ^ _T_1041;
  assign _T_1043 = _T_1038[3];
  assign _T_1044 = _T_1042 ^ _T_1043;
  assign _T_1045 = _T_1038[5];
  assign _T_1046 = _T_1044 ^ _T_1045;
  assign _T_1047 = _T_1038[15:1];
  assign _T_1048 = {_T_1046,_T_1047};
  assign _T_1051 = _T_1050 == 16'h0;
  assign _T_1052 = _T_1050[0];
  assign _T_1053 = _T_1050[2];
  assign _T_1054 = _T_1052 ^ _T_1053;
  assign _T_1055 = _T_1050[3];
  assign _T_1056 = _T_1054 ^ _T_1055;
  assign _T_1057 = _T_1050[5];
  assign _T_1058 = _T_1056 ^ _T_1057;
  assign _T_1059 = _T_1050[15:1];
  assign _T_1060 = {_T_1058,_T_1059};
  assign _T_1063 = _T_1062 == 16'h0;
  assign _T_1064 = _T_1062[0];
  assign _T_1065 = _T_1062[2];
  assign _T_1066 = _T_1064 ^ _T_1065;
  assign _T_1067 = _T_1062[3];
  assign _T_1068 = _T_1066 ^ _T_1067;
  assign _T_1069 = _T_1062[5];
  assign _T_1070 = _T_1068 ^ _T_1069;
  assign _T_1071 = _T_1062[15:1];
  assign _T_1072 = {_T_1070,_T_1071};
  assign _T_1075 = _T_1074 == 16'h0;
  assign _T_1076 = _T_1074[0];
  assign _T_1077 = _T_1074[2];
  assign _T_1078 = _T_1076 ^ _T_1077;
  assign _T_1079 = _T_1074[3];
  assign _T_1080 = _T_1078 ^ _T_1079;
  assign _T_1081 = _T_1074[5];
  assign _T_1082 = _T_1080 ^ _T_1081;
  assign _T_1083 = _T_1074[15:1];
  assign _T_1084 = {_T_1082,_T_1083};
  assign _T_1087 = _T_1086 == 16'h0;
  assign _T_1088 = _T_1086[0];
  assign _T_1089 = _T_1086[2];
  assign _T_1090 = _T_1088 ^ _T_1089;
  assign _T_1091 = _T_1086[3];
  assign _T_1092 = _T_1090 ^ _T_1091;
  assign _T_1093 = _T_1086[5];
  assign _T_1094 = _T_1092 ^ _T_1093;
  assign _T_1095 = _T_1086[15:1];
  assign _T_1096 = {_T_1094,_T_1095};
  assign _T_1099 = _T_1098 == 16'h0;
  assign _T_1100 = _T_1098[0];
  assign _T_1101 = _T_1098[2];
  assign _T_1102 = _T_1100 ^ _T_1101;
  assign _T_1103 = _T_1098[3];
  assign _T_1104 = _T_1102 ^ _T_1103;
  assign _T_1105 = _T_1098[5];
  assign _T_1106 = _T_1104 ^ _T_1105;
  assign _T_1107 = _T_1098[15:1];
  assign _T_1108 = {_T_1106,_T_1107};
  assign _T_1111 = _T_1110 == 16'h0;
  assign _T_1112 = _T_1110[0];
  assign _T_1113 = _T_1110[2];
  assign _T_1114 = _T_1112 ^ _T_1113;
  assign _T_1115 = _T_1110[3];
  assign _T_1116 = _T_1114 ^ _T_1115;
  assign _T_1117 = _T_1110[5];
  assign _T_1118 = _T_1116 ^ _T_1117;
  assign _T_1119 = _T_1110[15:1];
  assign _T_1120 = {_T_1118,_T_1119};
  assign _T_1123 = _T_1122 == 16'h0;
  assign _T_1124 = _T_1122[0];
  assign _T_1125 = _T_1122[2];
  assign _T_1126 = _T_1124 ^ _T_1125;
  assign _T_1127 = _T_1122[3];
  assign _T_1128 = _T_1126 ^ _T_1127;
  assign _T_1129 = _T_1122[5];
  assign _T_1130 = _T_1128 ^ _T_1129;
  assign _T_1131 = _T_1122[15:1];
  assign _T_1132 = {_T_1130,_T_1131};
  assign _T_1135 = _T_1134 == 16'h0;
  assign _T_1136 = _T_1134[0];
  assign _T_1137 = _T_1134[2];
  assign _T_1138 = _T_1136 ^ _T_1137;
  assign _T_1139 = _T_1134[3];
  assign _T_1140 = _T_1138 ^ _T_1139;
  assign _T_1141 = _T_1134[5];
  assign _T_1142 = _T_1140 ^ _T_1141;
  assign _T_1143 = _T_1134[15:1];
  assign _T_1144 = {_T_1142,_T_1143};
  assign _T_1147 = _T_1146 == 16'h0;
  assign _T_1148 = _T_1146[0];
  assign _T_1149 = _T_1146[2];
  assign _T_1150 = _T_1148 ^ _T_1149;
  assign _T_1151 = _T_1146[3];
  assign _T_1152 = _T_1150 ^ _T_1151;
  assign _T_1153 = _T_1146[5];
  assign _T_1154 = _T_1152 ^ _T_1153;
  assign _T_1155 = _T_1146[15:1];
  assign _T_1156 = {_T_1154,_T_1155};
  assign _T_1159 = _T_1158 == 16'h0;
  assign _T_1160 = _T_1158[0];
  assign _T_1161 = _T_1158[2];
  assign _T_1162 = _T_1160 ^ _T_1161;
  assign _T_1163 = _T_1158[3];
  assign _T_1164 = _T_1162 ^ _T_1163;
  assign _T_1165 = _T_1158[5];
  assign _T_1166 = _T_1164 ^ _T_1165;
  assign _T_1167 = _T_1158[15:1];
  assign _T_1168 = {_T_1166,_T_1167};
  assign _T_1171 = _T_1170 == 16'h0;
  assign _T_1172 = _T_1170[0];
  assign _T_1173 = _T_1170[2];
  assign _T_1174 = _T_1172 ^ _T_1173;
  assign _T_1175 = _T_1170[3];
  assign _T_1176 = _T_1174 ^ _T_1175;
  assign _T_1177 = _T_1170[5];
  assign _T_1178 = _T_1176 ^ _T_1177;
  assign _T_1179 = _T_1170[15:1];
  assign _T_1180 = {_T_1178,_T_1179};
  assign _T_1183 = _T_1182 == 16'h0;
  assign _T_1184 = _T_1182[0];
  assign _T_1185 = _T_1182[2];
  assign _T_1186 = _T_1184 ^ _T_1185;
  assign _T_1187 = _T_1182[3];
  assign _T_1188 = _T_1186 ^ _T_1187;
  assign _T_1189 = _T_1182[5];
  assign _T_1190 = _T_1188 ^ _T_1189;
  assign _T_1191 = _T_1182[15:1];
  assign _T_1192 = {_T_1190,_T_1191};
  assign _T_1195 = _T_1194 == 16'h0;
  assign _T_1196 = _T_1194[0];
  assign _T_1197 = _T_1194[2];
  assign _T_1198 = _T_1196 ^ _T_1197;
  assign _T_1199 = _T_1194[3];
  assign _T_1200 = _T_1198 ^ _T_1199;
  assign _T_1201 = _T_1194[5];
  assign _T_1202 = _T_1200 ^ _T_1201;
  assign _T_1203 = _T_1194[15:1];
  assign _T_1204 = {_T_1202,_T_1203};
  assign _T_1207 = _T_1206 == 16'h0;
  assign _T_1208 = _T_1206[0];
  assign _T_1209 = _T_1206[2];
  assign _T_1210 = _T_1208 ^ _T_1209;
  assign _T_1211 = _T_1206[3];
  assign _T_1212 = _T_1210 ^ _T_1211;
  assign _T_1213 = _T_1206[5];
  assign _T_1214 = _T_1212 ^ _T_1213;
  assign _T_1215 = _T_1206[15:1];
  assign _T_1216 = {_T_1214,_T_1215};
  assign _T_1219 = _T_1218 == 16'h0;
  assign _T_1220 = _T_1218[0];
  assign _T_1221 = _T_1218[2];
  assign _T_1222 = _T_1220 ^ _T_1221;
  assign _T_1223 = _T_1218[3];
  assign _T_1224 = _T_1222 ^ _T_1223;
  assign _T_1225 = _T_1218[5];
  assign _T_1226 = _T_1224 ^ _T_1225;
  assign _T_1227 = _T_1218[15:1];
  assign _T_1228 = {_T_1226,_T_1227};
  assign _T_1231 = _T_1230 == 16'h0;
  assign _T_1232 = _T_1230[0];
  assign _T_1233 = _T_1230[2];
  assign _T_1234 = _T_1232 ^ _T_1233;
  assign _T_1235 = _T_1230[3];
  assign _T_1236 = _T_1234 ^ _T_1235;
  assign _T_1237 = _T_1230[5];
  assign _T_1238 = _T_1236 ^ _T_1237;
  assign _T_1239 = _T_1230[15:1];
  assign _T_1240 = {_T_1238,_T_1239};
  assign _T_1243 = _T_1242 == 16'h0;
  assign _T_1244 = _T_1242[0];
  assign _T_1245 = _T_1242[2];
  assign _T_1246 = _T_1244 ^ _T_1245;
  assign _T_1247 = _T_1242[3];
  assign _T_1248 = _T_1246 ^ _T_1247;
  assign _T_1249 = _T_1242[5];
  assign _T_1250 = _T_1248 ^ _T_1249;
  assign _T_1251 = _T_1242[15:1];
  assign _T_1252 = {_T_1250,_T_1251};
  assign _T_1255 = _T_1254 == 16'h0;
  assign _T_1256 = _T_1254[0];
  assign _T_1257 = _T_1254[2];
  assign _T_1258 = _T_1256 ^ _T_1257;
  assign _T_1259 = _T_1254[3];
  assign _T_1260 = _T_1258 ^ _T_1259;
  assign _T_1261 = _T_1254[5];
  assign _T_1262 = _T_1260 ^ _T_1261;
  assign _T_1263 = _T_1254[15:1];
  assign _T_1264 = {_T_1262,_T_1263};
  assign _T_1267 = _T_1266 == 16'h0;
  assign _T_1268 = _T_1266[0];
  assign _T_1269 = _T_1266[2];
  assign _T_1270 = _T_1268 ^ _T_1269;
  assign _T_1271 = _T_1266[3];
  assign _T_1272 = _T_1270 ^ _T_1271;
  assign _T_1273 = _T_1266[5];
  assign _T_1274 = _T_1272 ^ _T_1273;
  assign _T_1275 = _T_1266[15:1];
  assign _T_1276 = {_T_1274,_T_1275};
  assign _T_1279 = _T_1278 == 16'h0;
  assign _T_1280 = _T_1278[0];
  assign _T_1281 = _T_1278[2];
  assign _T_1282 = _T_1280 ^ _T_1281;
  assign _T_1283 = _T_1278[3];
  assign _T_1284 = _T_1282 ^ _T_1283;
  assign _T_1285 = _T_1278[5];
  assign _T_1286 = _T_1284 ^ _T_1285;
  assign _T_1287 = _T_1278[15:1];
  assign _T_1288 = {_T_1286,_T_1287};
  assign _T_1291 = _T_1290 == 16'h0;
  assign _T_1292 = _T_1290[0];
  assign _T_1293 = _T_1290[2];
  assign _T_1294 = _T_1292 ^ _T_1293;
  assign _T_1295 = _T_1290[3];
  assign _T_1296 = _T_1294 ^ _T_1295;
  assign _T_1297 = _T_1290[5];
  assign _T_1298 = _T_1296 ^ _T_1297;
  assign _T_1299 = _T_1290[15:1];
  assign _T_1300 = {_T_1298,_T_1299};
  assign _T_1303 = _T_1302 == 16'h0;
  assign _T_1304 = _T_1302[0];
  assign _T_1305 = _T_1302[2];
  assign _T_1306 = _T_1304 ^ _T_1305;
  assign _T_1307 = _T_1302[3];
  assign _T_1308 = _T_1306 ^ _T_1307;
  assign _T_1309 = _T_1302[5];
  assign _T_1310 = _T_1308 ^ _T_1309;
  assign _T_1311 = _T_1302[15:1];
  assign _T_1312 = {_T_1310,_T_1311};
  assign _T_1315 = _T_1314 == 16'h0;
  assign _T_1316 = _T_1314[0];
  assign _T_1317 = _T_1314[2];
  assign _T_1318 = _T_1316 ^ _T_1317;
  assign _T_1319 = _T_1314[3];
  assign _T_1320 = _T_1318 ^ _T_1319;
  assign _T_1321 = _T_1314[5];
  assign _T_1322 = _T_1320 ^ _T_1321;
  assign _T_1323 = _T_1314[15:1];
  assign _T_1324 = {_T_1322,_T_1323};
  assign _T_1327 = _T_1326 == 16'h0;
  assign _T_1328 = _T_1326[0];
  assign _T_1329 = _T_1326[2];
  assign _T_1330 = _T_1328 ^ _T_1329;
  assign _T_1331 = _T_1326[3];
  assign _T_1332 = _T_1330 ^ _T_1331;
  assign _T_1333 = _T_1326[5];
  assign _T_1334 = _T_1332 ^ _T_1333;
  assign _T_1335 = _T_1326[15:1];
  assign _T_1336 = {_T_1334,_T_1335};
  assign _T_1339 = _T_1338 == 16'h0;
  assign _T_1340 = _T_1338[0];
  assign _T_1341 = _T_1338[2];
  assign _T_1342 = _T_1340 ^ _T_1341;
  assign _T_1343 = _T_1338[3];
  assign _T_1344 = _T_1342 ^ _T_1343;
  assign _T_1345 = _T_1338[5];
  assign _T_1346 = _T_1344 ^ _T_1345;
  assign _T_1347 = _T_1338[15:1];
  assign _T_1348 = {_T_1346,_T_1347};
  assign _T_1351 = _T_1350 == 16'h0;
  assign _T_1352 = _T_1350[0];
  assign _T_1353 = _T_1350[2];
  assign _T_1354 = _T_1352 ^ _T_1353;
  assign _T_1355 = _T_1350[3];
  assign _T_1356 = _T_1354 ^ _T_1355;
  assign _T_1357 = _T_1350[5];
  assign _T_1358 = _T_1356 ^ _T_1357;
  assign _T_1359 = _T_1350[15:1];
  assign _T_1360 = {_T_1358,_T_1359};
  assign _T_1363 = _T_1362 == 16'h0;
  assign _T_1364 = _T_1362[0];
  assign _T_1365 = _T_1362[2];
  assign _T_1366 = _T_1364 ^ _T_1365;
  assign _T_1367 = _T_1362[3];
  assign _T_1368 = _T_1366 ^ _T_1367;
  assign _T_1369 = _T_1362[5];
  assign _T_1370 = _T_1368 ^ _T_1369;
  assign _T_1371 = _T_1362[15:1];
  assign _T_1372 = {_T_1370,_T_1371};
  assign _T_1375 = _T_1374 == 16'h0;
  assign _T_1376 = _T_1374[0];
  assign _T_1377 = _T_1374[2];
  assign _T_1378 = _T_1376 ^ _T_1377;
  assign _T_1379 = _T_1374[3];
  assign _T_1380 = _T_1378 ^ _T_1379;
  assign _T_1381 = _T_1374[5];
  assign _T_1382 = _T_1380 ^ _T_1381;
  assign _T_1383 = _T_1374[15:1];
  assign _T_1384 = {_T_1382,_T_1383};
  assign _T_1387 = _T_1386 == 16'h0;
  assign _T_1388 = _T_1386[0];
  assign _T_1389 = _T_1386[2];
  assign _T_1390 = _T_1388 ^ _T_1389;
  assign _T_1391 = _T_1386[3];
  assign _T_1392 = _T_1390 ^ _T_1391;
  assign _T_1393 = _T_1386[5];
  assign _T_1394 = _T_1392 ^ _T_1393;
  assign _T_1395 = _T_1386[15:1];
  assign _T_1396 = {_T_1394,_T_1395};
  assign _T_1399 = _T_1398 == 16'h0;
  assign _T_1400 = _T_1398[0];
  assign _T_1401 = _T_1398[2];
  assign _T_1402 = _T_1400 ^ _T_1401;
  assign _T_1403 = _T_1398[3];
  assign _T_1404 = _T_1402 ^ _T_1403;
  assign _T_1405 = _T_1398[5];
  assign _T_1406 = _T_1404 ^ _T_1405;
  assign _T_1407 = _T_1398[15:1];
  assign _T_1408 = {_T_1406,_T_1407};
  assign _T_1411 = _T_1410 == 16'h0;
  assign _T_1412 = _T_1410[0];
  assign _T_1413 = _T_1410[2];
  assign _T_1414 = _T_1412 ^ _T_1413;
  assign _T_1415 = _T_1410[3];
  assign _T_1416 = _T_1414 ^ _T_1415;
  assign _T_1417 = _T_1410[5];
  assign _T_1418 = _T_1416 ^ _T_1417;
  assign _T_1419 = _T_1410[15:1];
  assign _T_1420 = {_T_1418,_T_1419};
  assign _T_1423 = _T_1422 == 16'h0;
  assign _T_1424 = _T_1422[0];
  assign _T_1425 = _T_1422[2];
  assign _T_1426 = _T_1424 ^ _T_1425;
  assign _T_1427 = _T_1422[3];
  assign _T_1428 = _T_1426 ^ _T_1427;
  assign _T_1429 = _T_1422[5];
  assign _T_1430 = _T_1428 ^ _T_1429;
  assign _T_1431 = _T_1422[15:1];
  assign _T_1432 = {_T_1430,_T_1431};
  assign _T_1435 = _T_1434 == 16'h0;
  assign _T_1436 = _T_1434[0];
  assign _T_1437 = _T_1434[2];
  assign _T_1438 = _T_1436 ^ _T_1437;
  assign _T_1439 = _T_1434[3];
  assign _T_1440 = _T_1438 ^ _T_1439;
  assign _T_1441 = _T_1434[5];
  assign _T_1442 = _T_1440 ^ _T_1441;
  assign _T_1443 = _T_1434[15:1];
  assign _T_1444 = {_T_1442,_T_1443};
  assign _T_1447 = _T_1446 == 16'h0;
  assign _T_1448 = _T_1446[0];
  assign _T_1449 = _T_1446[2];
  assign _T_1450 = _T_1448 ^ _T_1449;
  assign _T_1451 = _T_1446[3];
  assign _T_1452 = _T_1450 ^ _T_1451;
  assign _T_1453 = _T_1446[5];
  assign _T_1454 = _T_1452 ^ _T_1453;
  assign _T_1455 = _T_1446[15:1];
  assign _T_1456 = {_T_1454,_T_1455};
  assign _T_1459 = _T_1458 == 16'h0;
  assign _T_1460 = _T_1458[0];
  assign _T_1461 = _T_1458[2];
  assign _T_1462 = _T_1460 ^ _T_1461;
  assign _T_1463 = _T_1458[3];
  assign _T_1464 = _T_1462 ^ _T_1463;
  assign _T_1465 = _T_1458[5];
  assign _T_1466 = _T_1464 ^ _T_1465;
  assign _T_1467 = _T_1458[15:1];
  assign _T_1468 = {_T_1466,_T_1467};
  assign _T_1471 = _T_1470 == 16'h0;
  assign _T_1472 = _T_1470[0];
  assign _T_1473 = _T_1470[2];
  assign _T_1474 = _T_1472 ^ _T_1473;
  assign _T_1475 = _T_1470[3];
  assign _T_1476 = _T_1474 ^ _T_1475;
  assign _T_1477 = _T_1470[5];
  assign _T_1478 = _T_1476 ^ _T_1477;
  assign _T_1479 = _T_1470[15:1];
  assign _T_1480 = {_T_1478,_T_1479};
  assign _T_1483 = _T_1482 == 16'h0;
  assign _T_1484 = _T_1482[0];
  assign _T_1485 = _T_1482[2];
  assign _T_1486 = _T_1484 ^ _T_1485;
  assign _T_1487 = _T_1482[3];
  assign _T_1488 = _T_1486 ^ _T_1487;
  assign _T_1489 = _T_1482[5];
  assign _T_1490 = _T_1488 ^ _T_1489;
  assign _T_1491 = _T_1482[15:1];
  assign _T_1492 = {_T_1490,_T_1491};
  assign _T_1495 = _T_1494 == 16'h0;
  assign _T_1496 = _T_1494[0];
  assign _T_1497 = _T_1494[2];
  assign _T_1498 = _T_1496 ^ _T_1497;
  assign _T_1499 = _T_1494[3];
  assign _T_1500 = _T_1498 ^ _T_1499;
  assign _T_1501 = _T_1494[5];
  assign _T_1502 = _T_1500 ^ _T_1501;
  assign _T_1503 = _T_1494[15:1];
  assign _T_1504 = {_T_1502,_T_1503};
  assign _T_1507 = _T_1506 == 16'h0;
  assign _T_1508 = _T_1506[0];
  assign _T_1509 = _T_1506[2];
  assign _T_1510 = _T_1508 ^ _T_1509;
  assign _T_1511 = _T_1506[3];
  assign _T_1512 = _T_1510 ^ _T_1511;
  assign _T_1513 = _T_1506[5];
  assign _T_1514 = _T_1512 ^ _T_1513;
  assign _T_1515 = _T_1506[15:1];
  assign _T_1516 = {_T_1514,_T_1515};
  assign _T_1519 = _T_1518 == 16'h0;
  assign _T_1520 = _T_1518[0];
  assign _T_1521 = _T_1518[2];
  assign _T_1522 = _T_1520 ^ _T_1521;
  assign _T_1523 = _T_1518[3];
  assign _T_1524 = _T_1522 ^ _T_1523;
  assign _T_1525 = _T_1518[5];
  assign _T_1526 = _T_1524 ^ _T_1525;
  assign _T_1527 = _T_1518[15:1];
  assign _T_1528 = {_T_1526,_T_1527};
  assign _T_1531 = _T_1530 == 16'h0;
  assign _T_1532 = _T_1530[0];
  assign _T_1533 = _T_1530[2];
  assign _T_1534 = _T_1532 ^ _T_1533;
  assign _T_1535 = _T_1530[3];
  assign _T_1536 = _T_1534 ^ _T_1535;
  assign _T_1537 = _T_1530[5];
  assign _T_1538 = _T_1536 ^ _T_1537;
  assign _T_1539 = _T_1530[15:1];
  assign _T_1540 = {_T_1538,_T_1539};
  assign _T_1543 = _T_1542 == 16'h0;
  assign _T_1544 = _T_1542[0];
  assign _T_1545 = _T_1542[2];
  assign _T_1546 = _T_1544 ^ _T_1545;
  assign _T_1547 = _T_1542[3];
  assign _T_1548 = _T_1546 ^ _T_1547;
  assign _T_1549 = _T_1542[5];
  assign _T_1550 = _T_1548 ^ _T_1549;
  assign _T_1551 = _T_1542[15:1];
  assign _T_1552 = {_T_1550,_T_1551};
  assign _T_1555 = _T_1554 == 16'h0;
  assign _T_1556 = _T_1554[0];
  assign _T_1557 = _T_1554[2];
  assign _T_1558 = _T_1556 ^ _T_1557;
  assign _T_1559 = _T_1554[3];
  assign _T_1560 = _T_1558 ^ _T_1559;
  assign _T_1561 = _T_1554[5];
  assign _T_1562 = _T_1560 ^ _T_1561;
  assign _T_1563 = _T_1554[15:1];
  assign _T_1564 = {_T_1562,_T_1563};
  assign _T_1567 = _T_1566 == 16'h0;
  assign _T_1568 = _T_1566[0];
  assign _T_1569 = _T_1566[2];
  assign _T_1570 = _T_1568 ^ _T_1569;
  assign _T_1571 = _T_1566[3];
  assign _T_1572 = _T_1570 ^ _T_1571;
  assign _T_1573 = _T_1566[5];
  assign _T_1574 = _T_1572 ^ _T_1573;
  assign _T_1575 = _T_1566[15:1];
  assign _T_1576 = {_T_1574,_T_1575};
  assign _T_1579 = _T_1578 == 16'h0;
  assign _T_1580 = _T_1578[0];
  assign _T_1581 = _T_1578[2];
  assign _T_1582 = _T_1580 ^ _T_1581;
  assign _T_1583 = _T_1578[3];
  assign _T_1584 = _T_1582 ^ _T_1583;
  assign _T_1585 = _T_1578[5];
  assign _T_1586 = _T_1584 ^ _T_1585;
  assign _T_1587 = _T_1578[15:1];
  assign _T_1588 = {_T_1586,_T_1587};
  assign _T_1591 = _T_1590 == 16'h0;
  assign _T_1592 = _T_1590[0];
  assign _T_1593 = _T_1590[2];
  assign _T_1594 = _T_1592 ^ _T_1593;
  assign _T_1595 = _T_1590[3];
  assign _T_1596 = _T_1594 ^ _T_1595;
  assign _T_1597 = _T_1590[5];
  assign _T_1598 = _T_1596 ^ _T_1597;
  assign _T_1599 = _T_1590[15:1];
  assign _T_1600 = {_T_1598,_T_1599};
  assign _T_1603 = _T_1602 == 16'h0;
  assign _T_1604 = _T_1602[0];
  assign _T_1605 = _T_1602[2];
  assign _T_1606 = _T_1604 ^ _T_1605;
  assign _T_1607 = _T_1602[3];
  assign _T_1608 = _T_1606 ^ _T_1607;
  assign _T_1609 = _T_1602[5];
  assign _T_1610 = _T_1608 ^ _T_1609;
  assign _T_1611 = _T_1602[15:1];
  assign _T_1612 = {_T_1610,_T_1611};
  assign _T_1615 = _T_1614 == 16'h0;
  assign _T_1616 = _T_1614[0];
  assign _T_1617 = _T_1614[2];
  assign _T_1618 = _T_1616 ^ _T_1617;
  assign _T_1619 = _T_1614[3];
  assign _T_1620 = _T_1618 ^ _T_1619;
  assign _T_1621 = _T_1614[5];
  assign _T_1622 = _T_1620 ^ _T_1621;
  assign _T_1623 = _T_1614[15:1];
  assign _T_1624 = {_T_1622,_T_1623};
  assign _T_1627 = _T_1626 == 16'h0;
  assign _T_1628 = _T_1626[0];
  assign _T_1629 = _T_1626[2];
  assign _T_1630 = _T_1628 ^ _T_1629;
  assign _T_1631 = _T_1626[3];
  assign _T_1632 = _T_1630 ^ _T_1631;
  assign _T_1633 = _T_1626[5];
  assign _T_1634 = _T_1632 ^ _T_1633;
  assign _T_1635 = _T_1626[15:1];
  assign _T_1636 = {_T_1634,_T_1635};
  assign _T_1639 = _T_1638 == 16'h0;
  assign _T_1640 = _T_1638[0];
  assign _T_1641 = _T_1638[2];
  assign _T_1642 = _T_1640 ^ _T_1641;
  assign _T_1643 = _T_1638[3];
  assign _T_1644 = _T_1642 ^ _T_1643;
  assign _T_1645 = _T_1638[5];
  assign _T_1646 = _T_1644 ^ _T_1645;
  assign _T_1647 = _T_1638[15:1];
  assign _T_1648 = {_T_1646,_T_1647};
  assign _T_1651 = _T_1650 == 16'h0;
  assign _T_1652 = _T_1650[0];
  assign _T_1653 = _T_1650[2];
  assign _T_1654 = _T_1652 ^ _T_1653;
  assign _T_1655 = _T_1650[3];
  assign _T_1656 = _T_1654 ^ _T_1655;
  assign _T_1657 = _T_1650[5];
  assign _T_1658 = _T_1656 ^ _T_1657;
  assign _T_1659 = _T_1650[15:1];
  assign _T_1660 = {_T_1658,_T_1659};
  assign _T_1663 = _T_1662 == 16'h0;
  assign _T_1664 = _T_1662[0];
  assign _T_1665 = _T_1662[2];
  assign _T_1666 = _T_1664 ^ _T_1665;
  assign _T_1667 = _T_1662[3];
  assign _T_1668 = _T_1666 ^ _T_1667;
  assign _T_1669 = _T_1662[5];
  assign _T_1670 = _T_1668 ^ _T_1669;
  assign _T_1671 = _T_1662[15:1];
  assign _T_1672 = {_T_1670,_T_1671};
  assign _T_1675 = _T_1674 == 16'h0;
  assign _T_1676 = _T_1674[0];
  assign _T_1677 = _T_1674[2];
  assign _T_1678 = _T_1676 ^ _T_1677;
  assign _T_1679 = _T_1674[3];
  assign _T_1680 = _T_1678 ^ _T_1679;
  assign _T_1681 = _T_1674[5];
  assign _T_1682 = _T_1680 ^ _T_1681;
  assign _T_1683 = _T_1674[15:1];
  assign _T_1684 = {_T_1682,_T_1683};
  assign _T_1687 = _T_1686 == 16'h0;
  assign _T_1688 = _T_1686[0];
  assign _T_1689 = _T_1686[2];
  assign _T_1690 = _T_1688 ^ _T_1689;
  assign _T_1691 = _T_1686[3];
  assign _T_1692 = _T_1690 ^ _T_1691;
  assign _T_1693 = _T_1686[5];
  assign _T_1694 = _T_1692 ^ _T_1693;
  assign _T_1695 = _T_1686[15:1];
  assign _T_1696 = {_T_1694,_T_1695};
  assign _T_1699 = _T_1698 == 16'h0;
  assign _T_1700 = _T_1698[0];
  assign _T_1701 = _T_1698[2];
  assign _T_1702 = _T_1700 ^ _T_1701;
  assign _T_1703 = _T_1698[3];
  assign _T_1704 = _T_1702 ^ _T_1703;
  assign _T_1705 = _T_1698[5];
  assign _T_1706 = _T_1704 ^ _T_1705;
  assign _T_1707 = _T_1698[15:1];
  assign _T_1708 = {_T_1706,_T_1707};
  assign _T_1713 = _T_1712 == 16'h0;
  assign _T_1714 = _T_1712[0];
  assign _T_1715 = _T_1712[2];
  assign _T_1716 = _T_1714 ^ _T_1715;
  assign _T_1717 = _T_1712[3];
  assign _T_1718 = _T_1716 ^ _T_1717;
  assign _T_1719 = _T_1712[5];
  assign _T_1720 = _T_1718 ^ _T_1719;
  assign _T_1721 = _T_1712[15:1];
  assign _T_1722 = {_T_1720,_T_1721};
  assign _T_1725 = _T_1724 == 16'h0;
  assign _T_1726 = _T_1724[0];
  assign _T_1727 = _T_1724[2];
  assign _T_1728 = _T_1726 ^ _T_1727;
  assign _T_1729 = _T_1724[3];
  assign _T_1730 = _T_1728 ^ _T_1729;
  assign _T_1731 = _T_1724[5];
  assign _T_1732 = _T_1730 ^ _T_1731;
  assign _T_1733 = _T_1724[15:1];
  assign _T_1734 = {_T_1732,_T_1733};
  assign _T_1737 = _T_1736 == 16'h0;
  assign _T_1738 = _T_1736[0];
  assign _T_1739 = _T_1736[2];
  assign _T_1740 = _T_1738 ^ _T_1739;
  assign _T_1741 = _T_1736[3];
  assign _T_1742 = _T_1740 ^ _T_1741;
  assign _T_1743 = _T_1736[5];
  assign _T_1744 = _T_1742 ^ _T_1743;
  assign _T_1745 = _T_1736[15:1];
  assign _T_1746 = {_T_1744,_T_1745};
  assign _T_1749 = _T_1748 == 16'h0;
  assign _T_1750 = _T_1748[0];
  assign _T_1751 = _T_1748[2];
  assign _T_1752 = _T_1750 ^ _T_1751;
  assign _T_1753 = _T_1748[3];
  assign _T_1754 = _T_1752 ^ _T_1753;
  assign _T_1755 = _T_1748[5];
  assign _T_1756 = _T_1754 ^ _T_1755;
  assign _T_1757 = _T_1748[15:1];
  assign _T_1758 = {_T_1756,_T_1757};
  assign _T_1761 = _T_1760 == 16'h0;
  assign _T_1762 = _T_1760[0];
  assign _T_1763 = _T_1760[2];
  assign _T_1764 = _T_1762 ^ _T_1763;
  assign _T_1765 = _T_1760[3];
  assign _T_1766 = _T_1764 ^ _T_1765;
  assign _T_1767 = _T_1760[5];
  assign _T_1768 = _T_1766 ^ _T_1767;
  assign _T_1769 = _T_1760[15:1];
  assign _T_1770 = {_T_1768,_T_1769};
  assign _T_1773 = _T_1772 == 16'h0;
  assign _T_1774 = _T_1772[0];
  assign _T_1775 = _T_1772[2];
  assign _T_1776 = _T_1774 ^ _T_1775;
  assign _T_1777 = _T_1772[3];
  assign _T_1778 = _T_1776 ^ _T_1777;
  assign _T_1779 = _T_1772[5];
  assign _T_1780 = _T_1778 ^ _T_1779;
  assign _T_1781 = _T_1772[15:1];
  assign _T_1782 = {_T_1780,_T_1781};
  assign _T_1785 = _T_1784 == 16'h0;
  assign _T_1786 = _T_1784[0];
  assign _T_1787 = _T_1784[2];
  assign _T_1788 = _T_1786 ^ _T_1787;
  assign _T_1789 = _T_1784[3];
  assign _T_1790 = _T_1788 ^ _T_1789;
  assign _T_1791 = _T_1784[5];
  assign _T_1792 = _T_1790 ^ _T_1791;
  assign _T_1793 = _T_1784[15:1];
  assign _T_1794 = {_T_1792,_T_1793};
  assign _T_1797 = _T_1796 == 16'h0;
  assign _T_1798 = _T_1796[0];
  assign _T_1799 = _T_1796[2];
  assign _T_1800 = _T_1798 ^ _T_1799;
  assign _T_1801 = _T_1796[3];
  assign _T_1802 = _T_1800 ^ _T_1801;
  assign _T_1803 = _T_1796[5];
  assign _T_1804 = _T_1802 ^ _T_1803;
  assign _T_1805 = _T_1796[15:1];
  assign _T_1806 = {_T_1804,_T_1805};
  assign _T_1809 = _T_1808 == 16'h0;
  assign _T_1810 = _T_1808[0];
  assign _T_1811 = _T_1808[2];
  assign _T_1812 = _T_1810 ^ _T_1811;
  assign _T_1813 = _T_1808[3];
  assign _T_1814 = _T_1812 ^ _T_1813;
  assign _T_1815 = _T_1808[5];
  assign _T_1816 = _T_1814 ^ _T_1815;
  assign _T_1817 = _T_1808[15:1];
  assign _T_1818 = {_T_1816,_T_1817};
  assign _T_1821 = _T_1820 == 16'h0;
  assign _T_1822 = _T_1820[0];
  assign _T_1823 = _T_1820[2];
  assign _T_1824 = _T_1822 ^ _T_1823;
  assign _T_1825 = _T_1820[3];
  assign _T_1826 = _T_1824 ^ _T_1825;
  assign _T_1827 = _T_1820[5];
  assign _T_1828 = _T_1826 ^ _T_1827;
  assign _T_1829 = _T_1820[15:1];
  assign _T_1830 = {_T_1828,_T_1829};
  assign _T_1833 = _T_1832 == 16'h0;
  assign _T_1834 = _T_1832[0];
  assign _T_1835 = _T_1832[2];
  assign _T_1836 = _T_1834 ^ _T_1835;
  assign _T_1837 = _T_1832[3];
  assign _T_1838 = _T_1836 ^ _T_1837;
  assign _T_1839 = _T_1832[5];
  assign _T_1840 = _T_1838 ^ _T_1839;
  assign _T_1841 = _T_1832[15:1];
  assign _T_1842 = {_T_1840,_T_1841};
  assign _T_1845 = _T_1844 == 16'h0;
  assign _T_1846 = _T_1844[0];
  assign _T_1847 = _T_1844[2];
  assign _T_1848 = _T_1846 ^ _T_1847;
  assign _T_1849 = _T_1844[3];
  assign _T_1850 = _T_1848 ^ _T_1849;
  assign _T_1851 = _T_1844[5];
  assign _T_1852 = _T_1850 ^ _T_1851;
  assign _T_1853 = _T_1844[15:1];
  assign _T_1854 = {_T_1852,_T_1853};
  assign _T_1857 = _T_1856 == 16'h0;
  assign _T_1858 = _T_1856[0];
  assign _T_1859 = _T_1856[2];
  assign _T_1860 = _T_1858 ^ _T_1859;
  assign _T_1861 = _T_1856[3];
  assign _T_1862 = _T_1860 ^ _T_1861;
  assign _T_1863 = _T_1856[5];
  assign _T_1864 = _T_1862 ^ _T_1863;
  assign _T_1865 = _T_1856[15:1];
  assign _T_1866 = {_T_1864,_T_1865};
  assign _T_1869 = _T_1868 == 16'h0;
  assign _T_1870 = _T_1868[0];
  assign _T_1871 = _T_1868[2];
  assign _T_1872 = _T_1870 ^ _T_1871;
  assign _T_1873 = _T_1868[3];
  assign _T_1874 = _T_1872 ^ _T_1873;
  assign _T_1875 = _T_1868[5];
  assign _T_1876 = _T_1874 ^ _T_1875;
  assign _T_1877 = _T_1868[15:1];
  assign _T_1878 = {_T_1876,_T_1877};
  assign _T_1881 = _T_1880 == 16'h0;
  assign _T_1882 = _T_1880[0];
  assign _T_1883 = _T_1880[2];
  assign _T_1884 = _T_1882 ^ _T_1883;
  assign _T_1885 = _T_1880[3];
  assign _T_1886 = _T_1884 ^ _T_1885;
  assign _T_1887 = _T_1880[5];
  assign _T_1888 = _T_1886 ^ _T_1887;
  assign _T_1889 = _T_1880[15:1];
  assign _T_1890 = {_T_1888,_T_1889};
  assign _T_1893 = _T_1892 == 16'h0;
  assign _T_1894 = _T_1892[0];
  assign _T_1895 = _T_1892[2];
  assign _T_1896 = _T_1894 ^ _T_1895;
  assign _T_1897 = _T_1892[3];
  assign _T_1898 = _T_1896 ^ _T_1897;
  assign _T_1899 = _T_1892[5];
  assign _T_1900 = _T_1898 ^ _T_1899;
  assign _T_1901 = _T_1892[15:1];
  assign _T_1902 = {_T_1900,_T_1901};
  assign _T_1905 = _T_1904 == 16'h0;
  assign _T_1906 = _T_1904[0];
  assign _T_1907 = _T_1904[2];
  assign _T_1908 = _T_1906 ^ _T_1907;
  assign _T_1909 = _T_1904[3];
  assign _T_1910 = _T_1908 ^ _T_1909;
  assign _T_1911 = _T_1904[5];
  assign _T_1912 = _T_1910 ^ _T_1911;
  assign _T_1913 = _T_1904[15:1];
  assign _T_1914 = {_T_1912,_T_1913};
  assign _T_1917 = _T_1916 == 16'h0;
  assign _T_1918 = _T_1916[0];
  assign _T_1919 = _T_1916[2];
  assign _T_1920 = _T_1918 ^ _T_1919;
  assign _T_1921 = _T_1916[3];
  assign _T_1922 = _T_1920 ^ _T_1921;
  assign _T_1923 = _T_1916[5];
  assign _T_1924 = _T_1922 ^ _T_1923;
  assign _T_1925 = _T_1916[15:1];
  assign _T_1926 = {_T_1924,_T_1925};
  assign _T_1929 = _T_1928 == 16'h0;
  assign _T_1930 = _T_1928[0];
  assign _T_1931 = _T_1928[2];
  assign _T_1932 = _T_1930 ^ _T_1931;
  assign _T_1933 = _T_1928[3];
  assign _T_1934 = _T_1932 ^ _T_1933;
  assign _T_1935 = _T_1928[5];
  assign _T_1936 = _T_1934 ^ _T_1935;
  assign _T_1937 = _T_1928[15:1];
  assign _T_1938 = {_T_1936,_T_1937};
  assign _T_1941 = _T_1940 == 16'h0;
  assign _T_1942 = _T_1940[0];
  assign _T_1943 = _T_1940[2];
  assign _T_1944 = _T_1942 ^ _T_1943;
  assign _T_1945 = _T_1940[3];
  assign _T_1946 = _T_1944 ^ _T_1945;
  assign _T_1947 = _T_1940[5];
  assign _T_1948 = _T_1946 ^ _T_1947;
  assign _T_1949 = _T_1940[15:1];
  assign _T_1950 = {_T_1948,_T_1949};
  assign _T_1953 = _T_1952 == 16'h0;
  assign _T_1954 = _T_1952[0];
  assign _T_1955 = _T_1952[2];
  assign _T_1956 = _T_1954 ^ _T_1955;
  assign _T_1957 = _T_1952[3];
  assign _T_1958 = _T_1956 ^ _T_1957;
  assign _T_1959 = _T_1952[5];
  assign _T_1960 = _T_1958 ^ _T_1959;
  assign _T_1961 = _T_1952[15:1];
  assign _T_1962 = {_T_1960,_T_1961};
  assign _T_1965 = _T_1964 == 16'h0;
  assign _T_1966 = _T_1964[0];
  assign _T_1967 = _T_1964[2];
  assign _T_1968 = _T_1966 ^ _T_1967;
  assign _T_1969 = _T_1964[3];
  assign _T_1970 = _T_1968 ^ _T_1969;
  assign _T_1971 = _T_1964[5];
  assign _T_1972 = _T_1970 ^ _T_1971;
  assign _T_1973 = _T_1964[15:1];
  assign _T_1974 = {_T_1972,_T_1973};
  assign _T_1977 = _T_1976 == 16'h0;
  assign _T_1978 = _T_1976[0];
  assign _T_1979 = _T_1976[2];
  assign _T_1980 = _T_1978 ^ _T_1979;
  assign _T_1981 = _T_1976[3];
  assign _T_1982 = _T_1980 ^ _T_1981;
  assign _T_1983 = _T_1976[5];
  assign _T_1984 = _T_1982 ^ _T_1983;
  assign _T_1985 = _T_1976[15:1];
  assign _T_1986 = {_T_1984,_T_1985};
  assign _T_1989 = _T_1988 == 16'h0;
  assign _T_1990 = _T_1988[0];
  assign _T_1991 = _T_1988[2];
  assign _T_1992 = _T_1990 ^ _T_1991;
  assign _T_1993 = _T_1988[3];
  assign _T_1994 = _T_1992 ^ _T_1993;
  assign _T_1995 = _T_1988[5];
  assign _T_1996 = _T_1994 ^ _T_1995;
  assign _T_1997 = _T_1988[15:1];
  assign _T_1998 = {_T_1996,_T_1997};
  assign _T_2001 = _T_2000 == 16'h0;
  assign _T_2002 = _T_2000[0];
  assign _T_2003 = _T_2000[2];
  assign _T_2004 = _T_2002 ^ _T_2003;
  assign _T_2005 = _T_2000[3];
  assign _T_2006 = _T_2004 ^ _T_2005;
  assign _T_2007 = _T_2000[5];
  assign _T_2008 = _T_2006 ^ _T_2007;
  assign _T_2009 = _T_2000[15:1];
  assign _T_2010 = {_T_2008,_T_2009};
  assign _T_2013 = _T_2012 == 16'h0;
  assign _T_2014 = _T_2012[0];
  assign _T_2015 = _T_2012[2];
  assign _T_2016 = _T_2014 ^ _T_2015;
  assign _T_2017 = _T_2012[3];
  assign _T_2018 = _T_2016 ^ _T_2017;
  assign _T_2019 = _T_2012[5];
  assign _T_2020 = _T_2018 ^ _T_2019;
  assign _T_2021 = _T_2012[15:1];
  assign _T_2022 = {_T_2020,_T_2021};
  assign _T_2025 = _T_2024 == 16'h0;
  assign _T_2026 = _T_2024[0];
  assign _T_2027 = _T_2024[2];
  assign _T_2028 = _T_2026 ^ _T_2027;
  assign _T_2029 = _T_2024[3];
  assign _T_2030 = _T_2028 ^ _T_2029;
  assign _T_2031 = _T_2024[5];
  assign _T_2032 = _T_2030 ^ _T_2031;
  assign _T_2033 = _T_2024[15:1];
  assign _T_2034 = {_T_2032,_T_2033};
  assign _T_2037 = _T_2036 == 16'h0;
  assign _T_2038 = _T_2036[0];
  assign _T_2039 = _T_2036[2];
  assign _T_2040 = _T_2038 ^ _T_2039;
  assign _T_2041 = _T_2036[3];
  assign _T_2042 = _T_2040 ^ _T_2041;
  assign _T_2043 = _T_2036[5];
  assign _T_2044 = _T_2042 ^ _T_2043;
  assign _T_2045 = _T_2036[15:1];
  assign _T_2046 = {_T_2044,_T_2045};
  assign _T_2049 = _T_2048 == 16'h0;
  assign _T_2050 = _T_2048[0];
  assign _T_2051 = _T_2048[2];
  assign _T_2052 = _T_2050 ^ _T_2051;
  assign _T_2053 = _T_2048[3];
  assign _T_2054 = _T_2052 ^ _T_2053;
  assign _T_2055 = _T_2048[5];
  assign _T_2056 = _T_2054 ^ _T_2055;
  assign _T_2057 = _T_2048[15:1];
  assign _T_2058 = {_T_2056,_T_2057};
  assign _T_2061 = _T_2060 == 16'h0;
  assign _T_2062 = _T_2060[0];
  assign _T_2063 = _T_2060[2];
  assign _T_2064 = _T_2062 ^ _T_2063;
  assign _T_2065 = _T_2060[3];
  assign _T_2066 = _T_2064 ^ _T_2065;
  assign _T_2067 = _T_2060[5];
  assign _T_2068 = _T_2066 ^ _T_2067;
  assign _T_2069 = _T_2060[15:1];
  assign _T_2070 = {_T_2068,_T_2069};
  assign _T_2073 = _T_2072 == 16'h0;
  assign _T_2074 = _T_2072[0];
  assign _T_2075 = _T_2072[2];
  assign _T_2076 = _T_2074 ^ _T_2075;
  assign _T_2077 = _T_2072[3];
  assign _T_2078 = _T_2076 ^ _T_2077;
  assign _T_2079 = _T_2072[5];
  assign _T_2080 = _T_2078 ^ _T_2079;
  assign _T_2081 = _T_2072[15:1];
  assign _T_2082 = {_T_2080,_T_2081};
  assign _T_2085 = _T_2084 == 16'h0;
  assign _T_2086 = _T_2084[0];
  assign _T_2087 = _T_2084[2];
  assign _T_2088 = _T_2086 ^ _T_2087;
  assign _T_2089 = _T_2084[3];
  assign _T_2090 = _T_2088 ^ _T_2089;
  assign _T_2091 = _T_2084[5];
  assign _T_2092 = _T_2090 ^ _T_2091;
  assign _T_2093 = _T_2084[15:1];
  assign _T_2094 = {_T_2092,_T_2093};
  assign _T_2097 = _T_2096 == 16'h0;
  assign _T_2098 = _T_2096[0];
  assign _T_2099 = _T_2096[2];
  assign _T_2100 = _T_2098 ^ _T_2099;
  assign _T_2101 = _T_2096[3];
  assign _T_2102 = _T_2100 ^ _T_2101;
  assign _T_2103 = _T_2096[5];
  assign _T_2104 = _T_2102 ^ _T_2103;
  assign _T_2105 = _T_2096[15:1];
  assign _T_2106 = {_T_2104,_T_2105};
  assign _T_2109 = _T_2108 == 16'h0;
  assign _T_2110 = _T_2108[0];
  assign _T_2111 = _T_2108[2];
  assign _T_2112 = _T_2110 ^ _T_2111;
  assign _T_2113 = _T_2108[3];
  assign _T_2114 = _T_2112 ^ _T_2113;
  assign _T_2115 = _T_2108[5];
  assign _T_2116 = _T_2114 ^ _T_2115;
  assign _T_2117 = _T_2108[15:1];
  assign _T_2118 = {_T_2116,_T_2117};
  assign _T_2121 = _T_2120 == 16'h0;
  assign _T_2122 = _T_2120[0];
  assign _T_2123 = _T_2120[2];
  assign _T_2124 = _T_2122 ^ _T_2123;
  assign _T_2125 = _T_2120[3];
  assign _T_2126 = _T_2124 ^ _T_2125;
  assign _T_2127 = _T_2120[5];
  assign _T_2128 = _T_2126 ^ _T_2127;
  assign _T_2129 = _T_2120[15:1];
  assign _T_2130 = {_T_2128,_T_2129};
  assign _T_2133 = _T_2132 == 16'h0;
  assign _T_2134 = _T_2132[0];
  assign _T_2135 = _T_2132[2];
  assign _T_2136 = _T_2134 ^ _T_2135;
  assign _T_2137 = _T_2132[3];
  assign _T_2138 = _T_2136 ^ _T_2137;
  assign _T_2139 = _T_2132[5];
  assign _T_2140 = _T_2138 ^ _T_2139;
  assign _T_2141 = _T_2132[15:1];
  assign _T_2142 = {_T_2140,_T_2141};
  assign _T_2145 = _T_2144 == 16'h0;
  assign _T_2146 = _T_2144[0];
  assign _T_2147 = _T_2144[2];
  assign _T_2148 = _T_2146 ^ _T_2147;
  assign _T_2149 = _T_2144[3];
  assign _T_2150 = _T_2148 ^ _T_2149;
  assign _T_2151 = _T_2144[5];
  assign _T_2152 = _T_2150 ^ _T_2151;
  assign _T_2153 = _T_2144[15:1];
  assign _T_2154 = {_T_2152,_T_2153};
  assign _T_2157 = _T_2156 == 16'h0;
  assign _T_2158 = _T_2156[0];
  assign _T_2159 = _T_2156[2];
  assign _T_2160 = _T_2158 ^ _T_2159;
  assign _T_2161 = _T_2156[3];
  assign _T_2162 = _T_2160 ^ _T_2161;
  assign _T_2163 = _T_2156[5];
  assign _T_2164 = _T_2162 ^ _T_2163;
  assign _T_2165 = _T_2156[15:1];
  assign _T_2166 = {_T_2164,_T_2165};
  assign _T_2169 = _T_2168 == 16'h0;
  assign _T_2170 = _T_2168[0];
  assign _T_2171 = _T_2168[2];
  assign _T_2172 = _T_2170 ^ _T_2171;
  assign _T_2173 = _T_2168[3];
  assign _T_2174 = _T_2172 ^ _T_2173;
  assign _T_2175 = _T_2168[5];
  assign _T_2176 = _T_2174 ^ _T_2175;
  assign _T_2177 = _T_2168[15:1];
  assign _T_2178 = {_T_2176,_T_2177};
  assign _T_2181 = _T_2180 == 16'h0;
  assign _T_2182 = _T_2180[0];
  assign _T_2183 = _T_2180[2];
  assign _T_2184 = _T_2182 ^ _T_2183;
  assign _T_2185 = _T_2180[3];
  assign _T_2186 = _T_2184 ^ _T_2185;
  assign _T_2187 = _T_2180[5];
  assign _T_2188 = _T_2186 ^ _T_2187;
  assign _T_2189 = _T_2180[15:1];
  assign _T_2190 = {_T_2188,_T_2189};
  assign _T_2193 = _T_2192 == 16'h0;
  assign _T_2194 = _T_2192[0];
  assign _T_2195 = _T_2192[2];
  assign _T_2196 = _T_2194 ^ _T_2195;
  assign _T_2197 = _T_2192[3];
  assign _T_2198 = _T_2196 ^ _T_2197;
  assign _T_2199 = _T_2192[5];
  assign _T_2200 = _T_2198 ^ _T_2199;
  assign _T_2201 = _T_2192[15:1];
  assign _T_2202 = {_T_2200,_T_2201};
  assign _T_2205 = _T_2204 == 16'h0;
  assign _T_2206 = _T_2204[0];
  assign _T_2207 = _T_2204[2];
  assign _T_2208 = _T_2206 ^ _T_2207;
  assign _T_2209 = _T_2204[3];
  assign _T_2210 = _T_2208 ^ _T_2209;
  assign _T_2211 = _T_2204[5];
  assign _T_2212 = _T_2210 ^ _T_2211;
  assign _T_2213 = _T_2204[15:1];
  assign _T_2214 = {_T_2212,_T_2213};
  assign _T_2217 = _T_2216 == 16'h0;
  assign _T_2218 = _T_2216[0];
  assign _T_2219 = _T_2216[2];
  assign _T_2220 = _T_2218 ^ _T_2219;
  assign _T_2221 = _T_2216[3];
  assign _T_2222 = _T_2220 ^ _T_2221;
  assign _T_2223 = _T_2216[5];
  assign _T_2224 = _T_2222 ^ _T_2223;
  assign _T_2225 = _T_2216[15:1];
  assign _T_2226 = {_T_2224,_T_2225};
  assign _T_2229 = _T_2228 == 16'h0;
  assign _T_2230 = _T_2228[0];
  assign _T_2231 = _T_2228[2];
  assign _T_2232 = _T_2230 ^ _T_2231;
  assign _T_2233 = _T_2228[3];
  assign _T_2234 = _T_2232 ^ _T_2233;
  assign _T_2235 = _T_2228[5];
  assign _T_2236 = _T_2234 ^ _T_2235;
  assign _T_2237 = _T_2228[15:1];
  assign _T_2238 = {_T_2236,_T_2237};
  assign _T_2241 = _T_2240 == 16'h0;
  assign _T_2242 = _T_2240[0];
  assign _T_2243 = _T_2240[2];
  assign _T_2244 = _T_2242 ^ _T_2243;
  assign _T_2245 = _T_2240[3];
  assign _T_2246 = _T_2244 ^ _T_2245;
  assign _T_2247 = _T_2240[5];
  assign _T_2248 = _T_2246 ^ _T_2247;
  assign _T_2249 = _T_2240[15:1];
  assign _T_2250 = {_T_2248,_T_2249};
  assign _T_2253 = _T_2252 == 16'h0;
  assign _T_2254 = _T_2252[0];
  assign _T_2255 = _T_2252[2];
  assign _T_2256 = _T_2254 ^ _T_2255;
  assign _T_2257 = _T_2252[3];
  assign _T_2258 = _T_2256 ^ _T_2257;
  assign _T_2259 = _T_2252[5];
  assign _T_2260 = _T_2258 ^ _T_2259;
  assign _T_2261 = _T_2252[15:1];
  assign _T_2262 = {_T_2260,_T_2261};
  assign _T_2265 = _T_2264 == 16'h0;
  assign _T_2266 = _T_2264[0];
  assign _T_2267 = _T_2264[2];
  assign _T_2268 = _T_2266 ^ _T_2267;
  assign _T_2269 = _T_2264[3];
  assign _T_2270 = _T_2268 ^ _T_2269;
  assign _T_2271 = _T_2264[5];
  assign _T_2272 = _T_2270 ^ _T_2271;
  assign _T_2273 = _T_2264[15:1];
  assign _T_2274 = {_T_2272,_T_2273};
  assign _T_2277 = _T_2276 == 16'h0;
  assign _T_2278 = _T_2276[0];
  assign _T_2279 = _T_2276[2];
  assign _T_2280 = _T_2278 ^ _T_2279;
  assign _T_2281 = _T_2276[3];
  assign _T_2282 = _T_2280 ^ _T_2281;
  assign _T_2283 = _T_2276[5];
  assign _T_2284 = _T_2282 ^ _T_2283;
  assign _T_2285 = _T_2276[15:1];
  assign _T_2286 = {_T_2284,_T_2285};
  assign _T_2289 = _T_2288 == 16'h0;
  assign _T_2290 = _T_2288[0];
  assign _T_2291 = _T_2288[2];
  assign _T_2292 = _T_2290 ^ _T_2291;
  assign _T_2293 = _T_2288[3];
  assign _T_2294 = _T_2292 ^ _T_2293;
  assign _T_2295 = _T_2288[5];
  assign _T_2296 = _T_2294 ^ _T_2295;
  assign _T_2297 = _T_2288[15:1];
  assign _T_2298 = {_T_2296,_T_2297};
  assign _T_2301 = _T_2300 == 16'h0;
  assign _T_2302 = _T_2300[0];
  assign _T_2303 = _T_2300[2];
  assign _T_2304 = _T_2302 ^ _T_2303;
  assign _T_2305 = _T_2300[3];
  assign _T_2306 = _T_2304 ^ _T_2305;
  assign _T_2307 = _T_2300[5];
  assign _T_2308 = _T_2306 ^ _T_2307;
  assign _T_2309 = _T_2300[15:1];
  assign _T_2310 = {_T_2308,_T_2309};
  assign _T_2313 = _T_2312 == 16'h0;
  assign _T_2314 = _T_2312[0];
  assign _T_2315 = _T_2312[2];
  assign _T_2316 = _T_2314 ^ _T_2315;
  assign _T_2317 = _T_2312[3];
  assign _T_2318 = _T_2316 ^ _T_2317;
  assign _T_2319 = _T_2312[5];
  assign _T_2320 = _T_2318 ^ _T_2319;
  assign _T_2321 = _T_2312[15:1];
  assign _T_2322 = {_T_2320,_T_2321};
  assign _T_2325 = _T_2324 == 16'h0;
  assign _T_2326 = _T_2324[0];
  assign _T_2327 = _T_2324[2];
  assign _T_2328 = _T_2326 ^ _T_2327;
  assign _T_2329 = _T_2324[3];
  assign _T_2330 = _T_2328 ^ _T_2329;
  assign _T_2331 = _T_2324[5];
  assign _T_2332 = _T_2330 ^ _T_2331;
  assign _T_2333 = _T_2324[15:1];
  assign _T_2334 = {_T_2332,_T_2333};
  assign _T_2337 = _T_2336 == 16'h0;
  assign _T_2338 = _T_2336[0];
  assign _T_2339 = _T_2336[2];
  assign _T_2340 = _T_2338 ^ _T_2339;
  assign _T_2341 = _T_2336[3];
  assign _T_2342 = _T_2340 ^ _T_2341;
  assign _T_2343 = _T_2336[5];
  assign _T_2344 = _T_2342 ^ _T_2343;
  assign _T_2345 = _T_2336[15:1];
  assign _T_2346 = {_T_2344,_T_2345};
  assign _T_2349 = _T_2348 == 16'h0;
  assign _T_2350 = _T_2348[0];
  assign _T_2351 = _T_2348[2];
  assign _T_2352 = _T_2350 ^ _T_2351;
  assign _T_2353 = _T_2348[3];
  assign _T_2354 = _T_2352 ^ _T_2353;
  assign _T_2355 = _T_2348[5];
  assign _T_2356 = _T_2354 ^ _T_2355;
  assign _T_2357 = _T_2348[15:1];
  assign _T_2358 = {_T_2356,_T_2357};
  assign _T_2361 = _T_2360 == 16'h0;
  assign _T_2362 = _T_2360[0];
  assign _T_2363 = _T_2360[2];
  assign _T_2364 = _T_2362 ^ _T_2363;
  assign _T_2365 = _T_2360[3];
  assign _T_2366 = _T_2364 ^ _T_2365;
  assign _T_2367 = _T_2360[5];
  assign _T_2368 = _T_2366 ^ _T_2367;
  assign _T_2369 = _T_2360[15:1];
  assign _T_2370 = {_T_2368,_T_2369};
  assign _T_2373 = _T_2372 == 16'h0;
  assign _T_2374 = _T_2372[0];
  assign _T_2375 = _T_2372[2];
  assign _T_2376 = _T_2374 ^ _T_2375;
  assign _T_2377 = _T_2372[3];
  assign _T_2378 = _T_2376 ^ _T_2377;
  assign _T_2379 = _T_2372[5];
  assign _T_2380 = _T_2378 ^ _T_2379;
  assign _T_2381 = _T_2372[15:1];
  assign _T_2382 = {_T_2380,_T_2381};
  assign _T_2385 = _T_2384 == 16'h0;
  assign _T_2386 = _T_2384[0];
  assign _T_2387 = _T_2384[2];
  assign _T_2388 = _T_2386 ^ _T_2387;
  assign _T_2389 = _T_2384[3];
  assign _T_2390 = _T_2388 ^ _T_2389;
  assign _T_2391 = _T_2384[5];
  assign _T_2392 = _T_2390 ^ _T_2391;
  assign _T_2393 = _T_2384[15:1];
  assign _T_2394 = {_T_2392,_T_2393};
  assign _T_2397 = _T_2396 == 16'h0;
  assign _T_2398 = _T_2396[0];
  assign _T_2399 = _T_2396[2];
  assign _T_2400 = _T_2398 ^ _T_2399;
  assign _T_2401 = _T_2396[3];
  assign _T_2402 = _T_2400 ^ _T_2401;
  assign _T_2403 = _T_2396[5];
  assign _T_2404 = _T_2402 ^ _T_2403;
  assign _T_2405 = _T_2396[15:1];
  assign _T_2406 = {_T_2404,_T_2405};
  assign _T_2409 = _T_2408 == 16'h0;
  assign _T_2410 = _T_2408[0];
  assign _T_2411 = _T_2408[2];
  assign _T_2412 = _T_2410 ^ _T_2411;
  assign _T_2413 = _T_2408[3];
  assign _T_2414 = _T_2412 ^ _T_2413;
  assign _T_2415 = _T_2408[5];
  assign _T_2416 = _T_2414 ^ _T_2415;
  assign _T_2417 = _T_2408[15:1];
  assign _T_2418 = {_T_2416,_T_2417};
  assign _T_2421 = _T_2420 == 16'h0;
  assign _T_2422 = _T_2420[0];
  assign _T_2423 = _T_2420[2];
  assign _T_2424 = _T_2422 ^ _T_2423;
  assign _T_2425 = _T_2420[3];
  assign _T_2426 = _T_2424 ^ _T_2425;
  assign _T_2427 = _T_2420[5];
  assign _T_2428 = _T_2426 ^ _T_2427;
  assign _T_2429 = _T_2420[15:1];
  assign _T_2430 = {_T_2428,_T_2429};
  assign _T_2433 = _T_2432 == 16'h0;
  assign _T_2434 = _T_2432[0];
  assign _T_2435 = _T_2432[2];
  assign _T_2436 = _T_2434 ^ _T_2435;
  assign _T_2437 = _T_2432[3];
  assign _T_2438 = _T_2436 ^ _T_2437;
  assign _T_2439 = _T_2432[5];
  assign _T_2440 = _T_2438 ^ _T_2439;
  assign _T_2441 = _T_2432[15:1];
  assign _T_2442 = {_T_2440,_T_2441};
  assign _T_2445 = _T_2444 == 16'h0;
  assign _T_2446 = _T_2444[0];
  assign _T_2447 = _T_2444[2];
  assign _T_2448 = _T_2446 ^ _T_2447;
  assign _T_2449 = _T_2444[3];
  assign _T_2450 = _T_2448 ^ _T_2449;
  assign _T_2451 = _T_2444[5];
  assign _T_2452 = _T_2450 ^ _T_2451;
  assign _T_2453 = _T_2444[15:1];
  assign _T_2454 = {_T_2452,_T_2453};
  assign _T_2457 = _T_2456 == 16'h0;
  assign _T_2458 = _T_2456[0];
  assign _T_2459 = _T_2456[2];
  assign _T_2460 = _T_2458 ^ _T_2459;
  assign _T_2461 = _T_2456[3];
  assign _T_2462 = _T_2460 ^ _T_2461;
  assign _T_2463 = _T_2456[5];
  assign _T_2464 = _T_2462 ^ _T_2463;
  assign _T_2465 = _T_2456[15:1];
  assign _T_2466 = {_T_2464,_T_2465};
  assign _T_2469 = _T_2468 == 16'h0;
  assign _T_2470 = _T_2468[0];
  assign _T_2471 = _T_2468[2];
  assign _T_2472 = _T_2470 ^ _T_2471;
  assign _T_2473 = _T_2468[3];
  assign _T_2474 = _T_2472 ^ _T_2473;
  assign _T_2475 = _T_2468[5];
  assign _T_2476 = _T_2474 ^ _T_2475;
  assign _T_2477 = _T_2468[15:1];
  assign _T_2478 = {_T_2476,_T_2477};
  assign _T_2481 = _T_2480 == 16'h0;
  assign _T_2482 = _T_2480[0];
  assign _T_2483 = _T_2480[2];
  assign _T_2484 = _T_2482 ^ _T_2483;
  assign _T_2485 = _T_2480[3];
  assign _T_2486 = _T_2484 ^ _T_2485;
  assign _T_2487 = _T_2480[5];
  assign _T_2488 = _T_2486 ^ _T_2487;
  assign _T_2489 = _T_2480[15:1];
  assign _T_2490 = {_T_2488,_T_2489};
  assign _T_2493 = _T_2492 == 16'h0;
  assign _T_2494 = _T_2492[0];
  assign _T_2495 = _T_2492[2];
  assign _T_2496 = _T_2494 ^ _T_2495;
  assign _T_2497 = _T_2492[3];
  assign _T_2498 = _T_2496 ^ _T_2497;
  assign _T_2499 = _T_2492[5];
  assign _T_2500 = _T_2498 ^ _T_2499;
  assign _T_2501 = _T_2492[15:1];
  assign _T_2502 = {_T_2500,_T_2501};
  assign _T_2505 = _T_2504 == 16'h0;
  assign _T_2506 = _T_2504[0];
  assign _T_2507 = _T_2504[2];
  assign _T_2508 = _T_2506 ^ _T_2507;
  assign _T_2509 = _T_2504[3];
  assign _T_2510 = _T_2508 ^ _T_2509;
  assign _T_2511 = _T_2504[5];
  assign _T_2512 = _T_2510 ^ _T_2511;
  assign _T_2513 = _T_2504[15:1];
  assign _T_2514 = {_T_2512,_T_2513};
  assign _T_2517 = _T_2516 == 16'h0;
  assign _T_2518 = _T_2516[0];
  assign _T_2519 = _T_2516[2];
  assign _T_2520 = _T_2518 ^ _T_2519;
  assign _T_2521 = _T_2516[3];
  assign _T_2522 = _T_2520 ^ _T_2521;
  assign _T_2523 = _T_2516[5];
  assign _T_2524 = _T_2522 ^ _T_2523;
  assign _T_2525 = _T_2516[15:1];
  assign _T_2526 = {_T_2524,_T_2525};
  assign _T_2529 = _T_2528 == 16'h0;
  assign _T_2530 = _T_2528[0];
  assign _T_2531 = _T_2528[2];
  assign _T_2532 = _T_2530 ^ _T_2531;
  assign _T_2533 = _T_2528[3];
  assign _T_2534 = _T_2532 ^ _T_2533;
  assign _T_2535 = _T_2528[5];
  assign _T_2536 = _T_2534 ^ _T_2535;
  assign _T_2537 = _T_2528[15:1];
  assign _T_2538 = {_T_2536,_T_2537};
  assign _T_2541 = _T_2540 == 16'h0;
  assign _T_2542 = _T_2540[0];
  assign _T_2543 = _T_2540[2];
  assign _T_2544 = _T_2542 ^ _T_2543;
  assign _T_2545 = _T_2540[3];
  assign _T_2546 = _T_2544 ^ _T_2545;
  assign _T_2547 = _T_2540[5];
  assign _T_2548 = _T_2546 ^ _T_2547;
  assign _T_2549 = _T_2540[15:1];
  assign _T_2550 = {_T_2548,_T_2549};
  assign _T_2553 = _T_2552 == 16'h0;
  assign _T_2554 = _T_2552[0];
  assign _T_2555 = _T_2552[2];
  assign _T_2556 = _T_2554 ^ _T_2555;
  assign _T_2557 = _T_2552[3];
  assign _T_2558 = _T_2556 ^ _T_2557;
  assign _T_2559 = _T_2552[5];
  assign _T_2560 = _T_2558 ^ _T_2559;
  assign _T_2561 = _T_2552[15:1];
  assign _T_2562 = {_T_2560,_T_2561};
  assign _T_2565 = _T_2564 == 16'h0;
  assign _T_2566 = _T_2564[0];
  assign _T_2567 = _T_2564[2];
  assign _T_2568 = _T_2566 ^ _T_2567;
  assign _T_2569 = _T_2564[3];
  assign _T_2570 = _T_2568 ^ _T_2569;
  assign _T_2571 = _T_2564[5];
  assign _T_2572 = _T_2570 ^ _T_2571;
  assign _T_2573 = _T_2564[15:1];
  assign _T_2574 = {_T_2572,_T_2573};
  assign _T_2577 = _T_2576 == 16'h0;
  assign _T_2578 = _T_2576[0];
  assign _T_2579 = _T_2576[2];
  assign _T_2580 = _T_2578 ^ _T_2579;
  assign _T_2581 = _T_2576[3];
  assign _T_2582 = _T_2580 ^ _T_2581;
  assign _T_2583 = _T_2576[5];
  assign _T_2584 = _T_2582 ^ _T_2583;
  assign _T_2585 = _T_2576[15:1];
  assign _T_2586 = {_T_2584,_T_2585};
  assign _T_2589 = _T_2588 == 16'h0;
  assign _T_2590 = _T_2588[0];
  assign _T_2591 = _T_2588[2];
  assign _T_2592 = _T_2590 ^ _T_2591;
  assign _T_2593 = _T_2588[3];
  assign _T_2594 = _T_2592 ^ _T_2593;
  assign _T_2595 = _T_2588[5];
  assign _T_2596 = _T_2594 ^ _T_2595;
  assign _T_2597 = _T_2588[15:1];
  assign _T_2598 = {_T_2596,_T_2597};
  assign _T_2601 = _T_2600 == 16'h0;
  assign _T_2602 = _T_2600[0];
  assign _T_2603 = _T_2600[2];
  assign _T_2604 = _T_2602 ^ _T_2603;
  assign _T_2605 = _T_2600[3];
  assign _T_2606 = _T_2604 ^ _T_2605;
  assign _T_2607 = _T_2600[5];
  assign _T_2608 = _T_2606 ^ _T_2607;
  assign _T_2609 = _T_2600[15:1];
  assign _T_2610 = {_T_2608,_T_2609};
  assign _T_2613 = _T_2612 == 16'h0;
  assign _T_2614 = _T_2612[0];
  assign _T_2615 = _T_2612[2];
  assign _T_2616 = _T_2614 ^ _T_2615;
  assign _T_2617 = _T_2612[3];
  assign _T_2618 = _T_2616 ^ _T_2617;
  assign _T_2619 = _T_2612[5];
  assign _T_2620 = _T_2618 ^ _T_2619;
  assign _T_2621 = _T_2612[15:1];
  assign _T_2622 = {_T_2620,_T_2621};
  assign _T_2625 = _T_2624 == 16'h0;
  assign _T_2626 = _T_2624[0];
  assign _T_2627 = _T_2624[2];
  assign _T_2628 = _T_2626 ^ _T_2627;
  assign _T_2629 = _T_2624[3];
  assign _T_2630 = _T_2628 ^ _T_2629;
  assign _T_2631 = _T_2624[5];
  assign _T_2632 = _T_2630 ^ _T_2631;
  assign _T_2633 = _T_2624[15:1];
  assign _T_2634 = {_T_2632,_T_2633};
  assign _T_2637 = _T_2636 == 16'h0;
  assign _T_2638 = _T_2636[0];
  assign _T_2639 = _T_2636[2];
  assign _T_2640 = _T_2638 ^ _T_2639;
  assign _T_2641 = _T_2636[3];
  assign _T_2642 = _T_2640 ^ _T_2641;
  assign _T_2643 = _T_2636[5];
  assign _T_2644 = _T_2642 ^ _T_2643;
  assign _T_2645 = _T_2636[15:1];
  assign _T_2646 = {_T_2644,_T_2645};
  assign _T_2649 = _T_2648 == 16'h0;
  assign _T_2650 = _T_2648[0];
  assign _T_2651 = _T_2648[2];
  assign _T_2652 = _T_2650 ^ _T_2651;
  assign _T_2653 = _T_2648[3];
  assign _T_2654 = _T_2652 ^ _T_2653;
  assign _T_2655 = _T_2648[5];
  assign _T_2656 = _T_2654 ^ _T_2655;
  assign _T_2657 = _T_2648[15:1];
  assign _T_2658 = {_T_2656,_T_2657};
  assign _T_2661 = _T_2660 == 16'h0;
  assign _T_2662 = _T_2660[0];
  assign _T_2663 = _T_2660[2];
  assign _T_2664 = _T_2662 ^ _T_2663;
  assign _T_2665 = _T_2660[3];
  assign _T_2666 = _T_2664 ^ _T_2665;
  assign _T_2667 = _T_2660[5];
  assign _T_2668 = _T_2666 ^ _T_2667;
  assign _T_2669 = _T_2660[15:1];
  assign _T_2670 = {_T_2668,_T_2669};
  assign _T_2673 = _T_2672 == 16'h0;
  assign _T_2674 = _T_2672[0];
  assign _T_2675 = _T_2672[2];
  assign _T_2676 = _T_2674 ^ _T_2675;
  assign _T_2677 = _T_2672[3];
  assign _T_2678 = _T_2676 ^ _T_2677;
  assign _T_2679 = _T_2672[5];
  assign _T_2680 = _T_2678 ^ _T_2679;
  assign _T_2681 = _T_2672[15:1];
  assign _T_2682 = {_T_2680,_T_2681};
  assign _T_2685 = _T_2684 == 16'h0;
  assign _T_2686 = _T_2684[0];
  assign _T_2687 = _T_2684[2];
  assign _T_2688 = _T_2686 ^ _T_2687;
  assign _T_2689 = _T_2684[3];
  assign _T_2690 = _T_2688 ^ _T_2689;
  assign _T_2691 = _T_2684[5];
  assign _T_2692 = _T_2690 ^ _T_2691;
  assign _T_2693 = _T_2684[15:1];
  assign _T_2694 = {_T_2692,_T_2693};
  assign _T_2697 = _T_2696 == 16'h0;
  assign _T_2698 = _T_2696[0];
  assign _T_2699 = _T_2696[2];
  assign _T_2700 = _T_2698 ^ _T_2699;
  assign _T_2701 = _T_2696[3];
  assign _T_2702 = _T_2700 ^ _T_2701;
  assign _T_2703 = _T_2696[5];
  assign _T_2704 = _T_2702 ^ _T_2703;
  assign _T_2705 = _T_2696[15:1];
  assign _T_2706 = {_T_2704,_T_2705};
  assign _T_2709 = _T_2708 == 16'h0;
  assign _T_2710 = _T_2708[0];
  assign _T_2711 = _T_2708[2];
  assign _T_2712 = _T_2710 ^ _T_2711;
  assign _T_2713 = _T_2708[3];
  assign _T_2714 = _T_2712 ^ _T_2713;
  assign _T_2715 = _T_2708[5];
  assign _T_2716 = _T_2714 ^ _T_2715;
  assign _T_2717 = _T_2708[15:1];
  assign _T_2718 = {_T_2716,_T_2717};
  assign _T_2721 = _T_2720 == 16'h0;
  assign _T_2722 = _T_2720[0];
  assign _T_2723 = _T_2720[2];
  assign _T_2724 = _T_2722 ^ _T_2723;
  assign _T_2725 = _T_2720[3];
  assign _T_2726 = _T_2724 ^ _T_2725;
  assign _T_2727 = _T_2720[5];
  assign _T_2728 = _T_2726 ^ _T_2727;
  assign _T_2729 = _T_2720[15:1];
  assign _T_2730 = {_T_2728,_T_2729};
  assign _T_2733 = _T_2732 == 16'h0;
  assign _T_2734 = _T_2732[0];
  assign _T_2735 = _T_2732[2];
  assign _T_2736 = _T_2734 ^ _T_2735;
  assign _T_2737 = _T_2732[3];
  assign _T_2738 = _T_2736 ^ _T_2737;
  assign _T_2739 = _T_2732[5];
  assign _T_2740 = _T_2738 ^ _T_2739;
  assign _T_2741 = _T_2732[15:1];
  assign _T_2742 = {_T_2740,_T_2741};
  assign _T_2745 = _T_2744 == 16'h0;
  assign _T_2746 = _T_2744[0];
  assign _T_2747 = _T_2744[2];
  assign _T_2748 = _T_2746 ^ _T_2747;
  assign _T_2749 = _T_2744[3];
  assign _T_2750 = _T_2748 ^ _T_2749;
  assign _T_2751 = _T_2744[5];
  assign _T_2752 = _T_2750 ^ _T_2751;
  assign _T_2753 = _T_2744[15:1];
  assign _T_2754 = {_T_2752,_T_2753};
  assign _T_2757 = _T_2756 == 16'h0;
  assign _T_2758 = _T_2756[0];
  assign _T_2759 = _T_2756[2];
  assign _T_2760 = _T_2758 ^ _T_2759;
  assign _T_2761 = _T_2756[3];
  assign _T_2762 = _T_2760 ^ _T_2761;
  assign _T_2763 = _T_2756[5];
  assign _T_2764 = _T_2762 ^ _T_2763;
  assign _T_2765 = _T_2756[15:1];
  assign _T_2766 = {_T_2764,_T_2765};
  assign _T_2769 = _T_2768 == 16'h0;
  assign _T_2770 = _T_2768[0];
  assign _T_2771 = _T_2768[2];
  assign _T_2772 = _T_2770 ^ _T_2771;
  assign _T_2773 = _T_2768[3];
  assign _T_2774 = _T_2772 ^ _T_2773;
  assign _T_2775 = _T_2768[5];
  assign _T_2776 = _T_2774 ^ _T_2775;
  assign _T_2777 = _T_2768[15:1];
  assign _T_2778 = {_T_2776,_T_2777};
  assign _T_2781 = _T_2780 == 16'h0;
  assign _T_2782 = _T_2780[0];
  assign _T_2783 = _T_2780[2];
  assign _T_2784 = _T_2782 ^ _T_2783;
  assign _T_2785 = _T_2780[3];
  assign _T_2786 = _T_2784 ^ _T_2785;
  assign _T_2787 = _T_2780[5];
  assign _T_2788 = _T_2786 ^ _T_2787;
  assign _T_2789 = _T_2780[15:1];
  assign _T_2790 = {_T_2788,_T_2789};
  assign _T_2793 = _T_2792 == 16'h0;
  assign _T_2794 = _T_2792[0];
  assign _T_2795 = _T_2792[2];
  assign _T_2796 = _T_2794 ^ _T_2795;
  assign _T_2797 = _T_2792[3];
  assign _T_2798 = _T_2796 ^ _T_2797;
  assign _T_2799 = _T_2792[5];
  assign _T_2800 = _T_2798 ^ _T_2799;
  assign _T_2801 = _T_2792[15:1];
  assign _T_2802 = {_T_2800,_T_2801};
  assign _T_2805 = _T_2804 == 16'h0;
  assign _T_2806 = _T_2804[0];
  assign _T_2807 = _T_2804[2];
  assign _T_2808 = _T_2806 ^ _T_2807;
  assign _T_2809 = _T_2804[3];
  assign _T_2810 = _T_2808 ^ _T_2809;
  assign _T_2811 = _T_2804[5];
  assign _T_2812 = _T_2810 ^ _T_2811;
  assign _T_2813 = _T_2804[15:1];
  assign _T_2814 = {_T_2812,_T_2813};
  assign _T_2817 = _T_2816 == 16'h0;
  assign _T_2818 = _T_2816[0];
  assign _T_2819 = _T_2816[2];
  assign _T_2820 = _T_2818 ^ _T_2819;
  assign _T_2821 = _T_2816[3];
  assign _T_2822 = _T_2820 ^ _T_2821;
  assign _T_2823 = _T_2816[5];
  assign _T_2824 = _T_2822 ^ _T_2823;
  assign _T_2825 = _T_2816[15:1];
  assign _T_2826 = {_T_2824,_T_2825};
  assign _T_2829 = _T_2828 == 16'h0;
  assign _T_2830 = _T_2828[0];
  assign _T_2831 = _T_2828[2];
  assign _T_2832 = _T_2830 ^ _T_2831;
  assign _T_2833 = _T_2828[3];
  assign _T_2834 = _T_2832 ^ _T_2833;
  assign _T_2835 = _T_2828[5];
  assign _T_2836 = _T_2834 ^ _T_2835;
  assign _T_2837 = _T_2828[15:1];
  assign _T_2838 = {_T_2836,_T_2837};
  assign _T_2841 = _T_2840 == 16'h0;
  assign _T_2842 = _T_2840[0];
  assign _T_2843 = _T_2840[2];
  assign _T_2844 = _T_2842 ^ _T_2843;
  assign _T_2845 = _T_2840[3];
  assign _T_2846 = _T_2844 ^ _T_2845;
  assign _T_2847 = _T_2840[5];
  assign _T_2848 = _T_2846 ^ _T_2847;
  assign _T_2849 = _T_2840[15:1];
  assign _T_2850 = {_T_2848,_T_2849};
  assign _T_2853 = _T_2852 == 16'h0;
  assign _T_2854 = _T_2852[0];
  assign _T_2855 = _T_2852[2];
  assign _T_2856 = _T_2854 ^ _T_2855;
  assign _T_2857 = _T_2852[3];
  assign _T_2858 = _T_2856 ^ _T_2857;
  assign _T_2859 = _T_2852[5];
  assign _T_2860 = _T_2858 ^ _T_2859;
  assign _T_2861 = _T_2852[15:1];
  assign _T_2862 = {_T_2860,_T_2861};
  assign _T_2865 = _T_2864 == 16'h0;
  assign _T_2866 = _T_2864[0];
  assign _T_2867 = _T_2864[2];
  assign _T_2868 = _T_2866 ^ _T_2867;
  assign _T_2869 = _T_2864[3];
  assign _T_2870 = _T_2868 ^ _T_2869;
  assign _T_2871 = _T_2864[5];
  assign _T_2872 = _T_2870 ^ _T_2871;
  assign _T_2873 = _T_2864[15:1];
  assign _T_2874 = {_T_2872,_T_2873};
  assign _T_2877 = _T_2876 == 16'h0;
  assign _T_2878 = _T_2876[0];
  assign _T_2879 = _T_2876[2];
  assign _T_2880 = _T_2878 ^ _T_2879;
  assign _T_2881 = _T_2876[3];
  assign _T_2882 = _T_2880 ^ _T_2881;
  assign _T_2883 = _T_2876[5];
  assign _T_2884 = _T_2882 ^ _T_2883;
  assign _T_2885 = _T_2876[15:1];
  assign _T_2886 = {_T_2884,_T_2885};
  assign _T_2889 = _T_2888 == 16'h0;
  assign _T_2890 = _T_2888[0];
  assign _T_2891 = _T_2888[2];
  assign _T_2892 = _T_2890 ^ _T_2891;
  assign _T_2893 = _T_2888[3];
  assign _T_2894 = _T_2892 ^ _T_2893;
  assign _T_2895 = _T_2888[5];
  assign _T_2896 = _T_2894 ^ _T_2895;
  assign _T_2897 = _T_2888[15:1];
  assign _T_2898 = {_T_2896,_T_2897};
  assign _T_2901 = _T_2900 == 16'h0;
  assign _T_2902 = _T_2900[0];
  assign _T_2903 = _T_2900[2];
  assign _T_2904 = _T_2902 ^ _T_2903;
  assign _T_2905 = _T_2900[3];
  assign _T_2906 = _T_2904 ^ _T_2905;
  assign _T_2907 = _T_2900[5];
  assign _T_2908 = _T_2906 ^ _T_2907;
  assign _T_2909 = _T_2900[15:1];
  assign _T_2910 = {_T_2908,_T_2909};
  assign _T_2913 = _T_2912 == 16'h0;
  assign _T_2914 = _T_2912[0];
  assign _T_2915 = _T_2912[2];
  assign _T_2916 = _T_2914 ^ _T_2915;
  assign _T_2917 = _T_2912[3];
  assign _T_2918 = _T_2916 ^ _T_2917;
  assign _T_2919 = _T_2912[5];
  assign _T_2920 = _T_2918 ^ _T_2919;
  assign _T_2921 = _T_2912[15:1];
  assign _T_2922 = {_T_2920,_T_2921};
  assign _T_2925 = _T_2924 == 16'h0;
  assign _T_2926 = _T_2924[0];
  assign _T_2927 = _T_2924[2];
  assign _T_2928 = _T_2926 ^ _T_2927;
  assign _T_2929 = _T_2924[3];
  assign _T_2930 = _T_2928 ^ _T_2929;
  assign _T_2931 = _T_2924[5];
  assign _T_2932 = _T_2930 ^ _T_2931;
  assign _T_2933 = _T_2924[15:1];
  assign _T_2934 = {_T_2932,_T_2933};
  assign _T_2937 = _T_2936 == 16'h0;
  assign _T_2938 = _T_2936[0];
  assign _T_2939 = _T_2936[2];
  assign _T_2940 = _T_2938 ^ _T_2939;
  assign _T_2941 = _T_2936[3];
  assign _T_2942 = _T_2940 ^ _T_2941;
  assign _T_2943 = _T_2936[5];
  assign _T_2944 = _T_2942 ^ _T_2943;
  assign _T_2945 = _T_2936[15:1];
  assign _T_2946 = {_T_2944,_T_2945};
  assign _T_2949 = _T_2948 == 16'h0;
  assign _T_2950 = _T_2948[0];
  assign _T_2951 = _T_2948[2];
  assign _T_2952 = _T_2950 ^ _T_2951;
  assign _T_2953 = _T_2948[3];
  assign _T_2954 = _T_2952 ^ _T_2953;
  assign _T_2955 = _T_2948[5];
  assign _T_2956 = _T_2954 ^ _T_2955;
  assign _T_2957 = _T_2948[15:1];
  assign _T_2958 = {_T_2956,_T_2957};
  assign _T_2961 = _T_2960 == 16'h0;
  assign _T_2962 = _T_2960[0];
  assign _T_2963 = _T_2960[2];
  assign _T_2964 = _T_2962 ^ _T_2963;
  assign _T_2965 = _T_2960[3];
  assign _T_2966 = _T_2964 ^ _T_2965;
  assign _T_2967 = _T_2960[5];
  assign _T_2968 = _T_2966 ^ _T_2967;
  assign _T_2969 = _T_2960[15:1];
  assign _T_2970 = {_T_2968,_T_2969};
  assign _T_2973 = _T_2972 == 16'h0;
  assign _T_2974 = _T_2972[0];
  assign _T_2975 = _T_2972[2];
  assign _T_2976 = _T_2974 ^ _T_2975;
  assign _T_2977 = _T_2972[3];
  assign _T_2978 = _T_2976 ^ _T_2977;
  assign _T_2979 = _T_2972[5];
  assign _T_2980 = _T_2978 ^ _T_2979;
  assign _T_2981 = _T_2972[15:1];
  assign _T_2982 = {_T_2980,_T_2981};
  assign _T_2985 = _T_2984 == 16'h0;
  assign _T_2986 = _T_2984[0];
  assign _T_2987 = _T_2984[2];
  assign _T_2988 = _T_2986 ^ _T_2987;
  assign _T_2989 = _T_2984[3];
  assign _T_2990 = _T_2988 ^ _T_2989;
  assign _T_2991 = _T_2984[5];
  assign _T_2992 = _T_2990 ^ _T_2991;
  assign _T_2993 = _T_2984[15:1];
  assign _T_2994 = {_T_2992,_T_2993};
  assign _T_2997 = _T_2996 == 16'h0;
  assign _T_2998 = _T_2996[0];
  assign _T_2999 = _T_2996[2];
  assign _T_3000 = _T_2998 ^ _T_2999;
  assign _T_3001 = _T_2996[3];
  assign _T_3002 = _T_3000 ^ _T_3001;
  assign _T_3003 = _T_2996[5];
  assign _T_3004 = _T_3002 ^ _T_3003;
  assign _T_3005 = _T_2996[15:1];
  assign _T_3006 = {_T_3004,_T_3005};
  assign _T_3009 = _T_3008 == 16'h0;
  assign _T_3010 = _T_3008[0];
  assign _T_3011 = _T_3008[2];
  assign _T_3012 = _T_3010 ^ _T_3011;
  assign _T_3013 = _T_3008[3];
  assign _T_3014 = _T_3012 ^ _T_3013;
  assign _T_3015 = _T_3008[5];
  assign _T_3016 = _T_3014 ^ _T_3015;
  assign _T_3017 = _T_3008[15:1];
  assign _T_3018 = {_T_3016,_T_3017};
  assign _T_3021 = _T_3020 == 16'h0;
  assign _T_3022 = _T_3020[0];
  assign _T_3023 = _T_3020[2];
  assign _T_3024 = _T_3022 ^ _T_3023;
  assign _T_3025 = _T_3020[3];
  assign _T_3026 = _T_3024 ^ _T_3025;
  assign _T_3027 = _T_3020[5];
  assign _T_3028 = _T_3026 ^ _T_3027;
  assign _T_3029 = _T_3020[15:1];
  assign _T_3030 = {_T_3028,_T_3029};
  assign _T_3033 = _T_3032 == 16'h0;
  assign _T_3034 = _T_3032[0];
  assign _T_3035 = _T_3032[2];
  assign _T_3036 = _T_3034 ^ _T_3035;
  assign _T_3037 = _T_3032[3];
  assign _T_3038 = _T_3036 ^ _T_3037;
  assign _T_3039 = _T_3032[5];
  assign _T_3040 = _T_3038 ^ _T_3039;
  assign _T_3041 = _T_3032[15:1];
  assign _T_3042 = {_T_3040,_T_3041};
  assign _T_3045 = _T_3044 == 16'h0;
  assign _T_3046 = _T_3044[0];
  assign _T_3047 = _T_3044[2];
  assign _T_3048 = _T_3046 ^ _T_3047;
  assign _T_3049 = _T_3044[3];
  assign _T_3050 = _T_3048 ^ _T_3049;
  assign _T_3051 = _T_3044[5];
  assign _T_3052 = _T_3050 ^ _T_3051;
  assign _T_3053 = _T_3044[15:1];
  assign _T_3054 = {_T_3052,_T_3053};
  assign _T_3057 = _T_3056 == 16'h0;
  assign _T_3058 = _T_3056[0];
  assign _T_3059 = _T_3056[2];
  assign _T_3060 = _T_3058 ^ _T_3059;
  assign _T_3061 = _T_3056[3];
  assign _T_3062 = _T_3060 ^ _T_3061;
  assign _T_3063 = _T_3056[5];
  assign _T_3064 = _T_3062 ^ _T_3063;
  assign _T_3065 = _T_3056[15:1];
  assign _T_3066 = {_T_3064,_T_3065};
  assign _T_3069 = _T_3068 == 16'h0;
  assign _T_3070 = _T_3068[0];
  assign _T_3071 = _T_3068[2];
  assign _T_3072 = _T_3070 ^ _T_3071;
  assign _T_3073 = _T_3068[3];
  assign _T_3074 = _T_3072 ^ _T_3073;
  assign _T_3075 = _T_3068[5];
  assign _T_3076 = _T_3074 ^ _T_3075;
  assign _T_3077 = _T_3068[15:1];
  assign _T_3078 = {_T_3076,_T_3077};
  assign _T_3081 = _T_3080 == 16'h0;
  assign _T_3082 = _T_3080[0];
  assign _T_3083 = _T_3080[2];
  assign _T_3084 = _T_3082 ^ _T_3083;
  assign _T_3085 = _T_3080[3];
  assign _T_3086 = _T_3084 ^ _T_3085;
  assign _T_3087 = _T_3080[5];
  assign _T_3088 = _T_3086 ^ _T_3087;
  assign _T_3089 = _T_3080[15:1];
  assign _T_3090 = {_T_3088,_T_3089};
  assign _T_3093 = _T_3092 == 16'h0;
  assign _T_3094 = _T_3092[0];
  assign _T_3095 = _T_3092[2];
  assign _T_3096 = _T_3094 ^ _T_3095;
  assign _T_3097 = _T_3092[3];
  assign _T_3098 = _T_3096 ^ _T_3097;
  assign _T_3099 = _T_3092[5];
  assign _T_3100 = _T_3098 ^ _T_3099;
  assign _T_3101 = _T_3092[15:1];
  assign _T_3102 = {_T_3100,_T_3101};
  assign _T_3105 = _T_3104 == 16'h0;
  assign _T_3106 = _T_3104[0];
  assign _T_3107 = _T_3104[2];
  assign _T_3108 = _T_3106 ^ _T_3107;
  assign _T_3109 = _T_3104[3];
  assign _T_3110 = _T_3108 ^ _T_3109;
  assign _T_3111 = _T_3104[5];
  assign _T_3112 = _T_3110 ^ _T_3111;
  assign _T_3113 = _T_3104[15:1];
  assign _T_3114 = {_T_3112,_T_3113};
  assign _T_3117 = _T_3116 == 16'h0;
  assign _T_3118 = _T_3116[0];
  assign _T_3119 = _T_3116[2];
  assign _T_3120 = _T_3118 ^ _T_3119;
  assign _T_3121 = _T_3116[3];
  assign _T_3122 = _T_3120 ^ _T_3121;
  assign _T_3123 = _T_3116[5];
  assign _T_3124 = _T_3122 ^ _T_3123;
  assign _T_3125 = _T_3116[15:1];
  assign _T_3126 = {_T_3124,_T_3125};
  assign _T_3129 = _T_3128 == 16'h0;
  assign _T_3130 = _T_3128[0];
  assign _T_3131 = _T_3128[2];
  assign _T_3132 = _T_3130 ^ _T_3131;
  assign _T_3133 = _T_3128[3];
  assign _T_3134 = _T_3132 ^ _T_3133;
  assign _T_3135 = _T_3128[5];
  assign _T_3136 = _T_3134 ^ _T_3135;
  assign _T_3137 = _T_3128[15:1];
  assign _T_3138 = {_T_3136,_T_3137};
  assign _T_3141 = _T_3140 == 16'h0;
  assign _T_3142 = _T_3140[0];
  assign _T_3143 = _T_3140[2];
  assign _T_3144 = _T_3142 ^ _T_3143;
  assign _T_3145 = _T_3140[3];
  assign _T_3146 = _T_3144 ^ _T_3145;
  assign _T_3147 = _T_3140[5];
  assign _T_3148 = _T_3146 ^ _T_3147;
  assign _T_3149 = _T_3140[15:1];
  assign _T_3150 = {_T_3148,_T_3149};
  assign _T_3153 = _T_3152 == 16'h0;
  assign _T_3154 = _T_3152[0];
  assign _T_3155 = _T_3152[2];
  assign _T_3156 = _T_3154 ^ _T_3155;
  assign _T_3157 = _T_3152[3];
  assign _T_3158 = _T_3156 ^ _T_3157;
  assign _T_3159 = _T_3152[5];
  assign _T_3160 = _T_3158 ^ _T_3159;
  assign _T_3161 = _T_3152[15:1];
  assign _T_3162 = {_T_3160,_T_3161};
  assign _T_3165 = _T_3164 == 16'h0;
  assign _T_3166 = _T_3164[0];
  assign _T_3167 = _T_3164[2];
  assign _T_3168 = _T_3166 ^ _T_3167;
  assign _T_3169 = _T_3164[3];
  assign _T_3170 = _T_3168 ^ _T_3169;
  assign _T_3171 = _T_3164[5];
  assign _T_3172 = _T_3170 ^ _T_3171;
  assign _T_3173 = _T_3164[15:1];
  assign _T_3174 = {_T_3172,_T_3173};
  assign _T_3177 = _T_3176 == 16'h0;
  assign _T_3178 = _T_3176[0];
  assign _T_3179 = _T_3176[2];
  assign _T_3180 = _T_3178 ^ _T_3179;
  assign _T_3181 = _T_3176[3];
  assign _T_3182 = _T_3180 ^ _T_3181;
  assign _T_3183 = _T_3176[5];
  assign _T_3184 = _T_3182 ^ _T_3183;
  assign _T_3185 = _T_3176[15:1];
  assign _T_3186 = {_T_3184,_T_3185};
  assign _T_3189 = _T_3188 == 16'h0;
  assign _T_3190 = _T_3188[0];
  assign _T_3191 = _T_3188[2];
  assign _T_3192 = _T_3190 ^ _T_3191;
  assign _T_3193 = _T_3188[3];
  assign _T_3194 = _T_3192 ^ _T_3193;
  assign _T_3195 = _T_3188[5];
  assign _T_3196 = _T_3194 ^ _T_3195;
  assign _T_3197 = _T_3188[15:1];
  assign _T_3198 = {_T_3196,_T_3197};
  assign _T_3201 = _T_3200 == 16'h0;
  assign _T_3202 = _T_3200[0];
  assign _T_3203 = _T_3200[2];
  assign _T_3204 = _T_3202 ^ _T_3203;
  assign _T_3205 = _T_3200[3];
  assign _T_3206 = _T_3204 ^ _T_3205;
  assign _T_3207 = _T_3200[5];
  assign _T_3208 = _T_3206 ^ _T_3207;
  assign _T_3209 = _T_3200[15:1];
  assign _T_3210 = {_T_3208,_T_3209};
  assign _T_3213 = _T_3212 == 16'h0;
  assign _T_3214 = _T_3212[0];
  assign _T_3215 = _T_3212[2];
  assign _T_3216 = _T_3214 ^ _T_3215;
  assign _T_3217 = _T_3212[3];
  assign _T_3218 = _T_3216 ^ _T_3217;
  assign _T_3219 = _T_3212[5];
  assign _T_3220 = _T_3218 ^ _T_3219;
  assign _T_3221 = _T_3212[15:1];
  assign _T_3222 = {_T_3220,_T_3221};
  assign _T_3225 = _T_3224 == 16'h0;
  assign _T_3226 = _T_3224[0];
  assign _T_3227 = _T_3224[2];
  assign _T_3228 = _T_3226 ^ _T_3227;
  assign _T_3229 = _T_3224[3];
  assign _T_3230 = _T_3228 ^ _T_3229;
  assign _T_3231 = _T_3224[5];
  assign _T_3232 = _T_3230 ^ _T_3231;
  assign _T_3233 = _T_3224[15:1];
  assign _T_3234 = {_T_3232,_T_3233};
  assign _T_3243 = {_T_1786,_T_1774,_T_1762,_T_1750,_T_1738,_T_1726,_T_1714};
  assign _T_3251 = {_T_1882,_T_1870,_T_1858,_T_1846,_T_1834,_T_1822,_T_1810,_T_1798,_T_3243};
  assign _T_3258 = {_T_1978,_T_1966,_T_1954,_T_1942,_T_1930,_T_1918,_T_1906,_T_1894};
  assign _T_3267 = {_T_2074,_T_2062,_T_2050,_T_2038,_T_2026,_T_2014,_T_2002,_T_1990,_T_3258,_T_3251};
  assign _T_3274 = {_T_2170,_T_2158,_T_2146,_T_2134,_T_2122,_T_2110,_T_2098,_T_2086};
  assign _T_3282 = {_T_2266,_T_2254,_T_2242,_T_2230,_T_2218,_T_2206,_T_2194,_T_2182,_T_3274};
  assign _T_3289 = {_T_2362,_T_2350,_T_2338,_T_2326,_T_2314,_T_2302,_T_2290,_T_2278};
  assign _T_3298 = {_T_2458,_T_2446,_T_2434,_T_2422,_T_2410,_T_2398,_T_2386,_T_2374,_T_3289,_T_3282};
  assign _T_3306 = {_T_2554,_T_2542,_T_2530,_T_2518,_T_2506,_T_2494,_T_2482,_T_2470};
  assign _T_3314 = {_T_2650,_T_2638,_T_2626,_T_2614,_T_2602,_T_2590,_T_2578,_T_2566,_T_3306};
  assign _T_3321 = {_T_2746,_T_2734,_T_2722,_T_2710,_T_2698,_T_2686,_T_2674,_T_2662};
  assign _T_3330 = {_T_2842,_T_2830,_T_2818,_T_2806,_T_2794,_T_2782,_T_2770,_T_2758,_T_3321,_T_3314};
  assign _T_3337 = {_T_2938,_T_2926,_T_2914,_T_2902,_T_2890,_T_2878,_T_2866,_T_2854};
  assign _T_3345 = {_T_3034,_T_3022,_T_3010,_T_2998,_T_2986,_T_2974,_T_2962,_T_2950,_T_3337};
  assign _T_3352 = {_T_3130,_T_3118,_T_3106,_T_3094,_T_3082,_T_3070,_T_3058,_T_3046};
  assign _T_3361 = {_T_3226,_T_3214,_T_3202,_T_3190,_T_3178,_T_3166,_T_3154,_T_3142,_T_3352,_T_3345};
  assign _T_3363 = {_T_3361,_T_3330,_T_3298,_T_3267};
  assign _GEN_513 = _T_185 ? _T_3363 : 127'h0;
  assign _GEN_514 = _T_179 ? _T_184 : {{1'd0}, _GEN_513};
  assign _GEN_515 = _T_51 ? 128'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa : _GEN_514;
  assign _GEN_516 = _T_49 ? 128'h7fffffffffffffffffffffffffffffff : _GEN_515;
  assign _GEN_517 = _T_48 ? 128'h0 : _GEN_516;
  assign _GEN_518 = _T_34 == 1'h0;
  assign _GEN_519 = _T_35 == 1'h0;
  assign _GEN_520 = _GEN_518 & _GEN_519;
  assign _GEN_521 = _T_36 == 1'h0;
  assign _GEN_522 = _GEN_520 & _GEN_521;
  assign _GEN_523 = _T_37 == 1'h0;
  assign _GEN_524 = _GEN_522 & _GEN_523;
  assign _GEN_525 = _T_38 == 1'h0;
  assign _GEN_526 = _GEN_524 & _GEN_525;
  assign _GEN_527 = _T_39 == 1'h0;
  assign _GEN_528 = _GEN_526 & _GEN_527;
  assign _GEN_540 = _T_48 == 1'h0;
  assign _GEN_541 = _T_49 == 1'h0;
  assign _GEN_542 = _GEN_540 & _GEN_541;
  assign _GEN_543 = _T_51 == 1'h0;
  assign _GEN_544 = _GEN_542 & _GEN_543;
  assign _GEN_545 = _T_179 == 1'h0;
  assign _GEN_546 = _GEN_544 & _GEN_545;
  assign _GEN_547 = _T_185 == 1'h0;
  assign _GEN_548 = _GEN_546 & _GEN_547;
  assign io_success = 1'h0;
  assign system_clock = dpiClockGate_clock_out;
  assign system_reset = CountAndDriver_io_driven_value;
  assign system_debug_psd_test_mode = 1'h0;
  assign system_debug_psd_test_mode_reset = 1'h0;
  assign system_debug_systemjtag_jtag_TCK = DPIJTAGDriver_jtag_TCK;
  assign system_debug_systemjtag_jtag_TMS = DPIJTAGDriver_jtag_TMS;
  assign system_debug_systemjtag_jtag_TDI = DPIJTAGDriver_jtag_TDI;
  assign system_debug_systemjtag_reset = reset;
  assign system_debug_systemjtag_mfr_id = 11'h0;
  assign system_core_clock_0 = ClockSkew_clkout;
  assign system_reset_vector_0 = 32'h20000000;
  assign system_rtc_toggle = _T_1;
  assign system_global_interrupts = _GEN_517[126:0];
  assign system_mem_port_axi4_0_aw_ready = testRAM_2_io_axi4_0_aw_ready;
  assign system_mem_port_axi4_0_w_ready = testRAM_2_io_axi4_0_w_ready;
  assign system_mem_port_axi4_0_b_valid = testRAM_2_io_axi4_0_b_valid;
  assign system_mem_port_axi4_0_b_bits_id = testRAM_2_io_axi4_0_b_bits_id;
  assign system_mem_port_axi4_0_b_bits_resp = testRAM_2_io_axi4_0_b_bits_resp;
  assign system_mem_port_axi4_0_ar_ready = testRAM_2_io_axi4_0_ar_ready;
  assign system_mem_port_axi4_0_r_valid = testRAM_2_io_axi4_0_r_valid;
  assign system_mem_port_axi4_0_r_bits_id = testRAM_2_io_axi4_0_r_bits_id;
  assign system_mem_port_axi4_0_r_bits_data = testRAM_2_io_axi4_0_r_bits_data;
  assign system_mem_port_axi4_0_r_bits_resp = testRAM_2_io_axi4_0_r_bits_resp;
  assign system_mem_port_axi4_0_r_bits_last = testRAM_2_io_axi4_0_r_bits_last;
  assign system_sys_port_axi4_0_aw_ready = testRAM_1_io_axi4_0_aw_ready;
  assign system_sys_port_axi4_0_w_ready = testRAM_1_io_axi4_0_w_ready;
  assign system_sys_port_axi4_0_b_valid = testRAM_1_io_axi4_0_b_valid;
  assign system_sys_port_axi4_0_b_bits_id = testRAM_1_io_axi4_0_b_bits_id;
  assign system_sys_port_axi4_0_b_bits_resp = testRAM_1_io_axi4_0_b_bits_resp;
  assign system_sys_port_axi4_0_ar_ready = testRAM_1_io_axi4_0_ar_ready;
  assign system_sys_port_axi4_0_r_valid = testRAM_1_io_axi4_0_r_valid;
  assign system_sys_port_axi4_0_r_bits_id = testRAM_1_io_axi4_0_r_bits_id;
  assign system_sys_port_axi4_0_r_bits_data = testRAM_1_io_axi4_0_r_bits_data;
  assign system_sys_port_axi4_0_r_bits_resp = testRAM_1_io_axi4_0_r_bits_resp;
  assign system_sys_port_axi4_0_r_bits_last = testRAM_1_io_axi4_0_r_bits_last;
  assign system_periph_port_axi4_0_aw_ready = testRAM_io_axi4_0_aw_ready;
  assign system_periph_port_axi4_0_w_ready = testRAM_io_axi4_0_w_ready;
  assign system_periph_port_axi4_0_b_valid = testRAM_io_axi4_0_b_valid;
  assign system_periph_port_axi4_0_b_bits_id = testRAM_io_axi4_0_b_bits_id;
  assign system_periph_port_axi4_0_b_bits_resp = testRAM_io_axi4_0_b_bits_resp;
  assign system_periph_port_axi4_0_ar_ready = testRAM_io_axi4_0_ar_ready;
  assign system_periph_port_axi4_0_r_valid = testRAM_io_axi4_0_r_valid;
  assign system_periph_port_axi4_0_r_bits_id = testRAM_io_axi4_0_r_bits_id;
  assign system_periph_port_axi4_0_r_bits_data = testRAM_io_axi4_0_r_bits_data;
  assign system_periph_port_axi4_0_r_bits_resp = testRAM_io_axi4_0_r_bits_resp;
  assign system_periph_port_axi4_0_r_bits_last = testRAM_io_axi4_0_r_bits_last;
  assign system_front_port_axi4_0_aw_valid = 1'h0;
  assign system_front_port_axi4_0_aw_bits_id = 8'h0;
  assign system_front_port_axi4_0_aw_bits_addr = 32'h0;
  assign system_front_port_axi4_0_aw_bits_len = 8'h0;
  assign system_front_port_axi4_0_aw_bits_size = 3'h0;
  assign system_front_port_axi4_0_aw_bits_burst = 2'h0;
  assign system_front_port_axi4_0_aw_bits_lock = 1'h0;
  assign system_front_port_axi4_0_aw_bits_cache = 4'h0;
  assign system_front_port_axi4_0_aw_bits_prot = 3'h0;
  assign system_front_port_axi4_0_aw_bits_qos = 4'h0;
  assign system_front_port_axi4_0_w_valid = 1'h0;
  assign system_front_port_axi4_0_w_bits_data = 32'h0;
  assign system_front_port_axi4_0_w_bits_strb = 4'h0;
  assign system_front_port_axi4_0_w_bits_last = 1'h0;
  assign system_front_port_axi4_0_b_ready = 1'h0;
  assign system_front_port_axi4_0_ar_valid = 1'h0;
  assign system_front_port_axi4_0_ar_bits_id = 8'h0;
  assign system_front_port_axi4_0_ar_bits_addr = 32'h0;
  assign system_front_port_axi4_0_ar_bits_len = 8'h0;
  assign system_front_port_axi4_0_ar_bits_size = 3'h0;
  assign system_front_port_axi4_0_ar_bits_burst = 2'h0;
  assign system_front_port_axi4_0_ar_bits_lock = 1'h0;
  assign system_front_port_axi4_0_ar_bits_cache = 4'h0;
  assign system_front_port_axi4_0_ar_bits_prot = 3'h0;
  assign system_front_port_axi4_0_ar_bits_qos = 4'h0;
  assign system_front_port_axi4_0_r_ready = 1'h0;
  assign func_clock_clock = clock;
  assign ClockSkew_clkin = func_clock_io_clock_out;
  assign Pow2ClockDivider_clock = func_clock_io_clock_out;
  assign dpiClockGate_clock_in = Pow2ClockDivider_io_clock_out;
  assign c_core_reset_driver_clock = clock;
  assign testRAM_clock = system_clock;
  assign testRAM_reset = system_reset;
  assign testRAM_io_axi4_0_aw_valid = system_periph_port_axi4_0_aw_valid;
  assign testRAM_io_axi4_0_aw_bits_id = system_periph_port_axi4_0_aw_bits_id;
  assign testRAM_io_axi4_0_aw_bits_addr = system_periph_port_axi4_0_aw_bits_addr;
  assign testRAM_io_axi4_0_aw_bits_len = system_periph_port_axi4_0_aw_bits_len;
  assign testRAM_io_axi4_0_aw_bits_size = system_periph_port_axi4_0_aw_bits_size;
  assign testRAM_io_axi4_0_aw_bits_burst = system_periph_port_axi4_0_aw_bits_burst;
  assign testRAM_io_axi4_0_aw_bits_lock = system_periph_port_axi4_0_aw_bits_lock;
  assign testRAM_io_axi4_0_aw_bits_cache = system_periph_port_axi4_0_aw_bits_cache;
  assign testRAM_io_axi4_0_aw_bits_prot = system_periph_port_axi4_0_aw_bits_prot;
  assign testRAM_io_axi4_0_aw_bits_qos = system_periph_port_axi4_0_aw_bits_qos;
  assign testRAM_io_axi4_0_w_valid = system_periph_port_axi4_0_w_valid;
  assign testRAM_io_axi4_0_w_bits_data = system_periph_port_axi4_0_w_bits_data;
  assign testRAM_io_axi4_0_w_bits_strb = system_periph_port_axi4_0_w_bits_strb;
  assign testRAM_io_axi4_0_w_bits_last = system_periph_port_axi4_0_w_bits_last;
  assign testRAM_io_axi4_0_b_ready = system_periph_port_axi4_0_b_ready;
  assign testRAM_io_axi4_0_ar_valid = system_periph_port_axi4_0_ar_valid;
  assign testRAM_io_axi4_0_ar_bits_id = system_periph_port_axi4_0_ar_bits_id;
  assign testRAM_io_axi4_0_ar_bits_addr = system_periph_port_axi4_0_ar_bits_addr;
  assign testRAM_io_axi4_0_ar_bits_len = system_periph_port_axi4_0_ar_bits_len;
  assign testRAM_io_axi4_0_ar_bits_size = system_periph_port_axi4_0_ar_bits_size;
  assign testRAM_io_axi4_0_ar_bits_burst = system_periph_port_axi4_0_ar_bits_burst;
  assign testRAM_io_axi4_0_ar_bits_lock = system_periph_port_axi4_0_ar_bits_lock;
  assign testRAM_io_axi4_0_ar_bits_cache = system_periph_port_axi4_0_ar_bits_cache;
  assign testRAM_io_axi4_0_ar_bits_prot = system_periph_port_axi4_0_ar_bits_prot;
  assign testRAM_io_axi4_0_ar_bits_qos = system_periph_port_axi4_0_ar_bits_qos;
  assign testRAM_io_axi4_0_r_ready = system_periph_port_axi4_0_r_ready;
  assign testRAM_1_clock = system_clock;
  assign testRAM_1_reset = system_reset;
  assign testRAM_1_io_axi4_0_aw_valid = system_sys_port_axi4_0_aw_valid;
  assign testRAM_1_io_axi4_0_aw_bits_id = system_sys_port_axi4_0_aw_bits_id;
  assign testRAM_1_io_axi4_0_aw_bits_addr = system_sys_port_axi4_0_aw_bits_addr;
  assign testRAM_1_io_axi4_0_aw_bits_len = system_sys_port_axi4_0_aw_bits_len;
  assign testRAM_1_io_axi4_0_aw_bits_size = system_sys_port_axi4_0_aw_bits_size;
  assign testRAM_1_io_axi4_0_aw_bits_burst = system_sys_port_axi4_0_aw_bits_burst;
  assign testRAM_1_io_axi4_0_aw_bits_lock = system_sys_port_axi4_0_aw_bits_lock;
  assign testRAM_1_io_axi4_0_aw_bits_cache = system_sys_port_axi4_0_aw_bits_cache;
  assign testRAM_1_io_axi4_0_aw_bits_prot = system_sys_port_axi4_0_aw_bits_prot;
  assign testRAM_1_io_axi4_0_aw_bits_qos = system_sys_port_axi4_0_aw_bits_qos;
  assign testRAM_1_io_axi4_0_w_valid = system_sys_port_axi4_0_w_valid;
  assign testRAM_1_io_axi4_0_w_bits_data = system_sys_port_axi4_0_w_bits_data;
  assign testRAM_1_io_axi4_0_w_bits_strb = system_sys_port_axi4_0_w_bits_strb;
  assign testRAM_1_io_axi4_0_w_bits_last = system_sys_port_axi4_0_w_bits_last;
  assign testRAM_1_io_axi4_0_b_ready = system_sys_port_axi4_0_b_ready;
  assign testRAM_1_io_axi4_0_ar_valid = system_sys_port_axi4_0_ar_valid;
  assign testRAM_1_io_axi4_0_ar_bits_id = system_sys_port_axi4_0_ar_bits_id;
  assign testRAM_1_io_axi4_0_ar_bits_addr = system_sys_port_axi4_0_ar_bits_addr;
  assign testRAM_1_io_axi4_0_ar_bits_len = system_sys_port_axi4_0_ar_bits_len;
  assign testRAM_1_io_axi4_0_ar_bits_size = system_sys_port_axi4_0_ar_bits_size;
  assign testRAM_1_io_axi4_0_ar_bits_burst = system_sys_port_axi4_0_ar_bits_burst;
  assign testRAM_1_io_axi4_0_ar_bits_lock = system_sys_port_axi4_0_ar_bits_lock;
  assign testRAM_1_io_axi4_0_ar_bits_cache = system_sys_port_axi4_0_ar_bits_cache;
  assign testRAM_1_io_axi4_0_ar_bits_prot = system_sys_port_axi4_0_ar_bits_prot;
  assign testRAM_1_io_axi4_0_ar_bits_qos = system_sys_port_axi4_0_ar_bits_qos;
  assign testRAM_1_io_axi4_0_r_ready = system_sys_port_axi4_0_r_ready;
  assign testRAM_2_clock = system_clock;
  assign testRAM_2_reset = system_reset;
  assign testRAM_2_io_axi4_0_aw_valid = system_mem_port_axi4_0_aw_valid;
  assign testRAM_2_io_axi4_0_aw_bits_id = system_mem_port_axi4_0_aw_bits_id;
  assign testRAM_2_io_axi4_0_aw_bits_addr = system_mem_port_axi4_0_aw_bits_addr;
  assign testRAM_2_io_axi4_0_aw_bits_len = system_mem_port_axi4_0_aw_bits_len;
  assign testRAM_2_io_axi4_0_aw_bits_size = system_mem_port_axi4_0_aw_bits_size;
  assign testRAM_2_io_axi4_0_aw_bits_burst = system_mem_port_axi4_0_aw_bits_burst;
  assign testRAM_2_io_axi4_0_aw_bits_lock = system_mem_port_axi4_0_aw_bits_lock;
  assign testRAM_2_io_axi4_0_aw_bits_cache = system_mem_port_axi4_0_aw_bits_cache;
  assign testRAM_2_io_axi4_0_aw_bits_prot = system_mem_port_axi4_0_aw_bits_prot;
  assign testRAM_2_io_axi4_0_aw_bits_qos = system_mem_port_axi4_0_aw_bits_qos;
  assign testRAM_2_io_axi4_0_w_valid = system_mem_port_axi4_0_w_valid;
  assign testRAM_2_io_axi4_0_w_bits_data = system_mem_port_axi4_0_w_bits_data;
  assign testRAM_2_io_axi4_0_w_bits_strb = system_mem_port_axi4_0_w_bits_strb;
  assign testRAM_2_io_axi4_0_w_bits_last = system_mem_port_axi4_0_w_bits_last;
  assign testRAM_2_io_axi4_0_b_ready = system_mem_port_axi4_0_b_ready;
  assign testRAM_2_io_axi4_0_ar_valid = system_mem_port_axi4_0_ar_valid;
  assign testRAM_2_io_axi4_0_ar_bits_id = system_mem_port_axi4_0_ar_bits_id;
  assign testRAM_2_io_axi4_0_ar_bits_addr = system_mem_port_axi4_0_ar_bits_addr;
  assign testRAM_2_io_axi4_0_ar_bits_len = system_mem_port_axi4_0_ar_bits_len;
  assign testRAM_2_io_axi4_0_ar_bits_size = system_mem_port_axi4_0_ar_bits_size;
  assign testRAM_2_io_axi4_0_ar_bits_burst = system_mem_port_axi4_0_ar_bits_burst;
  assign testRAM_2_io_axi4_0_ar_bits_lock = system_mem_port_axi4_0_ar_bits_lock;
  assign testRAM_2_io_axi4_0_ar_bits_cache = system_mem_port_axi4_0_ar_bits_cache;
  assign testRAM_2_io_axi4_0_ar_bits_prot = system_mem_port_axi4_0_ar_bits_prot;
  assign testRAM_2_io_axi4_0_ar_bits_qos = system_mem_port_axi4_0_ar_bits_qos;
  assign testRAM_2_io_axi4_0_r_ready = system_mem_port_axi4_0_r_ready;
  assign DPIJTAGDriver_clock = clock;
  assign DPIJTAGDriver_reset = reset;
  assign DPIJTAGDriver_jtag_TDO_data = system_debug_systemjtag_jtag_TDO_data;
  assign DPIJTAGDriver_jtag_TDO_driven = system_debug_systemjtag_jtag_TDO_driven;
  assign system_reset_driver_clock = clock;
  assign CountAndDriver_clock = clock;
  assign CountAndDriver_reset = reset;
  assign CountAndDriver_io_default_value = ndm_reset | _T_28;
  assign CountAndDriver_io_count = plusarg_reader_out[15:0];
  assign core_reset_driver_clock = clock;
  assign core_monitor_m_0_clock = DataTap_5__0_clock;
  assign core_monitor_m_0_reset = DataTap_5__0_reset;
  assign core_monitor_m_0_hartid = DataTap_5__0_hartid;
  assign core_monitor_m_0_timer = DataTap_5__0_timer;
  assign core_monitor_m_0_valid = DataTap_5__0_valid;
  assign core_monitor_m_0_pc = DataTap_5__0_pc;
  assign core_monitor_m_0_wrdst = DataTap_5__0_wrdst;
  assign core_monitor_m_0_wrdata = DataTap_5__0_wrdata;
  assign core_monitor_m_0_wren = DataTap_5__0_wren;
  assign core_monitor_m_0_rd0src = DataTap_5__0_rd0src;
  assign core_monitor_m_0_rd0val = DataTap_5__0_rd0val;
  assign core_monitor_m_0_rd1src = DataTap_5__0_rd1src;
  assign core_monitor_m_0_rd1val = DataTap_5__0_rd1val;
  assign core_monitor_m_0_inst = DataTap_5__0_inst;
  assign core_monitor_m_1_clock = DataTap_5__1_clock;
  assign core_monitor_m_1_reset = DataTap_5__1_reset;
  assign core_monitor_m_1_hartid = DataTap_5__1_hartid;
  assign core_monitor_m_1_timer = DataTap_5__1_timer;
  assign core_monitor_m_1_valid = DataTap_5__1_valid;
  assign core_monitor_m_1_pc = DataTap_5__1_pc;
  assign core_monitor_m_1_wrdst = DataTap_5__1_wrdst;
  assign core_monitor_m_1_wrdata = DataTap_5__1_wrdata;
  assign core_monitor_m_1_wren = DataTap_5__1_wren;
  assign core_monitor_m_1_rd0src = DataTap_5__1_rd0src;
  assign core_monitor_m_1_rd0val = DataTap_5__1_rd0val;
  assign core_monitor_m_1_rd1src = DataTap_5__1_rd1src;
  assign core_monitor_m_1_rd1val = DataTap_5__1_rd1val;
  assign core_monitor_m_1_inst = DataTap_5__1_inst;
  assign InterruptsDriver_clock = 1'h0;
  assign InterruptsDriver_reset = 1'h0;
  assign dpitbh_clock = 1'h0;
  assign dpitbh_reset = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_186 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_198 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_210 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_222 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_234 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_246 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_258 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_270 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_282 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_294 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_306 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_318 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_330 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_342 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_354 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_366 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_378 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_390 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_402 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_414 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_426 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_438 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_450 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_462 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_474 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_486 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_498 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_510 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_522 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_534 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_546 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_558 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_570 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_582 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_594 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_606 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_618 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_630 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_642 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_654 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_666 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_678 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_690 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_702 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_714 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_726 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_738 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_750 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_762 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_774 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_786 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_798 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_810 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_822 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_834 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_846 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_858 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_870 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_882 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_894 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_906 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_918 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_930 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_942 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_954 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_966 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_978 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_990 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1002 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1014 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1026 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1038 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1050 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1062 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1074 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1086 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1098 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1110 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1122 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1134 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1146 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1158 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1170 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1182 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1194 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1206 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1218 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1230 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1242 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1254 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1266 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1278 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1290 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1302 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1314 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1326 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1338 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1350 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1362 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1374 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1386 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1398 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1410 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1422 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1434 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1446 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1458 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1470 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1482 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1494 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1506 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1518 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_1530 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_1542 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_1554 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_1566 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1578 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1590 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1602 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1614 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1626 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_1638 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1650 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1662 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1674 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1686 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1698 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1712 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1724 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_1736 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_1748 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_1760 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_1772 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_1784 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_1796 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_1808 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_1820 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_1832 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_1844 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_1856 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_1868 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_1880 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_1892 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_1904 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_1916 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_1928 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_1940 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_1952 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_1964 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_1976 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_1988 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_2000 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_2012 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_2024 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_2036 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_2048 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_2060 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_2072 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_2084 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_2096 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_2108 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_2120 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_2132 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_2144 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_2156 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_2168 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_2180 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_2192 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_2204 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_2216 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_2228 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_2240 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_2252 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_2264 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_2276 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_2288 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_2300 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_2312 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_2324 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_2336 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_2348 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_2360 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_2372 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_2384 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_2396 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_2408 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_2420 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_2432 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_2444 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_2456 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_2468 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_2480 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_2492 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_2504 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_2516 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_2528 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_2540 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_2552 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_2564 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_2576 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_2588 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_2600 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_2612 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_2624 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_2636 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_2648 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_2660 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_2672 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_2684 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_2696 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_2708 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_2720 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_2732 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_2744 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_2756 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_2768 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_2780 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_2792 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_2804 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_2816 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_2828 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_2840 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_2852 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_2864 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_2876 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_2888 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_2900 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_2912 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_2924 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_2936 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_2948 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_2960 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_2972 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_2984 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_2996 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3008 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3020 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3032 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3044 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3056 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3068 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3080 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3092 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3104 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3116 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3128 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3140 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3152 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3164 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3176 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3188 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3200 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3212 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3224 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge dpiClockGate_clock_out) begin
    if (reset) begin
      _T <= 5'h0;
    end else begin
      _T <= _T_3;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_4) begin
        _T_1 <= _T_5;
      end
    end
  end
  always @(posedge clock) begin
    if (reset) begin
      value_1 <= 7'h0;
    end else begin
      if (_T_45) begin
        value_1 <= 7'h0;
      end else begin
        value_1 <= _T_47;
      end
    end
    if (reset) begin
      value_2 <= 7'h0;
    end else begin
      if (_T_45) begin
        if (_T_180) begin
          value_2 <= 7'h0;
        end else begin
          value_2 <= _T_182;
        end
      end
    end
    if (_T_187) begin
      _T_186 <= 16'h1;
    end else begin
      _T_186 <= _T_196;
    end
    if (_T_199) begin
      _T_198 <= 16'h1;
    end else begin
      _T_198 <= _T_208;
    end
    if (_T_211) begin
      _T_210 <= 16'h1;
    end else begin
      _T_210 <= _T_220;
    end
    if (_T_223) begin
      _T_222 <= 16'h1;
    end else begin
      _T_222 <= _T_232;
    end
    if (_T_235) begin
      _T_234 <= 16'h1;
    end else begin
      _T_234 <= _T_244;
    end
    if (_T_247) begin
      _T_246 <= 16'h1;
    end else begin
      _T_246 <= _T_256;
    end
    if (_T_259) begin
      _T_258 <= 16'h1;
    end else begin
      _T_258 <= _T_268;
    end
    if (_T_271) begin
      _T_270 <= 16'h1;
    end else begin
      _T_270 <= _T_280;
    end
    if (_T_283) begin
      _T_282 <= 16'h1;
    end else begin
      _T_282 <= _T_292;
    end
    if (_T_295) begin
      _T_294 <= 16'h1;
    end else begin
      _T_294 <= _T_304;
    end
    if (_T_307) begin
      _T_306 <= 16'h1;
    end else begin
      _T_306 <= _T_316;
    end
    if (_T_319) begin
      _T_318 <= 16'h1;
    end else begin
      _T_318 <= _T_328;
    end
    if (_T_331) begin
      _T_330 <= 16'h1;
    end else begin
      _T_330 <= _T_340;
    end
    if (_T_343) begin
      _T_342 <= 16'h1;
    end else begin
      _T_342 <= _T_352;
    end
    if (_T_355) begin
      _T_354 <= 16'h1;
    end else begin
      _T_354 <= _T_364;
    end
    if (_T_367) begin
      _T_366 <= 16'h1;
    end else begin
      _T_366 <= _T_376;
    end
    if (_T_379) begin
      _T_378 <= 16'h1;
    end else begin
      _T_378 <= _T_388;
    end
    if (_T_391) begin
      _T_390 <= 16'h1;
    end else begin
      _T_390 <= _T_400;
    end
    if (_T_403) begin
      _T_402 <= 16'h1;
    end else begin
      _T_402 <= _T_412;
    end
    if (_T_415) begin
      _T_414 <= 16'h1;
    end else begin
      _T_414 <= _T_424;
    end
    if (_T_427) begin
      _T_426 <= 16'h1;
    end else begin
      _T_426 <= _T_436;
    end
    if (_T_439) begin
      _T_438 <= 16'h1;
    end else begin
      _T_438 <= _T_448;
    end
    if (_T_451) begin
      _T_450 <= 16'h1;
    end else begin
      _T_450 <= _T_460;
    end
    if (_T_463) begin
      _T_462 <= 16'h1;
    end else begin
      _T_462 <= _T_472;
    end
    if (_T_475) begin
      _T_474 <= 16'h1;
    end else begin
      _T_474 <= _T_484;
    end
    if (_T_487) begin
      _T_486 <= 16'h1;
    end else begin
      _T_486 <= _T_496;
    end
    if (_T_499) begin
      _T_498 <= 16'h1;
    end else begin
      _T_498 <= _T_508;
    end
    if (_T_511) begin
      _T_510 <= 16'h1;
    end else begin
      _T_510 <= _T_520;
    end
    if (_T_523) begin
      _T_522 <= 16'h1;
    end else begin
      _T_522 <= _T_532;
    end
    if (_T_535) begin
      _T_534 <= 16'h1;
    end else begin
      _T_534 <= _T_544;
    end
    if (_T_547) begin
      _T_546 <= 16'h1;
    end else begin
      _T_546 <= _T_556;
    end
    if (_T_559) begin
      _T_558 <= 16'h1;
    end else begin
      _T_558 <= _T_568;
    end
    if (_T_571) begin
      _T_570 <= 16'h1;
    end else begin
      _T_570 <= _T_580;
    end
    if (_T_583) begin
      _T_582 <= 16'h1;
    end else begin
      _T_582 <= _T_592;
    end
    if (_T_595) begin
      _T_594 <= 16'h1;
    end else begin
      _T_594 <= _T_604;
    end
    if (_T_607) begin
      _T_606 <= 16'h1;
    end else begin
      _T_606 <= _T_616;
    end
    if (_T_619) begin
      _T_618 <= 16'h1;
    end else begin
      _T_618 <= _T_628;
    end
    if (_T_631) begin
      _T_630 <= 16'h1;
    end else begin
      _T_630 <= _T_640;
    end
    if (_T_643) begin
      _T_642 <= 16'h1;
    end else begin
      _T_642 <= _T_652;
    end
    if (_T_655) begin
      _T_654 <= 16'h1;
    end else begin
      _T_654 <= _T_664;
    end
    if (_T_667) begin
      _T_666 <= 16'h1;
    end else begin
      _T_666 <= _T_676;
    end
    if (_T_679) begin
      _T_678 <= 16'h1;
    end else begin
      _T_678 <= _T_688;
    end
    if (_T_691) begin
      _T_690 <= 16'h1;
    end else begin
      _T_690 <= _T_700;
    end
    if (_T_703) begin
      _T_702 <= 16'h1;
    end else begin
      _T_702 <= _T_712;
    end
    if (_T_715) begin
      _T_714 <= 16'h1;
    end else begin
      _T_714 <= _T_724;
    end
    if (_T_727) begin
      _T_726 <= 16'h1;
    end else begin
      _T_726 <= _T_736;
    end
    if (_T_739) begin
      _T_738 <= 16'h1;
    end else begin
      _T_738 <= _T_748;
    end
    if (_T_751) begin
      _T_750 <= 16'h1;
    end else begin
      _T_750 <= _T_760;
    end
    if (_T_763) begin
      _T_762 <= 16'h1;
    end else begin
      _T_762 <= _T_772;
    end
    if (_T_775) begin
      _T_774 <= 16'h1;
    end else begin
      _T_774 <= _T_784;
    end
    if (_T_787) begin
      _T_786 <= 16'h1;
    end else begin
      _T_786 <= _T_796;
    end
    if (_T_799) begin
      _T_798 <= 16'h1;
    end else begin
      _T_798 <= _T_808;
    end
    if (_T_811) begin
      _T_810 <= 16'h1;
    end else begin
      _T_810 <= _T_820;
    end
    if (_T_823) begin
      _T_822 <= 16'h1;
    end else begin
      _T_822 <= _T_832;
    end
    if (_T_835) begin
      _T_834 <= 16'h1;
    end else begin
      _T_834 <= _T_844;
    end
    if (_T_847) begin
      _T_846 <= 16'h1;
    end else begin
      _T_846 <= _T_856;
    end
    if (_T_859) begin
      _T_858 <= 16'h1;
    end else begin
      _T_858 <= _T_868;
    end
    if (_T_871) begin
      _T_870 <= 16'h1;
    end else begin
      _T_870 <= _T_880;
    end
    if (_T_883) begin
      _T_882 <= 16'h1;
    end else begin
      _T_882 <= _T_892;
    end
    if (_T_895) begin
      _T_894 <= 16'h1;
    end else begin
      _T_894 <= _T_904;
    end
    if (_T_907) begin
      _T_906 <= 16'h1;
    end else begin
      _T_906 <= _T_916;
    end
    if (_T_919) begin
      _T_918 <= 16'h1;
    end else begin
      _T_918 <= _T_928;
    end
    if (_T_931) begin
      _T_930 <= 16'h1;
    end else begin
      _T_930 <= _T_940;
    end
    if (_T_943) begin
      _T_942 <= 16'h1;
    end else begin
      _T_942 <= _T_952;
    end
    if (_T_955) begin
      _T_954 <= 16'h1;
    end else begin
      _T_954 <= _T_964;
    end
    if (_T_967) begin
      _T_966 <= 16'h1;
    end else begin
      _T_966 <= _T_976;
    end
    if (_T_979) begin
      _T_978 <= 16'h1;
    end else begin
      _T_978 <= _T_988;
    end
    if (_T_991) begin
      _T_990 <= 16'h1;
    end else begin
      _T_990 <= _T_1000;
    end
    if (_T_1003) begin
      _T_1002 <= 16'h1;
    end else begin
      _T_1002 <= _T_1012;
    end
    if (_T_1015) begin
      _T_1014 <= 16'h1;
    end else begin
      _T_1014 <= _T_1024;
    end
    if (_T_1027) begin
      _T_1026 <= 16'h1;
    end else begin
      _T_1026 <= _T_1036;
    end
    if (_T_1039) begin
      _T_1038 <= 16'h1;
    end else begin
      _T_1038 <= _T_1048;
    end
    if (_T_1051) begin
      _T_1050 <= 16'h1;
    end else begin
      _T_1050 <= _T_1060;
    end
    if (_T_1063) begin
      _T_1062 <= 16'h1;
    end else begin
      _T_1062 <= _T_1072;
    end
    if (_T_1075) begin
      _T_1074 <= 16'h1;
    end else begin
      _T_1074 <= _T_1084;
    end
    if (_T_1087) begin
      _T_1086 <= 16'h1;
    end else begin
      _T_1086 <= _T_1096;
    end
    if (_T_1099) begin
      _T_1098 <= 16'h1;
    end else begin
      _T_1098 <= _T_1108;
    end
    if (_T_1111) begin
      _T_1110 <= 16'h1;
    end else begin
      _T_1110 <= _T_1120;
    end
    if (_T_1123) begin
      _T_1122 <= 16'h1;
    end else begin
      _T_1122 <= _T_1132;
    end
    if (_T_1135) begin
      _T_1134 <= 16'h1;
    end else begin
      _T_1134 <= _T_1144;
    end
    if (_T_1147) begin
      _T_1146 <= 16'h1;
    end else begin
      _T_1146 <= _T_1156;
    end
    if (_T_1159) begin
      _T_1158 <= 16'h1;
    end else begin
      _T_1158 <= _T_1168;
    end
    if (_T_1171) begin
      _T_1170 <= 16'h1;
    end else begin
      _T_1170 <= _T_1180;
    end
    if (_T_1183) begin
      _T_1182 <= 16'h1;
    end else begin
      _T_1182 <= _T_1192;
    end
    if (_T_1195) begin
      _T_1194 <= 16'h1;
    end else begin
      _T_1194 <= _T_1204;
    end
    if (_T_1207) begin
      _T_1206 <= 16'h1;
    end else begin
      _T_1206 <= _T_1216;
    end
    if (_T_1219) begin
      _T_1218 <= 16'h1;
    end else begin
      _T_1218 <= _T_1228;
    end
    if (_T_1231) begin
      _T_1230 <= 16'h1;
    end else begin
      _T_1230 <= _T_1240;
    end
    if (_T_1243) begin
      _T_1242 <= 16'h1;
    end else begin
      _T_1242 <= _T_1252;
    end
    if (_T_1255) begin
      _T_1254 <= 16'h1;
    end else begin
      _T_1254 <= _T_1264;
    end
    if (_T_1267) begin
      _T_1266 <= 16'h1;
    end else begin
      _T_1266 <= _T_1276;
    end
    if (_T_1279) begin
      _T_1278 <= 16'h1;
    end else begin
      _T_1278 <= _T_1288;
    end
    if (_T_1291) begin
      _T_1290 <= 16'h1;
    end else begin
      _T_1290 <= _T_1300;
    end
    if (_T_1303) begin
      _T_1302 <= 16'h1;
    end else begin
      _T_1302 <= _T_1312;
    end
    if (_T_1315) begin
      _T_1314 <= 16'h1;
    end else begin
      _T_1314 <= _T_1324;
    end
    if (_T_1327) begin
      _T_1326 <= 16'h1;
    end else begin
      _T_1326 <= _T_1336;
    end
    if (_T_1339) begin
      _T_1338 <= 16'h1;
    end else begin
      _T_1338 <= _T_1348;
    end
    if (_T_1351) begin
      _T_1350 <= 16'h1;
    end else begin
      _T_1350 <= _T_1360;
    end
    if (_T_1363) begin
      _T_1362 <= 16'h1;
    end else begin
      _T_1362 <= _T_1372;
    end
    if (_T_1375) begin
      _T_1374 <= 16'h1;
    end else begin
      _T_1374 <= _T_1384;
    end
    if (_T_1387) begin
      _T_1386 <= 16'h1;
    end else begin
      _T_1386 <= _T_1396;
    end
    if (_T_1399) begin
      _T_1398 <= 16'h1;
    end else begin
      _T_1398 <= _T_1408;
    end
    if (_T_1411) begin
      _T_1410 <= 16'h1;
    end else begin
      _T_1410 <= _T_1420;
    end
    if (_T_1423) begin
      _T_1422 <= 16'h1;
    end else begin
      _T_1422 <= _T_1432;
    end
    if (_T_1435) begin
      _T_1434 <= 16'h1;
    end else begin
      _T_1434 <= _T_1444;
    end
    if (_T_1447) begin
      _T_1446 <= 16'h1;
    end else begin
      _T_1446 <= _T_1456;
    end
    if (_T_1459) begin
      _T_1458 <= 16'h1;
    end else begin
      _T_1458 <= _T_1468;
    end
    if (_T_1471) begin
      _T_1470 <= 16'h1;
    end else begin
      _T_1470 <= _T_1480;
    end
    if (_T_1483) begin
      _T_1482 <= 16'h1;
    end else begin
      _T_1482 <= _T_1492;
    end
    if (_T_1495) begin
      _T_1494 <= 16'h1;
    end else begin
      _T_1494 <= _T_1504;
    end
    if (_T_1507) begin
      _T_1506 <= 16'h1;
    end else begin
      _T_1506 <= _T_1516;
    end
    if (_T_1519) begin
      _T_1518 <= 16'h1;
    end else begin
      _T_1518 <= _T_1528;
    end
    if (_T_1531) begin
      _T_1530 <= 16'h1;
    end else begin
      _T_1530 <= _T_1540;
    end
    if (_T_1543) begin
      _T_1542 <= 16'h1;
    end else begin
      _T_1542 <= _T_1552;
    end
    if (_T_1555) begin
      _T_1554 <= 16'h1;
    end else begin
      _T_1554 <= _T_1564;
    end
    if (_T_1567) begin
      _T_1566 <= 16'h1;
    end else begin
      _T_1566 <= _T_1576;
    end
    if (_T_1579) begin
      _T_1578 <= 16'h1;
    end else begin
      _T_1578 <= _T_1588;
    end
    if (_T_1591) begin
      _T_1590 <= 16'h1;
    end else begin
      _T_1590 <= _T_1600;
    end
    if (_T_1603) begin
      _T_1602 <= 16'h1;
    end else begin
      _T_1602 <= _T_1612;
    end
    if (_T_1615) begin
      _T_1614 <= 16'h1;
    end else begin
      _T_1614 <= _T_1624;
    end
    if (_T_1627) begin
      _T_1626 <= 16'h1;
    end else begin
      _T_1626 <= _T_1636;
    end
    if (_T_1639) begin
      _T_1638 <= 16'h1;
    end else begin
      _T_1638 <= _T_1648;
    end
    if (_T_1651) begin
      _T_1650 <= 16'h1;
    end else begin
      _T_1650 <= _T_1660;
    end
    if (_T_1663) begin
      _T_1662 <= 16'h1;
    end else begin
      _T_1662 <= _T_1672;
    end
    if (_T_1675) begin
      _T_1674 <= 16'h1;
    end else begin
      _T_1674 <= _T_1684;
    end
    if (_T_1687) begin
      _T_1686 <= 16'h1;
    end else begin
      _T_1686 <= _T_1696;
    end
    if (_T_1699) begin
      _T_1698 <= 16'h1;
    end else begin
      _T_1698 <= _T_1708;
    end
    if (_T_188) begin
      if (_T_1713) begin
        _T_1712 <= 16'h1;
      end else begin
        _T_1712 <= _T_1722;
      end
    end
    if (_T_200) begin
      if (_T_1725) begin
        _T_1724 <= 16'h1;
      end else begin
        _T_1724 <= _T_1734;
      end
    end
    if (_T_212) begin
      if (_T_1737) begin
        _T_1736 <= 16'h1;
      end else begin
        _T_1736 <= _T_1746;
      end
    end
    if (_T_224) begin
      if (_T_1749) begin
        _T_1748 <= 16'h1;
      end else begin
        _T_1748 <= _T_1758;
      end
    end
    if (_T_236) begin
      if (_T_1761) begin
        _T_1760 <= 16'h1;
      end else begin
        _T_1760 <= _T_1770;
      end
    end
    if (_T_248) begin
      if (_T_1773) begin
        _T_1772 <= 16'h1;
      end else begin
        _T_1772 <= _T_1782;
      end
    end
    if (_T_260) begin
      if (_T_1785) begin
        _T_1784 <= 16'h1;
      end else begin
        _T_1784 <= _T_1794;
      end
    end
    if (_T_272) begin
      if (_T_1797) begin
        _T_1796 <= 16'h1;
      end else begin
        _T_1796 <= _T_1806;
      end
    end
    if (_T_284) begin
      if (_T_1809) begin
        _T_1808 <= 16'h1;
      end else begin
        _T_1808 <= _T_1818;
      end
    end
    if (_T_296) begin
      if (_T_1821) begin
        _T_1820 <= 16'h1;
      end else begin
        _T_1820 <= _T_1830;
      end
    end
    if (_T_308) begin
      if (_T_1833) begin
        _T_1832 <= 16'h1;
      end else begin
        _T_1832 <= _T_1842;
      end
    end
    if (_T_320) begin
      if (_T_1845) begin
        _T_1844 <= 16'h1;
      end else begin
        _T_1844 <= _T_1854;
      end
    end
    if (_T_332) begin
      if (_T_1857) begin
        _T_1856 <= 16'h1;
      end else begin
        _T_1856 <= _T_1866;
      end
    end
    if (_T_344) begin
      if (_T_1869) begin
        _T_1868 <= 16'h1;
      end else begin
        _T_1868 <= _T_1878;
      end
    end
    if (_T_356) begin
      if (_T_1881) begin
        _T_1880 <= 16'h1;
      end else begin
        _T_1880 <= _T_1890;
      end
    end
    if (_T_368) begin
      if (_T_1893) begin
        _T_1892 <= 16'h1;
      end else begin
        _T_1892 <= _T_1902;
      end
    end
    if (_T_380) begin
      if (_T_1905) begin
        _T_1904 <= 16'h1;
      end else begin
        _T_1904 <= _T_1914;
      end
    end
    if (_T_392) begin
      if (_T_1917) begin
        _T_1916 <= 16'h1;
      end else begin
        _T_1916 <= _T_1926;
      end
    end
    if (_T_404) begin
      if (_T_1929) begin
        _T_1928 <= 16'h1;
      end else begin
        _T_1928 <= _T_1938;
      end
    end
    if (_T_416) begin
      if (_T_1941) begin
        _T_1940 <= 16'h1;
      end else begin
        _T_1940 <= _T_1950;
      end
    end
    if (_T_428) begin
      if (_T_1953) begin
        _T_1952 <= 16'h1;
      end else begin
        _T_1952 <= _T_1962;
      end
    end
    if (_T_440) begin
      if (_T_1965) begin
        _T_1964 <= 16'h1;
      end else begin
        _T_1964 <= _T_1974;
      end
    end
    if (_T_452) begin
      if (_T_1977) begin
        _T_1976 <= 16'h1;
      end else begin
        _T_1976 <= _T_1986;
      end
    end
    if (_T_464) begin
      if (_T_1989) begin
        _T_1988 <= 16'h1;
      end else begin
        _T_1988 <= _T_1998;
      end
    end
    if (_T_476) begin
      if (_T_2001) begin
        _T_2000 <= 16'h1;
      end else begin
        _T_2000 <= _T_2010;
      end
    end
    if (_T_488) begin
      if (_T_2013) begin
        _T_2012 <= 16'h1;
      end else begin
        _T_2012 <= _T_2022;
      end
    end
    if (_T_500) begin
      if (_T_2025) begin
        _T_2024 <= 16'h1;
      end else begin
        _T_2024 <= _T_2034;
      end
    end
    if (_T_512) begin
      if (_T_2037) begin
        _T_2036 <= 16'h1;
      end else begin
        _T_2036 <= _T_2046;
      end
    end
    if (_T_524) begin
      if (_T_2049) begin
        _T_2048 <= 16'h1;
      end else begin
        _T_2048 <= _T_2058;
      end
    end
    if (_T_536) begin
      if (_T_2061) begin
        _T_2060 <= 16'h1;
      end else begin
        _T_2060 <= _T_2070;
      end
    end
    if (_T_548) begin
      if (_T_2073) begin
        _T_2072 <= 16'h1;
      end else begin
        _T_2072 <= _T_2082;
      end
    end
    if (_T_560) begin
      if (_T_2085) begin
        _T_2084 <= 16'h1;
      end else begin
        _T_2084 <= _T_2094;
      end
    end
    if (_T_572) begin
      if (_T_2097) begin
        _T_2096 <= 16'h1;
      end else begin
        _T_2096 <= _T_2106;
      end
    end
    if (_T_584) begin
      if (_T_2109) begin
        _T_2108 <= 16'h1;
      end else begin
        _T_2108 <= _T_2118;
      end
    end
    if (_T_596) begin
      if (_T_2121) begin
        _T_2120 <= 16'h1;
      end else begin
        _T_2120 <= _T_2130;
      end
    end
    if (_T_608) begin
      if (_T_2133) begin
        _T_2132 <= 16'h1;
      end else begin
        _T_2132 <= _T_2142;
      end
    end
    if (_T_620) begin
      if (_T_2145) begin
        _T_2144 <= 16'h1;
      end else begin
        _T_2144 <= _T_2154;
      end
    end
    if (_T_632) begin
      if (_T_2157) begin
        _T_2156 <= 16'h1;
      end else begin
        _T_2156 <= _T_2166;
      end
    end
    if (_T_644) begin
      if (_T_2169) begin
        _T_2168 <= 16'h1;
      end else begin
        _T_2168 <= _T_2178;
      end
    end
    if (_T_656) begin
      if (_T_2181) begin
        _T_2180 <= 16'h1;
      end else begin
        _T_2180 <= _T_2190;
      end
    end
    if (_T_668) begin
      if (_T_2193) begin
        _T_2192 <= 16'h1;
      end else begin
        _T_2192 <= _T_2202;
      end
    end
    if (_T_680) begin
      if (_T_2205) begin
        _T_2204 <= 16'h1;
      end else begin
        _T_2204 <= _T_2214;
      end
    end
    if (_T_692) begin
      if (_T_2217) begin
        _T_2216 <= 16'h1;
      end else begin
        _T_2216 <= _T_2226;
      end
    end
    if (_T_704) begin
      if (_T_2229) begin
        _T_2228 <= 16'h1;
      end else begin
        _T_2228 <= _T_2238;
      end
    end
    if (_T_716) begin
      if (_T_2241) begin
        _T_2240 <= 16'h1;
      end else begin
        _T_2240 <= _T_2250;
      end
    end
    if (_T_728) begin
      if (_T_2253) begin
        _T_2252 <= 16'h1;
      end else begin
        _T_2252 <= _T_2262;
      end
    end
    if (_T_740) begin
      if (_T_2265) begin
        _T_2264 <= 16'h1;
      end else begin
        _T_2264 <= _T_2274;
      end
    end
    if (_T_752) begin
      if (_T_2277) begin
        _T_2276 <= 16'h1;
      end else begin
        _T_2276 <= _T_2286;
      end
    end
    if (_T_764) begin
      if (_T_2289) begin
        _T_2288 <= 16'h1;
      end else begin
        _T_2288 <= _T_2298;
      end
    end
    if (_T_776) begin
      if (_T_2301) begin
        _T_2300 <= 16'h1;
      end else begin
        _T_2300 <= _T_2310;
      end
    end
    if (_T_788) begin
      if (_T_2313) begin
        _T_2312 <= 16'h1;
      end else begin
        _T_2312 <= _T_2322;
      end
    end
    if (_T_800) begin
      if (_T_2325) begin
        _T_2324 <= 16'h1;
      end else begin
        _T_2324 <= _T_2334;
      end
    end
    if (_T_812) begin
      if (_T_2337) begin
        _T_2336 <= 16'h1;
      end else begin
        _T_2336 <= _T_2346;
      end
    end
    if (_T_824) begin
      if (_T_2349) begin
        _T_2348 <= 16'h1;
      end else begin
        _T_2348 <= _T_2358;
      end
    end
    if (_T_836) begin
      if (_T_2361) begin
        _T_2360 <= 16'h1;
      end else begin
        _T_2360 <= _T_2370;
      end
    end
    if (_T_848) begin
      if (_T_2373) begin
        _T_2372 <= 16'h1;
      end else begin
        _T_2372 <= _T_2382;
      end
    end
    if (_T_860) begin
      if (_T_2385) begin
        _T_2384 <= 16'h1;
      end else begin
        _T_2384 <= _T_2394;
      end
    end
    if (_T_872) begin
      if (_T_2397) begin
        _T_2396 <= 16'h1;
      end else begin
        _T_2396 <= _T_2406;
      end
    end
    if (_T_884) begin
      if (_T_2409) begin
        _T_2408 <= 16'h1;
      end else begin
        _T_2408 <= _T_2418;
      end
    end
    if (_T_896) begin
      if (_T_2421) begin
        _T_2420 <= 16'h1;
      end else begin
        _T_2420 <= _T_2430;
      end
    end
    if (_T_908) begin
      if (_T_2433) begin
        _T_2432 <= 16'h1;
      end else begin
        _T_2432 <= _T_2442;
      end
    end
    if (_T_920) begin
      if (_T_2445) begin
        _T_2444 <= 16'h1;
      end else begin
        _T_2444 <= _T_2454;
      end
    end
    if (_T_932) begin
      if (_T_2457) begin
        _T_2456 <= 16'h1;
      end else begin
        _T_2456 <= _T_2466;
      end
    end
    if (_T_944) begin
      if (_T_2469) begin
        _T_2468 <= 16'h1;
      end else begin
        _T_2468 <= _T_2478;
      end
    end
    if (_T_956) begin
      if (_T_2481) begin
        _T_2480 <= 16'h1;
      end else begin
        _T_2480 <= _T_2490;
      end
    end
    if (_T_968) begin
      if (_T_2493) begin
        _T_2492 <= 16'h1;
      end else begin
        _T_2492 <= _T_2502;
      end
    end
    if (_T_980) begin
      if (_T_2505) begin
        _T_2504 <= 16'h1;
      end else begin
        _T_2504 <= _T_2514;
      end
    end
    if (_T_992) begin
      if (_T_2517) begin
        _T_2516 <= 16'h1;
      end else begin
        _T_2516 <= _T_2526;
      end
    end
    if (_T_1004) begin
      if (_T_2529) begin
        _T_2528 <= 16'h1;
      end else begin
        _T_2528 <= _T_2538;
      end
    end
    if (_T_1016) begin
      if (_T_2541) begin
        _T_2540 <= 16'h1;
      end else begin
        _T_2540 <= _T_2550;
      end
    end
    if (_T_1028) begin
      if (_T_2553) begin
        _T_2552 <= 16'h1;
      end else begin
        _T_2552 <= _T_2562;
      end
    end
    if (_T_1040) begin
      if (_T_2565) begin
        _T_2564 <= 16'h1;
      end else begin
        _T_2564 <= _T_2574;
      end
    end
    if (_T_1052) begin
      if (_T_2577) begin
        _T_2576 <= 16'h1;
      end else begin
        _T_2576 <= _T_2586;
      end
    end
    if (_T_1064) begin
      if (_T_2589) begin
        _T_2588 <= 16'h1;
      end else begin
        _T_2588 <= _T_2598;
      end
    end
    if (_T_1076) begin
      if (_T_2601) begin
        _T_2600 <= 16'h1;
      end else begin
        _T_2600 <= _T_2610;
      end
    end
    if (_T_1088) begin
      if (_T_2613) begin
        _T_2612 <= 16'h1;
      end else begin
        _T_2612 <= _T_2622;
      end
    end
    if (_T_1100) begin
      if (_T_2625) begin
        _T_2624 <= 16'h1;
      end else begin
        _T_2624 <= _T_2634;
      end
    end
    if (_T_1112) begin
      if (_T_2637) begin
        _T_2636 <= 16'h1;
      end else begin
        _T_2636 <= _T_2646;
      end
    end
    if (_T_1124) begin
      if (_T_2649) begin
        _T_2648 <= 16'h1;
      end else begin
        _T_2648 <= _T_2658;
      end
    end
    if (_T_1136) begin
      if (_T_2661) begin
        _T_2660 <= 16'h1;
      end else begin
        _T_2660 <= _T_2670;
      end
    end
    if (_T_1148) begin
      if (_T_2673) begin
        _T_2672 <= 16'h1;
      end else begin
        _T_2672 <= _T_2682;
      end
    end
    if (_T_1160) begin
      if (_T_2685) begin
        _T_2684 <= 16'h1;
      end else begin
        _T_2684 <= _T_2694;
      end
    end
    if (_T_1172) begin
      if (_T_2697) begin
        _T_2696 <= 16'h1;
      end else begin
        _T_2696 <= _T_2706;
      end
    end
    if (_T_1184) begin
      if (_T_2709) begin
        _T_2708 <= 16'h1;
      end else begin
        _T_2708 <= _T_2718;
      end
    end
    if (_T_1196) begin
      if (_T_2721) begin
        _T_2720 <= 16'h1;
      end else begin
        _T_2720 <= _T_2730;
      end
    end
    if (_T_1208) begin
      if (_T_2733) begin
        _T_2732 <= 16'h1;
      end else begin
        _T_2732 <= _T_2742;
      end
    end
    if (_T_1220) begin
      if (_T_2745) begin
        _T_2744 <= 16'h1;
      end else begin
        _T_2744 <= _T_2754;
      end
    end
    if (_T_1232) begin
      if (_T_2757) begin
        _T_2756 <= 16'h1;
      end else begin
        _T_2756 <= _T_2766;
      end
    end
    if (_T_1244) begin
      if (_T_2769) begin
        _T_2768 <= 16'h1;
      end else begin
        _T_2768 <= _T_2778;
      end
    end
    if (_T_1256) begin
      if (_T_2781) begin
        _T_2780 <= 16'h1;
      end else begin
        _T_2780 <= _T_2790;
      end
    end
    if (_T_1268) begin
      if (_T_2793) begin
        _T_2792 <= 16'h1;
      end else begin
        _T_2792 <= _T_2802;
      end
    end
    if (_T_1280) begin
      if (_T_2805) begin
        _T_2804 <= 16'h1;
      end else begin
        _T_2804 <= _T_2814;
      end
    end
    if (_T_1292) begin
      if (_T_2817) begin
        _T_2816 <= 16'h1;
      end else begin
        _T_2816 <= _T_2826;
      end
    end
    if (_T_1304) begin
      if (_T_2829) begin
        _T_2828 <= 16'h1;
      end else begin
        _T_2828 <= _T_2838;
      end
    end
    if (_T_1316) begin
      if (_T_2841) begin
        _T_2840 <= 16'h1;
      end else begin
        _T_2840 <= _T_2850;
      end
    end
    if (_T_1328) begin
      if (_T_2853) begin
        _T_2852 <= 16'h1;
      end else begin
        _T_2852 <= _T_2862;
      end
    end
    if (_T_1340) begin
      if (_T_2865) begin
        _T_2864 <= 16'h1;
      end else begin
        _T_2864 <= _T_2874;
      end
    end
    if (_T_1352) begin
      if (_T_2877) begin
        _T_2876 <= 16'h1;
      end else begin
        _T_2876 <= _T_2886;
      end
    end
    if (_T_1364) begin
      if (_T_2889) begin
        _T_2888 <= 16'h1;
      end else begin
        _T_2888 <= _T_2898;
      end
    end
    if (_T_1376) begin
      if (_T_2901) begin
        _T_2900 <= 16'h1;
      end else begin
        _T_2900 <= _T_2910;
      end
    end
    if (_T_1388) begin
      if (_T_2913) begin
        _T_2912 <= 16'h1;
      end else begin
        _T_2912 <= _T_2922;
      end
    end
    if (_T_1400) begin
      if (_T_2925) begin
        _T_2924 <= 16'h1;
      end else begin
        _T_2924 <= _T_2934;
      end
    end
    if (_T_1412) begin
      if (_T_2937) begin
        _T_2936 <= 16'h1;
      end else begin
        _T_2936 <= _T_2946;
      end
    end
    if (_T_1424) begin
      if (_T_2949) begin
        _T_2948 <= 16'h1;
      end else begin
        _T_2948 <= _T_2958;
      end
    end
    if (_T_1436) begin
      if (_T_2961) begin
        _T_2960 <= 16'h1;
      end else begin
        _T_2960 <= _T_2970;
      end
    end
    if (_T_1448) begin
      if (_T_2973) begin
        _T_2972 <= 16'h1;
      end else begin
        _T_2972 <= _T_2982;
      end
    end
    if (_T_1460) begin
      if (_T_2985) begin
        _T_2984 <= 16'h1;
      end else begin
        _T_2984 <= _T_2994;
      end
    end
    if (_T_1472) begin
      if (_T_2997) begin
        _T_2996 <= 16'h1;
      end else begin
        _T_2996 <= _T_3006;
      end
    end
    if (_T_1484) begin
      if (_T_3009) begin
        _T_3008 <= 16'h1;
      end else begin
        _T_3008 <= _T_3018;
      end
    end
    if (_T_1496) begin
      if (_T_3021) begin
        _T_3020 <= 16'h1;
      end else begin
        _T_3020 <= _T_3030;
      end
    end
    if (_T_1508) begin
      if (_T_3033) begin
        _T_3032 <= 16'h1;
      end else begin
        _T_3032 <= _T_3042;
      end
    end
    if (_T_1520) begin
      if (_T_3045) begin
        _T_3044 <= 16'h1;
      end else begin
        _T_3044 <= _T_3054;
      end
    end
    if (_T_1532) begin
      if (_T_3057) begin
        _T_3056 <= 16'h1;
      end else begin
        _T_3056 <= _T_3066;
      end
    end
    if (_T_1544) begin
      if (_T_3069) begin
        _T_3068 <= 16'h1;
      end else begin
        _T_3068 <= _T_3078;
      end
    end
    if (_T_1556) begin
      if (_T_3081) begin
        _T_3080 <= 16'h1;
      end else begin
        _T_3080 <= _T_3090;
      end
    end
    if (_T_1568) begin
      if (_T_3093) begin
        _T_3092 <= 16'h1;
      end else begin
        _T_3092 <= _T_3102;
      end
    end
    if (_T_1580) begin
      if (_T_3105) begin
        _T_3104 <= 16'h1;
      end else begin
        _T_3104 <= _T_3114;
      end
    end
    if (_T_1592) begin
      if (_T_3117) begin
        _T_3116 <= 16'h1;
      end else begin
        _T_3116 <= _T_3126;
      end
    end
    if (_T_1604) begin
      if (_T_3129) begin
        _T_3128 <= 16'h1;
      end else begin
        _T_3128 <= _T_3138;
      end
    end
    if (_T_1616) begin
      if (_T_3141) begin
        _T_3140 <= 16'h1;
      end else begin
        _T_3140 <= _T_3150;
      end
    end
    if (_T_1628) begin
      if (_T_3153) begin
        _T_3152 <= 16'h1;
      end else begin
        _T_3152 <= _T_3162;
      end
    end
    if (_T_1640) begin
      if (_T_3165) begin
        _T_3164 <= 16'h1;
      end else begin
        _T_3164 <= _T_3174;
      end
    end
    if (_T_1652) begin
      if (_T_3177) begin
        _T_3176 <= 16'h1;
      end else begin
        _T_3176 <= _T_3186;
      end
    end
    if (_T_1664) begin
      if (_T_3189) begin
        _T_3188 <= 16'h1;
      end else begin
        _T_3188 <= _T_3198;
      end
    end
    if (_T_1676) begin
      if (_T_3201) begin
        _T_3200 <= 16'h1;
      end else begin
        _T_3200 <= _T_3210;
      end
    end
    if (_T_1688) begin
      if (_T_3213) begin
        _T_3212 <= 16'h1;
      end else begin
        _T_3212 <= _T_3222;
      end
    end
    if (_T_1700) begin
      if (_T_3225) begin
        _T_3224 <= 16'h1;
      end else begin
        _T_3224 <= _T_3234;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_528 & _T_43) begin
          $fwrite(32'h80000002,"Assertion failed: DriveInterruptType.%d not supported yet\n    at Interrupts.scala:195 assert(false.B, \"DriveInterruptType.%%d not supported yet\", drive_interrupt_type)\n",_T_30);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_528 & _T_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_548 & _T_43) begin
          $fwrite(32'h80000002,"Assertion failed: DriveInterruptType.%d not supported yet\n    at Interrupts.scala:222 assert(false.B, \"DriveInterruptType.%%d not supported yet\", drive_interrupt_type)\n",_T_44);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_548 & _T_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
