//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_28(
  output        _EVAL,
  input  [3:0]  _EVAL_0,
  output [7:0]  _EVAL_1,
  input         _EVAL_2,
  output [2:0]  _EVAL_3,
  output        _EVAL_4,
  input  [3:0]  _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  output [2:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input  [1:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [7:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  output [3:0]  _EVAL_21,
  output [31:0] _EVAL_22,
  output [1:0]  _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output        _EVAL_26,
  input  [2:0]  _EVAL_27,
  output        _EVAL_28,
  input  [3:0]  _EVAL_29,
  input         _EVAL_30,
  input  [2:0]  _EVAL_31,
  output        _EVAL_32,
  input  [30:0] _EVAL_33,
  input         _EVAL_34,
  input  [3:0]  _EVAL_35,
  output        _EVAL_36,
  input  [3:0]  _EVAL_37,
  output [3:0]  _EVAL_38,
  output [30:0] _EVAL_39,
  input  [2:0]  _EVAL_40,
  input  [2:0]  _EVAL_41,
  output [30:0] _EVAL_42,
  input         _EVAL_43,
  input  [1:0]  _EVAL_44,
  output [1:0]  _EVAL_45,
  input         _EVAL_46,
  input  [7:0]  _EVAL_47,
  output        _EVAL_48,
  output [1:0]  _EVAL_49,
  output [3:0]  _EVAL_50,
  input  [10:0] _EVAL_51,
  output [3:0]  _EVAL_52,
  input  [31:0] _EVAL_53,
  output        _EVAL_54,
  output [10:0] _EVAL_55,
  output        _EVAL_56,
  output [7:0]  _EVAL_57,
  input         _EVAL_58,
  output        _EVAL_59,
  input  [10:0] _EVAL_60,
  input  [30:0] _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  input  [31:0] _EVAL_64,
  input         _EVAL_65,
  output [31:0] _EVAL_66,
  output        _EVAL_67,
  output [2:0]  _EVAL_68,
  input  [3:0]  _EVAL_69,
  output [3:0]  _EVAL_70,
  output [3:0]  _EVAL_71,
  output [3:0]  _EVAL_72,
  output [2:0]  _EVAL_73,
  output [3:0]  _EVAL_74,
  output [3:0]  _EVAL_75,
  output        _EVAL_76,
  output [10:0] _EVAL_77,
  output [1:0]  _EVAL_78
);
  wire  Queue_15__EVAL;
  wire  Queue_15__EVAL_0;
  wire  Queue_15__EVAL_1;
  wire  Queue_15__EVAL_2;
  wire  Queue_15__EVAL_3;
  wire [10:0] Queue_15__EVAL_4;
  wire  Queue_15__EVAL_5;
  wire [10:0] Queue_15__EVAL_6;
  wire  Queue_3__EVAL;
  wire  Queue_3__EVAL_0;
  wire  Queue_3__EVAL_1;
  wire [10:0] Queue_3__EVAL_2;
  wire [10:0] Queue_3__EVAL_3;
  wire  Queue_3__EVAL_4;
  wire  Queue_3__EVAL_5;
  wire  Queue_3__EVAL_6;
  wire  Queue__EVAL;
  wire  Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire [10:0] Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire [10:0] Queue__EVAL_6;
  wire  Queue_6__EVAL;
  wire  Queue_6__EVAL_0;
  wire  Queue_6__EVAL_1;
  wire [10:0] Queue_6__EVAL_2;
  wire [10:0] Queue_6__EVAL_3;
  wire  Queue_6__EVAL_4;
  wire  Queue_6__EVAL_5;
  wire  Queue_6__EVAL_6;
  wire  Queue_13__EVAL;
  wire  Queue_13__EVAL_0;
  wire  Queue_13__EVAL_1;
  wire [10:0] Queue_13__EVAL_2;
  wire [10:0] Queue_13__EVAL_3;
  wire  Queue_13__EVAL_4;
  wire  Queue_13__EVAL_5;
  wire  Queue_13__EVAL_6;
  wire  Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire [10:0] Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire [10:0] Queue_1__EVAL_6;
  wire  Queue_11__EVAL;
  wire  Queue_11__EVAL_0;
  wire  Queue_11__EVAL_1;
  wire [10:0] Queue_11__EVAL_2;
  wire [10:0] Queue_11__EVAL_3;
  wire  Queue_11__EVAL_4;
  wire  Queue_11__EVAL_5;
  wire  Queue_11__EVAL_6;
  wire  Queue_9__EVAL;
  wire  Queue_9__EVAL_0;
  wire  Queue_9__EVAL_1;
  wire  Queue_9__EVAL_2;
  wire  Queue_9__EVAL_3;
  wire [10:0] Queue_9__EVAL_4;
  wire  Queue_9__EVAL_5;
  wire [10:0] Queue_9__EVAL_6;
  wire  Queue_2__EVAL;
  wire  Queue_2__EVAL_0;
  wire  Queue_2__EVAL_1;
  wire [10:0] Queue_2__EVAL_2;
  wire  Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire [10:0] Queue_2__EVAL_5;
  wire  Queue_2__EVAL_6;
  wire  Queue_5__EVAL;
  wire  Queue_5__EVAL_0;
  wire  Queue_5__EVAL_1;
  wire [10:0] Queue_5__EVAL_2;
  wire [10:0] Queue_5__EVAL_3;
  wire  Queue_5__EVAL_4;
  wire  Queue_5__EVAL_5;
  wire  Queue_5__EVAL_6;
  wire  Queue_8__EVAL;
  wire  Queue_8__EVAL_0;
  wire  Queue_8__EVAL_1;
  wire  Queue_8__EVAL_2;
  wire  Queue_8__EVAL_3;
  wire [10:0] Queue_8__EVAL_4;
  wire  Queue_8__EVAL_5;
  wire [10:0] Queue_8__EVAL_6;
  wire  Queue_12__EVAL;
  wire  Queue_12__EVAL_0;
  wire  Queue_12__EVAL_1;
  wire [10:0] Queue_12__EVAL_2;
  wire [10:0] Queue_12__EVAL_3;
  wire  Queue_12__EVAL_4;
  wire  Queue_12__EVAL_5;
  wire  Queue_12__EVAL_6;
  wire  Queue_4__EVAL;
  wire  Queue_4__EVAL_0;
  wire  Queue_4__EVAL_1;
  wire [10:0] Queue_4__EVAL_2;
  wire [10:0] Queue_4__EVAL_3;
  wire  Queue_4__EVAL_4;
  wire  Queue_4__EVAL_5;
  wire  Queue_4__EVAL_6;
  wire  Queue_14__EVAL;
  wire  Queue_14__EVAL_0;
  wire  Queue_14__EVAL_1;
  wire [10:0] Queue_14__EVAL_2;
  wire [10:0] Queue_14__EVAL_3;
  wire  Queue_14__EVAL_4;
  wire  Queue_14__EVAL_5;
  wire  Queue_14__EVAL_6;
  wire  Queue_7__EVAL;
  wire  Queue_7__EVAL_0;
  wire  Queue_7__EVAL_1;
  wire  Queue_7__EVAL_2;
  wire  Queue_7__EVAL_3;
  wire [10:0] Queue_7__EVAL_4;
  wire  Queue_7__EVAL_5;
  wire [10:0] Queue_7__EVAL_6;
  wire  Queue_10__EVAL;
  wire  Queue_10__EVAL_0;
  wire  Queue_10__EVAL_1;
  wire [10:0] Queue_10__EVAL_2;
  wire  Queue_10__EVAL_3;
  wire  Queue_10__EVAL_4;
  wire [10:0] Queue_10__EVAL_5;
  wire  Queue_10__EVAL_6;
  wire  _EVAL_269;
  wire  _EVAL_129;
  wire  _EVAL_240;
  wire  _EVAL_103;
  wire  _EVAL_164;
  wire  _EVAL_263;
  wire  _EVAL_213;
  wire  _EVAL_257;
  wire  _EVAL_204;
  wire  _EVAL_202;
  wire  _EVAL_195;
  wire  _EVAL_212;
  wire  _EVAL_153;
  wire  _EVAL_180;
  wire  _EVAL_225;
  wire  _EVAL_231;
  wire  _EVAL_186;
  wire  _EVAL_168;
  wire  _EVAL_185;
  wire  _EVAL_182;
  wire  _EVAL_170;
  wire  _EVAL_142;
  wire  _EVAL_245;
  wire  _EVAL_100;
  wire  _EVAL_94;
  wire  _EVAL_84;
  wire  _EVAL_179;
  wire  _EVAL_205;
  wire  _EVAL_172;
  wire  _EVAL_159;
  wire  _EVAL_206;
  wire  _EVAL_115;
  wire  _EVAL_117;
  wire  _EVAL_266;
  wire  _EVAL_260;
  wire  _EVAL_194;
  wire  _EVAL_224;
  wire  _EVAL_96;
  wire  _EVAL_259;
  wire  _EVAL_251;
  wire  _EVAL_219;
  wire  _EVAL_89;
  wire  _EVAL_101;
  wire  _EVAL_141;
  wire  _EVAL_145;
  wire [15:0] _EVAL_208;
  wire  _EVAL_169;
  wire  _EVAL_230;
  wire [15:0] _EVAL_110;
  wire  _EVAL_250;
  wire  _EVAL_97;
  wire [15:0] _EVAL_234;
  wire  _EVAL_121;
  wire [10:0] _EVAL_166;
  wire [10:0] _EVAL_178;
  wire [10:0] _EVAL_244;
  wire [10:0] _EVAL_241;
  wire [10:0] _EVAL_150;
  wire  _EVAL_134;
  wire  _EVAL_183;
  wire [10:0] _EVAL_126;
  wire [10:0] _EVAL_132;
  wire [10:0] _EVAL_181;
  wire [10:0] _EVAL_270;
  wire [10:0] _EVAL_220;
  wire [10:0] _EVAL_239;
  wire [10:0] _EVAL_154;
  wire [10:0] _EVAL_207;
  wire [10:0] _EVAL_198;
  wire [10:0] _EVAL_151;
  wire  _EVAL_80;
  wire  _EVAL_254;
  wire [10:0] _EVAL_156;
  wire [10:0] _EVAL_265;
  wire [10:0] _EVAL_221;
  wire [10:0] _EVAL_255;
  wire [10:0] _EVAL_146;
  wire [10:0] _EVAL_167;
  wire [10:0] _EVAL_165;
  wire [10:0] _EVAL_268;
  wire [10:0] _EVAL_138;
  wire [10:0] _EVAL_247;
  wire [10:0] _EVAL_106;
  wire [10:0] _EVAL_201;
  wire [10:0] _EVAL_92;
  wire [10:0] _EVAL_218;
  wire [10:0] _EVAL_229;
  wire [10:0] _EVAL_99;
  wire [10:0] _EVAL_114;
  wire [10:0] _EVAL_139;
  wire [15:0] _EVAL_226;
  wire  _EVAL_249;
  wire [10:0] _EVAL_95;
  wire [10:0] _EVAL_187;
  wire [10:0] _EVAL_203;
  wire  _EVAL_144;
  wire  _EVAL_124;
  wire  _EVAL_123;
  wire  _EVAL_261;
  wire  _EVAL_258;
  wire  _EVAL_122;
  wire [10:0] _EVAL_211;
  wire [10:0] _EVAL_191;
  wire  _EVAL_171;
  wire  _EVAL_111;
  wire  _EVAL_87;
  wire  _EVAL_112;
  wire  _EVAL_192;
  wire  _EVAL_256;
  wire [10:0] _EVAL_217;
  wire [10:0] _EVAL_238;
  wire  _EVAL_242;
  wire  _EVAL_130;
  wire  _EVAL_160;
  wire [10:0] _EVAL_158;
  wire  _EVAL_119;
  wire  _EVAL_199;
  wire  _EVAL_91;
  wire [10:0] _EVAL_90;
  wire  _EVAL_125;
  wire  _EVAL_210;
  wire  _EVAL_140;
  wire  _EVAL_135;
  wire [10:0] _EVAL_128;
  wire  _EVAL_85;
  wire  _EVAL_107;
  wire  _EVAL_200;
  wire  _EVAL_223;
  wire  _EVAL_161;
  wire  _EVAL_216;
  wire  _EVAL_196;
  wire [10:0] _EVAL_86;
  wire  _EVAL_148;
  wire  _EVAL_131;
  wire  _EVAL_79;
  wire  _EVAL_232;
  wire  _EVAL_109;
  wire  _EVAL_93;
  SiFive__EVAL_25 Queue_15 (
    ._EVAL(Queue_15__EVAL),
    ._EVAL_0(Queue_15__EVAL_0),
    ._EVAL_1(Queue_15__EVAL_1),
    ._EVAL_2(Queue_15__EVAL_2),
    ._EVAL_3(Queue_15__EVAL_3),
    ._EVAL_4(Queue_15__EVAL_4),
    ._EVAL_5(Queue_15__EVAL_5),
    ._EVAL_6(Queue_15__EVAL_6)
  );
  SiFive__EVAL_27 Queue_3 (
    ._EVAL(Queue_3__EVAL),
    ._EVAL_0(Queue_3__EVAL_0),
    ._EVAL_1(Queue_3__EVAL_1),
    ._EVAL_2(Queue_3__EVAL_2),
    ._EVAL_3(Queue_3__EVAL_3),
    ._EVAL_4(Queue_3__EVAL_4),
    ._EVAL_5(Queue_3__EVAL_5),
    ._EVAL_6(Queue_3__EVAL_6)
  );
  SiFive__EVAL_25 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6)
  );
  SiFive__EVAL_27 Queue_6 (
    ._EVAL(Queue_6__EVAL),
    ._EVAL_0(Queue_6__EVAL_0),
    ._EVAL_1(Queue_6__EVAL_1),
    ._EVAL_2(Queue_6__EVAL_2),
    ._EVAL_3(Queue_6__EVAL_3),
    ._EVAL_4(Queue_6__EVAL_4),
    ._EVAL_5(Queue_6__EVAL_5),
    ._EVAL_6(Queue_6__EVAL_6)
  );
  SiFive__EVAL_27 Queue_13 (
    ._EVAL(Queue_13__EVAL),
    ._EVAL_0(Queue_13__EVAL_0),
    ._EVAL_1(Queue_13__EVAL_1),
    ._EVAL_2(Queue_13__EVAL_2),
    ._EVAL_3(Queue_13__EVAL_3),
    ._EVAL_4(Queue_13__EVAL_4),
    ._EVAL_5(Queue_13__EVAL_5),
    ._EVAL_6(Queue_13__EVAL_6)
  );
  SiFive__EVAL_25 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6)
  );
  SiFive__EVAL_27 Queue_11 (
    ._EVAL(Queue_11__EVAL),
    ._EVAL_0(Queue_11__EVAL_0),
    ._EVAL_1(Queue_11__EVAL_1),
    ._EVAL_2(Queue_11__EVAL_2),
    ._EVAL_3(Queue_11__EVAL_3),
    ._EVAL_4(Queue_11__EVAL_4),
    ._EVAL_5(Queue_11__EVAL_5),
    ._EVAL_6(Queue_11__EVAL_6)
  );
  SiFive__EVAL_25 Queue_9 (
    ._EVAL(Queue_9__EVAL),
    ._EVAL_0(Queue_9__EVAL_0),
    ._EVAL_1(Queue_9__EVAL_1),
    ._EVAL_2(Queue_9__EVAL_2),
    ._EVAL_3(Queue_9__EVAL_3),
    ._EVAL_4(Queue_9__EVAL_4),
    ._EVAL_5(Queue_9__EVAL_5),
    ._EVAL_6(Queue_9__EVAL_6)
  );
  SiFive__EVAL_26 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6)
  );
  SiFive__EVAL_27 Queue_5 (
    ._EVAL(Queue_5__EVAL),
    ._EVAL_0(Queue_5__EVAL_0),
    ._EVAL_1(Queue_5__EVAL_1),
    ._EVAL_2(Queue_5__EVAL_2),
    ._EVAL_3(Queue_5__EVAL_3),
    ._EVAL_4(Queue_5__EVAL_4),
    ._EVAL_5(Queue_5__EVAL_5),
    ._EVAL_6(Queue_5__EVAL_6)
  );
  SiFive__EVAL_25 Queue_8 (
    ._EVAL(Queue_8__EVAL),
    ._EVAL_0(Queue_8__EVAL_0),
    ._EVAL_1(Queue_8__EVAL_1),
    ._EVAL_2(Queue_8__EVAL_2),
    ._EVAL_3(Queue_8__EVAL_3),
    ._EVAL_4(Queue_8__EVAL_4),
    ._EVAL_5(Queue_8__EVAL_5),
    ._EVAL_6(Queue_8__EVAL_6)
  );
  SiFive__EVAL_27 Queue_12 (
    ._EVAL(Queue_12__EVAL),
    ._EVAL_0(Queue_12__EVAL_0),
    ._EVAL_1(Queue_12__EVAL_1),
    ._EVAL_2(Queue_12__EVAL_2),
    ._EVAL_3(Queue_12__EVAL_3),
    ._EVAL_4(Queue_12__EVAL_4),
    ._EVAL_5(Queue_12__EVAL_5),
    ._EVAL_6(Queue_12__EVAL_6)
  );
  SiFive__EVAL_27 Queue_4 (
    ._EVAL(Queue_4__EVAL),
    ._EVAL_0(Queue_4__EVAL_0),
    ._EVAL_1(Queue_4__EVAL_1),
    ._EVAL_2(Queue_4__EVAL_2),
    ._EVAL_3(Queue_4__EVAL_3),
    ._EVAL_4(Queue_4__EVAL_4),
    ._EVAL_5(Queue_4__EVAL_5),
    ._EVAL_6(Queue_4__EVAL_6)
  );
  SiFive__EVAL_27 Queue_14 (
    ._EVAL(Queue_14__EVAL),
    ._EVAL_0(Queue_14__EVAL_0),
    ._EVAL_1(Queue_14__EVAL_1),
    ._EVAL_2(Queue_14__EVAL_2),
    ._EVAL_3(Queue_14__EVAL_3),
    ._EVAL_4(Queue_14__EVAL_4),
    ._EVAL_5(Queue_14__EVAL_5),
    ._EVAL_6(Queue_14__EVAL_6)
  );
  SiFive__EVAL_25 Queue_7 (
    ._EVAL(Queue_7__EVAL),
    ._EVAL_0(Queue_7__EVAL_0),
    ._EVAL_1(Queue_7__EVAL_1),
    ._EVAL_2(Queue_7__EVAL_2),
    ._EVAL_3(Queue_7__EVAL_3),
    ._EVAL_4(Queue_7__EVAL_4),
    ._EVAL_5(Queue_7__EVAL_5),
    ._EVAL_6(Queue_7__EVAL_6)
  );
  SiFive__EVAL_26 Queue_10 (
    ._EVAL(Queue_10__EVAL),
    ._EVAL_0(Queue_10__EVAL_0),
    ._EVAL_1(Queue_10__EVAL_1),
    ._EVAL_2(Queue_10__EVAL_2),
    ._EVAL_3(Queue_10__EVAL_3),
    ._EVAL_4(Queue_10__EVAL_4),
    ._EVAL_5(Queue_10__EVAL_5),
    ._EVAL_6(Queue_10__EVAL_6)
  );
  assign _EVAL_269 = Queue_13__EVAL_4;
  assign _EVAL_129 = Queue_2__EVAL_3;
  assign _EVAL_240 = Queue_1__EVAL_1;
  assign _EVAL_103 = Queue__EVAL_1;
  assign _EVAL_164 = 4'h1 == _EVAL_69 ? _EVAL_240 : _EVAL_103;
  assign _EVAL_263 = 4'h2 == _EVAL_69 ? _EVAL_129 : _EVAL_164;
  assign _EVAL_213 = Queue_7__EVAL_1;
  assign _EVAL_257 = Queue_6__EVAL_4;
  assign _EVAL_204 = Queue_5__EVAL_4;
  assign _EVAL_202 = Queue_4__EVAL_4;
  assign _EVAL_195 = Queue_3__EVAL_4;
  assign _EVAL_212 = 4'h3 == _EVAL_69 ? _EVAL_195 : _EVAL_263;
  assign _EVAL_153 = 4'h4 == _EVAL_69 ? _EVAL_202 : _EVAL_212;
  assign _EVAL_180 = 4'h5 == _EVAL_69 ? _EVAL_204 : _EVAL_153;
  assign _EVAL_225 = 4'h6 == _EVAL_69 ? _EVAL_257 : _EVAL_180;
  assign _EVAL_231 = 4'h7 == _EVAL_69 ? _EVAL_213 : _EVAL_225;
  assign _EVAL_186 = 4'h8 == _EVAL_69 ? 1'h0 : _EVAL_231;
  assign _EVAL_168 = 4'h9 == _EVAL_69 ? 1'h0 : _EVAL_186;
  assign _EVAL_185 = 4'ha == _EVAL_69 ? 1'h0 : _EVAL_168;
  assign _EVAL_182 = 4'hb == _EVAL_69 ? 1'h0 : _EVAL_185;
  assign _EVAL_170 = 4'hc == _EVAL_69 ? 1'h0 : _EVAL_182;
  assign _EVAL_142 = 4'hd == _EVAL_69 ? 1'h0 : _EVAL_170;
  assign _EVAL_245 = 4'he == _EVAL_69 ? 1'h0 : _EVAL_142;
  assign _EVAL_100 = 4'hf == _EVAL_69 ? 1'h0 : _EVAL_245;
  assign _EVAL_94 = Queue_15__EVAL_1;
  assign _EVAL_84 = Queue_14__EVAL_4;
  assign _EVAL_179 = Queue_12__EVAL_4;
  assign _EVAL_205 = Queue_11__EVAL_4;
  assign _EVAL_172 = Queue_10__EVAL_3;
  assign _EVAL_159 = Queue_9__EVAL_1;
  assign _EVAL_206 = Queue_8__EVAL_1;
  assign _EVAL_115 = 4'h1 == _EVAL_18 ? _EVAL_159 : _EVAL_206;
  assign _EVAL_117 = 4'h2 == _EVAL_18 ? _EVAL_172 : _EVAL_115;
  assign _EVAL_266 = 4'h3 == _EVAL_18 ? _EVAL_205 : _EVAL_117;
  assign _EVAL_260 = 4'h4 == _EVAL_18 ? _EVAL_179 : _EVAL_266;
  assign _EVAL_194 = 4'h5 == _EVAL_18 ? _EVAL_269 : _EVAL_260;
  assign _EVAL_224 = 4'h6 == _EVAL_18 ? _EVAL_84 : _EVAL_194;
  assign _EVAL_96 = 4'h7 == _EVAL_18 ? _EVAL_94 : _EVAL_224;
  assign _EVAL_259 = 4'h8 == _EVAL_18 ? 1'h0 : _EVAL_96;
  assign _EVAL_251 = 4'h9 == _EVAL_18 ? 1'h0 : _EVAL_259;
  assign _EVAL_219 = 4'ha == _EVAL_18 ? 1'h0 : _EVAL_251;
  assign _EVAL_89 = 4'hb == _EVAL_18 ? 1'h0 : _EVAL_219;
  assign _EVAL_101 = 4'hc == _EVAL_18 ? 1'h0 : _EVAL_89;
  assign _EVAL_141 = 4'hd == _EVAL_18 ? 1'h0 : _EVAL_101;
  assign _EVAL_145 = 4'he == _EVAL_18 ? 1'h0 : _EVAL_141;
  assign _EVAL_208 = 16'h1 << _EVAL_18;
  assign _EVAL_169 = _EVAL_208[4];
  assign _EVAL_230 = _EVAL_17 & _EVAL_62;
  assign _EVAL_110 = 16'h1 << _EVAL_35;
  assign _EVAL_250 = _EVAL_110[6];
  assign _EVAL_97 = _EVAL_230 & _EVAL_250;
  assign _EVAL_234 = 16'h1 << _EVAL_69;
  assign _EVAL_121 = _EVAL_234[0];
  assign _EVAL_166 = Queue_10__EVAL_2;
  assign _EVAL_178 = Queue_9__EVAL_6;
  assign _EVAL_244 = Queue_8__EVAL_6;
  assign _EVAL_241 = 4'h1 == _EVAL_29 ? _EVAL_178 : _EVAL_244;
  assign _EVAL_150 = 4'h2 == _EVAL_29 ? _EVAL_166 : _EVAL_241;
  assign _EVAL_134 = _EVAL_30 & _EVAL_6;
  assign _EVAL_183 = _EVAL_234[4];
  assign _EVAL_126 = Queue_15__EVAL_6;
  assign _EVAL_132 = Queue_14__EVAL_3;
  assign _EVAL_181 = Queue_13__EVAL_3;
  assign _EVAL_270 = Queue_12__EVAL_3;
  assign _EVAL_220 = Queue_11__EVAL_3;
  assign _EVAL_239 = 4'h3 == _EVAL_29 ? _EVAL_220 : _EVAL_150;
  assign _EVAL_154 = 4'h4 == _EVAL_29 ? _EVAL_270 : _EVAL_239;
  assign _EVAL_207 = 4'h5 == _EVAL_29 ? _EVAL_181 : _EVAL_154;
  assign _EVAL_198 = 4'h6 == _EVAL_29 ? _EVAL_132 : _EVAL_207;
  assign _EVAL_151 = 4'h7 == _EVAL_29 ? _EVAL_126 : _EVAL_198;
  assign _EVAL_80 = _EVAL_110[7];
  assign _EVAL_254 = _EVAL_230 & _EVAL_80;
  assign _EVAL_156 = Queue_7__EVAL_6;
  assign _EVAL_265 = Queue_6__EVAL_3;
  assign _EVAL_221 = Queue_5__EVAL_3;
  assign _EVAL_255 = Queue_4__EVAL_3;
  assign _EVAL_146 = Queue_3__EVAL_3;
  assign _EVAL_167 = Queue_2__EVAL_2;
  assign _EVAL_165 = Queue_1__EVAL_6;
  assign _EVAL_268 = Queue__EVAL_6;
  assign _EVAL_138 = 4'h1 == _EVAL_35 ? _EVAL_165 : _EVAL_268;
  assign _EVAL_247 = 4'h2 == _EVAL_35 ? _EVAL_167 : _EVAL_138;
  assign _EVAL_106 = 4'h3 == _EVAL_35 ? _EVAL_146 : _EVAL_247;
  assign _EVAL_201 = 4'h4 == _EVAL_35 ? _EVAL_255 : _EVAL_106;
  assign _EVAL_92 = 4'h5 == _EVAL_35 ? _EVAL_221 : _EVAL_201;
  assign _EVAL_218 = 4'h6 == _EVAL_35 ? _EVAL_265 : _EVAL_92;
  assign _EVAL_229 = 4'h7 == _EVAL_35 ? _EVAL_156 : _EVAL_218;
  assign _EVAL_99 = 4'h8 == _EVAL_35 ? 11'h0 : _EVAL_229;
  assign _EVAL_114 = 4'h9 == _EVAL_35 ? 11'h0 : _EVAL_99;
  assign _EVAL_139 = 4'ha == _EVAL_35 ? 11'h0 : _EVAL_114;
  assign _EVAL_226 = 16'h1 << _EVAL_29;
  assign _EVAL_249 = _EVAL_226[2];
  assign _EVAL_95 = 4'hb == _EVAL_35 ? 11'h0 : _EVAL_139;
  assign _EVAL_187 = 4'hc == _EVAL_35 ? 11'h0 : _EVAL_95;
  assign _EVAL_203 = 4'hd == _EVAL_35 ? 11'h0 : _EVAL_187;
  assign _EVAL_144 = _EVAL_226[4];
  assign _EVAL_124 = _EVAL_2 & _EVAL_12;
  assign _EVAL_123 = _EVAL_208[6];
  assign _EVAL_261 = _EVAL_226[6];
  assign _EVAL_258 = _EVAL_110[1];
  assign _EVAL_122 = _EVAL_230 & _EVAL_258;
  assign _EVAL_211 = 4'h8 == _EVAL_29 ? 11'h0 : _EVAL_151;
  assign _EVAL_191 = 4'h9 == _EVAL_29 ? 11'h0 : _EVAL_211;
  assign _EVAL_171 = _EVAL_234[2];
  assign _EVAL_111 = 4'hf == _EVAL_18 ? 1'h0 : _EVAL_145;
  assign _EVAL_87 = _EVAL_110[2];
  assign _EVAL_112 = _EVAL_230 & _EVAL_87;
  assign _EVAL_192 = _EVAL_226[5];
  assign _EVAL_256 = _EVAL_226[3];
  assign _EVAL_217 = 4'ha == _EVAL_29 ? 11'h0 : _EVAL_191;
  assign _EVAL_238 = 4'hb == _EVAL_29 ? 11'h0 : _EVAL_217;
  assign _EVAL_242 = _EVAL_110[5];
  assign _EVAL_130 = _EVAL_230 & _EVAL_242;
  assign _EVAL_160 = _EVAL_208[3];
  assign _EVAL_158 = 4'hc == _EVAL_29 ? 11'h0 : _EVAL_238;
  assign _EVAL_119 = _EVAL_110[0];
  assign _EVAL_199 = _EVAL_230 & _EVAL_119;
  assign _EVAL_91 = _EVAL_234[6];
  assign _EVAL_90 = 4'hd == _EVAL_29 ? 11'h0 : _EVAL_158;
  assign _EVAL_125 = _EVAL_234[5];
  assign _EVAL_210 = _EVAL_226[1];
  assign _EVAL_140 = _EVAL_208[2];
  assign _EVAL_135 = _EVAL_208[0];
  assign _EVAL_128 = 4'he == _EVAL_29 ? 11'h0 : _EVAL_90;
  assign _EVAL_85 = _EVAL_226[7];
  assign _EVAL_107 = _EVAL_208[5];
  assign _EVAL_200 = _EVAL_234[1];
  assign _EVAL_223 = _EVAL_63 & _EVAL_25;
  assign _EVAL_161 = _EVAL_234[3];
  assign _EVAL_216 = _EVAL_110[4];
  assign _EVAL_196 = _EVAL_110[3];
  assign _EVAL_86 = 4'he == _EVAL_35 ? 11'h0 : _EVAL_203;
  assign _EVAL_148 = _EVAL_208[7];
  assign _EVAL_131 = _EVAL_230 & _EVAL_216;
  assign _EVAL_79 = _EVAL_226[0];
  assign _EVAL_232 = _EVAL_230 & _EVAL_196;
  assign _EVAL_109 = _EVAL_234[7];
  assign _EVAL_93 = _EVAL_208[1];
  assign _EVAL_22 = _EVAL_64;
  assign Queue_9__EVAL_5 = _EVAL_124 & _EVAL_93;
  assign Queue_3__EVAL_1 = _EVAL_34;
  assign Queue_7__EVAL_3 = _EVAL_46;
  assign Queue_1__EVAL_3 = _EVAL_46;
  assign Queue_15__EVAL_2 = _EVAL_134 & _EVAL_85;
  assign Queue_10__EVAL = _EVAL_124 & _EVAL_140;
  assign Queue_2__EVAL_4 = _EVAL_112 & _EVAL_24;
  assign Queue_15__EVAL_3 = _EVAL_46;
  assign Queue_5__EVAL_2 = _EVAL_60;
  assign Queue_3__EVAL_5 = _EVAL_46;
  assign Queue_13__EVAL_2 = _EVAL_51;
  assign Queue_5__EVAL = _EVAL_130 & _EVAL_24;
  assign Queue_13__EVAL_1 = _EVAL_34;
  assign Queue_13__EVAL_0 = _EVAL_124 & _EVAL_107;
  assign Queue_11__EVAL_1 = _EVAL_34;
  assign _EVAL_52 = _EVAL_5;
  assign _EVAL_71 = _EVAL_69;
  assign _EVAL_3 = _EVAL_40;
  assign _EVAL_39 = _EVAL_61;
  assign Queue_14__EVAL_5 = _EVAL_46;
  assign Queue__EVAL = _EVAL_34;
  assign _EVAL_26 = _EVAL_65;
  assign Queue_1__EVAL_5 = _EVAL_223 & _EVAL_200;
  assign _EVAL_21 = _EVAL_14;
  assign Queue_7__EVAL_5 = _EVAL_223 & _EVAL_109;
  assign Queue_8__EVAL_3 = _EVAL_46;
  assign Queue_10__EVAL_1 = _EVAL_46;
  assign _EVAL_42 = _EVAL_33;
  assign _EVAL_49 = _EVAL_11;
  assign Queue_4__EVAL_2 = _EVAL_60;
  assign Queue_14__EVAL = _EVAL_134 & _EVAL_261;
  assign Queue_4__EVAL_1 = _EVAL_34;
  assign _EVAL_10 = _EVAL_41;
  assign _EVAL_76 = _EVAL_62;
  assign Queue_14__EVAL_2 = _EVAL_51;
  assign _EVAL_48 = _EVAL_9;
  assign Queue_14__EVAL_1 = _EVAL_34;
  assign Queue__EVAL_3 = _EVAL_46;
  assign Queue_9__EVAL_2 = _EVAL_134 & _EVAL_210;
  assign _EVAL_45 = _EVAL_8;
  assign Queue_13__EVAL = _EVAL_134 & _EVAL_192;
  assign Queue_2__EVAL_5 = _EVAL_60;
  assign Queue_12__EVAL_1 = _EVAL_34;
  assign _EVAL_32 = _EVAL_17;
  assign _EVAL_66 = _EVAL_53;
  assign Queue_11__EVAL_0 = _EVAL_124 & _EVAL_160;
  assign Queue_14__EVAL_0 = _EVAL_124 & _EVAL_123;
  assign Queue__EVAL_4 = _EVAL_60;
  assign Queue_15__EVAL = _EVAL_34;
  assign Queue_6__EVAL = _EVAL_97 & _EVAL_24;
  assign Queue_5__EVAL_5 = _EVAL_46;
  assign _EVAL_67 = _EVAL_30;
  assign Queue__EVAL_2 = _EVAL_199 & _EVAL_24;
  assign Queue_9__EVAL_4 = _EVAL_51;
  assign _EVAL_28 = _EVAL_43;
  assign _EVAL_50 = _EVAL_35;
  assign Queue_3__EVAL_0 = _EVAL_223 & _EVAL_161;
  assign Queue_2__EVAL_1 = _EVAL_46;
  assign Queue_6__EVAL_5 = _EVAL_46;
  assign Queue_3__EVAL = _EVAL_232 & _EVAL_24;
  assign Queue_12__EVAL_2 = _EVAL_51;
  assign Queue_11__EVAL_2 = _EVAL_51;
  assign Queue_10__EVAL_0 = _EVAL_34;
  assign Queue_8__EVAL_5 = _EVAL_124 & _EVAL_135;
  assign Queue_5__EVAL_0 = _EVAL_223 & _EVAL_125;
  assign Queue_9__EVAL_3 = _EVAL_46;
  assign _EVAL_78 = _EVAL_13;
  assign _EVAL_59 = _EVAL_2 & _EVAL_111;
  assign Queue_1__EVAL_4 = _EVAL_60;
  assign _EVAL_36 = _EVAL_58;
  assign Queue_9__EVAL = _EVAL_34;
  assign _EVAL_73 = _EVAL_27;
  assign Queue_5__EVAL_1 = _EVAL_34;
  assign _EVAL_75 = _EVAL_16;
  assign _EVAL_77 = 4'hf == _EVAL_29 ? 11'h0 : _EVAL_128;
  assign _EVAL_4 = _EVAL_6;
  assign _EVAL_56 = _EVAL_24;
  assign _EVAL_68 = _EVAL_31;
  assign Queue_4__EVAL_0 = _EVAL_223 & _EVAL_183;
  assign Queue_12__EVAL = _EVAL_134 & _EVAL_144;
  assign Queue_6__EVAL_2 = _EVAL_60;
  assign Queue_7__EVAL_2 = _EVAL_254 & _EVAL_24;
  assign Queue_1__EVAL_2 = _EVAL_122 & _EVAL_24;
  assign _EVAL = _EVAL_12 & _EVAL_111;
  assign _EVAL_7 = _EVAL_19;
  assign Queue_12__EVAL_0 = _EVAL_124 & _EVAL_169;
  assign Queue_3__EVAL_2 = _EVAL_60;
  assign Queue_7__EVAL = _EVAL_34;
  assign Queue_1__EVAL = _EVAL_34;
  assign _EVAL_54 = _EVAL_25 & _EVAL_100;
  assign Queue_4__EVAL_5 = _EVAL_46;
  assign _EVAL_55 = 4'hf == _EVAL_35 ? 11'h0 : _EVAL_86;
  assign Queue_6__EVAL_1 = _EVAL_34;
  assign Queue_8__EVAL_2 = _EVAL_134 & _EVAL_79;
  assign Queue_15__EVAL_5 = _EVAL_124 & _EVAL_148;
  assign Queue_8__EVAL_4 = _EVAL_51;
  assign Queue_6__EVAL_0 = _EVAL_223 & _EVAL_91;
  assign _EVAL_57 = _EVAL_47;
  assign _EVAL_23 = _EVAL_44;
  assign Queue__EVAL_5 = _EVAL_223 & _EVAL_121;
  assign Queue_11__EVAL_5 = _EVAL_46;
  assign Queue_8__EVAL = _EVAL_34;
  assign Queue_12__EVAL_5 = _EVAL_46;
  assign Queue_10__EVAL_4 = _EVAL_134 & _EVAL_249;
  assign _EVAL_74 = _EVAL_29;
  assign _EVAL_38 = _EVAL_18;
  assign Queue_7__EVAL_4 = _EVAL_60;
  assign Queue_10__EVAL_5 = _EVAL_51;
  assign Queue_2__EVAL_0 = _EVAL_34;
  assign Queue_11__EVAL = _EVAL_134 & _EVAL_256;
  assign Queue_15__EVAL_4 = _EVAL_51;
  assign _EVAL_72 = _EVAL_37;
  assign _EVAL_70 = _EVAL_0;
  assign Queue_13__EVAL_5 = _EVAL_46;
  assign _EVAL_1 = _EVAL_15;
  assign Queue_4__EVAL = _EVAL_131 & _EVAL_24;
  assign _EVAL_20 = _EVAL_63 & _EVAL_100;
  assign Queue_2__EVAL = _EVAL_223 & _EVAL_171;
endmodule
