//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_86_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [7:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_23;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_47;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_87;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_92;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_97;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_126;
  reg [31:0] _RAND_5;
  reg  _EVAL_142;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_145;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_197;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_198;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_206;
  reg [31:0] _RAND_10;
  reg  _EVAL_212;
  reg [31:0] _RAND_11;
  reg  _EVAL_234;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_252;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_261;
  reg [31:0] _RAND_14;
  wire  _EVAL_18;
  wire  _EVAL_46;
  wire  _EVAL_192;
  wire  _EVAL_30;
  wire [1:0] _EVAL_179;
  wire [3:0] _EVAL_210;
  wire [2:0] _EVAL_49;
  wire [2:0] _EVAL_72;
  wire  _EVAL_240;
  wire  _EVAL_111;
  wire  _EVAL_242;
  wire  _EVAL_257;
  wire  _EVAL_102;
  wire  _EVAL_154;
  wire  _EVAL_159;
  wire  _EVAL_259;
  wire  _EVAL_129;
  wire  _EVAL_229;
  wire  _EVAL_139;
  wire  _EVAL_223;
  wire  _EVAL_90;
  wire  _EVAL_185;
  wire  _EVAL_36;
  wire  _EVAL_100;
  wire  _EVAL_41;
  wire  _EVAL_224;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_160;
  wire  _EVAL_150;
  wire  _EVAL_54;
  wire  _EVAL_233;
  wire  _EVAL_101;
  wire  _EVAL_162;
  wire  _EVAL_120;
  wire  _EVAL_71;
  wire  _EVAL_253;
  wire [1:0] _EVAL_177;
  wire  _EVAL_79;
  wire  _EVAL_98;
  wire  _EVAL_196;
  wire  _EVAL_201;
  wire  _EVAL_271;
  wire  _EVAL_117;
  wire  _EVAL_125;
  wire  _EVAL_272;
  wire  _EVAL_121;
  wire  _EVAL_64;
  wire  _EVAL_67;
  wire  _EVAL_176;
  wire  _EVAL_124;
  wire  _EVAL_204;
  wire  _EVAL_108;
  wire  _EVAL_84;
  wire  _EVAL_169;
  wire  _EVAL_17;
  wire  _EVAL_24;
  wire  _EVAL_237;
  wire  _EVAL_94;
  wire  _EVAL_219;
  wire  _EVAL_274;
  wire  _EVAL_255;
  wire  _EVAL_109;
  wire  _EVAL_221;
  wire  _EVAL_115;
  wire  _EVAL_265;
  wire  _EVAL_32;
  wire  _EVAL_172;
  wire  _EVAL_33;
  wire  _EVAL_56;
  wire [7:0] _EVAL_44;
  wire [7:0] _EVAL_215;
  wire [7:0] _EVAL_93;
  wire  _EVAL_258;
  wire  _EVAL_29;
  wire  _EVAL_280;
  wire  _EVAL_217;
  wire  _EVAL_170;
  wire  _EVAL_110;
  wire  _EVAL_218;
  wire  _EVAL_195;
  wire  _EVAL_22;
  wire  _EVAL_144;
  wire  _EVAL_194;
  wire [12:0] _EVAL_42;
  wire [5:0] _EVAL_184;
  wire  _EVAL_208;
  wire  _EVAL_188;
  wire  _EVAL_245;
  wire  _EVAL_264;
  wire  _EVAL_151;
  wire [5:0] _EVAL_66;
  wire [31:0] _EVAL_116;
  wire [31:0] _EVAL_279;
  wire  _EVAL_85;
  wire  _EVAL_99;
  wire [2:0] _EVAL_35;
  wire  _EVAL_112;
  wire  _EVAL_130;
  wire [12:0] _EVAL_189;
  wire [5:0] _EVAL_105;
  wire [5:0] _EVAL_248;
  wire [2:0] _EVAL_25;
  wire [31:0] _EVAL_267;
  wire [32:0] _EVAL_131;
  wire [32:0] _EVAL_173;
  wire [32:0] _EVAL_239;
  wire  _EVAL_104;
  wire  _EVAL_163;
  wire  _EVAL_183;
  wire  _EVAL_69;
  wire  _EVAL_205;
  wire  _EVAL_149;
  wire  _EVAL_53;
  wire [1:0] _EVAL_134;
  wire [1:0] _EVAL_96;
  wire  _EVAL_40;
  wire  _EVAL_281;
  wire  _EVAL_244;
  wire  _EVAL_37;
  wire  _EVAL_180;
  wire [7:0] _EVAL_199;
  wire  _EVAL_55;
  wire  _EVAL_76;
  wire  _EVAL_246;
  wire  _EVAL_278;
  wire  _EVAL_62;
  wire  _EVAL_138;
  wire  _EVAL_152;
  wire [1:0] _EVAL_157;
  wire [1:0] _EVAL_262;
  wire [1:0] _EVAL_59;
  wire [1:0] _EVAL_166;
  wire  _EVAL_45;
  wire  _EVAL_203;
  wire  _EVAL_20;
  wire [31:0] _EVAL_103;
  wire  _EVAL_282;
  wire  _EVAL_164;
  wire  _EVAL_228;
  wire  _EVAL_27;
  wire  _EVAL_168;
  wire  _EVAL_236;
  wire [1:0] _EVAL_119;
  wire [1:0] _EVAL_226;
  wire [1:0] _EVAL_275;
  wire  _EVAL_65;
  wire  _EVAL_82;
  wire [2:0] _EVAL_114;
  wire [2:0] _EVAL_60;
  wire [2:0] _EVAL_238;
  wire  _EVAL_283;
  wire  _EVAL_182;
  wire  _EVAL_39;
  wire  _EVAL_128;
  wire  _EVAL_175;
  wire  _EVAL_141;
  wire  _EVAL_222;
  wire  _EVAL_91;
  wire [2:0] _EVAL_250;
  wire  _EVAL_123;
  wire  _EVAL_19;
  wire  _EVAL_187;
  wire  _EVAL_256;
  wire  _EVAL_147;
  wire  _EVAL_106;
  wire  _EVAL_48;
  wire  _EVAL_107;
  wire  _EVAL_51;
  wire  _EVAL_178;
  wire  _EVAL_207;
  wire  _EVAL_146;
  wire  _EVAL_95;
  wire  _EVAL_73;
  wire  _EVAL_52;
  wire  _EVAL_61;
  wire  _EVAL_83;
  wire  _EVAL_135;
  wire  _EVAL_270;
  wire  _EVAL_57;
  wire  _EVAL_28;
  wire  _EVAL_133;
  wire  _EVAL_273;
  wire  _EVAL_63;
  wire  _EVAL_21;
  wire  _EVAL_153;
  wire  _EVAL_161;
  wire  _EVAL_77;
  wire  _EVAL_155;
  wire  _EVAL_171;
  wire  _EVAL_186;
  wire  _EVAL_249;
  wire  _EVAL_181;
  wire  _EVAL_81;
  wire  _EVAL_193;
  wire  _EVAL_31;
  wire  _EVAL_78;
  wire  _EVAL_225;
  wire  _EVAL_80;
  wire  _EVAL_118;
  wire  _EVAL_167;
  wire  _EVAL_216;
  wire  _EVAL_232;
  wire  _EVAL_43;
  wire  _EVAL_276;
  wire  _EVAL_140;
  wire  _EVAL_211;
  wire  _EVAL_235;
  wire  _EVAL_266;
  wire  _EVAL_70;
  wire  _EVAL_214;
  wire  _EVAL_34;
  wire  _EVAL_127;
  wire  _EVAL_254;
  wire  _EVAL_122;
  wire  _EVAL_251;
  wire  _EVAL_165;
  wire  _EVAL_132;
  wire  _EVAL_58;
  wire  _EVAL_231;
  wire  _EVAL_26;
  wire  _EVAL_260;
  wire  _EVAL_269;
  wire  _EVAL_227;
  wire  _EVAL_191;
  wire  _EVAL_68;
  wire  _EVAL_213;
  wire  _EVAL_137;
  wire  _EVAL_263;
  wire  _EVAL_277;
  wire  _EVAL_200;
  wire  _EVAL_202;
  wire  _EVAL_209;
  wire  _EVAL_220;
  wire  _EVAL_113;
  wire  _EVAL_74;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_18 = _EVAL_14 == 1'h0;
  assign _EVAL_46 = _EVAL_18 | _EVAL_11;
  assign _EVAL_192 = _EVAL_126 == 3'h0;
  assign _EVAL_30 = _EVAL_15 >= 3'h3;
  assign _EVAL_179 = _EVAL_15[1:0];
  assign _EVAL_210 = 4'h1 << _EVAL_179;
  assign _EVAL_49 = _EVAL_210[2:0];
  assign _EVAL_72 = _EVAL_49 | 3'h1;
  assign _EVAL_240 = _EVAL_72[2];
  assign _EVAL_111 = _EVAL_1[2];
  assign _EVAL_242 = _EVAL_111 == 1'h0;
  assign _EVAL_257 = _EVAL_240 & _EVAL_242;
  assign _EVAL_102 = _EVAL_30 | _EVAL_257;
  assign _EVAL_154 = _EVAL_72[1];
  assign _EVAL_159 = _EVAL_1[1];
  assign _EVAL_259 = _EVAL_242 & _EVAL_159;
  assign _EVAL_129 = _EVAL_154 & _EVAL_259;
  assign _EVAL_229 = _EVAL_102 | _EVAL_129;
  assign _EVAL_139 = _EVAL_72[0];
  assign _EVAL_223 = _EVAL_1[0];
  assign _EVAL_90 = _EVAL_223 == 1'h0;
  assign _EVAL_185 = _EVAL_259 & _EVAL_90;
  assign _EVAL_36 = _EVAL_139 & _EVAL_185;
  assign _EVAL_100 = _EVAL_229 | _EVAL_36;
  assign _EVAL_41 = _EVAL_9 != 3'h0;
  assign _EVAL_224 = _EVAL_41 | _EVAL_11;
  assign _EVAL_88 = _EVAL_224 == 1'h0;
  assign _EVAL_89 = _EVAL_159 == 1'h0;
  assign _EVAL_160 = _EVAL_111 & _EVAL_89;
  assign _EVAL_150 = _EVAL_1 == _EVAL_47;
  assign _EVAL_54 = _EVAL_150 | _EVAL_11;
  assign _EVAL_233 = _EVAL_111 & _EVAL_159;
  assign _EVAL_101 = _EVAL_233 & _EVAL_223;
  assign _EVAL_162 = _EVAL_5 == _EVAL_87;
  assign _EVAL_120 = _EVAL_162 | _EVAL_11;
  assign _EVAL_71 = _EVAL_120 == 1'h0;
  assign _EVAL_253 = _EVAL_3 == 3'h3;
  assign _EVAL_177 = _EVAL_197 >> _EVAL_12;
  assign _EVAL_79 = _EVAL_177[0];
  assign _EVAL_98 = _EVAL_79 == 1'h0;
  assign _EVAL_196 = _EVAL_3 == 3'h6;
  assign _EVAL_201 = _EVAL_240 & _EVAL_111;
  assign _EVAL_271 = _EVAL_30 | _EVAL_201;
  assign _EVAL_117 = _EVAL_154 & _EVAL_233;
  assign _EVAL_125 = _EVAL_271 | _EVAL_117;
  assign _EVAL_272 = _EVAL_139 & _EVAL_101;
  assign _EVAL_121 = _EVAL_125 | _EVAL_272;
  assign _EVAL_64 = _EVAL_233 & _EVAL_90;
  assign _EVAL_67 = _EVAL_139 & _EVAL_64;
  assign _EVAL_176 = _EVAL_125 | _EVAL_67;
  assign _EVAL_124 = _EVAL_154 & _EVAL_160;
  assign _EVAL_204 = _EVAL_271 | _EVAL_124;
  assign _EVAL_108 = _EVAL_160 & _EVAL_223;
  assign _EVAL_84 = _EVAL_139 & _EVAL_108;
  assign _EVAL_169 = _EVAL_204 | _EVAL_84;
  assign _EVAL_17 = _EVAL_160 & _EVAL_90;
  assign _EVAL_24 = _EVAL_139 & _EVAL_17;
  assign _EVAL_237 = _EVAL_204 | _EVAL_24;
  assign _EVAL_94 = _EVAL_259 & _EVAL_223;
  assign _EVAL_219 = _EVAL_139 & _EVAL_94;
  assign _EVAL_274 = _EVAL_229 | _EVAL_219;
  assign _EVAL_255 = _EVAL_242 & _EVAL_89;
  assign _EVAL_109 = _EVAL_154 & _EVAL_255;
  assign _EVAL_221 = _EVAL_102 | _EVAL_109;
  assign _EVAL_115 = _EVAL_255 & _EVAL_223;
  assign _EVAL_265 = _EVAL_139 & _EVAL_115;
  assign _EVAL_32 = _EVAL_221 | _EVAL_265;
  assign _EVAL_172 = _EVAL_255 & _EVAL_90;
  assign _EVAL_33 = _EVAL_139 & _EVAL_172;
  assign _EVAL_56 = _EVAL_221 | _EVAL_33;
  assign _EVAL_44 = {_EVAL_121,_EVAL_176,_EVAL_169,_EVAL_237,_EVAL_274,_EVAL_100,_EVAL_32,_EVAL_56};
  assign _EVAL_215 = ~ _EVAL_44;
  assign _EVAL_93 = _EVAL_10 & _EVAL_215;
  assign _EVAL_258 = _EVAL_93 == 8'h0;
  assign _EVAL_29 = _EVAL_258 | _EVAL_11;
  assign _EVAL_280 = _EVAL_29 == 1'h0;
  assign _EVAL_217 = _EVAL_15 == _EVAL_206;
  assign _EVAL_170 = _EVAL_217 | _EVAL_11;
  assign _EVAL_110 = _EVAL_170 == 1'h0;
  assign _EVAL_218 = _EVAL_30 | _EVAL_11;
  assign _EVAL_195 = _EVAL_13 & _EVAL;
  assign _EVAL_22 = _EVAL_97 == 3'h0;
  assign _EVAL_144 = _EVAL_195 & _EVAL_22;
  assign _EVAL_194 = _EVAL_3 == 3'h5;
  assign _EVAL_42 = 13'h3f << _EVAL_15;
  assign _EVAL_184 = _EVAL_42[5:0];
  assign _EVAL_208 = _EVAL_5 <= 3'h6;
  assign _EVAL_188 = _EVAL_3 == 3'h7;
  assign _EVAL_245 = _EVAL & _EVAL_188;
  assign _EVAL_264 = _EVAL_9 == _EVAL_261;
  assign _EVAL_151 = _EVAL & _EVAL_253;
  assign _EVAL_66 = ~ _EVAL_184;
  assign _EVAL_116 = {{26'd0}, _EVAL_66};
  assign _EVAL_279 = _EVAL_1 & _EVAL_116;
  assign _EVAL_85 = _EVAL_279 == 32'h0;
  assign _EVAL_99 = _EVAL_85 | _EVAL_11;
  assign _EVAL_35 = _EVAL_23 - 3'h1;
  assign _EVAL_112 = _EVAL_23 == 3'h0;
  assign _EVAL_130 = _EVAL_5[0];
  assign _EVAL_189 = 13'h3f << _EVAL_0;
  assign _EVAL_105 = _EVAL_189[5:0];
  assign _EVAL_248 = ~ _EVAL_105;
  assign _EVAL_25 = _EVAL_248[5:3];
  assign _EVAL_267 = _EVAL_1 ^ 32'h80000000;
  assign _EVAL_131 = {1'b0,$signed(_EVAL_267)};
  assign _EVAL_173 = $signed(_EVAL_131) & $signed(-33'sh20000);
  assign _EVAL_239 = $signed(_EVAL_173);
  assign _EVAL_104 = _EVAL_3 == 3'h2;
  assign _EVAL_163 = _EVAL & _EVAL_104;
  assign _EVAL_183 = _EVAL_7 & _EVAL_6;
  assign _EVAL_69 = _EVAL_183 & _EVAL_112;
  assign _EVAL_205 = _EVAL_5 == 3'h6;
  assign _EVAL_149 = _EVAL_205 == 1'h0;
  assign _EVAL_53 = _EVAL_69 & _EVAL_149;
  assign _EVAL_134 = 2'h1 << _EVAL_16;
  assign _EVAL_96 = _EVAL_53 ? _EVAL_134 : 2'h0;
  assign _EVAL_40 = _EVAL_2 == 1'h0;
  assign _EVAL_281 = _EVAL_40 | _EVAL_11;
  assign _EVAL_244 = _EVAL_9 <= 3'h3;
  assign _EVAL_37 = _EVAL_244 | _EVAL_11;
  assign _EVAL_180 = _EVAL_37 == 1'h0;
  assign _EVAL_199 = ~ _EVAL_10;
  assign _EVAL_55 = _EVAL_199 == 8'h0;
  assign _EVAL_76 = _EVAL_16 == _EVAL_234;
  assign _EVAL_246 = _EVAL_92 == 3'h0;
  assign _EVAL_278 = _EVAL_195 & _EVAL_246;
  assign _EVAL_62 = _EVAL_0 == _EVAL_198;
  assign _EVAL_138 = _EVAL_62 | _EVAL_11;
  assign _EVAL_152 = _EVAL_138 == 1'h0;
  assign _EVAL_157 = 2'h1 << _EVAL_12;
  assign _EVAL_262 = _EVAL_278 ? _EVAL_157 : 2'h0;
  assign _EVAL_59 = _EVAL_262 | _EVAL_197;
  assign _EVAL_166 = _EVAL_59 >> _EVAL_16;
  assign _EVAL_45 = _EVAL_166[0];
  assign _EVAL_203 = _EVAL_45 | _EVAL_11;
  assign _EVAL_20 = _EVAL_203 == 1'h0;
  assign _EVAL_103 = _EVAL_252 + 32'h1;
  assign _EVAL_282 = _EVAL_262 != _EVAL_96;
  assign _EVAL_164 = _EVAL_262 != 2'h0;
  assign _EVAL_228 = _EVAL_164 == 1'h0;
  assign _EVAL_27 = _EVAL_282 | _EVAL_228;
  assign _EVAL_168 = _EVAL_9 == 3'h0;
  assign _EVAL_236 = _EVAL_168 | _EVAL_11;
  assign _EVAL_119 = _EVAL_197 | _EVAL_262;
  assign _EVAL_226 = ~ _EVAL_96;
  assign _EVAL_275 = _EVAL_119 & _EVAL_226;
  assign _EVAL_65 = _EVAL_3[2];
  assign _EVAL_82 = _EVAL_65 == 1'h0;
  assign _EVAL_114 = _EVAL_66[5:3];
  assign _EVAL_60 = _EVAL_97 - 3'h1;
  assign _EVAL_238 = _EVAL_126 - 3'h1;
  assign _EVAL_283 = _EVAL_192 == 1'h0;
  assign _EVAL_182 = _EVAL_3 == 3'h1;
  assign _EVAL_39 = _EVAL & _EVAL_182;
  assign _EVAL_128 = _EVAL_15 <= 3'h6;
  assign _EVAL_175 = $signed(_EVAL_239) == $signed(33'sh0);
  assign _EVAL_141 = _EVAL_128 & _EVAL_175;
  assign _EVAL_222 = _EVAL & _EVAL_194;
  assign _EVAL_91 = _EVAL_195 | _EVAL_183;
  assign _EVAL_250 = _EVAL_92 - 3'h1;
  assign _EVAL_123 = _EVAL_197 != 2'h0;
  assign _EVAL_19 = _EVAL_123 == 1'h0;
  assign _EVAL_187 = plusarg_reader_out == 32'h0;
  assign _EVAL_256 = _EVAL_19 | _EVAL_187;
  assign _EVAL_147 = _EVAL_252 < plusarg_reader_out;
  assign _EVAL_106 = _EVAL_256 | _EVAL_147;
  assign _EVAL_48 = _EVAL_106 | _EVAL_11;
  assign _EVAL_107 = _EVAL_10 == _EVAL_44;
  assign _EVAL_51 = _EVAL_3 == 3'h4;
  assign _EVAL_178 = _EVAL_107 | _EVAL_11;
  assign _EVAL_207 = _EVAL_178 == 1'h0;
  assign _EVAL_146 = _EVAL_3 == _EVAL_145;
  assign _EVAL_95 = _EVAL_146 | _EVAL_11;
  assign _EVAL_73 = _EVAL_95 == 1'h0;
  assign _EVAL_52 = _EVAL_9 <= 3'h4;
  assign _EVAL_61 = _EVAL_264 | _EVAL_11;
  assign _EVAL_83 = _EVAL_5 == 3'h4;
  assign _EVAL_135 = _EVAL_6 & _EVAL_83;
  assign _EVAL_270 = _EVAL_14 == _EVAL_142;
  assign _EVAL_57 = _EVAL_270 | _EVAL_11;
  assign _EVAL_28 = _EVAL_57 == 1'h0;
  assign _EVAL_133 = _EVAL_9 <= 3'h2;
  assign _EVAL_273 = _EVAL_133 | _EVAL_11;
  assign _EVAL_63 = _EVAL_5 == 3'h1;
  assign _EVAL_21 = _EVAL_6 & _EVAL_63;
  assign _EVAL_153 = _EVAL_55 | _EVAL_11;
  assign _EVAL_161 = _EVAL_153 == 1'h0;
  assign _EVAL_77 = _EVAL_8 == 1'h0;
  assign _EVAL_155 = _EVAL_52 | _EVAL_11;
  assign _EVAL_171 = _EVAL_236 == 1'h0;
  assign _EVAL_186 = _EVAL_0 >= 3'h3;
  assign _EVAL_249 = _EVAL_186 | _EVAL_11;
  assign _EVAL_181 = _EVAL_249 == 1'h0;
  assign _EVAL_81 = _EVAL_76 | _EVAL_11;
  assign _EVAL_193 = _EVAL_81 == 1'h0;
  assign _EVAL_31 = _EVAL_5 == 3'h2;
  assign _EVAL_78 = _EVAL_6 & _EVAL_31;
  assign _EVAL_225 = _EVAL_5 == 3'h5;
  assign _EVAL_80 = _EVAL_5 == 3'h0;
  assign _EVAL_118 = _EVAL_6 & _EVAL_80;
  assign _EVAL_167 = _EVAL_141 | _EVAL_11;
  assign _EVAL_216 = _EVAL_208 | _EVAL_11;
  assign _EVAL_232 = _EVAL_216 == 1'h0;
  assign _EVAL_43 = _EVAL_98 | _EVAL_11;
  assign _EVAL_276 = _EVAL_43 == 1'h0;
  assign _EVAL_140 = _EVAL_18 | _EVAL_8;
  assign _EVAL_211 = _EVAL_140 | _EVAL_11;
  assign _EVAL_235 = _EVAL_211 == 1'h0;
  assign _EVAL_266 = _EVAL_218 == 1'h0;
  assign _EVAL_70 = _EVAL_3 == 3'h0;
  assign _EVAL_214 = _EVAL & _EVAL_70;
  assign _EVAL_34 = _EVAL_6 & _EVAL_283;
  assign _EVAL_127 = _EVAL_54 == 1'h0;
  assign _EVAL_254 = _EVAL_27 | _EVAL_11;
  assign _EVAL_122 = _EVAL_11 == 1'h0;
  assign _EVAL_251 = _EVAL_99 == 1'h0;
  assign _EVAL_165 = _EVAL_12 == _EVAL_212;
  assign _EVAL_132 = _EVAL_165 | _EVAL_11;
  assign _EVAL_58 = _EVAL_77 | _EVAL_11;
  assign _EVAL_231 = _EVAL_58 == 1'h0;
  assign _EVAL_26 = _EVAL_281 == 1'h0;
  assign _EVAL_260 = _EVAL_155 == 1'h0;
  assign _EVAL_269 = _EVAL_6 & _EVAL_225;
  assign _EVAL_227 = _EVAL_22 == 1'h0;
  assign _EVAL_191 = _EVAL_61 == 1'h0;
  assign _EVAL_68 = _EVAL_167 == 1'h0;
  assign _EVAL_213 = _EVAL & _EVAL_51;
  assign _EVAL_137 = _EVAL & _EVAL_227;
  assign _EVAL_263 = _EVAL_6 & _EVAL_205;
  assign _EVAL_277 = _EVAL_48 == 1'h0;
  assign _EVAL_200 = _EVAL_183 & _EVAL_192;
  assign _EVAL_202 = _EVAL_132 == 1'h0;
  assign _EVAL_209 = _EVAL_254 == 1'h0;
  assign _EVAL_220 = _EVAL & _EVAL_196;
  assign _EVAL_113 = _EVAL_273 == 1'h0;
  assign _EVAL_74 = _EVAL_46 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_47 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_87 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_92 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_97 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_126 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_142 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_145 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_197 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_198 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_206 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_212 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_234 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_252 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_261 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_11) begin
      _EVAL_23 <= 3'h0;
    end else begin
      if (_EVAL_183) begin
        if (_EVAL_112) begin
          if (_EVAL_130) begin
            _EVAL_23 <= _EVAL_25;
          end else begin
            _EVAL_23 <= 3'h0;
          end
        end else begin
          _EVAL_23 <= _EVAL_35;
        end
      end
    end
    if (_EVAL_144) begin
      _EVAL_47 <= _EVAL_1;
    end
    if (_EVAL_200) begin
      _EVAL_87 <= _EVAL_5;
    end
    if (_EVAL_11) begin
      _EVAL_92 <= 3'h0;
    end else begin
      if (_EVAL_195) begin
        if (_EVAL_246) begin
          if (_EVAL_82) begin
            _EVAL_92 <= _EVAL_114;
          end else begin
            _EVAL_92 <= 3'h0;
          end
        end else begin
          _EVAL_92 <= _EVAL_250;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_97 <= 3'h0;
    end else begin
      if (_EVAL_195) begin
        if (_EVAL_22) begin
          if (_EVAL_82) begin
            _EVAL_97 <= _EVAL_114;
          end else begin
            _EVAL_97 <= 3'h0;
          end
        end else begin
          _EVAL_97 <= _EVAL_60;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_126 <= 3'h0;
    end else begin
      if (_EVAL_183) begin
        if (_EVAL_192) begin
          if (_EVAL_130) begin
            _EVAL_126 <= _EVAL_25;
          end else begin
            _EVAL_126 <= 3'h0;
          end
        end else begin
          _EVAL_126 <= _EVAL_238;
        end
      end
    end
    if (_EVAL_200) begin
      _EVAL_142 <= _EVAL_14;
    end
    if (_EVAL_144) begin
      _EVAL_145 <= _EVAL_3;
    end
    if (_EVAL_11) begin
      _EVAL_197 <= 2'h0;
    end else begin
      _EVAL_197 <= _EVAL_275;
    end
    if (_EVAL_200) begin
      _EVAL_198 <= _EVAL_0;
    end
    if (_EVAL_144) begin
      _EVAL_206 <= _EVAL_15;
    end
    if (_EVAL_144) begin
      _EVAL_212 <= _EVAL_12;
    end
    if (_EVAL_200) begin
      _EVAL_234 <= _EVAL_16;
    end
    if (_EVAL_11) begin
      _EVAL_252 <= 32'h0;
    end else begin
      if (_EVAL_91) begin
        _EVAL_252 <= 32'h0;
      end else begin
        _EVAL_252 <= _EVAL_103;
      end
    end
    if (_EVAL_144) begin
      _EVAL_261 <= _EVAL_9;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(757cd941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d1d407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f6c8d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9301317)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34829bb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a72214c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6618f884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f1cfa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(925571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0321069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dfd192a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3896813)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0d71cd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a81aa1b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e664da64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97d7e3a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cc965d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4eab5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c802fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac3bf095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7692c77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c42e96fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5ec70a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba6474f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27a1d181)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f89e183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b11db30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5ab765a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43ca8df8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1312dd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b15eb2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93bd7a10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac66f4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cc728cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a289d278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bc97d04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d70d05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f9ae626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(710fe105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ed040f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bb8609a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afe0c019)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e4acac0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0ecb700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c24c8837)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c90ac999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54d12b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6960d4a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e4c20e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d489177f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3777fa8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6097ef0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9f721d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e16be20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9421a40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81450337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55f7467c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d2616af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(613e5455)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e79067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f096302)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5246ffcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4992ed43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(308d6e68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(766738a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb11eabb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
