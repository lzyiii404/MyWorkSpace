//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_51_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [4:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [4:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [1:0] _EVAL_21;
  reg [31:0] _RAND_0;
  reg [4:0] _EVAL_106;
  reg [31:0] _RAND_1;
  reg [31:0] _EVAL_139;
  reg [31:0] _RAND_2;
  reg [4:0] _EVAL_152;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_180;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_193;
  reg [31:0] _RAND_5;
  reg [31:0] _EVAL_196;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_233;
  reg [31:0] _RAND_7;
  reg [5:0] _EVAL_258;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_306;
  reg [31:0] _RAND_9;
  reg  _EVAL_320;
  reg [31:0] _RAND_10;
  reg [5:0] _EVAL_323;
  reg [31:0] _RAND_11;
  reg  _EVAL_325;
  reg [31:0] _RAND_12;
  reg [5:0] _EVAL_341;
  reg [31:0] _RAND_13;
  reg [5:0] _EVAL_347;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_351;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_357;
  reg [31:0] _RAND_16;
  wire  _EVAL_276;
  wire  _EVAL_292;
  wire  _EVAL_197;
  wire  _EVAL_82;
  wire  _EVAL_85;
  wire [3:0] _EVAL_309;
  wire  _EVAL_348;
  wire  _EVAL_287;
  wire  _EVAL_54;
  wire  _EVAL_70;
  wire  _EVAL_46;
  wire  _EVAL_281;
  wire  _EVAL_262;
  wire  _EVAL_286;
  wire  _EVAL_231;
  wire  _EVAL_184;
  wire [31:0] _EVAL_263;
  wire [32:0] _EVAL_211;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_33;
  wire  _EVAL_328;
  wire [22:0] _EVAL_135;
  wire [7:0] _EVAL_343;
  wire [7:0] _EVAL_76;
  wire [31:0] _EVAL_169;
  wire  _EVAL_95;
  wire [31:0] _EVAL_22;
  wire [32:0] _EVAL_108;
  wire [32:0] _EVAL_295;
  wire [32:0] _EVAL_223;
  wire  _EVAL_125;
  wire  _EVAL_153;
  wire  _EVAL_317;
  wire  _EVAL_356;
  wire [1:0] _EVAL_313;
  wire [1:0] _EVAL_352;
  wire  _EVAL_148;
  wire  _EVAL_307;
  wire  _EVAL_111;
  wire  _EVAL_183;
  wire  _EVAL_246;
  wire  _EVAL_140;
  wire  _EVAL_342;
  wire  _EVAL_207;
  wire  _EVAL_141;
  wire  _EVAL_302;
  wire  _EVAL_122;
  wire  _EVAL_267;
  wire  _EVAL_336;
  wire  _EVAL_298;
  wire  _EVAL_100;
  wire  _EVAL_327;
  wire  _EVAL_282;
  wire  _EVAL_144;
  wire  _EVAL_168;
  wire  _EVAL_319;
  wire  _EVAL_132;
  wire  _EVAL_94;
  wire [3:0] _EVAL_208;
  wire [3:0] _EVAL_29;
  wire [3:0] _EVAL_47;
  wire  _EVAL_142;
  wire [1:0] _EVAL_93;
  wire  _EVAL_155;
  wire  _EVAL_56;
  wire  _EVAL_165;
  wire  _EVAL_92;
  wire  _EVAL_252;
  wire  _EVAL_151;
  wire  _EVAL_202;
  wire [31:0] _EVAL_237;
  wire [32:0] _EVAL_273;
  wire [32:0] _EVAL_41;
  wire [32:0] _EVAL_296;
  wire [31:0] _EVAL_51;
  wire [32:0] _EVAL_43;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_102;
  wire  _EVAL_290;
  wire  _EVAL_264;
  wire  _EVAL_161;
  wire [32:0] _EVAL_175;
  wire [32:0] _EVAL_222;
  wire [32:0] _EVAL_84;
  wire  _EVAL_185;
  wire  _EVAL_162;
  wire [31:0] _EVAL_304;
  wire [32:0] _EVAL_189;
  wire [32:0] _EVAL_133;
  wire [32:0] _EVAL_24;
  wire  _EVAL_114;
  wire  _EVAL_335;
  wire [31:0] _EVAL_52;
  wire [32:0] _EVAL_34;
  wire [32:0] _EVAL_32;
  wire [32:0] _EVAL_186;
  wire  _EVAL_120;
  wire  _EVAL_40;
  wire [31:0] _EVAL_340;
  wire [32:0] _EVAL_105;
  wire [32:0] _EVAL_48;
  wire [32:0] _EVAL_271;
  wire  _EVAL_293;
  wire  _EVAL_128;
  wire  _EVAL_269;
  wire  _EVAL_121;
  wire  _EVAL_265;
  wire [5:0] _EVAL_158;
  wire [5:0] _EVAL_49;
  wire  _EVAL_55;
  wire  _EVAL_154;
  wire  _EVAL_30;
  wire [31:0] _EVAL_159;
  wire [31:0] _EVAL_318;
  wire [31:0] _EVAL_194;
  wire  _EVAL_322;
  wire [31:0] _EVAL_213;
  wire [32:0] _EVAL_31;
  wire [32:0] _EVAL_88;
  wire [32:0] _EVAL_28;
  wire  _EVAL_127;
  wire  _EVAL_115;
  wire [1:0] _EVAL_72;
  wire  _EVAL_355;
  wire  _EVAL_270;
  wire  _EVAL_353;
  wire  _EVAL_134;
  wire  _EVAL_236;
  wire  _EVAL_249;
  wire  _EVAL_245;
  wire  _EVAL_79;
  wire  _EVAL_203;
  wire  _EVAL_294;
  wire  _EVAL_23;
  wire  _EVAL_260;
  wire  _EVAL_173;
  wire  _EVAL_230;
  wire  _EVAL_75;
  wire  _EVAL_349;
  wire  _EVAL_218;
  wire [5:0] _EVAL_239;
  wire  _EVAL_204;
  wire  _EVAL_113;
  wire  _EVAL_177;
  wire  _EVAL_164;
  wire  _EVAL_179;
  wire  _EVAL_280;
  wire  _EVAL_358;
  wire  _EVAL_181;
  wire  _EVAL_209;
  wire [31:0] _EVAL_244;
  wire [31:0] _EVAL_195;
  wire  _EVAL_63;
  wire  _EVAL_61;
  wire  _EVAL_107;
  wire  _EVAL_316;
  wire  _EVAL_224;
  wire  _EVAL_42;
  wire  _EVAL_337;
  wire  _EVAL_35;
  wire [31:0] _EVAL_266;
  wire  _EVAL_57;
  wire  _EVAL_321;
  wire  _EVAL_101;
  wire  _EVAL_274;
  wire  _EVAL_279;
  wire  _EVAL_330;
  wire  _EVAL_45;
  wire  _EVAL_126;
  wire  _EVAL_27;
  wire  _EVAL_227;
  wire  _EVAL_205;
  wire [22:0] _EVAL_261;
  wire [7:0] _EVAL_117;
  wire [7:0] _EVAL_272;
  wire [5:0] _EVAL_240;
  wire  _EVAL_283;
  wire [5:0] _EVAL_332;
  wire  _EVAL_78;
  wire  _EVAL_344;
  wire  _EVAL_301;
  wire  _EVAL_87;
  wire  _EVAL_71;
  wire  _EVAL_38;
  wire  _EVAL_345;
  wire  _EVAL_138;
  wire  _EVAL_253;
  wire  _EVAL_324;
  wire  _EVAL_53;
  wire  _EVAL_257;
  wire  _EVAL_39;
  wire  _EVAL_214;
  wire  _EVAL_346;
  wire  _EVAL_86;
  wire  _EVAL_220;
  wire  _EVAL_229;
  wire  _EVAL_145;
  wire  _EVAL_90;
  wire [31:0] _EVAL_187;
  wire [31:0] _EVAL_188;
  wire  _EVAL_123;
  wire  _EVAL_277;
  wire  _EVAL_110;
  wire [31:0] _EVAL_190;
  wire  _EVAL_217;
  wire  _EVAL_228;
  wire  _EVAL_216;
  wire  _EVAL_291;
  wire  _EVAL_97;
  wire  _EVAL_64;
  wire  _EVAL_297;
  wire  _EVAL_89;
  wire  _EVAL_234;
  wire  _EVAL_178;
  wire  _EVAL_212;
  wire  _EVAL_167;
  wire  _EVAL_338;
  wire  _EVAL_235;
  wire  _EVAL_104;
  wire  _EVAL_232;
  wire  _EVAL_112;
  wire  _EVAL_109;
  wire  _EVAL_130;
  wire  _EVAL_243;
  wire  _EVAL_80;
  wire  _EVAL_334;
  wire  _EVAL_299;
  wire  _EVAL_226;
  wire  _EVAL_147;
  wire  _EVAL_314;
  wire  _EVAL_20;
  wire  _EVAL_312;
  wire  _EVAL_254;
  wire  _EVAL_124;
  wire [5:0] _EVAL_69;
  wire  _EVAL_242;
  wire  _EVAL_60;
  wire  _EVAL_96;
  wire  _EVAL_354;
  wire  _EVAL_198;
  wire  _EVAL_149;
  wire  _EVAL_26;
  wire  _EVAL_201;
  wire  _EVAL_25;
  wire  _EVAL_129;
  wire  _EVAL_200;
  wire [31:0] _EVAL_103;
  wire [31:0] _EVAL_176;
  wire  _EVAL_50;
  wire  _EVAL_278;
  wire  _EVAL_136;
  wire  _EVAL_131;
  wire  _EVAL_118;
  wire  _EVAL_160;
  wire  _EVAL_98;
  wire  _EVAL_288;
  wire  _EVAL_215;
  wire  _EVAL_171;
  wire  _EVAL_268;
  wire  _EVAL_137;
  wire  _EVAL_219;
  wire  _EVAL_44;
  wire  _EVAL_166;
  wire  _EVAL_143;
  wire  _EVAL_191;
  wire  _EVAL_331;
  wire  _EVAL_199;
  wire  _EVAL_37;
  wire  _EVAL_326;
  wire  _EVAL_66;
  wire  _EVAL_329;
  wire  _EVAL_256;
  wire  _EVAL_59;
  wire  _EVAL_67;
  wire  _EVAL_305;
  wire  _EVAL_119;
  wire  _EVAL_116;
  wire  _EVAL_300;
  wire  _EVAL_150;
  wire  _EVAL_275;
  wire  _EVAL_36;
  wire  _EVAL_315;
  wire  _EVAL_210;
  wire  _EVAL_146;
  wire  _EVAL_310;
  wire  _EVAL_192;
  wire  _EVAL_170;
  wire  _EVAL_62;
  wire  _EVAL_174;
  wire  _EVAL_247;
  wire  _EVAL_289;
  wire  _EVAL_221;
  wire  _EVAL_81;
  wire  _EVAL_65;
  wire  _EVAL_333;
  wire  _EVAL_99;
  wire  _EVAL_259;
  wire [31:0] _EVAL_225;
  wire  _EVAL_285;
  wire  _EVAL_19;
  wire  _EVAL_308;
  wire  _EVAL_251;
  wire  _EVAL_58;
  wire  _EVAL_83;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_68;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_276 = _EVAL_18 & _EVAL;
  assign _EVAL_292 = _EVAL_5 & _EVAL_3;
  assign _EVAL_197 = _EVAL_276 | _EVAL_292;
  assign _EVAL_82 = _EVAL_2 == 3'h2;
  assign _EVAL_85 = _EVAL & _EVAL_82;
  assign _EVAL_309 = ~ _EVAL_8;
  assign _EVAL_348 = _EVAL_309 == 4'h0;
  assign _EVAL_287 = _EVAL_348 | _EVAL_11;
  assign _EVAL_54 = _EVAL_196 != 32'h0;
  assign _EVAL_70 = _EVAL_54 == 1'h0;
  assign _EVAL_46 = plusarg_reader_out == 32'h0;
  assign _EVAL_281 = _EVAL_70 | _EVAL_46;
  assign _EVAL_262 = _EVAL_139 < plusarg_reader_out;
  assign _EVAL_286 = _EVAL_281 | _EVAL_262;
  assign _EVAL_231 = _EVAL_286 | _EVAL_11;
  assign _EVAL_184 = _EVAL_231 == 1'h0;
  assign _EVAL_263 = _EVAL_13 ^ 32'h2000000;
  assign _EVAL_211 = {1'b0,$signed(_EVAL_263)};
  assign _EVAL_163 = $signed(_EVAL_211) & $signed(-33'sh10000);
  assign _EVAL_33 = $signed(_EVAL_163);
  assign _EVAL_328 = $signed(_EVAL_33) == $signed(33'sh0);
  assign _EVAL_135 = 23'hff << _EVAL_6;
  assign _EVAL_343 = _EVAL_135[7:0];
  assign _EVAL_76 = ~ _EVAL_343;
  assign _EVAL_169 = {{24'd0}, _EVAL_76};
  assign _EVAL_95 = _EVAL_6 <= 4'h8;
  assign _EVAL_22 = _EVAL_13 ^ 32'h3000;
  assign _EVAL_108 = {1'b0,$signed(_EVAL_22)};
  assign _EVAL_295 = $signed(_EVAL_108) & $signed(-33'sh1000);
  assign _EVAL_223 = $signed(_EVAL_295);
  assign _EVAL_125 = $signed(_EVAL_223) == $signed(33'sh0);
  assign _EVAL_153 = _EVAL_95 & _EVAL_125;
  assign _EVAL_317 = _EVAL_6 >= 4'h2;
  assign _EVAL_356 = _EVAL_6[0];
  assign _EVAL_313 = 2'h1 << _EVAL_356;
  assign _EVAL_352 = _EVAL_313 | 2'h1;
  assign _EVAL_148 = _EVAL_352[1];
  assign _EVAL_307 = _EVAL_13[1];
  assign _EVAL_111 = _EVAL_148 & _EVAL_307;
  assign _EVAL_183 = _EVAL_317 | _EVAL_111;
  assign _EVAL_246 = _EVAL_352[0];
  assign _EVAL_140 = _EVAL_13[0];
  assign _EVAL_342 = _EVAL_307 & _EVAL_140;
  assign _EVAL_207 = _EVAL_246 & _EVAL_342;
  assign _EVAL_141 = _EVAL_183 | _EVAL_207;
  assign _EVAL_302 = _EVAL_140 == 1'h0;
  assign _EVAL_122 = _EVAL_307 & _EVAL_302;
  assign _EVAL_267 = _EVAL_246 & _EVAL_122;
  assign _EVAL_336 = _EVAL_183 | _EVAL_267;
  assign _EVAL_298 = _EVAL_307 == 1'h0;
  assign _EVAL_100 = _EVAL_148 & _EVAL_298;
  assign _EVAL_327 = _EVAL_317 | _EVAL_100;
  assign _EVAL_282 = _EVAL_298 & _EVAL_140;
  assign _EVAL_144 = _EVAL_246 & _EVAL_282;
  assign _EVAL_168 = _EVAL_327 | _EVAL_144;
  assign _EVAL_319 = _EVAL_298 & _EVAL_302;
  assign _EVAL_132 = _EVAL_246 & _EVAL_319;
  assign _EVAL_94 = _EVAL_327 | _EVAL_132;
  assign _EVAL_208 = {_EVAL_141,_EVAL_336,_EVAL_168,_EVAL_94};
  assign _EVAL_29 = ~ _EVAL_208;
  assign _EVAL_47 = _EVAL_8 & _EVAL_29;
  assign _EVAL_142 = _EVAL_47 == 4'h0;
  assign _EVAL_93 = _EVAL_9[4:3];
  assign _EVAL_155 = _EVAL_93 == 2'h0;
  assign _EVAL_56 = _EVAL_93 == 2'h1;
  assign _EVAL_165 = _EVAL_155 | _EVAL_56;
  assign _EVAL_92 = _EVAL_93 == 2'h2;
  assign _EVAL_252 = _EVAL_165 | _EVAL_92;
  assign _EVAL_151 = _EVAL_93 == 2'h3;
  assign _EVAL_202 = _EVAL_252 | _EVAL_151;
  assign _EVAL_237 = _EVAL_13 ^ 32'h40000000;
  assign _EVAL_273 = {1'b0,$signed(_EVAL_237)};
  assign _EVAL_41 = $signed(_EVAL_273) & $signed(-33'sh2000);
  assign _EVAL_296 = $signed(_EVAL_41);
  assign _EVAL_51 = _EVAL_13 ^ 32'hc000000;
  assign _EVAL_43 = {1'b0,$signed(_EVAL_51)};
  assign _EVAL_172 = $signed(_EVAL_43) & $signed(-33'sh4000000);
  assign _EVAL_102 = $signed(_EVAL_172);
  assign _EVAL_290 = $signed(_EVAL_102) == $signed(33'sh0);
  assign _EVAL_264 = _EVAL_125 | _EVAL_290;
  assign _EVAL_161 = _EVAL_264 | _EVAL_328;
  assign _EVAL_175 = {1'b0,$signed(_EVAL_13)};
  assign _EVAL_222 = $signed(_EVAL_175) & $signed(-33'sh5000);
  assign _EVAL_84 = $signed(_EVAL_222);
  assign _EVAL_185 = $signed(_EVAL_84) == $signed(33'sh0);
  assign _EVAL_162 = _EVAL_161 | _EVAL_185;
  assign _EVAL_304 = _EVAL_13 ^ 32'h1800000;
  assign _EVAL_189 = {1'b0,$signed(_EVAL_304)};
  assign _EVAL_133 = $signed(_EVAL_189) & $signed(-33'sh8000);
  assign _EVAL_24 = $signed(_EVAL_133);
  assign _EVAL_114 = $signed(_EVAL_24) == $signed(33'sh0);
  assign _EVAL_335 = _EVAL_162 | _EVAL_114;
  assign _EVAL_52 = _EVAL_13 ^ 32'h1900000;
  assign _EVAL_34 = {1'b0,$signed(_EVAL_52)};
  assign _EVAL_32 = $signed(_EVAL_34) & $signed(-33'sh2000);
  assign _EVAL_186 = $signed(_EVAL_32);
  assign _EVAL_120 = $signed(_EVAL_186) == $signed(33'sh0);
  assign _EVAL_40 = _EVAL_335 | _EVAL_120;
  assign _EVAL_340 = _EVAL_13 ^ 32'h20000000;
  assign _EVAL_105 = {1'b0,$signed(_EVAL_340)};
  assign _EVAL_48 = $signed(_EVAL_105) & $signed(-33'sh2000);
  assign _EVAL_271 = $signed(_EVAL_48);
  assign _EVAL_293 = $signed(_EVAL_271) == $signed(33'sh0);
  assign _EVAL_128 = _EVAL_40 | _EVAL_293;
  assign _EVAL_269 = _EVAL_323 == 6'h0;
  assign _EVAL_121 = _EVAL_2[2];
  assign _EVAL_265 = _EVAL_121 == 1'h0;
  assign _EVAL_158 = _EVAL_76[7:2];
  assign _EVAL_49 = _EVAL_323 - 6'h1;
  assign _EVAL_55 = _EVAL_2 == 3'h4;
  assign _EVAL_154 = _EVAL_258 == 6'h0;
  assign _EVAL_30 = _EVAL_276 & _EVAL_154;
  assign _EVAL_159 = 32'h1 << _EVAL_16;
  assign _EVAL_318 = _EVAL_30 ? _EVAL_159 : 32'h0;
  assign _EVAL_194 = _EVAL_196 | _EVAL_318;
  assign _EVAL_322 = _EVAL_6 <= 4'h6;
  assign _EVAL_213 = _EVAL_13 ^ 32'h80000000;
  assign _EVAL_31 = {1'b0,$signed(_EVAL_213)};
  assign _EVAL_88 = $signed(_EVAL_31) & $signed(-33'sh20000);
  assign _EVAL_28 = $signed(_EVAL_88);
  assign _EVAL_127 = $signed(_EVAL_28) == $signed(33'sh0);
  assign _EVAL_115 = _EVAL_322 & _EVAL_127;
  assign _EVAL_72 = _EVAL_16[4:3];
  assign _EVAL_355 = _EVAL_72 == 2'h1;
  assign _EVAL_270 = _EVAL_2 == 3'h1;
  assign _EVAL_353 = _EVAL & _EVAL_270;
  assign _EVAL_134 = _EVAL_6 <= 4'h2;
  assign _EVAL_236 = _EVAL_134 & _EVAL_128;
  assign _EVAL_249 = _EVAL_17 == 3'h0;
  assign _EVAL_245 = _EVAL_249 | _EVAL_11;
  assign _EVAL_79 = $signed(_EVAL_296) == $signed(33'sh0);
  assign _EVAL_203 = _EVAL_79 | _EVAL_127;
  assign _EVAL_294 = _EVAL_203 | _EVAL_290;
  assign _EVAL_23 = _EVAL_294 | _EVAL_328;
  assign _EVAL_260 = _EVAL_15 >= 4'h2;
  assign _EVAL_173 = _EVAL_260 | _EVAL_11;
  assign _EVAL_230 = _EVAL_173 == 1'h0;
  assign _EVAL_75 = _EVAL_2 == 3'h6;
  assign _EVAL_349 = _EVAL_72 == 2'h3;
  assign _EVAL_218 = _EVAL_17 <= 3'h2;
  assign _EVAL_239 = _EVAL_347 - 6'h1;
  assign _EVAL_204 = _EVAL_1 == 1'h0;
  assign _EVAL_113 = _EVAL_204 | _EVAL_11;
  assign _EVAL_177 = _EVAL_14 == _EVAL_325;
  assign _EVAL_164 = _EVAL_177 | _EVAL_11;
  assign _EVAL_179 = _EVAL_341 == 6'h0;
  assign _EVAL_280 = _EVAL_292 & _EVAL_179;
  assign _EVAL_358 = _EVAL_10 == 3'h6;
  assign _EVAL_181 = _EVAL_358 == 1'h0;
  assign _EVAL_209 = _EVAL_280 & _EVAL_181;
  assign _EVAL_244 = 32'h1 << _EVAL_9;
  assign _EVAL_195 = _EVAL_209 ? _EVAL_244 : 32'h0;
  assign _EVAL_63 = _EVAL_14 == 1'h0;
  assign _EVAL_61 = _EVAL_63 | _EVAL_12;
  assign _EVAL_107 = _EVAL_61 | _EVAL_11;
  assign _EVAL_316 = _EVAL_107 == 1'h0;
  assign _EVAL_224 = _EVAL_17 <= 3'h4;
  assign _EVAL_42 = _EVAL_224 | _EVAL_11;
  assign _EVAL_337 = _EVAL_42 == 1'h0;
  assign _EVAL_35 = _EVAL_218 | _EVAL_11;
  assign _EVAL_266 = _EVAL_196 >> _EVAL_16;
  assign _EVAL_57 = _EVAL_266[0];
  assign _EVAL_321 = _EVAL_12 == 1'h0;
  assign _EVAL_101 = _EVAL_321 | _EVAL_11;
  assign _EVAL_274 = _EVAL_101 == 1'h0;
  assign _EVAL_279 = _EVAL_10 == 3'h0;
  assign _EVAL_330 = _EVAL_57 == 1'h0;
  assign _EVAL_45 = _EVAL_330 | _EVAL_11;
  assign _EVAL_126 = _EVAL_45 == 1'h0;
  assign _EVAL_27 = _EVAL_6 == _EVAL_357;
  assign _EVAL_227 = _EVAL_27 | _EVAL_11;
  assign _EVAL_205 = _EVAL_10[0];
  assign _EVAL_261 = 23'hff << _EVAL_15;
  assign _EVAL_117 = _EVAL_261[7:0];
  assign _EVAL_272 = ~ _EVAL_117;
  assign _EVAL_240 = _EVAL_272[7:2];
  assign _EVAL_283 = _EVAL & _EVAL_75;
  assign _EVAL_332 = _EVAL_258 - 6'h1;
  assign _EVAL_78 = _EVAL_317 | _EVAL_11;
  assign _EVAL_344 = _EVAL_78 == 1'h0;
  assign _EVAL_301 = _EVAL_2 == 3'h5;
  assign _EVAL_87 = _EVAL_347 == 6'h0;
  assign _EVAL_71 = _EVAL_87 == 1'h0;
  assign _EVAL_38 = _EVAL_2 == _EVAL_233;
  assign _EVAL_345 = _EVAL_38 | _EVAL_11;
  assign _EVAL_138 = _EVAL_23 | _EVAL_185;
  assign _EVAL_253 = _EVAL_138 | _EVAL_114;
  assign _EVAL_324 = _EVAL_318 != _EVAL_195;
  assign _EVAL_53 = _EVAL_318 != 32'h0;
  assign _EVAL_257 = _EVAL_53 == 1'h0;
  assign _EVAL_39 = _EVAL_324 | _EVAL_257;
  assign _EVAL_214 = _EVAL_39 | _EVAL_11;
  assign _EVAL_346 = _EVAL_72 == 2'h0;
  assign _EVAL_86 = _EVAL_346 | _EVAL_355;
  assign _EVAL_220 = _EVAL_72 == 2'h2;
  assign _EVAL_229 = _EVAL_86 | _EVAL_220;
  assign _EVAL_145 = _EVAL_229 | _EVAL_349;
  assign _EVAL_90 = _EVAL & _EVAL_301;
  assign _EVAL_187 = ~ _EVAL_195;
  assign _EVAL_188 = _EVAL_13 & _EVAL_169;
  assign _EVAL_123 = _EVAL_188 == 32'h0;
  assign _EVAL_277 = _EVAL_10 == 3'h1;
  assign _EVAL_110 = _EVAL_3 & _EVAL_277;
  assign _EVAL_190 = _EVAL_139 + 32'h1;
  assign _EVAL_217 = _EVAL_17 != 3'h0;
  assign _EVAL_228 = _EVAL_217 | _EVAL_11;
  assign _EVAL_216 = _EVAL_227 == 1'h0;
  assign _EVAL_291 = _EVAL_10 == _EVAL_306;
  assign _EVAL_97 = _EVAL_291 | _EVAL_11;
  assign _EVAL_64 = _EVAL_228 == 1'h0;
  assign _EVAL_297 = _EVAL_269 == 1'h0;
  assign _EVAL_89 = _EVAL_145 | _EVAL_11;
  assign _EVAL_234 = _EVAL_89 == 1'h0;
  assign _EVAL_178 = _EVAL_0 == 2'h0;
  assign _EVAL_212 = _EVAL_178 | _EVAL_11;
  assign _EVAL_167 = _EVAL_212 == 1'h0;
  assign _EVAL_338 = _EVAL_9 == _EVAL_152;
  assign _EVAL_235 = _EVAL_245 == 1'h0;
  assign _EVAL_104 = _EVAL_15 == _EVAL_193;
  assign _EVAL_232 = _EVAL_104 | _EVAL_11;
  assign _EVAL_112 = _EVAL & _EVAL_297;
  assign _EVAL_109 = _EVAL_0 <= 2'h2;
  assign _EVAL_130 = _EVAL_109 | _EVAL_11;
  assign _EVAL_243 = _EVAL_130 == 1'h0;
  assign _EVAL_80 = _EVAL_3 & _EVAL_279;
  assign _EVAL_334 = _EVAL_236 | _EVAL_11;
  assign _EVAL_299 = _EVAL_142 | _EVAL_11;
  assign _EVAL_226 = _EVAL_2 == 3'h3;
  assign _EVAL_147 = _EVAL & _EVAL_226;
  assign _EVAL_314 = _EVAL_287 == 1'h0;
  assign _EVAL_20 = _EVAL_16 == _EVAL_106;
  assign _EVAL_312 = _EVAL_20 | _EVAL_11;
  assign _EVAL_254 = _EVAL_312 == 1'h0;
  assign _EVAL_124 = _EVAL_4 == _EVAL_320;
  assign _EVAL_69 = _EVAL_341 - 6'h1;
  assign _EVAL_242 = _EVAL_202 | _EVAL_11;
  assign _EVAL_60 = _EVAL_10 == 3'h2;
  assign _EVAL_96 = _EVAL_164 == 1'h0;
  assign _EVAL_354 = _EVAL_2 == 3'h0;
  assign _EVAL_198 = _EVAL_292 & _EVAL_87;
  assign _EVAL_149 = _EVAL_11 == 1'h0;
  assign _EVAL_26 = _EVAL_3 & _EVAL_71;
  assign _EVAL_201 = _EVAL_10 <= 3'h6;
  assign _EVAL_25 = _EVAL_201 | _EVAL_11;
  assign _EVAL_129 = _EVAL_25 == 1'h0;
  assign _EVAL_200 = _EVAL_242 == 1'h0;
  assign _EVAL_103 = _EVAL_318 | _EVAL_196;
  assign _EVAL_176 = _EVAL_103 >> _EVAL_9;
  assign _EVAL_50 = _EVAL_176[0];
  assign _EVAL_278 = _EVAL_50 | _EVAL_11;
  assign _EVAL_136 = _EVAL_278 == 1'h0;
  assign _EVAL_131 = _EVAL_17 == _EVAL_351;
  assign _EVAL_118 = _EVAL_131 | _EVAL_11;
  assign _EVAL_160 = _EVAL_118 == 1'h0;
  assign _EVAL_98 = _EVAL_13 == _EVAL_180;
  assign _EVAL_288 = _EVAL_98 | _EVAL_11;
  assign _EVAL_215 = _EVAL_288 == 1'h0;
  assign _EVAL_171 = _EVAL_63 | _EVAL_11;
  assign _EVAL_268 = _EVAL_115 | _EVAL_11;
  assign _EVAL_137 = _EVAL_124 | _EVAL_11;
  assign _EVAL_219 = _EVAL_137 == 1'h0;
  assign _EVAL_44 = _EVAL_253 | _EVAL_120;
  assign _EVAL_166 = _EVAL_44 | _EVAL_293;
  assign _EVAL_143 = _EVAL_322 & _EVAL_166;
  assign _EVAL_191 = _EVAL_10 == 3'h5;
  assign _EVAL_331 = _EVAL_113 == 1'h0;
  assign _EVAL_199 = _EVAL_8 == _EVAL_208;
  assign _EVAL_37 = _EVAL_199 | _EVAL_11;
  assign _EVAL_326 = _EVAL_299 == 1'h0;
  assign _EVAL_66 = _EVAL_338 | _EVAL_11;
  assign _EVAL_329 = _EVAL_66 == 1'h0;
  assign _EVAL_256 = _EVAL_0 == _EVAL_21;
  assign _EVAL_59 = _EVAL_256 | _EVAL_11;
  assign _EVAL_67 = _EVAL_59 == 1'h0;
  assign _EVAL_305 = _EVAL_2 == 3'h7;
  assign _EVAL_119 = _EVAL & _EVAL_305;
  assign _EVAL_116 = _EVAL & _EVAL_55;
  assign _EVAL_300 = _EVAL_143 | _EVAL_153;
  assign _EVAL_150 = _EVAL_0 != 2'h2;
  assign _EVAL_275 = _EVAL_150 | _EVAL_11;
  assign _EVAL_36 = _EVAL_275 == 1'h0;
  assign _EVAL_315 = _EVAL_300 | _EVAL_11;
  assign _EVAL_210 = _EVAL_345 == 1'h0;
  assign _EVAL_146 = _EVAL & _EVAL_354;
  assign _EVAL_310 = _EVAL_171 == 1'h0;
  assign _EVAL_192 = _EVAL_153 | _EVAL_11;
  assign _EVAL_170 = _EVAL_17 <= 3'h3;
  assign _EVAL_62 = _EVAL_170 | _EVAL_11;
  assign _EVAL_174 = _EVAL_62 == 1'h0;
  assign _EVAL_247 = _EVAL_3 & _EVAL_191;
  assign _EVAL_289 = _EVAL_315 == 1'h0;
  assign _EVAL_221 = _EVAL_268 == 1'h0;
  assign _EVAL_81 = _EVAL_334 == 1'h0;
  assign _EVAL_65 = _EVAL_276 & _EVAL_269;
  assign _EVAL_333 = _EVAL_232 == 1'h0;
  assign _EVAL_99 = _EVAL_214 == 1'h0;
  assign _EVAL_259 = _EVAL_3 & _EVAL_60;
  assign _EVAL_225 = _EVAL_194 & _EVAL_187;
  assign _EVAL_285 = _EVAL_97 == 1'h0;
  assign _EVAL_19 = _EVAL_37 == 1'h0;
  assign _EVAL_308 = _EVAL_192 == 1'h0;
  assign _EVAL_251 = _EVAL_10 == 3'h4;
  assign _EVAL_58 = _EVAL_3 & _EVAL_251;
  assign _EVAL_83 = _EVAL_35 == 1'h0;
  assign _EVAL_156 = _EVAL_123 | _EVAL_11;
  assign _EVAL_157 = _EVAL_3 & _EVAL_358;
  assign _EVAL_68 = _EVAL_156 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_21 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_106 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_139 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_152 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_180 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_193 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_196 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_233 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_258 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_306 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_320 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_323 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_325 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_341 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_347 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_351 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_357 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_7) begin
    if (_EVAL_198) begin
      _EVAL_21 <= _EVAL_0;
    end
    if (_EVAL_65) begin
      _EVAL_106 <= _EVAL_16;
    end
    if (_EVAL_11) begin
      _EVAL_139 <= 32'h0;
    end else begin
      if (_EVAL_197) begin
        _EVAL_139 <= 32'h0;
      end else begin
        _EVAL_139 <= _EVAL_190;
      end
    end
    if (_EVAL_198) begin
      _EVAL_152 <= _EVAL_9;
    end
    if (_EVAL_65) begin
      _EVAL_180 <= _EVAL_13;
    end
    if (_EVAL_198) begin
      _EVAL_193 <= _EVAL_15;
    end
    if (_EVAL_11) begin
      _EVAL_196 <= 32'h0;
    end else begin
      _EVAL_196 <= _EVAL_225;
    end
    if (_EVAL_65) begin
      _EVAL_233 <= _EVAL_2;
    end
    if (_EVAL_11) begin
      _EVAL_258 <= 6'h0;
    end else begin
      if (_EVAL_276) begin
        if (_EVAL_154) begin
          if (_EVAL_265) begin
            _EVAL_258 <= _EVAL_158;
          end else begin
            _EVAL_258 <= 6'h0;
          end
        end else begin
          _EVAL_258 <= _EVAL_332;
        end
      end
    end
    if (_EVAL_198) begin
      _EVAL_306 <= _EVAL_10;
    end
    if (_EVAL_198) begin
      _EVAL_320 <= _EVAL_4;
    end
    if (_EVAL_11) begin
      _EVAL_323 <= 6'h0;
    end else begin
      if (_EVAL_276) begin
        if (_EVAL_269) begin
          if (_EVAL_265) begin
            _EVAL_323 <= _EVAL_158;
          end else begin
            _EVAL_323 <= 6'h0;
          end
        end else begin
          _EVAL_323 <= _EVAL_49;
        end
      end
    end
    if (_EVAL_198) begin
      _EVAL_325 <= _EVAL_14;
    end
    if (_EVAL_11) begin
      _EVAL_341 <= 6'h0;
    end else begin
      if (_EVAL_292) begin
        if (_EVAL_179) begin
          if (_EVAL_205) begin
            _EVAL_341 <= _EVAL_240;
          end else begin
            _EVAL_341 <= 6'h0;
          end
        end else begin
          _EVAL_341 <= _EVAL_69;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_347 <= 6'h0;
    end else begin
      if (_EVAL_292) begin
        if (_EVAL_87) begin
          if (_EVAL_205) begin
            _EVAL_347 <= _EVAL_240;
          end else begin
            _EVAL_347 <= 6'h0;
          end
        end else begin
          _EVAL_347 <= _EVAL_239;
        end
      end
    end
    if (_EVAL_65) begin
      _EVAL_351 <= _EVAL_17;
    end
    if (_EVAL_65) begin
      _EVAL_357 <= _EVAL_6;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74db03c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_329) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(962d759c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82d7a034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59789c6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(558776fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5df99af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fa6f74d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ae247e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(145aab47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75e70d47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25a50a15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4329642d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4df54c08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53d908e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f95c90e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d10a15d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffc0635d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_337) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d7b074f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b57f039)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_333) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d8efed1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3c2b4d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8080103d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67067536)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89c5a392)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1e61337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dbb9507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef58725c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa75cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b09e6aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccc5ad20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54ecac37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae777c29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee02a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d277dee8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddd85367)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(605b583a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6b51c2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ed8fbca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7372fc00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2e1961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0c4e820)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe2ed2f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6c4a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6eed756)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4ffdf11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b155c999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_310) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15862e73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cd77937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88ab9ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d8b3a9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30f39ccf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ae3f55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57fd17bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff9b1253)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bba8db1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_333) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68f78eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(697c890e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_310) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38cd54cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fed96f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d14dbdea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d227dcf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa2c54f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42220f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56170f0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed03ca9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a13b679f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_329) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a856154d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72b639d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb8ffbdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dc16c3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e83381)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46a30c0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9c70d5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd7759d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e5cacf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3803e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d556c663)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6994f50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82383f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f737ac6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5f7af5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88180a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54764ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbbfb924)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(697ce0bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2e038b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e4bc5e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42908a27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
