//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_47(
  input  [1:0]  _EVAL,
  output [3:0]  _EVAL_0,
  input  [5:0]  _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output [1:0]  _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  output        _EVAL_11,
  output [5:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [63:0] _EVAL_14,
  output [3:0]  _EVAL_15,
  output [5:0]  _EVAL_16,
  input  [3:0]  _EVAL_17,
  input  [2:0]  _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  input  [5:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output [2:0]  _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  output [2:0]  _EVAL_28,
  input         _EVAL_29,
  input  [3:0]  _EVAL_30,
  output [7:0]  _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input  [31:0] _EVAL_34,
  output [31:0] _EVAL_35,
  output        _EVAL_36,
  input         _EVAL_37,
  output [63:0] _EVAL_38,
  output [31:0] _EVAL_39,
  output        _EVAL_40
);
  wire [3:0] Repeater__EVAL;
  wire  Repeater__EVAL_0;
  wire [5:0] Repeater__EVAL_1;
  wire  Repeater__EVAL_2;
  wire [1:0] Repeater__EVAL_3;
  wire  Repeater__EVAL_4;
  wire [2:0] Repeater__EVAL_5;
  wire [1:0] Repeater__EVAL_6;
  wire [2:0] Repeater__EVAL_7;
  wire  Repeater__EVAL_8;
  wire  Repeater__EVAL_9;
  wire  Repeater__EVAL_10;
  wire  Repeater__EVAL_11;
  wire [5:0] Repeater__EVAL_12;
  wire [3:0] Repeater__EVAL_13;
  wire  Repeater__EVAL_14;
  wire  Repeater__EVAL_15;
  wire  Repeater__EVAL_16;
  wire [63:0] Repeater__EVAL_17;
  wire  Repeater__EVAL_18;
  wire  Repeater__EVAL_19;
  wire  Repeater__EVAL_20;
  wire [63:0] Repeater__EVAL_21;
  reg  _EVAL_42;
  reg [31:0] _RAND_0;
  reg  _EVAL_43;
  reg [31:0] _RAND_1;
  reg  _EVAL_45;
  reg [31:0] _RAND_2;
  reg  _EVAL_50;
  reg [31:0] _RAND_3;
  reg  _EVAL_52;
  reg [31:0] _RAND_4;
  reg  _EVAL_58;
  reg [31:0] _RAND_5;
  reg  _EVAL_77;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_80;
  reg [31:0] _RAND_7;
  reg  _EVAL_91;
  reg [31:0] _RAND_8;
  reg  _EVAL_92;
  reg [31:0] _RAND_9;
  reg  _EVAL_96;
  reg [31:0] _RAND_10;
  reg  _EVAL_104;
  reg [31:0] _RAND_11;
  reg  _EVAL_113;
  reg [31:0] _RAND_12;
  reg  _EVAL_116;
  reg [31:0] _RAND_13;
  reg  _EVAL_126;
  reg [31:0] _RAND_14;
  reg  _EVAL_127;
  reg [31:0] _RAND_15;
  reg  _EVAL_129;
  reg [31:0] _RAND_16;
  reg  _EVAL_142;
  reg [31:0] _RAND_17;
  reg  _EVAL_148;
  reg [31:0] _RAND_18;
  reg  _EVAL_149;
  reg [31:0] _RAND_19;
  reg  _EVAL_150;
  reg [31:0] _RAND_20;
  reg  _EVAL_159;
  reg [31:0] _RAND_21;
  reg  _EVAL_169;
  reg [31:0] _RAND_22;
  reg  _EVAL_172;
  reg [31:0] _RAND_23;
  reg  _EVAL_175;
  reg [31:0] _RAND_24;
  reg  _EVAL_177;
  reg [31:0] _RAND_25;
  reg  _EVAL_180;
  reg [31:0] _RAND_26;
  reg  _EVAL_199;
  reg [31:0] _RAND_27;
  reg [31:0] _EVAL_201;
  reg [31:0] _RAND_28;
  reg  _EVAL_204;
  reg [31:0] _RAND_29;
  reg  _EVAL_208;
  reg [31:0] _RAND_30;
  reg  _EVAL_216;
  reg [31:0] _RAND_31;
  reg  _EVAL_225;
  reg [31:0] _RAND_32;
  reg  _EVAL_232;
  reg [31:0] _RAND_33;
  reg  _EVAL_235;
  reg [31:0] _RAND_34;
  reg  _EVAL_237;
  reg [31:0] _RAND_35;
  reg  _EVAL_241;
  reg [31:0] _RAND_36;
  reg  _EVAL_243;
  reg [31:0] _RAND_37;
  reg  _EVAL_244;
  reg [31:0] _RAND_38;
  wire  _EVAL_160;
  wire [5:0] _EVAL_118;
  wire  _EVAL_81;
  wire  _EVAL_210;
  wire  _EVAL_207;
  wire  _EVAL_193;
  wire  _EVAL_109;
  wire  _EVAL_176;
  wire  _EVAL_230;
  wire  _EVAL_236;
  wire  _EVAL_56;
  wire  _EVAL_87;
  wire  _EVAL_137;
  wire  _EVAL_222;
  wire  _EVAL_112;
  wire  _EVAL_200;
  wire  _EVAL_212;
  wire  _EVAL_97;
  wire  _EVAL_74;
  wire  _EVAL_78;
  wire  _EVAL_60;
  wire  _EVAL_164;
  wire  _EVAL_102;
  wire  _EVAL_144;
  wire  _EVAL_107;
  wire  _EVAL_228;
  wire  _EVAL_55;
  wire  _EVAL_182;
  wire  _EVAL_188;
  wire  _EVAL_66;
  wire  _EVAL_95;
  wire  _EVAL_145;
  wire  _EVAL_125;
  wire  _EVAL_248;
  wire  _EVAL_90;
  wire  _EVAL_53;
  wire [1:0] _EVAL_46;
  wire [3:0] _EVAL_233;
  wire [2:0] _EVAL_124;
  wire [2:0] _EVAL_73;
  wire  _EVAL_114;
  wire  _EVAL_198;
  wire  _EVAL_111;
  wire  _EVAL_86;
  wire  _EVAL_245;
  wire  _EVAL_101;
  wire  _EVAL_183;
  wire  _EVAL_223;
  wire  _EVAL_231;
  wire  _EVAL_179;
  wire  _EVAL_168;
  wire  _EVAL_132;
  wire  _EVAL_63;
  wire  _EVAL_221;
  wire [2:0] _EVAL_246;
  wire  _EVAL_65;
  wire  _EVAL_57;
  wire  _EVAL_249;
  wire  _EVAL_121;
  wire  _EVAL_110;
  wire  _EVAL_185;
  wire  _EVAL_234;
  wire [31:0] _EVAL_156;
  wire [31:0] _EVAL_224;
  wire [63:0] _EVAL_173;
  wire [31:0] _EVAL_123;
  wire [3:0] _EVAL_171;
  wire [17:0] _EVAL_202;
  wire [2:0] _EVAL_158;
  wire [2:0] _EVAL_59;
  wire  _EVAL_136;
  wire  _EVAL_184;
  wire  _EVAL_214;
  wire  _EVAL_120;
  wire  _EVAL_240;
  wire [17:0] _EVAL_88;
  wire [2:0] _EVAL_106;
  wire [2:0] _EVAL_68;
  wire  _EVAL_227;
  wire  _EVAL_197;
  wire  _EVAL_94;
  wire [31:0] _EVAL_48;
  wire  _EVAL_213;
  wire  _EVAL_161;
  wire  _EVAL_247;
  wire  _EVAL_252;
  wire  _EVAL_49;
  wire  _EVAL_82;
  wire  _EVAL_203;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_75;
  wire [3:0] _EVAL_157;
  wire [7:0] _EVAL_154;
  wire [7:0] _EVAL_205;
  wire  _EVAL_181;
  wire  _EVAL_128;
  wire  _EVAL_147;
  wire  _EVAL_79;
  wire  _EVAL_250;
  wire  _EVAL_217;
  wire  _EVAL_47;
  wire  _EVAL_117;
  wire  _EVAL_69;
  wire  _EVAL_85;
  wire  _EVAL_220;
  wire  _EVAL_194;
  wire  _EVAL_84;
  wire  _EVAL_54;
  wire  _EVAL_146;
  wire  _EVAL_72;
  wire  _EVAL_71;
  wire  _EVAL_174;
  wire  _EVAL_51;
  wire  _EVAL_219;
  wire  _EVAL_191;
  wire  _EVAL_41;
  wire  _EVAL_152;
  wire  _EVAL_170;
  wire  _EVAL_215;
  wire  _EVAL_251;
  wire  _EVAL_135;
  wire [7:0] _EVAL_209;
  wire [31:0] _EVAL_133;
  wire  _EVAL_226;
  wire  _EVAL_178;
  wire  _EVAL_134;
  wire  _EVAL_108;
  wire  _EVAL_122;
  wire  _EVAL_44;
  wire  _EVAL_83;
  wire  _EVAL_190;
  SiFive__EVAL_46 Repeater (
    ._EVAL(Repeater__EVAL),
    ._EVAL_0(Repeater__EVAL_0),
    ._EVAL_1(Repeater__EVAL_1),
    ._EVAL_2(Repeater__EVAL_2),
    ._EVAL_3(Repeater__EVAL_3),
    ._EVAL_4(Repeater__EVAL_4),
    ._EVAL_5(Repeater__EVAL_5),
    ._EVAL_6(Repeater__EVAL_6),
    ._EVAL_7(Repeater__EVAL_7),
    ._EVAL_8(Repeater__EVAL_8),
    ._EVAL_9(Repeater__EVAL_9),
    ._EVAL_10(Repeater__EVAL_10),
    ._EVAL_11(Repeater__EVAL_11),
    ._EVAL_12(Repeater__EVAL_12),
    ._EVAL_13(Repeater__EVAL_13),
    ._EVAL_14(Repeater__EVAL_14),
    ._EVAL_15(Repeater__EVAL_15),
    ._EVAL_16(Repeater__EVAL_16),
    ._EVAL_17(Repeater__EVAL_17),
    ._EVAL_18(Repeater__EVAL_18),
    ._EVAL_19(Repeater__EVAL_19),
    ._EVAL_20(Repeater__EVAL_20),
    ._EVAL_21(Repeater__EVAL_21)
  );
  assign _EVAL_160 = _EVAL_104 == 1'h0;
  assign _EVAL_118 = Repeater__EVAL_1;
  assign _EVAL_81 = 6'h1 == _EVAL_118 ? _EVAL_175 : _EVAL_225;
  assign _EVAL_210 = 6'h2 == _EVAL_118 ? _EVAL_113 : _EVAL_81;
  assign _EVAL_207 = 6'h3 == _EVAL_118 ? _EVAL_180 : _EVAL_210;
  assign _EVAL_193 = 6'h4 == _EVAL_118 ? _EVAL_45 : _EVAL_207;
  assign _EVAL_109 = 6'h5 == _EVAL_118 ? _EVAL_232 : _EVAL_193;
  assign _EVAL_176 = 6'h6 == _EVAL_118 ? _EVAL_91 : _EVAL_109;
  assign _EVAL_230 = 6'h7 == _EVAL_118 ? _EVAL_52 : _EVAL_176;
  assign _EVAL_236 = 6'h8 == _EVAL_118 ? _EVAL_129 : _EVAL_230;
  assign _EVAL_56 = 6'h9 == _EVAL_118 ? _EVAL_237 : _EVAL_236;
  assign _EVAL_87 = 6'ha == _EVAL_118 ? _EVAL_43 : _EVAL_56;
  assign _EVAL_137 = 6'hb == _EVAL_118 ? _EVAL_244 : _EVAL_87;
  assign _EVAL_222 = 6'hc == _EVAL_118 ? _EVAL_142 : _EVAL_137;
  assign _EVAL_112 = 6'hd == _EVAL_118 ? _EVAL_172 : _EVAL_222;
  assign _EVAL_200 = 6'he == _EVAL_118 ? _EVAL_169 : _EVAL_112;
  assign _EVAL_212 = 6'hf == _EVAL_118 ? _EVAL_241 : _EVAL_200;
  assign _EVAL_97 = 6'h10 == _EVAL_118 ? _EVAL_126 : _EVAL_212;
  assign _EVAL_74 = 6'h11 == _EVAL_118 ? _EVAL_149 : _EVAL_97;
  assign _EVAL_78 = 6'h12 == _EVAL_118 ? _EVAL_150 : _EVAL_74;
  assign _EVAL_60 = 6'h13 == _EVAL_118 ? _EVAL_177 : _EVAL_78;
  assign _EVAL_164 = 6'h14 == _EVAL_118 ? _EVAL_159 : _EVAL_60;
  assign _EVAL_102 = 6'h15 == _EVAL_118 ? _EVAL_42 : _EVAL_164;
  assign _EVAL_144 = 6'h16 == _EVAL_118 ? _EVAL_208 : _EVAL_102;
  assign _EVAL_107 = 6'h17 == _EVAL_118 ? _EVAL_58 : _EVAL_144;
  assign _EVAL_228 = 6'h18 == _EVAL_118 ? _EVAL_199 : _EVAL_107;
  assign _EVAL_55 = 6'h19 == _EVAL_118 ? _EVAL_216 : _EVAL_228;
  assign _EVAL_182 = 6'h1a == _EVAL_118 ? _EVAL_116 : _EVAL_55;
  assign _EVAL_188 = 6'h1b == _EVAL_118 ? _EVAL_235 : _EVAL_182;
  assign _EVAL_66 = 6'h1c == _EVAL_118 ? _EVAL_148 : _EVAL_188;
  assign _EVAL_95 = 6'h1d == _EVAL_118 ? _EVAL_127 : _EVAL_66;
  assign _EVAL_145 = 6'h1e == _EVAL_118 ? _EVAL_204 : _EVAL_95;
  assign _EVAL_125 = 6'h1f == _EVAL_118 ? _EVAL_243 : _EVAL_145;
  assign _EVAL_248 = 6'h20 == _EVAL_118 ? _EVAL_92 : _EVAL_125;
  assign _EVAL_90 = _EVAL_160 ? _EVAL_248 : _EVAL_50;
  assign _EVAL_53 = _EVAL_17 >= 4'h3;
  assign _EVAL_46 = _EVAL_17[1:0];
  assign _EVAL_233 = 4'h1 << _EVAL_46;
  assign _EVAL_124 = _EVAL_233[2:0];
  assign _EVAL_73 = _EVAL_124 | 3'h1;
  assign _EVAL_114 = _EVAL_73[2];
  assign _EVAL_198 = _EVAL_34[2];
  assign _EVAL_111 = _EVAL_114 & _EVAL_198;
  assign _EVAL_86 = _EVAL_53 | _EVAL_111;
  assign _EVAL_245 = _EVAL_73[1];
  assign _EVAL_101 = _EVAL_34[1];
  assign _EVAL_183 = _EVAL_198 & _EVAL_101;
  assign _EVAL_223 = _EVAL_245 & _EVAL_183;
  assign _EVAL_231 = _EVAL_86 | _EVAL_223;
  assign _EVAL_179 = _EVAL_73[0];
  assign _EVAL_168 = _EVAL_34[0];
  assign _EVAL_132 = _EVAL_183 & _EVAL_168;
  assign _EVAL_63 = _EVAL_179 & _EVAL_132;
  assign _EVAL_221 = _EVAL_231 | _EVAL_63;
  assign _EVAL_246 = Repeater__EVAL_7;
  assign _EVAL_65 = _EVAL_246[0];
  assign _EVAL_57 = _EVAL_101 == 1'h0;
  assign _EVAL_249 = _EVAL_198 & _EVAL_57;
  assign _EVAL_121 = _EVAL_249 & _EVAL_168;
  assign _EVAL_110 = _EVAL_179 & _EVAL_121;
  assign _EVAL_185 = _EVAL_18[2];
  assign _EVAL_234 = _EVAL_185 == 1'h0;
  assign _EVAL_156 = Repeater__EVAL_17[63:32];
  assign _EVAL_224 = _EVAL_14[31:0];
  assign _EVAL_173 = {_EVAL_156,_EVAL_224};
  assign _EVAL_123 = _EVAL_173[31:0];
  assign _EVAL_171 = Repeater__EVAL;
  assign _EVAL_202 = 18'h7 << _EVAL_171;
  assign _EVAL_158 = _EVAL_202[2:0];
  assign _EVAL_59 = ~ _EVAL_158;
  assign _EVAL_136 = _EVAL_59[2:2];
  assign _EVAL_184 = _EVAL_104 == _EVAL_136;
  assign _EVAL_214 = _EVAL_65 == 1'h0;
  assign _EVAL_120 = _EVAL_184 | _EVAL_214;
  assign _EVAL_240 = ~ _EVAL_136;
  assign _EVAL_88 = 18'h7 << _EVAL_17;
  assign _EVAL_106 = _EVAL_88[2:0];
  assign _EVAL_68 = ~ _EVAL_106;
  assign _EVAL_227 = _EVAL_68[2:2];
  assign _EVAL_197 = _EVAL_96 & _EVAL_227;
  assign _EVAL_94 = _EVAL_197 == 1'h0;
  assign _EVAL_48 = _EVAL_94 ? _EVAL_7 : _EVAL_201;
  assign _EVAL_213 = _EVAL_168 == 1'h0;
  assign _EVAL_161 = _EVAL_183 & _EVAL_213;
  assign _EVAL_247 = _EVAL_179 & _EVAL_161;
  assign _EVAL_252 = _EVAL_231 | _EVAL_247;
  assign _EVAL_49 = _EVAL_249 & _EVAL_213;
  assign _EVAL_82 = _EVAL_96 == _EVAL_227;
  assign _EVAL_203 = _EVAL_234 == 1'h0;
  assign _EVAL_238 = _EVAL_82 | _EVAL_203;
  assign _EVAL_239 = _EVAL_23 | _EVAL_77;
  assign _EVAL_75 = _EVAL_90 & _EVAL_240;
  assign _EVAL_157 = _EVAL_94 ? _EVAL_30 : _EVAL_80;
  assign _EVAL_154 = {_EVAL_30,_EVAL_157};
  assign _EVAL_205 = _EVAL_234 ? _EVAL_154 : 8'hff;
  assign _EVAL_181 = Repeater__EVAL_11;
  assign _EVAL_128 = _EVAL_179 & _EVAL_49;
  assign _EVAL_147 = _EVAL_198 == 1'h0;
  assign _EVAL_79 = _EVAL_147 & _EVAL_101;
  assign _EVAL_250 = _EVAL_79 & _EVAL_168;
  assign _EVAL_217 = _EVAL_179 & _EVAL_250;
  assign _EVAL_47 = _EVAL_147 & _EVAL_57;
  assign _EVAL_117 = _EVAL_47 & _EVAL_168;
  assign _EVAL_69 = _EVAL_179 & _EVAL_117;
  assign _EVAL_85 = _EVAL_245 & _EVAL_249;
  assign _EVAL_220 = _EVAL_86 | _EVAL_85;
  assign _EVAL_194 = _EVAL_220 | _EVAL_110;
  assign _EVAL_84 = _EVAL_220 | _EVAL_128;
  assign _EVAL_54 = _EVAL_114 & _EVAL_147;
  assign _EVAL_146 = _EVAL_53 | _EVAL_54;
  assign _EVAL_72 = _EVAL_245 & _EVAL_79;
  assign _EVAL_71 = _EVAL_146 | _EVAL_72;
  assign _EVAL_174 = _EVAL_71 | _EVAL_217;
  assign _EVAL_51 = _EVAL_79 & _EVAL_213;
  assign _EVAL_219 = _EVAL_179 & _EVAL_51;
  assign _EVAL_191 = _EVAL_71 | _EVAL_219;
  assign _EVAL_41 = _EVAL_245 & _EVAL_47;
  assign _EVAL_152 = _EVAL_146 | _EVAL_41;
  assign _EVAL_170 = _EVAL_152 | _EVAL_69;
  assign _EVAL_215 = _EVAL_47 & _EVAL_213;
  assign _EVAL_251 = _EVAL_179 & _EVAL_215;
  assign _EVAL_135 = _EVAL_152 | _EVAL_251;
  assign _EVAL_209 = {_EVAL_221,_EVAL_252,_EVAL_194,_EVAL_84,_EVAL_174,_EVAL_191,_EVAL_170,_EVAL_135};
  assign _EVAL_133 = _EVAL_173[63:32];
  assign _EVAL_226 = _EVAL_104 + 1'h1;
  assign _EVAL_178 = _EVAL_238 == 1'h0;
  assign _EVAL_134 = _EVAL_33 | _EVAL_178;
  assign _EVAL_108 = _EVAL_96 + 1'h1;
  assign _EVAL_122 = _EVAL_134 & _EVAL_19;
  assign _EVAL_44 = _EVAL_4 & _EVAL_181;
  assign _EVAL_83 = _EVAL_122 & _EVAL_178;
  assign _EVAL_190 = _EVAL_75 | _EVAL_104;
  assign _EVAL_15 = _EVAL_17;
  assign Repeater__EVAL_13 = _EVAL_13;
  assign _EVAL_31 = _EVAL_209 & _EVAL_205;
  assign _EVAL_35 = _EVAL_34;
  assign Repeater__EVAL_15 = _EVAL_120 == 1'h0;
  assign Repeater__EVAL_10 = _EVAL_24;
  assign Repeater__EVAL_3 = _EVAL;
  assign _EVAL_26 = _EVAL_19 & _EVAL_238;
  assign _EVAL_22 = _EVAL_18;
  assign Repeater__EVAL_0 = _EVAL_8;
  assign _EVAL_11 = Repeater__EVAL_19;
  assign _EVAL_39 = _EVAL_190 ? _EVAL_133 : _EVAL_123;
  assign Repeater__EVAL_4 = _EVAL_37;
  assign _EVAL_0 = Repeater__EVAL;
  assign _EVAL_27 = _EVAL_33 | _EVAL_178;
  assign Repeater__EVAL_21 = _EVAL_14;
  assign _EVAL_3 = Repeater__EVAL_11;
  assign Repeater__EVAL_8 = _EVAL_32;
  assign Repeater__EVAL_2 = _EVAL_29;
  assign _EVAL_16 = _EVAL_1;
  assign _EVAL_38 = {_EVAL_7,_EVAL_48};
  assign _EVAL_25 = Repeater__EVAL_7;
  assign Repeater__EVAL_12 = _EVAL_21;
  assign _EVAL_28 = _EVAL_9;
  assign _EVAL_36 = Repeater__EVAL_14;
  assign _EVAL_2 = Repeater__EVAL_20;
  assign Repeater__EVAL_5 = _EVAL_10;
  assign _EVAL_20 = Repeater__EVAL_9;
  assign _EVAL_6 = Repeater__EVAL_6;
  assign _EVAL_12 = Repeater__EVAL_1;
  assign _EVAL_40 = _EVAL_23 | _EVAL_77;
  assign Repeater__EVAL_18 = _EVAL_4;
  assign Repeater__EVAL_16 = _EVAL_5;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_42 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_43 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_45 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_50 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_52 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_58 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_77 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_80 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_91 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_92 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_96 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_104 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_113 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_116 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_126 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_127 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_129 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_142 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_148 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_149 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_150 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_159 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_169 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_172 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_175 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_177 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_180 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_199 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_201 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_204 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_208 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_216 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_225 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_232 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_235 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_237 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_241 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_243 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_244 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_5) begin
    if (_EVAL_122) begin
      if (6'h15 == _EVAL_1) begin
        _EVAL_42 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'ha == _EVAL_1) begin
        _EVAL_43 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h4 == _EVAL_1) begin
        _EVAL_45 <= _EVAL_198;
      end
    end
    if (_EVAL_160) begin
      if (6'h20 == _EVAL_118) begin
        _EVAL_50 <= _EVAL_92;
      end else begin
        if (6'h1f == _EVAL_118) begin
          _EVAL_50 <= _EVAL_243;
        end else begin
          if (6'h1e == _EVAL_118) begin
            _EVAL_50 <= _EVAL_204;
          end else begin
            if (6'h1d == _EVAL_118) begin
              _EVAL_50 <= _EVAL_127;
            end else begin
              if (6'h1c == _EVAL_118) begin
                _EVAL_50 <= _EVAL_148;
              end else begin
                if (6'h1b == _EVAL_118) begin
                  _EVAL_50 <= _EVAL_235;
                end else begin
                  if (6'h1a == _EVAL_118) begin
                    _EVAL_50 <= _EVAL_116;
                  end else begin
                    if (6'h19 == _EVAL_118) begin
                      _EVAL_50 <= _EVAL_216;
                    end else begin
                      if (6'h18 == _EVAL_118) begin
                        _EVAL_50 <= _EVAL_199;
                      end else begin
                        if (6'h17 == _EVAL_118) begin
                          _EVAL_50 <= _EVAL_58;
                        end else begin
                          if (6'h16 == _EVAL_118) begin
                            _EVAL_50 <= _EVAL_208;
                          end else begin
                            if (6'h15 == _EVAL_118) begin
                              _EVAL_50 <= _EVAL_42;
                            end else begin
                              if (6'h14 == _EVAL_118) begin
                                _EVAL_50 <= _EVAL_159;
                              end else begin
                                if (6'h13 == _EVAL_118) begin
                                  _EVAL_50 <= _EVAL_177;
                                end else begin
                                  if (6'h12 == _EVAL_118) begin
                                    _EVAL_50 <= _EVAL_150;
                                  end else begin
                                    if (6'h11 == _EVAL_118) begin
                                      _EVAL_50 <= _EVAL_149;
                                    end else begin
                                      if (6'h10 == _EVAL_118) begin
                                        _EVAL_50 <= _EVAL_126;
                                      end else begin
                                        if (6'hf == _EVAL_118) begin
                                          _EVAL_50 <= _EVAL_241;
                                        end else begin
                                          if (6'he == _EVAL_118) begin
                                            _EVAL_50 <= _EVAL_169;
                                          end else begin
                                            if (6'hd == _EVAL_118) begin
                                              _EVAL_50 <= _EVAL_172;
                                            end else begin
                                              if (6'hc == _EVAL_118) begin
                                                _EVAL_50 <= _EVAL_142;
                                              end else begin
                                                if (6'hb == _EVAL_118) begin
                                                  _EVAL_50 <= _EVAL_244;
                                                end else begin
                                                  if (6'ha == _EVAL_118) begin
                                                    _EVAL_50 <= _EVAL_43;
                                                  end else begin
                                                    if (6'h9 == _EVAL_118) begin
                                                      _EVAL_50 <= _EVAL_237;
                                                    end else begin
                                                      if (6'h8 == _EVAL_118) begin
                                                        _EVAL_50 <= _EVAL_129;
                                                      end else begin
                                                        if (6'h7 == _EVAL_118) begin
                                                          _EVAL_50 <= _EVAL_52;
                                                        end else begin
                                                          if (6'h6 == _EVAL_118) begin
                                                            _EVAL_50 <= _EVAL_91;
                                                          end else begin
                                                            if (6'h5 == _EVAL_118) begin
                                                              _EVAL_50 <= _EVAL_232;
                                                            end else begin
                                                              if (6'h4 == _EVAL_118) begin
                                                                _EVAL_50 <= _EVAL_45;
                                                              end else begin
                                                                if (6'h3 == _EVAL_118) begin
                                                                  _EVAL_50 <= _EVAL_180;
                                                                end else begin
                                                                  if (6'h2 == _EVAL_118) begin
                                                                    _EVAL_50 <= _EVAL_113;
                                                                  end else begin
                                                                    if (6'h1 == _EVAL_118) begin
                                                                      _EVAL_50 <= _EVAL_175;
                                                                    end else begin
                                                                      _EVAL_50 <= _EVAL_225;
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_122) begin
      if (6'h7 == _EVAL_1) begin
        _EVAL_52 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h17 == _EVAL_1) begin
        _EVAL_58 <= _EVAL_198;
      end
    end
    if (_EVAL_32) begin
      _EVAL_77 <= 1'h0;
    end else begin
      if (_EVAL_122) begin
        if (_EVAL_238) begin
          _EVAL_77 <= 1'h0;
        end else begin
          _EVAL_77 <= _EVAL_239;
        end
      end
    end
    if (_EVAL_83) begin
      if (_EVAL_94) begin
        _EVAL_80 <= _EVAL_30;
      end
    end
    if (_EVAL_122) begin
      if (6'h6 == _EVAL_1) begin
        _EVAL_91 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h20 == _EVAL_1) begin
        _EVAL_92 <= _EVAL_198;
      end
    end
    if (_EVAL_32) begin
      _EVAL_96 <= 1'h0;
    end else begin
      if (_EVAL_122) begin
        if (_EVAL_238) begin
          _EVAL_96 <= 1'h0;
        end else begin
          _EVAL_96 <= _EVAL_108;
        end
      end
    end
    if (_EVAL_32) begin
      _EVAL_104 <= 1'h0;
    end else begin
      if (_EVAL_44) begin
        if (_EVAL_120) begin
          _EVAL_104 <= 1'h0;
        end else begin
          _EVAL_104 <= _EVAL_226;
        end
      end
    end
    if (_EVAL_122) begin
      if (6'h2 == _EVAL_1) begin
        _EVAL_113 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h1a == _EVAL_1) begin
        _EVAL_116 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h10 == _EVAL_1) begin
        _EVAL_126 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h1d == _EVAL_1) begin
        _EVAL_127 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h8 == _EVAL_1) begin
        _EVAL_129 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'hc == _EVAL_1) begin
        _EVAL_142 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h1c == _EVAL_1) begin
        _EVAL_148 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h11 == _EVAL_1) begin
        _EVAL_149 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h12 == _EVAL_1) begin
        _EVAL_150 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h14 == _EVAL_1) begin
        _EVAL_159 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'he == _EVAL_1) begin
        _EVAL_169 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'hd == _EVAL_1) begin
        _EVAL_172 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h1 == _EVAL_1) begin
        _EVAL_175 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h13 == _EVAL_1) begin
        _EVAL_177 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h3 == _EVAL_1) begin
        _EVAL_180 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h18 == _EVAL_1) begin
        _EVAL_199 <= _EVAL_198;
      end
    end
    if (_EVAL_83) begin
      if (_EVAL_94) begin
        _EVAL_201 <= _EVAL_7;
      end
    end
    if (_EVAL_122) begin
      if (6'h1e == _EVAL_1) begin
        _EVAL_204 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h16 == _EVAL_1) begin
        _EVAL_208 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h19 == _EVAL_1) begin
        _EVAL_216 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h0 == _EVAL_1) begin
        _EVAL_225 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h5 == _EVAL_1) begin
        _EVAL_232 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h1b == _EVAL_1) begin
        _EVAL_235 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h9 == _EVAL_1) begin
        _EVAL_237 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'hf == _EVAL_1) begin
        _EVAL_241 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'h1f == _EVAL_1) begin
        _EVAL_243 <= _EVAL_198;
      end
    end
    if (_EVAL_122) begin
      if (6'hb == _EVAL_1) begin
        _EVAL_244 <= _EVAL_198;
      end
    end
  end
endmodule
