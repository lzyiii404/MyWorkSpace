//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_41_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [6:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [6:0]  _EVAL_7,
  input  [29:0] _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input  [7:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_34;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_35;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_45;
  reg [31:0] _RAND_2;
  reg [6:0] _EVAL_82;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_99;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_104;
  reg [31:0] _RAND_5;
  reg  _EVAL_127;
  reg [31:0] _RAND_6;
  reg [72:0] _EVAL_179;
  reg [95:0] _RAND_7;
  reg  _EVAL_185;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_245;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_254;
  reg [31:0] _RAND_10;
  reg [29:0] _EVAL_255;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_261;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_279;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_299;
  reg [31:0] _RAND_14;
  reg [4:0] _EVAL_301;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_387;
  reg [31:0] _RAND_16;
  wire [1:0] _EVAL_353;
  wire [3:0] _EVAL_399;
  wire [2:0] _EVAL_222;
  wire [2:0] _EVAL_216;
  wire  _EVAL_206;
  wire  _EVAL_123;
  wire  _EVAL_170;
  wire  _EVAL_282;
  wire  _EVAL_164;
  wire  _EVAL_152;
  wire [3:0] _EVAL_325;
  wire  _EVAL_109;
  wire [2:0] _EVAL_390;
  wire  _EVAL_329;
  wire  _EVAL_260;
  wire  _EVAL_81;
  wire  _EVAL_307;
  wire  _EVAL_246;
  wire  _EVAL_113;
  wire [3:0] _EVAL_73;
  wire  _EVAL_252;
  wire [2:0] _EVAL_225;
  wire  _EVAL_314;
  wire  _EVAL_76;
  wire  _EVAL_309;
  wire  _EVAL_150;
  wire  _EVAL_50;
  wire  _EVAL_328;
  wire  _EVAL_358;
  wire  _EVAL_343;
  wire  _EVAL_98;
  wire [29:0] _EVAL_258;
  wire [30:0] _EVAL_338;
  wire [30:0] _EVAL_223;
  wire [30:0] _EVAL_121;
  wire  _EVAL_384;
  wire [29:0] _EVAL_80;
  wire [30:0] _EVAL_288;
  wire [30:0] _EVAL_21;
  wire [30:0] _EVAL_286;
  wire  _EVAL_162;
  wire  _EVAL_93;
  wire  _EVAL_171;
  wire  _EVAL_268;
  wire  _EVAL_62;
  wire  _EVAL_32;
  wire  _EVAL_217;
  wire  _EVAL_350;
  wire  _EVAL_176;
  wire  _EVAL_290;
  wire  _EVAL_108;
  wire  _EVAL_332;
  wire  _EVAL_110;
  wire  _EVAL_116;
  wire  _EVAL_38;
  wire  _EVAL_364;
  wire  _EVAL_120;
  wire  _EVAL_351;
  wire  _EVAL_370;
  wire  _EVAL_348;
  wire  _EVAL_237;
  wire  _EVAL_41;
  wire  _EVAL_131;
  wire  _EVAL_231;
  wire  _EVAL_42;
  wire [31:0] _EVAL_167;
  wire  _EVAL_210;
  wire  _EVAL_197;
  wire [127:0] _EVAL_89;
  wire [127:0] _EVAL_235;
  wire  _EVAL_129;
  wire  _EVAL_29;
  wire  _EVAL_95;
  wire  _EVAL_155;
  wire  _EVAL_79;
  wire  _EVAL_320;
  wire [72:0] _EVAL_308;
  wire  _EVAL_385;
  wire  _EVAL_336;
  wire  _EVAL_111;
  wire  _EVAL_168;
  wire  _EVAL_190;
  wire [127:0] _EVAL_345;
  wire [127:0] _EVAL_24;
  wire [72:0] _EVAL_230;
  wire  _EVAL_367;
  wire  _EVAL_102;
  wire  _EVAL_36;
  wire  _EVAL_55;
  wire  _EVAL_23;
  wire  _EVAL_122;
  wire  _EVAL_228;
  wire [29:0] _EVAL_376;
  wire [30:0] _EVAL_146;
  wire [30:0] _EVAL_356;
  wire [30:0] _EVAL_54;
  wire  _EVAL_334;
  wire  _EVAL_377;
  wire  _EVAL_149;
  wire  _EVAL_67;
  wire  _EVAL_47;
  wire  _EVAL_58;
  wire [29:0] _EVAL_212;
  wire [30:0] _EVAL_224;
  wire [30:0] _EVAL_53;
  wire [30:0] _EVAL_335;
  wire  _EVAL_148;
  wire  _EVAL_74;
  wire [30:0] _EVAL_92;
  wire [30:0] _EVAL_219;
  wire [30:0] _EVAL_277;
  wire  _EVAL_101;
  wire  _EVAL_145;
  wire [29:0] _EVAL_291;
  wire [30:0] _EVAL_208;
  wire [30:0] _EVAL_227;
  wire [30:0] _EVAL_310;
  wire  _EVAL_397;
  wire  _EVAL_26;
  wire  _EVAL_161;
  wire [29:0] _EVAL_144;
  wire [30:0] _EVAL_214;
  wire [30:0] _EVAL_163;
  wire [30:0] _EVAL_315;
  wire  _EVAL_52;
  wire  _EVAL_209;
  wire  _EVAL_359;
  wire  _EVAL_28;
  wire  _EVAL_361;
  wire  _EVAL_139;
  wire  _EVAL_289;
  wire  _EVAL_262;
  wire  _EVAL_257;
  wire  _EVAL_340;
  wire  _EVAL_360;
  wire  _EVAL_259;
  wire  _EVAL_372;
  wire  _EVAL_31;
  wire  _EVAL_363;
  wire  _EVAL_203;
  wire  _EVAL_382;
  wire  _EVAL_135;
  wire  _EVAL_267;
  wire  _EVAL_349;
  wire  _EVAL_178;
  wire  _EVAL_199;
  wire  _EVAL_341;
  wire  _EVAL_147;
  wire  _EVAL_319;
  wire  _EVAL_19;
  wire  _EVAL_25;
  wire  _EVAL_201;
  wire  _EVAL_221;
  wire  _EVAL_300;
  wire  _EVAL_240;
  wire  _EVAL_69;
  wire  _EVAL_27;
  wire  _EVAL_243;
  wire  _EVAL_362;
  wire  _EVAL_174;
  wire  _EVAL_77;
  wire  _EVAL_193;
  wire [7:0] _EVAL_138;
  wire [7:0] _EVAL_192;
  wire [7:0] _EVAL_157;
  wire  _EVAL_215;
  wire  _EVAL_133;
  wire  _EVAL_40;
  wire  _EVAL_78;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_70;
  wire [7:0] _EVAL_295;
  wire  _EVAL_303;
  wire  _EVAL_182;
  wire [72:0] _EVAL_322;
  wire  _EVAL_87;
  wire  _EVAL_247;
  wire  _EVAL_323;
  wire  _EVAL_72;
  wire [22:0] _EVAL_60;
  wire [7:0] _EVAL_253;
  wire [7:0] _EVAL_158;
  wire [4:0] _EVAL_166;
  wire [4:0] _EVAL_248;
  wire  _EVAL_125;
  wire  _EVAL_103;
  wire  _EVAL_43;
  wire  _EVAL_180;
  wire  _EVAL_226;
  wire  _EVAL_177;
  wire  _EVAL_218;
  wire  _EVAL_313;
  wire  _EVAL_234;
  wire  _EVAL_107;
  wire  _EVAL_251;
  wire  _EVAL_250;
  wire  _EVAL_165;
  wire  _EVAL_275;
  wire  _EVAL_269;
  wire  _EVAL_241;
  wire  _EVAL_284;
  wire  _EVAL_388;
  wire  _EVAL_281;
  wire  _EVAL_142;
  wire  _EVAL_151;
  wire  _EVAL_86;
  wire  _EVAL_112;
  wire  _EVAL_172;
  wire  _EVAL_270;
  wire  _EVAL_294;
  wire  _EVAL_46;
  wire [72:0] _EVAL_375;
  wire [72:0] _EVAL_64;
  wire  _EVAL_369;
  wire  _EVAL_395;
  wire  _EVAL_383;
  wire  _EVAL_97;
  wire  _EVAL_276;
  wire  _EVAL_265;
  wire  _EVAL_141;
  wire  _EVAL_37;
  wire  _EVAL_140;
  wire [22:0] _EVAL_169;
  wire [7:0] _EVAL_344;
  wire [7:0] _EVAL_327;
  wire [4:0] _EVAL_287;
  wire  _EVAL_324;
  wire  _EVAL_88;
  wire  _EVAL_333;
  wire  _EVAL_83;
  wire [4:0] _EVAL_119;
  wire  _EVAL_393;
  wire  _EVAL_274;
  wire  _EVAL_159;
  wire  _EVAL_191;
  wire  _EVAL_196;
  wire  _EVAL_337;
  wire  _EVAL_202;
  wire  _EVAL_391;
  wire  _EVAL_293;
  wire  _EVAL_207;
  wire [4:0] _EVAL_188;
  wire  _EVAL_381;
  wire  _EVAL_66;
  wire  _EVAL_63;
  wire  _EVAL_154;
  wire  _EVAL_195;
  wire  _EVAL_352;
  wire  _EVAL_94;
  wire  _EVAL_379;
  wire  _EVAL_56;
  wire  _EVAL_184;
  wire [4:0] _EVAL_239;
  wire  _EVAL_136;
  wire  _EVAL_160;
  wire  _EVAL_392;
  wire  _EVAL_48;
  wire  _EVAL_143;
  wire  _EVAL_238;
  wire  _EVAL_321;
  wire  _EVAL_91;
  wire  _EVAL_306;
  wire  _EVAL_249;
  wire  _EVAL_124;
  wire  _EVAL_368;
  wire  _EVAL_132;
  wire  _EVAL_330;
  wire  _EVAL_204;
  wire  _EVAL_292;
  wire [29:0] _EVAL_312;
  wire  _EVAL_232;
  wire  _EVAL_374;
  wire  _EVAL_398;
  wire  _EVAL_355;
  wire  _EVAL_114;
  wire  _EVAL_200;
  wire  _EVAL_198;
  wire  _EVAL_90;
  wire  _EVAL_126;
  wire [29:0] _EVAL_357;
  wire  _EVAL_304;
  wire  _EVAL_39;
  wire  _EVAL_298;
  wire  _EVAL_59;
  wire  _EVAL_65;
  wire  _EVAL_242;
  wire  _EVAL_394;
  wire  _EVAL_285;
  wire  _EVAL_305;
  wire  _EVAL_220;
  wire  _EVAL_331;
  wire  _EVAL_205;
  wire  _EVAL_57;
  wire  _EVAL_100;
  wire  _EVAL_233;
  wire  _EVAL_68;
  wire  _EVAL_386;
  wire  _EVAL_96;
  wire  _EVAL_264;
  wire  _EVAL_365;
  wire  _EVAL_380;
  wire [72:0] _EVAL_266;
  wire  _EVAL_134;
  wire  _EVAL_311;
  wire  _EVAL_389;
  wire  _EVAL_106;
  wire  _EVAL_211;
  wire  _EVAL_346;
  wire  _EVAL_297;
  wire  _EVAL_186;
  wire  _EVAL_181;
  wire  _EVAL_278;
  wire  _EVAL_130;
  wire  _EVAL_118;
  wire  _EVAL_173;
  wire  _EVAL_280;
  wire  _EVAL_30;
  wire  _EVAL_396;
  wire  _EVAL_44;
  wire [72:0] _EVAL_354;
  wire [72:0] _EVAL_371;
  wire  _EVAL_85;
  wire  _EVAL_105;
  wire  _EVAL_117;
  wire  _EVAL_317;
  wire  _EVAL_256;
  wire  _EVAL_366;
  wire  _EVAL_189;
  wire  _EVAL_71;
  wire  _EVAL_244;
  wire  _EVAL_20;
  wire  _EVAL_302;
  wire  _EVAL_229;
  wire  _EVAL_84;
  wire  _EVAL_115;
  wire  _EVAL_283;
  wire  _EVAL_187;
  wire  _EVAL_373;
  wire  _EVAL_263;
  wire  _EVAL_194;
  wire  _EVAL_61;
  wire  _EVAL_175;
  wire  _EVAL_339;
  wire  _EVAL_183;
  wire  _EVAL_213;
  wire  _EVAL_156;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_353 = _EVAL_6[1:0];
  assign _EVAL_399 = 4'h1 << _EVAL_353;
  assign _EVAL_222 = _EVAL_399[2:0];
  assign _EVAL_216 = _EVAL_222 | 3'h1;
  assign _EVAL_206 = _EVAL_216[2];
  assign _EVAL_123 = _EVAL_8[2];
  assign _EVAL_170 = _EVAL_206 & _EVAL_123;
  assign _EVAL_282 = _EVAL_1 == 7'h48;
  assign _EVAL_164 = _EVAL_1 == 7'h40;
  assign _EVAL_152 = _EVAL_282 | _EVAL_164;
  assign _EVAL_325 = _EVAL_1[6:3];
  assign _EVAL_109 = _EVAL_325 == 4'h8;
  assign _EVAL_390 = _EVAL_1[2:0];
  assign _EVAL_329 = 3'h1 <= _EVAL_390;
  assign _EVAL_260 = _EVAL_109 & _EVAL_329;
  assign _EVAL_81 = _EVAL_152 | _EVAL_260;
  assign _EVAL_307 = _EVAL_7 == 7'h48;
  assign _EVAL_246 = _EVAL_7 == 7'h40;
  assign _EVAL_113 = _EVAL_307 | _EVAL_246;
  assign _EVAL_73 = _EVAL_7[6:3];
  assign _EVAL_252 = _EVAL_73 == 4'h8;
  assign _EVAL_225 = _EVAL_7[2:0];
  assign _EVAL_314 = 3'h1 <= _EVAL_225;
  assign _EVAL_76 = _EVAL_252 & _EVAL_314;
  assign _EVAL_309 = _EVAL_113 | _EVAL_76;
  assign _EVAL_150 = _EVAL_7 == 7'h20;
  assign _EVAL_50 = _EVAL_309 | _EVAL_150;
  assign _EVAL_328 = _EVAL_73 == 4'h0;
  assign _EVAL_358 = _EVAL_50 | _EVAL_328;
  assign _EVAL_343 = _EVAL_73 == 4'h1;
  assign _EVAL_98 = _EVAL_358 | _EVAL_343;
  assign _EVAL_258 = _EVAL_8 ^ 30'h3000;
  assign _EVAL_338 = {1'b0,$signed(_EVAL_258)};
  assign _EVAL_223 = $signed(_EVAL_338) & $signed(-31'sh1000);
  assign _EVAL_121 = $signed(_EVAL_223);
  assign _EVAL_384 = $signed(_EVAL_121) == $signed(31'sh0);
  assign _EVAL_80 = _EVAL_8 ^ 30'h1900000;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_80)};
  assign _EVAL_21 = $signed(_EVAL_288) & $signed(-31'sh2000);
  assign _EVAL_286 = $signed(_EVAL_21);
  assign _EVAL_162 = $signed(_EVAL_286) == $signed(31'sh0);
  assign _EVAL_93 = _EVAL_73 == 4'h2;
  assign _EVAL_171 = _EVAL_98 | _EVAL_93;
  assign _EVAL_268 = _EVAL_216[0];
  assign _EVAL_62 = _EVAL_123 == 1'h0;
  assign _EVAL_32 = _EVAL_8[1];
  assign _EVAL_217 = _EVAL_32 == 1'h0;
  assign _EVAL_350 = _EVAL_62 & _EVAL_217;
  assign _EVAL_176 = _EVAL_8[0];
  assign _EVAL_290 = _EVAL_350 & _EVAL_176;
  assign _EVAL_108 = _EVAL_268 & _EVAL_290;
  assign _EVAL_332 = _EVAL_123 & _EVAL_32;
  assign _EVAL_110 = _EVAL_332 & _EVAL_176;
  assign _EVAL_116 = _EVAL_6 >= 4'h3;
  assign _EVAL_38 = _EVAL_206 & _EVAL_62;
  assign _EVAL_364 = _EVAL_116 | _EVAL_38;
  assign _EVAL_120 = _EVAL_216[1];
  assign _EVAL_351 = _EVAL_120 & _EVAL_350;
  assign _EVAL_370 = _EVAL_364 | _EVAL_351;
  assign _EVAL_348 = _EVAL_4 == _EVAL_185;
  assign _EVAL_237 = _EVAL_348 | _EVAL_2;
  assign _EVAL_41 = _EVAL_237 == 1'h0;
  assign _EVAL_131 = _EVAL_18 & _EVAL_13;
  assign _EVAL_231 = _EVAL_5 & _EVAL;
  assign _EVAL_42 = _EVAL_131 | _EVAL_231;
  assign _EVAL_167 = _EVAL_34 + 32'h1;
  assign _EVAL_210 = _EVAL_254 == 5'h0;
  assign _EVAL_197 = _EVAL_131 & _EVAL_210;
  assign _EVAL_89 = 128'h1 << _EVAL_7;
  assign _EVAL_235 = _EVAL_197 ? _EVAL_89 : 128'h0;
  assign _EVAL_129 = _EVAL_62 & _EVAL_32;
  assign _EVAL_29 = _EVAL_129 & _EVAL_176;
  assign _EVAL_95 = _EVAL_268 & _EVAL_29;
  assign _EVAL_155 = _EVAL_10 != 3'h0;
  assign _EVAL_79 = _EVAL_12 == _EVAL_279;
  assign _EVAL_320 = _EVAL_79 | _EVAL_2;
  assign _EVAL_308 = _EVAL_235[72:0];
  assign _EVAL_385 = _EVAL_104 == 5'h0;
  assign _EVAL_336 = _EVAL_231 & _EVAL_385;
  assign _EVAL_111 = _EVAL_0 == 3'h6;
  assign _EVAL_168 = _EVAL_111 == 1'h0;
  assign _EVAL_190 = _EVAL_336 & _EVAL_168;
  assign _EVAL_345 = 128'h1 << _EVAL_1;
  assign _EVAL_24 = _EVAL_190 ? _EVAL_345 : 128'h0;
  assign _EVAL_230 = _EVAL_24[72:0];
  assign _EVAL_367 = _EVAL_308 != _EVAL_230;
  assign _EVAL_102 = _EVAL_308 != 73'h0;
  assign _EVAL_36 = _EVAL_102 == 1'h0;
  assign _EVAL_55 = _EVAL_367 | _EVAL_36;
  assign _EVAL_23 = _EVAL_12 == 2'h0;
  assign _EVAL_122 = _EVAL_23 | _EVAL_2;
  assign _EVAL_228 = _EVAL_122 == 1'h0;
  assign _EVAL_376 = _EVAL_8 ^ 30'hc000000;
  assign _EVAL_146 = {1'b0,$signed(_EVAL_376)};
  assign _EVAL_356 = $signed(_EVAL_146) & $signed(-31'sh4000000);
  assign _EVAL_54 = $signed(_EVAL_356);
  assign _EVAL_334 = $signed(_EVAL_54) == $signed(31'sh0);
  assign _EVAL_377 = _EVAL_384 | _EVAL_334;
  assign _EVAL_149 = _EVAL_45 == 5'h0;
  assign _EVAL_67 = _EVAL_149 == 1'h0;
  assign _EVAL_47 = _EVAL & _EVAL_67;
  assign _EVAL_58 = _EVAL_325 == 4'h0;
  assign _EVAL_212 = _EVAL_8 ^ 30'h2000000;
  assign _EVAL_224 = {1'b0,$signed(_EVAL_212)};
  assign _EVAL_53 = $signed(_EVAL_224) & $signed(-31'sh10000);
  assign _EVAL_335 = $signed(_EVAL_53);
  assign _EVAL_148 = $signed(_EVAL_335) == $signed(31'sh0);
  assign _EVAL_74 = _EVAL_334 | _EVAL_148;
  assign _EVAL_92 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_219 = $signed(_EVAL_92) & $signed(-31'sh5000);
  assign _EVAL_277 = $signed(_EVAL_219);
  assign _EVAL_101 = $signed(_EVAL_277) == $signed(31'sh0);
  assign _EVAL_145 = _EVAL_74 | _EVAL_101;
  assign _EVAL_291 = _EVAL_8 ^ 30'h1800000;
  assign _EVAL_208 = {1'b0,$signed(_EVAL_291)};
  assign _EVAL_227 = $signed(_EVAL_208) & $signed(-31'sh8000);
  assign _EVAL_310 = $signed(_EVAL_227);
  assign _EVAL_397 = $signed(_EVAL_310) == $signed(31'sh0);
  assign _EVAL_26 = _EVAL_145 | _EVAL_397;
  assign _EVAL_161 = _EVAL_26 | _EVAL_162;
  assign _EVAL_144 = _EVAL_8 ^ 30'h20000000;
  assign _EVAL_214 = {1'b0,$signed(_EVAL_144)};
  assign _EVAL_163 = $signed(_EVAL_214) & $signed(-31'sh2000);
  assign _EVAL_315 = $signed(_EVAL_163);
  assign _EVAL_52 = $signed(_EVAL_315) == $signed(31'sh0);
  assign _EVAL_209 = _EVAL_161 | _EVAL_52;
  assign _EVAL_359 = _EVAL_9 == 3'h3;
  assign _EVAL_28 = _EVAL_13 & _EVAL_359;
  assign _EVAL_361 = _EVAL_179 != 73'h0;
  assign _EVAL_139 = _EVAL_361 == 1'h0;
  assign _EVAL_289 = plusarg_reader_out == 32'h0;
  assign _EVAL_262 = _EVAL_139 | _EVAL_289;
  assign _EVAL_257 = _EVAL_34 < plusarg_reader_out;
  assign _EVAL_340 = _EVAL_262 | _EVAL_257;
  assign _EVAL_360 = _EVAL_116 | _EVAL_170;
  assign _EVAL_259 = _EVAL_120 & _EVAL_332;
  assign _EVAL_372 = _EVAL_360 | _EVAL_259;
  assign _EVAL_31 = _EVAL_268 & _EVAL_110;
  assign _EVAL_363 = _EVAL_372 | _EVAL_31;
  assign _EVAL_203 = _EVAL_176 == 1'h0;
  assign _EVAL_382 = _EVAL_332 & _EVAL_203;
  assign _EVAL_135 = _EVAL_268 & _EVAL_382;
  assign _EVAL_267 = _EVAL_372 | _EVAL_135;
  assign _EVAL_349 = _EVAL_123 & _EVAL_217;
  assign _EVAL_178 = _EVAL_120 & _EVAL_349;
  assign _EVAL_199 = _EVAL_360 | _EVAL_178;
  assign _EVAL_341 = _EVAL_349 & _EVAL_176;
  assign _EVAL_147 = _EVAL_268 & _EVAL_341;
  assign _EVAL_319 = _EVAL_199 | _EVAL_147;
  assign _EVAL_19 = _EVAL_349 & _EVAL_203;
  assign _EVAL_25 = _EVAL_268 & _EVAL_19;
  assign _EVAL_201 = _EVAL_199 | _EVAL_25;
  assign _EVAL_221 = _EVAL_120 & _EVAL_129;
  assign _EVAL_300 = _EVAL_364 | _EVAL_221;
  assign _EVAL_240 = _EVAL_300 | _EVAL_95;
  assign _EVAL_69 = _EVAL_129 & _EVAL_203;
  assign _EVAL_27 = _EVAL_268 & _EVAL_69;
  assign _EVAL_243 = _EVAL_300 | _EVAL_27;
  assign _EVAL_362 = _EVAL_370 | _EVAL_108;
  assign _EVAL_174 = _EVAL_350 & _EVAL_203;
  assign _EVAL_77 = _EVAL_268 & _EVAL_174;
  assign _EVAL_193 = _EVAL_370 | _EVAL_77;
  assign _EVAL_138 = {_EVAL_363,_EVAL_267,_EVAL_319,_EVAL_201,_EVAL_240,_EVAL_243,_EVAL_362,_EVAL_193};
  assign _EVAL_192 = ~ _EVAL_138;
  assign _EVAL_157 = _EVAL_14 & _EVAL_192;
  assign _EVAL_215 = _EVAL_157 == 8'h0;
  assign _EVAL_133 = _EVAL_215 | _EVAL_2;
  assign _EVAL_40 = _EVAL_133 == 1'h0;
  assign _EVAL_78 = _EVAL_6 <= 4'h6;
  assign _EVAL_271 = _EVAL_10 <= 3'h3;
  assign _EVAL_272 = _EVAL_6 == _EVAL_245;
  assign _EVAL_273 = _EVAL_272 | _EVAL_2;
  assign _EVAL_70 = _EVAL_273 == 1'h0;
  assign _EVAL_295 = ~ _EVAL_14;
  assign _EVAL_303 = _EVAL_295 == 8'h0;
  assign _EVAL_182 = _EVAL_9 == 3'h4;
  assign _EVAL_322 = _EVAL_179 >> _EVAL_7;
  assign _EVAL_87 = _EVAL_322[0];
  assign _EVAL_247 = _EVAL_301 == 5'h0;
  assign _EVAL_323 = _EVAL_9[2];
  assign _EVAL_72 = _EVAL_323 == 1'h0;
  assign _EVAL_60 = 23'hff << _EVAL_6;
  assign _EVAL_253 = _EVAL_60[7:0];
  assign _EVAL_158 = ~ _EVAL_253;
  assign _EVAL_166 = _EVAL_158[7:3];
  assign _EVAL_248 = _EVAL_301 - 5'h1;
  assign _EVAL_125 = _EVAL_9 == 3'h2;
  assign _EVAL_103 = _EVAL_10 == 3'h0;
  assign _EVAL_43 = _EVAL_103 | _EVAL_2;
  assign _EVAL_180 = _EVAL_9 == 3'h6;
  assign _EVAL_226 = _EVAL_13 & _EVAL_180;
  assign _EVAL_177 = _EVAL_9 == 3'h7;
  assign _EVAL_218 = _EVAL_6 <= 4'h8;
  assign _EVAL_313 = _EVAL_218 & _EVAL_384;
  assign _EVAL_234 = _EVAL_313 | _EVAL_2;
  assign _EVAL_107 = _EVAL_234 == 1'h0;
  assign _EVAL_251 = _EVAL_155 | _EVAL_2;
  assign _EVAL_250 = _EVAL_7 == _EVAL_35;
  assign _EVAL_165 = _EVAL_250 | _EVAL_2;
  assign _EVAL_275 = _EVAL_165 == 1'h0;
  assign _EVAL_269 = _EVAL_16 == 1'h0;
  assign _EVAL_241 = _EVAL_269 | _EVAL_11;
  assign _EVAL_284 = _EVAL_241 | _EVAL_2;
  assign _EVAL_388 = _EVAL_377 | _EVAL_148;
  assign _EVAL_281 = _EVAL_388 | _EVAL_101;
  assign _EVAL_142 = _EVAL_281 | _EVAL_397;
  assign _EVAL_151 = _EVAL_142 | _EVAL_162;
  assign _EVAL_86 = _EVAL_151 | _EVAL_52;
  assign _EVAL_112 = _EVAL_78 & _EVAL_209;
  assign _EVAL_172 = _EVAL_313 | _EVAL_112;
  assign _EVAL_270 = _EVAL_172 | _EVAL_2;
  assign _EVAL_294 = _EVAL_303 | _EVAL_2;
  assign _EVAL_46 = _EVAL_294 == 1'h0;
  assign _EVAL_375 = _EVAL_308 | _EVAL_179;
  assign _EVAL_64 = _EVAL_375 >> _EVAL_1;
  assign _EVAL_369 = _EVAL_64[0];
  assign _EVAL_395 = _EVAL_369 | _EVAL_2;
  assign _EVAL_383 = _EVAL_395 == 1'h0;
  assign _EVAL_97 = _EVAL_8 == _EVAL_255;
  assign _EVAL_276 = _EVAL_97 | _EVAL_2;
  assign _EVAL_265 = _EVAL_12 != 2'h2;
  assign _EVAL_141 = _EVAL_265 | _EVAL_2;
  assign _EVAL_37 = _EVAL_141 == 1'h0;
  assign _EVAL_140 = _EVAL_0[0];
  assign _EVAL_169 = 23'hff << _EVAL_17;
  assign _EVAL_344 = _EVAL_169[7:0];
  assign _EVAL_327 = ~ _EVAL_344;
  assign _EVAL_287 = _EVAL_327[7:3];
  assign _EVAL_324 = _EVAL_14 == _EVAL_138;
  assign _EVAL_88 = _EVAL_10 == _EVAL_387;
  assign _EVAL_333 = _EVAL_88 | _EVAL_2;
  assign _EVAL_83 = _EVAL_333 == 1'h0;
  assign _EVAL_119 = _EVAL_254 - 5'h1;
  assign _EVAL_393 = _EVAL_1 == 7'h20;
  assign _EVAL_274 = _EVAL_81 | _EVAL_393;
  assign _EVAL_159 = _EVAL_274 | _EVAL_58;
  assign _EVAL_191 = _EVAL_325 == 4'h1;
  assign _EVAL_196 = _EVAL_159 | _EVAL_191;
  assign _EVAL_337 = _EVAL_325 == 4'h2;
  assign _EVAL_202 = _EVAL_196 | _EVAL_337;
  assign _EVAL_391 = _EVAL_325 == 4'h3;
  assign _EVAL_293 = _EVAL_202 | _EVAL_391;
  assign _EVAL_207 = _EVAL_276 == 1'h0;
  assign _EVAL_188 = _EVAL_45 - 5'h1;
  assign _EVAL_381 = _EVAL_6 <= 4'h2;
  assign _EVAL_66 = _EVAL_381 & _EVAL_86;
  assign _EVAL_63 = _EVAL_66 | _EVAL_2;
  assign _EVAL_154 = _EVAL_9 == 3'h0;
  assign _EVAL_195 = _EVAL_13 & _EVAL_154;
  assign _EVAL_352 = _EVAL_1 == _EVAL_82;
  assign _EVAL_94 = _EVAL_352 | _EVAL_2;
  assign _EVAL_379 = _EVAL_17 >= 4'h3;
  assign _EVAL_56 = _EVAL_379 | _EVAL_2;
  assign _EVAL_184 = _EVAL_0 == _EVAL_99;
  assign _EVAL_239 = _EVAL_104 - 5'h1;
  assign _EVAL_136 = _EVAL_293 | _EVAL_2;
  assign _EVAL_160 = _EVAL_136 == 1'h0;
  assign _EVAL_392 = 4'h6 == _EVAL_6;
  assign _EVAL_48 = _EVAL_94 == 1'h0;
  assign _EVAL_143 = _EVAL_55 | _EVAL_2;
  assign _EVAL_238 = _EVAL_143 == 1'h0;
  assign _EVAL_321 = _EVAL_0 == 3'h2;
  assign _EVAL_91 = _EVAL & _EVAL_111;
  assign _EVAL_306 = _EVAL_324 | _EVAL_2;
  assign _EVAL_249 = _EVAL_306 == 1'h0;
  assign _EVAL_124 = _EVAL_10 <= 3'h4;
  assign _EVAL_368 = _EVAL_124 | _EVAL_2;
  assign _EVAL_132 = _EVAL_368 == 1'h0;
  assign _EVAL_330 = _EVAL_13 & _EVAL_125;
  assign _EVAL_204 = _EVAL_63 == 1'h0;
  assign _EVAL_292 = _EVAL_0 == 3'h0;
  assign _EVAL_312 = {{22'd0}, _EVAL_158};
  assign _EVAL_232 = _EVAL_340 | _EVAL_2;
  assign _EVAL_374 = _EVAL_10 <= 3'h2;
  assign _EVAL_398 = _EVAL_374 | _EVAL_2;
  assign _EVAL_355 = _EVAL_398 == 1'h0;
  assign _EVAL_114 = _EVAL_231 & _EVAL_149;
  assign _EVAL_200 = _EVAL_56 == 1'h0;
  assign _EVAL_198 = _EVAL_12 <= 2'h2;
  assign _EVAL_90 = _EVAL_198 | _EVAL_2;
  assign _EVAL_126 = _EVAL_90 == 1'h0;
  assign _EVAL_357 = _EVAL_8 & _EVAL_312;
  assign _EVAL_304 = _EVAL_357 == 30'h0;
  assign _EVAL_39 = _EVAL_304 | _EVAL_2;
  assign _EVAL_298 = _EVAL_184 | _EVAL_2;
  assign _EVAL_59 = _EVAL_298 == 1'h0;
  assign _EVAL_65 = _EVAL_0 == 3'h4;
  assign _EVAL_242 = _EVAL & _EVAL_65;
  assign _EVAL_394 = _EVAL_17 == _EVAL_299;
  assign _EVAL_285 = _EVAL_73 == 4'h3;
  assign _EVAL_305 = _EVAL_171 | _EVAL_285;
  assign _EVAL_220 = _EVAL_305 | _EVAL_2;
  assign _EVAL_331 = _EVAL_220 == 1'h0;
  assign _EVAL_205 = _EVAL & _EVAL_321;
  assign _EVAL_57 = _EVAL_320 == 1'h0;
  assign _EVAL_100 = _EVAL_9 == 3'h1;
  assign _EVAL_233 = _EVAL_13 & _EVAL_177;
  assign _EVAL_68 = _EVAL_284 == 1'h0;
  assign _EVAL_386 = _EVAL_246 ? _EVAL_392 : 1'h0;
  assign _EVAL_96 = _EVAL_386 | _EVAL_2;
  assign _EVAL_264 = _EVAL_96 == 1'h0;
  assign _EVAL_365 = _EVAL_15 == 1'h0;
  assign _EVAL_380 = _EVAL_87 == 1'h0;
  assign _EVAL_266 = ~ _EVAL_230;
  assign _EVAL_134 = _EVAL_11 == 1'h0;
  assign _EVAL_311 = _EVAL_9 == _EVAL_261;
  assign _EVAL_389 = _EVAL_311 | _EVAL_2;
  assign _EVAL_106 = _EVAL_251 == 1'h0;
  assign _EVAL_211 = _EVAL_0 == 3'h5;
  assign _EVAL_346 = _EVAL_380 | _EVAL_2;
  assign _EVAL_297 = _EVAL_346 == 1'h0;
  assign _EVAL_186 = _EVAL & _EVAL_292;
  assign _EVAL_181 = _EVAL_365 | _EVAL_2;
  assign _EVAL_278 = _EVAL_2 == 1'h0;
  assign _EVAL_130 = _EVAL_0 <= 3'h6;
  assign _EVAL_118 = _EVAL_130 | _EVAL_2;
  assign _EVAL_173 = _EVAL_389 == 1'h0;
  assign _EVAL_280 = _EVAL_270 == 1'h0;
  assign _EVAL_30 = _EVAL_269 | _EVAL_2;
  assign _EVAL_396 = _EVAL_30 == 1'h0;
  assign _EVAL_44 = _EVAL_271 | _EVAL_2;
  assign _EVAL_354 = _EVAL_179 | _EVAL_308;
  assign _EVAL_371 = _EVAL_354 & _EVAL_266;
  assign _EVAL_85 = _EVAL & _EVAL_211;
  assign _EVAL_105 = _EVAL_116 | _EVAL_2;
  assign _EVAL_117 = _EVAL_247 == 1'h0;
  assign _EVAL_317 = _EVAL_13 & _EVAL_117;
  assign _EVAL_256 = _EVAL_44 == 1'h0;
  assign _EVAL_366 = _EVAL_232 == 1'h0;
  assign _EVAL_189 = _EVAL_9 == 3'h5;
  assign _EVAL_71 = _EVAL_16 == _EVAL_127;
  assign _EVAL_244 = _EVAL_13 & _EVAL_182;
  assign _EVAL_20 = _EVAL_134 | _EVAL_2;
  assign _EVAL_302 = _EVAL_105 == 1'h0;
  assign _EVAL_229 = _EVAL_71 | _EVAL_2;
  assign _EVAL_84 = _EVAL_229 == 1'h0;
  assign _EVAL_115 = _EVAL_13 & _EVAL_100;
  assign _EVAL_283 = _EVAL_181 == 1'h0;
  assign _EVAL_187 = _EVAL_13 & _EVAL_189;
  assign _EVAL_373 = _EVAL_0 == 3'h1;
  assign _EVAL_263 = _EVAL & _EVAL_373;
  assign _EVAL_194 = _EVAL_394 | _EVAL_2;
  assign _EVAL_61 = _EVAL_194 == 1'h0;
  assign _EVAL_175 = _EVAL_43 == 1'h0;
  assign _EVAL_339 = _EVAL_118 == 1'h0;
  assign _EVAL_183 = _EVAL_131 & _EVAL_247;
  assign _EVAL_213 = _EVAL_20 == 1'h0;
  assign _EVAL_156 = _EVAL_39 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_34 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_45 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_82 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_99 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_104 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_127 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  _EVAL_179 = _RAND_7[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_185 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_245 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_254 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_255 = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_261 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_279 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_299 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_301 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_387 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_2) begin
      _EVAL_34 <= 32'h0;
    end else begin
      if (_EVAL_42) begin
        _EVAL_34 <= 32'h0;
      end else begin
        _EVAL_34 <= _EVAL_167;
      end
    end
    if (_EVAL_183) begin
      _EVAL_35 <= _EVAL_7;
    end
    if (_EVAL_2) begin
      _EVAL_45 <= 5'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_149) begin
          if (_EVAL_140) begin
            _EVAL_45 <= _EVAL_287;
          end else begin
            _EVAL_45 <= 5'h0;
          end
        end else begin
          _EVAL_45 <= _EVAL_188;
        end
      end
    end
    if (_EVAL_114) begin
      _EVAL_82 <= _EVAL_1;
    end
    if (_EVAL_114) begin
      _EVAL_99 <= _EVAL_0;
    end
    if (_EVAL_2) begin
      _EVAL_104 <= 5'h0;
    end else begin
      if (_EVAL_231) begin
        if (_EVAL_385) begin
          if (_EVAL_140) begin
            _EVAL_104 <= _EVAL_287;
          end else begin
            _EVAL_104 <= 5'h0;
          end
        end else begin
          _EVAL_104 <= _EVAL_239;
        end
      end
    end
    if (_EVAL_114) begin
      _EVAL_127 <= _EVAL_16;
    end
    if (_EVAL_2) begin
      _EVAL_179 <= 73'h0;
    end else begin
      _EVAL_179 <= _EVAL_371;
    end
    if (_EVAL_114) begin
      _EVAL_185 <= _EVAL_4;
    end
    if (_EVAL_183) begin
      _EVAL_245 <= _EVAL_6;
    end
    if (_EVAL_2) begin
      _EVAL_254 <= 5'h0;
    end else begin
      if (_EVAL_131) begin
        if (_EVAL_210) begin
          if (_EVAL_72) begin
            _EVAL_254 <= _EVAL_166;
          end else begin
            _EVAL_254 <= 5'h0;
          end
        end else begin
          _EVAL_254 <= _EVAL_119;
        end
      end
    end
    if (_EVAL_183) begin
      _EVAL_255 <= _EVAL_8;
    end
    if (_EVAL_183) begin
      _EVAL_261 <= _EVAL_9;
    end
    if (_EVAL_114) begin
      _EVAL_279 <= _EVAL_12;
    end
    if (_EVAL_114) begin
      _EVAL_299 <= _EVAL_17;
    end
    if (_EVAL_2) begin
      _EVAL_301 <= 5'h0;
    end else begin
      if (_EVAL_131) begin
        if (_EVAL_247) begin
          if (_EVAL_72) begin
            _EVAL_301 <= _EVAL_166;
          end else begin
            _EVAL_301 <= 5'h0;
          end
        end else begin
          _EVAL_301 <= _EVAL_248;
        end
      end
    end
    if (_EVAL_183) begin
      _EVAL_387 <= _EVAL_10;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17f3da19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d673b6b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b2f22aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6116b5c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d74706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdc4eb7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da48e53a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93411d67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4471e030)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8c3882c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59f72d92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c1d6de6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f6d8c19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5341c13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9187a35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e019781)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_339) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26b56dcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efe9c350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df9dd6b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41f1c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a73850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a753262)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(675d10b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1a76e7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_339) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(399a3d89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(244b0db7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27a77bb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7435d774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d1ad0d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_396) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fd9fa08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3316527)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bda0bf8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(995c9503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a87044f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1934dc57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14f46b05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e207368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a7c93c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(723680fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6cefb6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d94d4c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db4c8b89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1f526b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffe0a457)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e64073ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bed14de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89f89999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea3175f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_396) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9803612a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35bcf518)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a66f9ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3479da0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59be64af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a24c046)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e92dcc07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c378380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e123aac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_383) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c04a8f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78a0ad58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(459ad225)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b46b95c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66d05123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e479c9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(121fc043)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c316e4da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b642b530)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a54462f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7056dcd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af4ae2b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cd01c5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffc9f94c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bebebf6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fbeae33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4e09378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35791d46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca002ad5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4f8f7aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f14b347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7477cee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f5a4b1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44b836e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1ce142c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e533b999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c8ed7e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32974b58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4b2b337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35fe6db9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_383) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(944a946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90a69ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d8750bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
