//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_267_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [31:0] _EVAL_6,
  input  [7:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [31:0] _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input  [3:0]  _EVAL_19,
  input         _EVAL_20,
  input  [3:0]  _EVAL_21,
  input         _EVAL_22,
  input  [1:0]  _EVAL_23,
  input         _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  input  [3:0]  _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input  [3:0]  _EVAL_31,
  input  [3:0]  _EVAL_32,
  input         _EVAL_33
);
  wire [31:0] plusarg_reader_out;
  reg [4:0] _EVAL_148;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_162;
  reg [31:0] _RAND_1;
  reg [1:0] _EVAL_167;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_173;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_183;
  reg [31:0] _RAND_4;
  reg [8:0] _EVAL_197;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_232;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_245;
  reg [31:0] _RAND_7;
  reg  _EVAL_311;
  reg [31:0] _RAND_8;
  reg [31:0] _EVAL_316;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_369;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_370;
  reg [31:0] _RAND_11;
  reg [4:0] _EVAL_411;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_420;
  reg [31:0] _RAND_13;
  reg [31:0] _EVAL_439;
  reg [31:0] _RAND_14;
  reg  _EVAL_471;
  reg [31:0] _RAND_15;
  reg [31:0] _EVAL_488;
  reg [31:0] _RAND_16;
  reg [4:0] _EVAL_495;
  reg [31:0] _RAND_17;
  reg [4:0] _EVAL_503;
  reg [31:0] _RAND_18;
  reg [2:0] _EVAL_512;
  reg [31:0] _RAND_19;
  reg [1:0] _EVAL_530;
  reg [31:0] _RAND_20;
  reg [3:0] _EVAL_551;
  reg [31:0] _RAND_21;
  reg [4:0] _EVAL_567;
  reg [31:0] _RAND_22;
  reg [3:0] _EVAL_615;
  reg [31:0] _RAND_23;
  reg [2:0] _EVAL_631;
  reg [31:0] _RAND_24;
  reg [3:0] _EVAL_641;
  reg [31:0] _RAND_25;
  reg [4:0] _EVAL_651;
  reg [31:0] _RAND_26;
  reg [1:0] _EVAL_667;
  reg [31:0] _RAND_27;
  wire [31:0] _EVAL_85;
  wire  _EVAL_84;
  wire  _EVAL_359;
  wire [32:0] _EVAL_367;
  wire  _EVAL_485;
  wire  _EVAL_123;
  wire  _EVAL_540;
  wire  _EVAL_494;
  wire  _EVAL_110;
  wire  _EVAL_440;
  wire  _EVAL_48;
  wire  _EVAL_621;
  wire  _EVAL_630;
  wire [22:0] _EVAL_671;
  wire [7:0] _EVAL_206;
  wire [7:0] _EVAL_347;
  wire [4:0] _EVAL_544;
  wire  _EVAL_138;
  wire  _EVAL_653;
  wire [1:0] _EVAL_386;
  wire [3:0] _EVAL_135;
  wire [2:0] _EVAL_204;
  wire [2:0] _EVAL_83;
  wire  _EVAL_254;
  wire  _EVAL_617;
  wire  _EVAL_288;
  wire  _EVAL_287;
  wire  _EVAL_121;
  wire  _EVAL_153;
  wire  _EVAL_672;
  wire  _EVAL_76;
  wire  _EVAL_293;
  wire  _EVAL_374;
  wire  _EVAL_114;
  wire [32:0] _EVAL_100;
  wire [32:0] _EVAL_161;
  wire  _EVAL_209;
  wire [31:0] _EVAL_483;
  wire [32:0] _EVAL_230;
  wire [32:0] _EVAL_225;
  wire [32:0] _EVAL_189;
  wire  _EVAL_213;
  wire  _EVAL_658;
  wire [2:0] _EVAL_180;
  wire  _EVAL_125;
  wire  _EVAL_41;
  wire  _EVAL_97;
  wire  _EVAL_36;
  wire [31:0] _EVAL_136;
  wire [32:0] _EVAL_429;
  wire  _EVAL_649;
  wire  _EVAL_270;
  wire  _EVAL_305;
  wire  _EVAL_575;
  wire  _EVAL_317;
  wire  _EVAL_492;
  wire  _EVAL_645;
  wire  _EVAL_201;
  wire  _EVAL_496;
  wire  _EVAL_406;
  wire  _EVAL_486;
  wire  _EVAL_82;
  wire  _EVAL_389;
  wire  _EVAL_468;
  wire  _EVAL_396;
  wire  _EVAL_461;
  wire  _EVAL_354;
  wire  _EVAL_43;
  wire  _EVAL_555;
  wire  _EVAL_79;
  wire  _EVAL_68;
  wire  _EVAL_527;
  wire  _EVAL_554;
  wire  _EVAL_453;
  wire  _EVAL_480;
  wire  _EVAL_533;
  wire  _EVAL_647;
  wire  _EVAL_301;
  wire  _EVAL_561;
  wire  _EVAL_280;
  wire  _EVAL_164;
  wire  _EVAL_509;
  wire  _EVAL_50;
  wire  _EVAL_81;
  wire  _EVAL_170;
  wire  _EVAL_178;
  wire  _EVAL_580;
  wire  _EVAL_390;
  wire  _EVAL_579;
  wire [7:0] _EVAL_410;
  wire [7:0] _EVAL_636;
  wire [7:0] _EVAL_310;
  wire [4:0] _EVAL_140;
  wire  _EVAL_147;
  wire  _EVAL_477;
  wire  _EVAL_395;
  wire [22:0] _EVAL_376;
  wire [7:0] _EVAL_332;
  wire [7:0] _EVAL_200;
  wire [31:0] _EVAL_150;
  wire [31:0] _EVAL_434;
  wire [8:0] _EVAL_40;
  wire [31:0] _EVAL_257;
  wire [32:0] _EVAL_426;
  wire [32:0] _EVAL_600;
  wire [32:0] _EVAL_212;
  wire  _EVAL_432;
  wire [32:0] _EVAL_571;
  wire [32:0] _EVAL_193;
  wire  _EVAL_93;
  wire  _EVAL_563;
  wire [31:0] _EVAL_656;
  wire [32:0] _EVAL_442;
  wire [32:0] _EVAL_60;
  wire [32:0] _EVAL_623;
  wire  _EVAL_325;
  wire  _EVAL_65;
  wire  _EVAL_654;
  wire  _EVAL_111;
  wire  _EVAL_522;
  wire [15:0] _EVAL_472;
  wire [15:0] _EVAL_402;
  wire [8:0] _EVAL_628;
  wire [8:0] _EVAL_543;
  wire [8:0] _EVAL_497;
  wire  _EVAL_393;
  wire  _EVAL_505;
  wire [4:0] _EVAL_523;
  wire [31:0] _EVAL_326;
  wire [32:0] _EVAL_286;
  wire [32:0] _EVAL_602;
  wire  _EVAL_604;
  wire  _EVAL_279;
  wire  _EVAL_158;
  wire  _EVAL_514;
  wire [22:0] _EVAL_487;
  wire [7:0] _EVAL_320;
  wire [7:0] _EVAL_86;
  wire [31:0] _EVAL_626;
  wire  _EVAL_236;
  wire [31:0] _EVAL_360;
  wire [32:0] _EVAL_582;
  wire [32:0] _EVAL_205;
  wire [32:0] _EVAL_223;
  wire  _EVAL_217;
  wire  _EVAL_581;
  wire [31:0] _EVAL_648;
  wire [32:0] _EVAL_156;
  wire [32:0] _EVAL_45;
  wire [32:0] _EVAL_122;
  wire  _EVAL_560;
  wire  _EVAL_511;
  wire [31:0] _EVAL_260;
  wire [32:0] _EVAL_235;
  wire [32:0] _EVAL_454;
  wire [32:0] _EVAL_104;
  wire  _EVAL_566;
  wire  _EVAL_504;
  wire [31:0] _EVAL_233;
  wire [32:0] _EVAL_365;
  wire [32:0] _EVAL_620;
  wire [32:0] _EVAL_226;
  wire  _EVAL_549;
  wire  _EVAL_242;
  wire [32:0] _EVAL_625;
  wire [32:0] _EVAL_271;
  wire [32:0] _EVAL_329;
  wire  _EVAL_663;
  wire  _EVAL_253;
  wire [32:0] _EVAL_427;
  wire  _EVAL_349;
  wire  _EVAL_565;
  wire  _EVAL_457;
  wire  _EVAL_146;
  wire  _EVAL_474;
  wire [2:0] _EVAL_534;
  wire  _EVAL_95;
  wire  _EVAL_52;
  wire  _EVAL_394;
  wire  _EVAL_669;
  wire  _EVAL_264;
  wire [31:0] _EVAL_650;
  wire [32:0] _EVAL_587;
  wire [32:0] _EVAL_598;
  wire [32:0] _EVAL_415;
  wire  _EVAL_456;
  wire  _EVAL_53;
  wire [31:0] _EVAL_606;
  wire [32:0] _EVAL_56;
  wire  _EVAL_520;
  wire  _EVAL_149;
  wire  _EVAL_218;
  wire  _EVAL_577;
  wire  _EVAL_315;
  wire [2:0] _EVAL_609;
  wire  _EVAL_282;
  wire  _EVAL_256;
  wire  _EVAL_416;
  wire  _EVAL_518;
  wire [32:0] _EVAL_339;
  wire [32:0] _EVAL_412;
  wire  _EVAL_69;
  wire  _EVAL_601;
  wire [31:0] _EVAL_614;
  wire [32:0] _EVAL_240;
  wire [32:0] _EVAL_421;
  wire  _EVAL_510;
  wire  _EVAL_352;
  wire  _EVAL_448;
  wire  _EVAL_436;
  wire  _EVAL_186;
  wire  _EVAL_576;
  wire [31:0] _EVAL_476;
  wire [32:0] _EVAL_344;
  wire [32:0] _EVAL_313;
  wire  _EVAL_531;
  wire  _EVAL_536;
  wire  _EVAL_552;
  wire  _EVAL_489;
  wire  _EVAL_371;
  wire  _EVAL_589;
  wire [31:0] _EVAL_398;
  wire [32:0] _EVAL_72;
  wire [32:0] _EVAL_277;
  wire  _EVAL_478;
  wire  _EVAL_333;
  wire  _EVAL_224;
  wire [31:0] _EVAL_662;
  wire [32:0] _EVAL_661;
  wire [32:0] _EVAL_238;
  wire [31:0] _EVAL_348;
  wire  _EVAL_392;
  wire  _EVAL_583;
  wire [31:0] _EVAL_263;
  wire [32:0] _EVAL_283;
  wire [32:0] _EVAL_55;
  wire [32:0] _EVAL_537;
  wire  _EVAL_608;
  wire  _EVAL_517;
  wire  _EVAL_265;
  wire  _EVAL_475;
  wire  _EVAL_408;
  wire  _EVAL_187;
  wire [31:0] _EVAL_239;
  wire [32:0] _EVAL_116;
  wire [32:0] _EVAL_603;
  wire [32:0] _EVAL_78;
  wire  _EVAL_372;
  wire  _EVAL_249;
  wire [32:0] _EVAL_447;
  wire  _EVAL_450;
  wire  _EVAL_105;
  wire [32:0] _EVAL_124;
  wire  _EVAL_585;
  wire  _EVAL_595;
  wire  _EVAL_159;
  wire [31:0] _EVAL_479;
  wire [32:0] _EVAL_203;
  wire [32:0] _EVAL_573;
  wire [32:0] _EVAL_227;
  wire  _EVAL_296;
  wire [32:0] _EVAL_462;
  wire  _EVAL_613;
  wire  _EVAL_521;
  wire  _EVAL_89;
  wire  _EVAL_548;
  wire  _EVAL_538;
  wire [31:0] _EVAL_592;
  wire [32:0] _EVAL_80;
  wire [32:0] _EVAL_557;
  wire [32:0] _EVAL_190;
  wire  _EVAL_130;
  wire  _EVAL_291;
  wire  _EVAL_665;
  wire [32:0] _EVAL_337;
  wire  _EVAL_199;
  wire  _EVAL_119;
  wire [31:0] _EVAL_166;
  wire [32:0] _EVAL_659;
  wire [32:0] _EVAL_616;
  wire [32:0] _EVAL_126;
  wire  _EVAL_430;
  wire  _EVAL_145;
  wire [31:0] _EVAL_532;
  wire [32:0] _EVAL_361;
  wire [32:0] _EVAL_611;
  wire [32:0] _EVAL_545;
  wire  _EVAL_177;
  wire  _EVAL_290;
  wire  _EVAL_473;
  wire  _EVAL_118;
  wire [32:0] _EVAL_449;
  wire [32:0] _EVAL_252;
  wire  _EVAL_655;
  wire  _EVAL_168;
  wire  _EVAL_605;
  wire [1:0] _EVAL_493;
  wire  _EVAL_335;
  wire  _EVAL_446;
  wire  _EVAL_44;
  wire  _EVAL_258;
  wire  _EVAL_62;
  wire  _EVAL_171;
  wire  _EVAL_535;
  wire  _EVAL_364;
  wire  _EVAL_338;
  wire  _EVAL_38;
  wire  _EVAL_129;
  wire  _EVAL_507;
  wire  _EVAL_646;
  wire  _EVAL_163;
  wire  _EVAL_157;
  wire  _EVAL_334;
  wire  _EVAL_101;
  wire  _EVAL_237;
  wire  _EVAL_572;
  wire [15:0] _EVAL_466;
  wire [15:0] _EVAL_425;
  wire [8:0] _EVAL_463;
  wire  _EVAL_102;
  wire  _EVAL_342;
  wire  _EVAL_482;
  wire  _EVAL_377;
  wire  _EVAL_528;
  wire  _EVAL_35;
  wire  _EVAL_564;
  wire  _EVAL_500;
  wire  _EVAL_399;
  wire  _EVAL_165;
  wire [7:0] _EVAL_596;
  wire  _EVAL_350;
  wire  _EVAL_216;
  wire  _EVAL_635;
  wire [4:0] _EVAL_622;
  wire  _EVAL_590;
  wire  _EVAL_292;
  wire  _EVAL_137;
  wire  _EVAL_366;
  wire [4:0] _EVAL_49;
  wire  _EVAL_134;
  wire  _EVAL_599;
  wire [32:0] _EVAL_34;
  wire  _EVAL_381;
  wire  _EVAL_192;
  wire  _EVAL_214;
  wire  _EVAL_87;
  wire  _EVAL_324;
  wire [1:0] _EVAL_194;
  wire [1:0] _EVAL_433;
  wire [1:0] _EVAL_642;
  wire [31:0] _EVAL_99;
  wire [32:0] _EVAL_272;
  wire [31:0] _EVAL_175;
  wire  _EVAL_184;
  wire  _EVAL_417;
  wire  _EVAL_441;
  wire  _EVAL_139;
  wire  _EVAL_574;
  wire [32:0] _EVAL_98;
  wire  _EVAL_586;
  wire  _EVAL_559;
  wire  _EVAL_553;
  wire  _EVAL_524;
  wire [31:0] _EVAL_47;
  wire [32:0] _EVAL_46;
  wire [32:0] _EVAL_319;
  wire  _EVAL_231;
  wire  _EVAL_444;
  wire  _EVAL_490;
  wire  _EVAL_244;
  wire  _EVAL_673;
  wire  _EVAL_303;
  wire [31:0] _EVAL_73;
  wire [32:0] _EVAL_391;
  wire [32:0] _EVAL_368;
  wire [32:0] _EVAL_299;
  wire  _EVAL_529;
  wire  _EVAL_90;
  wire  _EVAL_413;
  wire  _EVAL_414;
  wire  _EVAL_593;
  wire [4:0] _EVAL_401;
  wire  _EVAL_211;
  wire  _EVAL_597;
  wire  _EVAL_397;
  wire  _EVAL_318;
  wire  _EVAL_51;
  wire  _EVAL_546;
  wire  _EVAL_103;
  wire [31:0] _EVAL_556;
  wire [32:0] _EVAL_269;
  wire [32:0] _EVAL_465;
  wire [32:0] _EVAL_37;
  wire  _EVAL_638;
  wire [1:0] _EVAL_558;
  wire [1:0] _EVAL_77;
  wire [4:0] _EVAL_141;
  wire [1:0] _EVAL_154;
  wire  _EVAL_424;
  wire  _EVAL_562;
  wire  _EVAL_351;
  wire  _EVAL_356;
  wire  _EVAL_67;
  wire [1:0] _EVAL_314;
  wire  _EVAL_70;
  wire  _EVAL_308;
  wire  _EVAL_255;
  wire  _EVAL_131;
  wire  _EVAL_327;
  wire  _EVAL_63;
  wire  _EVAL_619;
  wire  _EVAL_498;
  wire  _EVAL_208;
  wire  _EVAL_246;
  wire [32:0] _EVAL_343;
  wire  _EVAL_152;
  wire  _EVAL_578;
  wire [32:0] _EVAL_250;
  wire [32:0] _EVAL_169;
  wire  _EVAL_380;
  wire  _EVAL_215;
  wire [32:0] _EVAL_484;
  wire  _EVAL_353;
  wire  _EVAL_285;
  wire  _EVAL_451;
  wire  _EVAL_176;
  wire  _EVAL_261;
  wire  _EVAL_312;
  wire  _EVAL_407;
  wire  _EVAL_328;
  wire  _EVAL_428;
  wire  _EVAL_437;
  wire  _EVAL_435;
  wire  _EVAL_58;
  wire  _EVAL_248;
  wire  _EVAL_382;
  wire  _EVAL_357;
  wire  _EVAL_542;
  wire  _EVAL_634;
  wire [4:0] _EVAL_666;
  wire  _EVAL_132;
  wire  _EVAL_657;
  wire  _EVAL_422;
  wire  _EVAL_174;
  wire  _EVAL_142;
  wire  _EVAL_185;
  wire  _EVAL_610;
  wire  _EVAL_273;
  wire  _EVAL_516;
  wire [4:0] _EVAL_196;
  wire [32:0] _EVAL_275;
  wire  _EVAL_639;
  wire  _EVAL_222;
  wire  _EVAL_547;
  wire  _EVAL_207;
  wire  _EVAL_133;
  wire  _EVAL_243;
  wire  _EVAL_526;
  wire  _EVAL_550;
  wire  _EVAL_307;
  wire  _EVAL_336;
  wire  _EVAL_637;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_75;
  wire  _EVAL_191;
  wire  _EVAL_584;
  wire  _EVAL_61;
  wire  _EVAL_251;
  wire  _EVAL_458;
  wire  _EVAL_388;
  wire [1:0] _EVAL_71;
  wire  _EVAL_355;
  wire  _EVAL_670;
  wire  _EVAL_66;
  wire  _EVAL_375;
  wire  _EVAL_228;
  wire  _EVAL_607;
  wire  _EVAL_127;
  wire  _EVAL_385;
  wire  _EVAL_96;
  wire  _EVAL_321;
  wire  _EVAL_469;
  wire  _EVAL_373;
  wire  _EVAL_241;
  wire  _EVAL_74;
  wire  _EVAL_181;
  wire  _EVAL_627;
  wire  _EVAL_506;
  wire  _EVAL_117;
  wire  _EVAL_501;
  wire  _EVAL_229;
  wire  _EVAL_267;
  wire  _EVAL_91;
  wire  _EVAL_618;
  wire  _EVAL_297;
  wire  _EVAL_640;
  wire  _EVAL_455;
  wire  _EVAL_644;
  wire  _EVAL_107;
  wire  _EVAL_594;
  wire  _EVAL_160;
  wire [4:0] _EVAL_358;
  wire  _EVAL_128;
  wire  _EVAL_404;
  wire  _EVAL_220;
  wire  _EVAL_304;
  wire  _EVAL_400;
  wire  _EVAL_464;
  wire  _EVAL_262;
  wire  _EVAL_508;
  wire  _EVAL_569;
  wire  _EVAL_384;
  wire  _EVAL_541;
  wire  _EVAL_276;
  wire  _EVAL_491;
  wire  _EVAL_403;
  wire  _EVAL_668;
  wire  _EVAL_298;
  wire  _EVAL_179;
  wire  _EVAL_88;
  wire  _EVAL_284;
  wire [1:0] _EVAL_341;
  wire  _EVAL_443;
  wire  _EVAL_115;
  wire  _EVAL_247;
  wire  _EVAL_570;
  wire  _EVAL_302;
  wire  _EVAL_431;
  wire  _EVAL_664;
  wire  _EVAL_525;
  wire  _EVAL_59;
  wire  _EVAL_331;
  wire  _EVAL_64;
  wire  _EVAL_234;
  wire  _EVAL_445;
  wire  _EVAL_383;
  wire  _EVAL_345;
  wire  _EVAL_460;
  wire  _EVAL_652;
  wire  _EVAL_182;
  wire  _EVAL_281;
  wire  _EVAL_306;
  wire [8:0] _EVAL_588;
  wire  _EVAL_109;
  wire  _EVAL_362;
  wire  _EVAL_346;
  wire  _EVAL_502;
  wire  _EVAL_405;
  wire  _EVAL_452;
  wire  _EVAL_423;
  wire  _EVAL_195;
  wire  _EVAL_210;
  wire [31:0] _EVAL_155;
  wire  _EVAL_660;
  wire  _EVAL_378;
  wire  _EVAL_106;
  wire  _EVAL_268;
  wire  _EVAL_459;
  wire  _EVAL_151;
  wire  _EVAL_591;
  wire  _EVAL_143;
  wire  _EVAL_643;
  wire  _EVAL_54;
  wire  _EVAL_278;
  wire  _EVAL_120;
  wire  _EVAL_42;
  wire  _EVAL_632;
  wire  _EVAL_539;
  wire  _EVAL_266;
  wire  _EVAL_633;
  wire  _EVAL_419;
  wire  _EVAL_330;
  wire  _EVAL_309;
  wire [8:0] _EVAL_387;
  wire [8:0] _EVAL_295;
  wire  _EVAL_467;
  wire  _EVAL_202;
  wire  _EVAL_274;
  wire  _EVAL_363;
  wire  _EVAL_289;
  wire  _EVAL_219;
  wire  _EVAL_470;
  wire  _EVAL_221;
  wire  _EVAL_513;
  wire  _EVAL_94;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_85 = _EVAL_12 ^ 32'h40000000;
  assign _EVAL_84 = _EVAL_11 == 3'h4;
  assign _EVAL_359 = _EVAL_26 & _EVAL_84;
  assign _EVAL_367 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_485 = _EVAL_16 & _EVAL_33;
  assign _EVAL_123 = _EVAL_503 == 5'h0;
  assign _EVAL_540 = _EVAL_485 & _EVAL_123;
  assign _EVAL_494 = _EVAL_9 == 3'h4;
  assign _EVAL_110 = _EVAL_33 & _EVAL_494;
  assign _EVAL_440 = _EVAL_11 == _EVAL_512;
  assign _EVAL_48 = _EVAL_440 | _EVAL_28;
  assign _EVAL_621 = _EVAL_48 == 1'h0;
  assign _EVAL_630 = _EVAL_14[0];
  assign _EVAL_671 = 23'hff << _EVAL_32;
  assign _EVAL_206 = _EVAL_671[7:0];
  assign _EVAL_347 = ~ _EVAL_206;
  assign _EVAL_544 = _EVAL_347[7:3];
  assign _EVAL_138 = _EVAL_12[0];
  assign _EVAL_653 = _EVAL_138 == 1'h0;
  assign _EVAL_386 = _EVAL_21[1:0];
  assign _EVAL_135 = 4'h1 << _EVAL_386;
  assign _EVAL_204 = _EVAL_135[2:0];
  assign _EVAL_83 = _EVAL_204 | 3'h1;
  assign _EVAL_254 = _EVAL_83[0];
  assign _EVAL_617 = _EVAL_12[2];
  assign _EVAL_288 = _EVAL_617 == 1'h0;
  assign _EVAL_287 = _EVAL_12[1];
  assign _EVAL_121 = _EVAL_288 & _EVAL_287;
  assign _EVAL_153 = _EVAL_121 & _EVAL_653;
  assign _EVAL_672 = _EVAL_254 & _EVAL_153;
  assign _EVAL_76 = _EVAL_9[2];
  assign _EVAL_293 = _EVAL_19 == _EVAL_551;
  assign _EVAL_374 = _EVAL_293 | _EVAL_28;
  assign _EVAL_114 = _EVAL_374 == 1'h0;
  assign _EVAL_100 = $signed(_EVAL_367) & $signed(-33'sh5000);
  assign _EVAL_161 = $signed(_EVAL_100);
  assign _EVAL_209 = $signed(_EVAL_161) == $signed(33'sh0);
  assign _EVAL_483 = _EVAL_15 ^ 32'h40000000;
  assign _EVAL_230 = {1'b0,$signed(_EVAL_483)};
  assign _EVAL_225 = $signed(_EVAL_230) & $signed(-33'sh2000);
  assign _EVAL_189 = $signed(_EVAL_225);
  assign _EVAL_213 = _EVAL_31[3:3];
  assign _EVAL_658 = _EVAL_213 == 1'h0;
  assign _EVAL_180 = _EVAL_31[2:0];
  assign _EVAL_125 = 3'h1 <= _EVAL_180;
  assign _EVAL_41 = _EVAL_658 & _EVAL_125;
  assign _EVAL_97 = _EVAL_287 == 1'h0;
  assign _EVAL_36 = _EVAL_288 & _EVAL_97;
  assign _EVAL_136 = _EVAL_6 ^ 32'h80000000;
  assign _EVAL_429 = {1'b0,$signed(_EVAL_136)};
  assign _EVAL_649 = _EVAL_21 >= 4'h3;
  assign _EVAL_270 = _EVAL_83[2];
  assign _EVAL_305 = _EVAL_270 & _EVAL_617;
  assign _EVAL_575 = _EVAL_649 | _EVAL_305;
  assign _EVAL_317 = _EVAL_83[1];
  assign _EVAL_492 = _EVAL_617 & _EVAL_287;
  assign _EVAL_645 = _EVAL_317 & _EVAL_492;
  assign _EVAL_201 = _EVAL_575 | _EVAL_645;
  assign _EVAL_496 = _EVAL_492 & _EVAL_138;
  assign _EVAL_406 = _EVAL_254 & _EVAL_496;
  assign _EVAL_486 = _EVAL_201 | _EVAL_406;
  assign _EVAL_82 = _EVAL_492 & _EVAL_653;
  assign _EVAL_389 = _EVAL_254 & _EVAL_82;
  assign _EVAL_468 = _EVAL_201 | _EVAL_389;
  assign _EVAL_396 = _EVAL_617 & _EVAL_97;
  assign _EVAL_461 = _EVAL_317 & _EVAL_396;
  assign _EVAL_354 = _EVAL_575 | _EVAL_461;
  assign _EVAL_43 = _EVAL_396 & _EVAL_138;
  assign _EVAL_555 = _EVAL_254 & _EVAL_43;
  assign _EVAL_79 = _EVAL_354 | _EVAL_555;
  assign _EVAL_68 = _EVAL_396 & _EVAL_653;
  assign _EVAL_527 = _EVAL_254 & _EVAL_68;
  assign _EVAL_554 = _EVAL_354 | _EVAL_527;
  assign _EVAL_453 = _EVAL_270 & _EVAL_288;
  assign _EVAL_480 = _EVAL_649 | _EVAL_453;
  assign _EVAL_533 = _EVAL_317 & _EVAL_121;
  assign _EVAL_647 = _EVAL_480 | _EVAL_533;
  assign _EVAL_301 = _EVAL_121 & _EVAL_138;
  assign _EVAL_561 = _EVAL_254 & _EVAL_301;
  assign _EVAL_280 = _EVAL_647 | _EVAL_561;
  assign _EVAL_164 = _EVAL_647 | _EVAL_672;
  assign _EVAL_509 = _EVAL_317 & _EVAL_36;
  assign _EVAL_50 = _EVAL_480 | _EVAL_509;
  assign _EVAL_81 = _EVAL_36 & _EVAL_138;
  assign _EVAL_170 = _EVAL_254 & _EVAL_81;
  assign _EVAL_178 = _EVAL_50 | _EVAL_170;
  assign _EVAL_580 = _EVAL_36 & _EVAL_653;
  assign _EVAL_390 = _EVAL_254 & _EVAL_580;
  assign _EVAL_579 = _EVAL_50 | _EVAL_390;
  assign _EVAL_410 = {_EVAL_486,_EVAL_468,_EVAL_79,_EVAL_554,_EVAL_280,_EVAL_164,_EVAL_178,_EVAL_579};
  assign _EVAL_636 = ~ _EVAL_410;
  assign _EVAL_310 = _EVAL_7 & _EVAL_636;
  assign _EVAL_140 = _EVAL_503 - 5'h1;
  assign _EVAL_147 = _EVAL_15 == _EVAL_316;
  assign _EVAL_477 = _EVAL_7 == _EVAL_410;
  assign _EVAL_395 = _EVAL_477 | _EVAL_28;
  assign _EVAL_376 = 23'hff << _EVAL_21;
  assign _EVAL_332 = _EVAL_376[7:0];
  assign _EVAL_200 = ~ _EVAL_332;
  assign _EVAL_150 = {{24'd0}, _EVAL_200};
  assign _EVAL_434 = _EVAL_12 & _EVAL_150;
  assign _EVAL_40 = _EVAL_197 >> _EVAL_5;
  assign _EVAL_257 = _EVAL_6 ^ 32'h40000000;
  assign _EVAL_426 = {1'b0,$signed(_EVAL_257)};
  assign _EVAL_600 = $signed(_EVAL_426) & $signed(-33'sh2000);
  assign _EVAL_212 = $signed(_EVAL_600);
  assign _EVAL_432 = $signed(_EVAL_212) == $signed(33'sh0);
  assign _EVAL_571 = $signed(_EVAL_429) & $signed(-33'sh20000);
  assign _EVAL_193 = $signed(_EVAL_571);
  assign _EVAL_93 = $signed(_EVAL_193) == $signed(33'sh0);
  assign _EVAL_563 = _EVAL_432 | _EVAL_93;
  assign _EVAL_656 = _EVAL_6 ^ 32'h3000;
  assign _EVAL_442 = {1'b0,$signed(_EVAL_656)};
  assign _EVAL_60 = $signed(_EVAL_442) & $signed(-33'sh1000);
  assign _EVAL_623 = $signed(_EVAL_60);
  assign _EVAL_325 = $signed(_EVAL_623) == $signed(33'sh0);
  assign _EVAL_65 = _EVAL_563 | _EVAL_325;
  assign _EVAL_654 = _EVAL_11 == 3'h0;
  assign _EVAL_111 = _EVAL_651 == 5'h0;
  assign _EVAL_522 = _EVAL_485 & _EVAL_111;
  assign _EVAL_472 = 16'h1 << _EVAL_5;
  assign _EVAL_402 = _EVAL_522 ? _EVAL_472 : 16'h0;
  assign _EVAL_628 = _EVAL_402[8:0];
  assign _EVAL_543 = _EVAL_628 | _EVAL_197;
  assign _EVAL_497 = _EVAL_543 >> _EVAL_19;
  assign _EVAL_393 = _EVAL_497[0];
  assign _EVAL_505 = _EVAL_76 == 1'h0;
  assign _EVAL_523 = _EVAL_200[7:3];
  assign _EVAL_326 = _EVAL_6 ^ 32'h1900000;
  assign _EVAL_286 = {1'b0,$signed(_EVAL_326)};
  assign _EVAL_602 = $signed(_EVAL_286) & $signed(-33'sh2000);
  assign _EVAL_604 = _EVAL_395 == 1'h0;
  assign _EVAL_279 = _EVAL_8 == 2'h0;
  assign _EVAL_158 = _EVAL_279 | _EVAL_28;
  assign _EVAL_514 = _EVAL_158 == 1'h0;
  assign _EVAL_487 = 23'hff << _EVAL_27;
  assign _EVAL_320 = _EVAL_487[7:0];
  assign _EVAL_86 = ~ _EVAL_320;
  assign _EVAL_626 = {{24'd0}, _EVAL_86};
  assign _EVAL_236 = $signed(_EVAL_189) == $signed(33'sh0);
  assign _EVAL_360 = _EVAL_15 ^ 32'h80000000;
  assign _EVAL_582 = {1'b0,$signed(_EVAL_360)};
  assign _EVAL_205 = $signed(_EVAL_582) & $signed(-33'sh20000);
  assign _EVAL_223 = $signed(_EVAL_205);
  assign _EVAL_217 = $signed(_EVAL_223) == $signed(33'sh0);
  assign _EVAL_581 = _EVAL_236 | _EVAL_217;
  assign _EVAL_648 = _EVAL_15 ^ 32'h3000;
  assign _EVAL_156 = {1'b0,$signed(_EVAL_648)};
  assign _EVAL_45 = $signed(_EVAL_156) & $signed(-33'sh1000);
  assign _EVAL_122 = $signed(_EVAL_45);
  assign _EVAL_560 = $signed(_EVAL_122) == $signed(33'sh0);
  assign _EVAL_511 = _EVAL_581 | _EVAL_560;
  assign _EVAL_260 = _EVAL_15 ^ 32'hc000000;
  assign _EVAL_235 = {1'b0,$signed(_EVAL_260)};
  assign _EVAL_454 = $signed(_EVAL_235) & $signed(-33'sh4000000);
  assign _EVAL_104 = $signed(_EVAL_454);
  assign _EVAL_566 = $signed(_EVAL_104) == $signed(33'sh0);
  assign _EVAL_504 = _EVAL_511 | _EVAL_566;
  assign _EVAL_233 = _EVAL_15 ^ 32'h2000000;
  assign _EVAL_365 = {1'b0,$signed(_EVAL_233)};
  assign _EVAL_620 = $signed(_EVAL_365) & $signed(-33'sh10000);
  assign _EVAL_226 = $signed(_EVAL_620);
  assign _EVAL_549 = $signed(_EVAL_226) == $signed(33'sh0);
  assign _EVAL_242 = _EVAL_504 | _EVAL_549;
  assign _EVAL_625 = {1'b0,$signed(_EVAL_15)};
  assign _EVAL_271 = $signed(_EVAL_625) & $signed(-33'sh1000);
  assign _EVAL_329 = $signed(_EVAL_271);
  assign _EVAL_663 = $signed(_EVAL_329) == $signed(33'sh0);
  assign _EVAL_253 = _EVAL_242 | _EVAL_663;
  assign _EVAL_427 = {1'b0,$signed(_EVAL_6)};
  assign _EVAL_349 = _EVAL_5 == 4'h8;
  assign _EVAL_565 = _EVAL_5 == 4'h0;
  assign _EVAL_457 = _EVAL_349 | _EVAL_565;
  assign _EVAL_146 = _EVAL_5[3:3];
  assign _EVAL_474 = _EVAL_146 == 1'h0;
  assign _EVAL_534 = _EVAL_5[2:0];
  assign _EVAL_95 = 3'h1 <= _EVAL_534;
  assign _EVAL_52 = _EVAL_474 & _EVAL_95;
  assign _EVAL_394 = _EVAL_457 | _EVAL_52;
  assign _EVAL_669 = _EVAL_394 | _EVAL_28;
  assign _EVAL_264 = _EVAL_8 != 2'h2;
  assign _EVAL_650 = _EVAL_12 ^ 32'hc000000;
  assign _EVAL_587 = {1'b0,$signed(_EVAL_650)};
  assign _EVAL_598 = $signed(_EVAL_587) & $signed(-33'sh4000000);
  assign _EVAL_415 = $signed(_EVAL_598);
  assign _EVAL_456 = _EVAL_31 == _EVAL_370;
  assign _EVAL_53 = _EVAL_14 == 3'h2;
  assign _EVAL_606 = _EVAL_12 ^ 32'h3000;
  assign _EVAL_56 = {1'b0,$signed(_EVAL_606)};
  assign _EVAL_520 = _EVAL_25 != 3'h0;
  assign _EVAL_149 = _EVAL_520 | _EVAL_28;
  assign _EVAL_218 = _EVAL_149 == 1'h0;
  assign _EVAL_577 = _EVAL_19[3:3];
  assign _EVAL_315 = _EVAL_577 == 1'h0;
  assign _EVAL_609 = _EVAL_19[2:0];
  assign _EVAL_282 = 3'h1 <= _EVAL_609;
  assign _EVAL_256 = _EVAL_315 & _EVAL_282;
  assign _EVAL_416 = 4'h6 == _EVAL_27;
  assign _EVAL_518 = _EVAL_264 | _EVAL_28;
  assign _EVAL_339 = {1'b0,$signed(_EVAL_85)};
  assign _EVAL_412 = $signed(_EVAL_339) & $signed(-33'sh2000);
  assign _EVAL_69 = _EVAL_420 == 5'h0;
  assign _EVAL_601 = _EVAL_69 == 1'h0;
  assign _EVAL_614 = _EVAL_6 ^ 32'h1800000;
  assign _EVAL_240 = {1'b0,$signed(_EVAL_614)};
  assign _EVAL_421 = $signed(_EVAL_240) & $signed(-33'sh8000);
  assign _EVAL_510 = _EVAL_30 & _EVAL_22;
  assign _EVAL_352 = _EVAL_567 == 5'h0;
  assign _EVAL_448 = _EVAL_510 & _EVAL_352;
  assign _EVAL_436 = _EVAL_23 == _EVAL_167;
  assign _EVAL_186 = _EVAL_436 | _EVAL_28;
  assign _EVAL_576 = _EVAL_186 == 1'h0;
  assign _EVAL_476 = _EVAL_12 ^ 32'h1800000;
  assign _EVAL_344 = {1'b0,$signed(_EVAL_476)};
  assign _EVAL_313 = $signed(_EVAL_344) & $signed(-33'sh8000);
  assign _EVAL_531 = _EVAL_19 == 4'h8;
  assign _EVAL_536 = _EVAL_19 == 4'h0;
  assign _EVAL_552 = _EVAL_531 | _EVAL_536;
  assign _EVAL_489 = _EVAL_552 | _EVAL_256;
  assign _EVAL_371 = _EVAL_489 | _EVAL_28;
  assign _EVAL_589 = _EVAL_371 == 1'h0;
  assign _EVAL_398 = _EVAL_6 ^ 32'h2000000;
  assign _EVAL_72 = {1'b0,$signed(_EVAL_398)};
  assign _EVAL_277 = $signed(_EVAL_72) & $signed(-33'sh10000);
  assign _EVAL_478 = _EVAL_9 == _EVAL_369;
  assign _EVAL_333 = _EVAL_478 | _EVAL_28;
  assign _EVAL_224 = _EVAL_333 == 1'h0;
  assign _EVAL_662 = _EVAL_15 ^ 32'h1900000;
  assign _EVAL_661 = {1'b0,$signed(_EVAL_662)};
  assign _EVAL_238 = $signed(_EVAL_661) & $signed(-33'sh2000);
  assign _EVAL_348 = _EVAL_6 & _EVAL_626;
  assign _EVAL_392 = _EVAL_9 == 3'h2;
  assign _EVAL_583 = _EVAL_33 & _EVAL_392;
  assign _EVAL_263 = _EVAL_6 ^ 32'h4000;
  assign _EVAL_283 = {1'b0,$signed(_EVAL_263)};
  assign _EVAL_55 = $signed(_EVAL_283) & $signed(-33'sh1000);
  assign _EVAL_537 = $signed(_EVAL_55);
  assign _EVAL_608 = 4'h6 == _EVAL_21;
  assign _EVAL_517 = _EVAL_148 == 5'h0;
  assign _EVAL_265 = _EVAL_517 == 1'h0;
  assign _EVAL_475 = _EVAL_4 & _EVAL_265;
  assign _EVAL_408 = _EVAL_310 == 8'h0;
  assign _EVAL_187 = _EVAL_408 | _EVAL_28;
  assign _EVAL_239 = _EVAL_6 ^ 32'hc000000;
  assign _EVAL_116 = {1'b0,$signed(_EVAL_239)};
  assign _EVAL_603 = $signed(_EVAL_116) & $signed(-33'sh4000000);
  assign _EVAL_78 = $signed(_EVAL_603);
  assign _EVAL_372 = $signed(_EVAL_78) == $signed(33'sh0);
  assign _EVAL_249 = _EVAL_65 | _EVAL_372;
  assign _EVAL_447 = $signed(_EVAL_277);
  assign _EVAL_450 = $signed(_EVAL_447) == $signed(33'sh0);
  assign _EVAL_105 = _EVAL_249 | _EVAL_450;
  assign _EVAL_124 = $signed(_EVAL_421);
  assign _EVAL_585 = _EVAL_25 <= 3'h4;
  assign _EVAL_595 = _EVAL_585 | _EVAL_28;
  assign _EVAL_159 = _EVAL_595 == 1'h0;
  assign _EVAL_479 = _EVAL_12 ^ 32'h80000000;
  assign _EVAL_203 = {1'b0,$signed(_EVAL_479)};
  assign _EVAL_573 = $signed(_EVAL_203) & $signed(-33'sh20000);
  assign _EVAL_227 = $signed(_EVAL_573);
  assign _EVAL_296 = _EVAL_21 <= 4'h6;
  assign _EVAL_462 = $signed(_EVAL_412);
  assign _EVAL_613 = $signed(_EVAL_462) == $signed(33'sh0);
  assign _EVAL_521 = $signed(_EVAL_227) == $signed(33'sh0);
  assign _EVAL_89 = _EVAL_613 | _EVAL_521;
  assign _EVAL_548 = $signed(_EVAL_415) == $signed(33'sh0);
  assign _EVAL_538 = _EVAL_89 | _EVAL_548;
  assign _EVAL_592 = _EVAL_12 ^ 32'h2000000;
  assign _EVAL_80 = {1'b0,$signed(_EVAL_592)};
  assign _EVAL_557 = $signed(_EVAL_80) & $signed(-33'sh10000);
  assign _EVAL_190 = $signed(_EVAL_557);
  assign _EVAL_130 = $signed(_EVAL_190) == $signed(33'sh0);
  assign _EVAL_291 = _EVAL_538 | _EVAL_130;
  assign _EVAL_665 = _EVAL_291 | _EVAL_209;
  assign _EVAL_337 = $signed(_EVAL_313);
  assign _EVAL_199 = $signed(_EVAL_337) == $signed(33'sh0);
  assign _EVAL_119 = _EVAL_665 | _EVAL_199;
  assign _EVAL_166 = _EVAL_12 ^ 32'h1900000;
  assign _EVAL_659 = {1'b0,$signed(_EVAL_166)};
  assign _EVAL_616 = $signed(_EVAL_659) & $signed(-33'sh2000);
  assign _EVAL_126 = $signed(_EVAL_616);
  assign _EVAL_430 = $signed(_EVAL_126) == $signed(33'sh0);
  assign _EVAL_145 = _EVAL_119 | _EVAL_430;
  assign _EVAL_532 = _EVAL_12 ^ 32'h20000000;
  assign _EVAL_361 = {1'b0,$signed(_EVAL_532)};
  assign _EVAL_611 = $signed(_EVAL_361) & $signed(-33'sh2000);
  assign _EVAL_545 = $signed(_EVAL_611);
  assign _EVAL_177 = $signed(_EVAL_545) == $signed(33'sh0);
  assign _EVAL_290 = _EVAL_145 | _EVAL_177;
  assign _EVAL_473 = _EVAL_296 & _EVAL_290;
  assign _EVAL_118 = _EVAL_21 <= 4'h8;
  assign _EVAL_449 = $signed(_EVAL_56) & $signed(-33'sh1000);
  assign _EVAL_252 = $signed(_EVAL_449);
  assign _EVAL_655 = $signed(_EVAL_252) == $signed(33'sh0);
  assign _EVAL_168 = _EVAL_118 & _EVAL_655;
  assign _EVAL_605 = _EVAL_473 | _EVAL_168;
  assign _EVAL_493 = _EVAL_667 >> _EVAL_13;
  assign _EVAL_335 = _EVAL_493[0];
  assign _EVAL_446 = _EVAL_335 == 1'h0;
  assign _EVAL_44 = _EVAL_446 | _EVAL_28;
  assign _EVAL_258 = _EVAL_296 & _EVAL_521;
  assign _EVAL_62 = _EVAL_258 | _EVAL_28;
  assign _EVAL_171 = _EVAL_649 | _EVAL_28;
  assign _EVAL_535 = _EVAL_18 == 1'h0;
  assign _EVAL_364 = _EVAL_535 | _EVAL_28;
  assign _EVAL_338 = _EVAL_364 == 1'h0;
  assign _EVAL_38 = _EVAL_25 <= 3'h2;
  assign _EVAL_129 = _EVAL_38 | _EVAL_28;
  assign _EVAL_507 = _EVAL_129 == 1'h0;
  assign _EVAL_646 = _EVAL_393 | _EVAL_28;
  assign _EVAL_163 = _EVAL_646 == 1'h0;
  assign _EVAL_157 = _EVAL_411 == 5'h0;
  assign _EVAL_334 = _EVAL_510 & _EVAL_157;
  assign _EVAL_101 = _EVAL_14 == 3'h6;
  assign _EVAL_237 = _EVAL_101 == 1'h0;
  assign _EVAL_572 = _EVAL_334 & _EVAL_237;
  assign _EVAL_466 = 16'h1 << _EVAL_19;
  assign _EVAL_425 = _EVAL_572 ? _EVAL_466 : 16'h0;
  assign _EVAL_463 = _EVAL_425[8:0];
  assign _EVAL_102 = _EVAL_628 != _EVAL_463;
  assign _EVAL_342 = _EVAL_628 != 9'h0;
  assign _EVAL_482 = _EVAL_342 == 1'h0;
  assign _EVAL_377 = _EVAL_102 | _EVAL_482;
  assign _EVAL_528 = _EVAL_377 | _EVAL_28;
  assign _EVAL_35 = _EVAL_510 & _EVAL_69;
  assign _EVAL_564 = _EVAL_25 <= 3'h3;
  assign _EVAL_500 = _EVAL_564 | _EVAL_28;
  assign _EVAL_399 = _EVAL_14 == 3'h0;
  assign _EVAL_165 = _EVAL_22 & _EVAL_399;
  assign _EVAL_596 = ~ _EVAL_7;
  assign _EVAL_350 = _EVAL_27 <= 4'h6;
  assign _EVAL_216 = _EVAL_350 & _EVAL_93;
  assign _EVAL_635 = _EVAL_216 | _EVAL_28;
  assign _EVAL_622 = _EVAL_567 - 5'h1;
  assign _EVAL_590 = _EVAL_25 == 3'h0;
  assign _EVAL_292 = _EVAL_590 | _EVAL_28;
  assign _EVAL_137 = _EVAL_292 == 1'h0;
  assign _EVAL_366 = _EVAL_1 == 1'h0;
  assign _EVAL_49 = _EVAL_148 - 5'h1;
  assign _EVAL_134 = _EVAL_29 == 1'h0;
  assign _EVAL_599 = _EVAL_134 | _EVAL_28;
  assign _EVAL_34 = $signed(_EVAL_427) & $signed(-33'sh1000);
  assign _EVAL_381 = _EVAL_14[2];
  assign _EVAL_192 = _EVAL_14[1];
  assign _EVAL_214 = _EVAL_192 == 1'h0;
  assign _EVAL_87 = _EVAL_381 & _EVAL_214;
  assign _EVAL_324 = _EVAL_448 & _EVAL_87;
  assign _EVAL_194 = 2'h1 << _EVAL_13;
  assign _EVAL_433 = _EVAL_324 ? _EVAL_194 : 2'h0;
  assign _EVAL_642 = _EVAL_667 | _EVAL_433;
  assign _EVAL_99 = _EVAL_15 ^ 32'h4000;
  assign _EVAL_272 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_175 = _EVAL_15 & 32'h3f;
  assign _EVAL_184 = _EVAL_175 == 32'h0;
  assign _EVAL_417 = _EVAL_184 | _EVAL_28;
  assign _EVAL_441 = _EVAL_12 == _EVAL_439;
  assign _EVAL_139 = _EVAL_441 | _EVAL_28;
  assign _EVAL_574 = _EVAL_139 == 1'h0;
  assign _EVAL_98 = $signed(_EVAL_34);
  assign _EVAL_586 = $signed(_EVAL_98) == $signed(33'sh0);
  assign _EVAL_559 = _EVAL_31 == 4'h0;
  assign _EVAL_553 = _EVAL_1 == _EVAL_311;
  assign _EVAL_524 = _EVAL_553 | _EVAL_28;
  assign _EVAL_47 = _EVAL_15 ^ 32'h20000000;
  assign _EVAL_46 = {1'b0,$signed(_EVAL_47)};
  assign _EVAL_319 = $signed(_EVAL_46) & $signed(-33'sh2000);
  assign _EVAL_231 = _EVAL_171 == 1'h0;
  assign _EVAL_444 = _EVAL_14 <= 3'h6;
  assign _EVAL_490 = _EVAL_5 == _EVAL_641;
  assign _EVAL_244 = _EVAL_490 | _EVAL_28;
  assign _EVAL_673 = _EVAL_244 == 1'h0;
  assign _EVAL_303 = $signed(_EVAL_537) == $signed(33'sh0);
  assign _EVAL_73 = _EVAL_15 ^ 32'h1800000;
  assign _EVAL_391 = {1'b0,$signed(_EVAL_73)};
  assign _EVAL_368 = $signed(_EVAL_391) & $signed(-33'sh8000);
  assign _EVAL_299 = $signed(_EVAL_368);
  assign _EVAL_529 = _EVAL_25 == _EVAL_183;
  assign _EVAL_90 = $signed(_EVAL_124) == $signed(33'sh0);
  assign _EVAL_413 = _EVAL_14 == 3'h1;
  assign _EVAL_414 = _EVAL_444 | _EVAL_28;
  assign _EVAL_593 = _EVAL_414 == 1'h0;
  assign _EVAL_401 = _EVAL_411 - 5'h1;
  assign _EVAL_211 = _EVAL_565 ? _EVAL_608 : 1'h0;
  assign _EVAL_597 = _EVAL_211 | _EVAL_28;
  assign _EVAL_397 = _EVAL_597 == 1'h0;
  assign _EVAL_318 = _EVAL_31 == 4'h8;
  assign _EVAL_51 = _EVAL_318 | _EVAL_559;
  assign _EVAL_546 = _EVAL_51 | _EVAL_41;
  assign _EVAL_103 = _EVAL_546 | _EVAL_28;
  assign _EVAL_556 = _EVAL_6 ^ 32'h20000000;
  assign _EVAL_269 = {1'b0,$signed(_EVAL_556)};
  assign _EVAL_465 = $signed(_EVAL_269) & $signed(-33'sh2000);
  assign _EVAL_37 = $signed(_EVAL_465);
  assign _EVAL_638 = _EVAL_10 & _EVAL_2;
  assign _EVAL_558 = 2'h1 << _EVAL_17;
  assign _EVAL_77 = _EVAL_638 ? _EVAL_558 : 2'h0;
  assign _EVAL_141 = _EVAL_86[7:3];
  assign _EVAL_154 = ~ _EVAL_77;
  assign _EVAL_424 = _EVAL_13 == _EVAL_471;
  assign _EVAL_562 = _EVAL_424 | _EVAL_28;
  assign _EVAL_351 = _EVAL_147 | _EVAL_28;
  assign _EVAL_356 = _EVAL_351 == 1'h0;
  assign _EVAL_67 = _EVAL_21 <= 4'h2;
  assign _EVAL_314 = _EVAL_433 | _EVAL_667;
  assign _EVAL_70 = _EVAL_529 | _EVAL_28;
  assign _EVAL_308 = _EVAL_70 == 1'h0;
  assign _EVAL_255 = _EVAL_26 & _EVAL_654;
  assign _EVAL_131 = _EVAL_366 | _EVAL_28;
  assign _EVAL_327 = _EVAL_131 == 1'h0;
  assign _EVAL_63 = _EVAL_11[0];
  assign _EVAL_619 = _EVAL_23 <= 2'h2;
  assign _EVAL_498 = _EVAL_619 | _EVAL_28;
  assign _EVAL_208 = $signed(_EVAL_299) == $signed(33'sh0);
  assign _EVAL_246 = _EVAL_253 | _EVAL_208;
  assign _EVAL_343 = $signed(_EVAL_238);
  assign _EVAL_152 = $signed(_EVAL_343) == $signed(33'sh0);
  assign _EVAL_578 = _EVAL_246 | _EVAL_152;
  assign _EVAL_250 = $signed(_EVAL_272) & $signed(-33'sh1000);
  assign _EVAL_169 = $signed(_EVAL_250);
  assign _EVAL_380 = $signed(_EVAL_169) == $signed(33'sh0);
  assign _EVAL_215 = _EVAL_578 | _EVAL_380;
  assign _EVAL_484 = $signed(_EVAL_319);
  assign _EVAL_353 = $signed(_EVAL_484) == $signed(33'sh0);
  assign _EVAL_285 = _EVAL_215 | _EVAL_353;
  assign _EVAL_451 = _EVAL_197 != 9'h0;
  assign _EVAL_176 = _EVAL_451 == 1'h0;
  assign _EVAL_261 = plusarg_reader_out == 32'h0;
  assign _EVAL_312 = _EVAL_176 | _EVAL_261;
  assign _EVAL_407 = _EVAL_488 < plusarg_reader_out;
  assign _EVAL_328 = _EVAL_312 | _EVAL_407;
  assign _EVAL_428 = _EVAL_40[0];
  assign _EVAL_437 = _EVAL_428 == 1'h0;
  assign _EVAL_435 = _EVAL_32 == _EVAL_245;
  assign _EVAL_58 = _EVAL_3 & _EVAL_26;
  assign _EVAL_248 = _EVAL_123 == 1'h0;
  assign _EVAL_382 = _EVAL_33 & _EVAL_248;
  assign _EVAL_357 = _EVAL_105 | _EVAL_586;
  assign _EVAL_542 = _EVAL_357 | _EVAL_90;
  assign _EVAL_634 = _EVAL_495 == 5'h0;
  assign _EVAL_666 = _EVAL_495 - 5'h1;
  assign _EVAL_132 = _EVAL_328 | _EVAL_28;
  assign _EVAL_657 = _EVAL_132 == 1'h0;
  assign _EVAL_422 = _EVAL == _EVAL_631;
  assign _EVAL_174 = _EVAL_422 | _EVAL_28;
  assign _EVAL_142 = _EVAL_22 & _EVAL_601;
  assign _EVAL_185 = _EVAL_8 == _EVAL_530;
  assign _EVAL_610 = _EVAL_185 | _EVAL_28;
  assign _EVAL_273 = _EVAL_11 == 3'h6;
  assign _EVAL_516 = _EVAL_26 & _EVAL_273;
  assign _EVAL_196 = _EVAL_651 - 5'h1;
  assign _EVAL_275 = $signed(_EVAL_602);
  assign _EVAL_639 = $signed(_EVAL_275) == $signed(33'sh0);
  assign _EVAL_222 = _EVAL_542 | _EVAL_639;
  assign _EVAL_547 = _EVAL_222 | _EVAL_303;
  assign _EVAL_207 = $signed(_EVAL_37) == $signed(33'sh0);
  assign _EVAL_133 = _EVAL_547 | _EVAL_207;
  assign _EVAL_243 = _EVAL_133 | _EVAL_28;
  assign _EVAL_526 = _EVAL_243 == 1'h0;
  assign _EVAL_550 = _EVAL_456 | _EVAL_28;
  assign _EVAL_307 = _EVAL_550 == 1'h0;
  assign _EVAL_336 = _EVAL_348 == 32'h0;
  assign _EVAL_637 = _EVAL_336 | _EVAL_28;
  assign _EVAL_322 = _EVAL_655 | _EVAL_548;
  assign _EVAL_323 = _EVAL_8 <= 2'h2;
  assign _EVAL_75 = _EVAL_323 | _EVAL_28;
  assign _EVAL_191 = _EVAL_14 == 3'h5;
  assign _EVAL_584 = _EVAL_22 & _EVAL_191;
  assign _EVAL_61 = _EVAL <= 3'h5;
  assign _EVAL_251 = _EVAL_596 == 8'h0;
  assign _EVAL_458 = _EVAL_251 | _EVAL_28;
  assign _EVAL_388 = _EVAL_9 == 3'h5;
  assign _EVAL_71 = _EVAL_314 >> _EVAL_17;
  assign _EVAL_355 = _EVAL_71[0];
  assign _EVAL_670 = _EVAL_355 | _EVAL_28;
  assign _EVAL_66 = _EVAL_9 == 3'h6;
  assign _EVAL_375 = _EVAL_33 & _EVAL_66;
  assign _EVAL_228 = _EVAL_6 == _EVAL_173;
  assign _EVAL_607 = _EVAL_228 | _EVAL_28;
  assign _EVAL_127 = _EVAL_607 == 1'h0;
  assign _EVAL_385 = _EVAL_21 == _EVAL_615;
  assign _EVAL_96 = _EVAL_417 == 1'h0;
  assign _EVAL_321 = _EVAL_20 & _EVAL_4;
  assign _EVAL_469 = _EVAL_321 & _EVAL_517;
  assign _EVAL_373 = _EVAL_24 == 1'h0;
  assign _EVAL_241 = _EVAL_373 | _EVAL_28;
  assign _EVAL_74 = _EVAL_241 == 1'h0;
  assign _EVAL_181 = _EVAL_168 | _EVAL_28;
  assign _EVAL_627 = _EVAL_75 == 1'h0;
  assign _EVAL_506 = _EVAL_9 == 3'h1;
  assign _EVAL_117 = _EVAL_434 == 32'h0;
  assign _EVAL_501 = _EVAL_637 == 1'h0;
  assign _EVAL_229 = _EVAL_22 & _EVAL_101;
  assign _EVAL_267 = _EVAL_500 == 1'h0;
  assign _EVAL_91 = _EVAL <= 3'h2;
  assign _EVAL_618 = _EVAL_91 | _EVAL_28;
  assign _EVAL_297 = _EVAL_618 == 1'h0;
  assign _EVAL_640 = _EVAL_22 & _EVAL_53;
  assign _EVAL_455 = _EVAL_14 == _EVAL_232;
  assign _EVAL_644 = _EVAL_27 >= 4'h3;
  assign _EVAL_107 = _EVAL_644 | _EVAL_28;
  assign _EVAL_594 = _EVAL_11 == 3'h1;
  assign _EVAL_160 = _EVAL_435 | _EVAL_28;
  assign _EVAL_358 = _EVAL_420 - 5'h1;
  assign _EVAL_128 = _EVAL_524 == 1'h0;
  assign _EVAL_404 = _EVAL == 3'h0;
  assign _EVAL_220 = _EVAL_366 | _EVAL_29;
  assign _EVAL_304 = _EVAL_220 | _EVAL_28;
  assign _EVAL_400 = _EVAL_44 == 1'h0;
  assign _EVAL_464 = _EVAL_610 == 1'h0;
  assign _EVAL_262 = _EVAL_9 == 3'h0;
  assign _EVAL_508 = _EVAL_33 & _EVAL_262;
  assign _EVAL_569 = _EVAL_634 == 1'h0;
  assign _EVAL_384 = _EVAL_26 & _EVAL_569;
  assign _EVAL_541 = _EVAL_58 & _EVAL_634;
  assign _EVAL_276 = _EVAL_27 == _EVAL_162;
  assign _EVAL_491 = _EVAL_276 | _EVAL_28;
  assign _EVAL_403 = _EVAL_491 == 1'h0;
  assign _EVAL_668 = _EVAL_322 | _EVAL_130;
  assign _EVAL_298 = _EVAL_668 | _EVAL_209;
  assign _EVAL_179 = _EVAL_298 | _EVAL_199;
  assign _EVAL_88 = _EVAL_179 | _EVAL_430;
  assign _EVAL_284 = _EVAL_11 == 3'h7;
  assign _EVAL_341 = _EVAL_642 & _EVAL_154;
  assign _EVAL_443 = _EVAL_26 & _EVAL_594;
  assign _EVAL_115 = _EVAL_160 == 1'h0;
  assign _EVAL_247 = _EVAL_437 | _EVAL_28;
  assign _EVAL_570 = _EVAL_455 | _EVAL_28;
  assign _EVAL_302 = _EVAL_117 | _EVAL_28;
  assign _EVAL_431 = _EVAL_302 == 1'h0;
  assign _EVAL_664 = _EVAL_485 | _EVAL_510;
  assign _EVAL_525 = _EVAL_669 == 1'h0;
  assign _EVAL_59 = _EVAL_385 | _EVAL_28;
  assign _EVAL_331 = _EVAL_62 == 1'h0;
  assign _EVAL_64 = _EVAL_304 == 1'h0;
  assign _EVAL_234 = _EVAL_11 == 3'h5;
  assign _EVAL_445 = _EVAL_26 & _EVAL_234;
  assign _EVAL_383 = _EVAL_88 | _EVAL_177;
  assign _EVAL_345 = _EVAL_67 & _EVAL_383;
  assign _EVAL_460 = _EVAL_14 == 3'h4;
  assign _EVAL_652 = _EVAL_59 == 1'h0;
  assign _EVAL_182 = _EVAL_9 == 3'h7;
  assign _EVAL_281 = _EVAL_345 | _EVAL_28;
  assign _EVAL_306 = _EVAL_562 == 1'h0;
  assign _EVAL_588 = ~ _EVAL_463;
  assign _EVAL_109 = _EVAL_61 | _EVAL_28;
  assign _EVAL_362 = _EVAL_109 == 1'h0;
  assign _EVAL_346 = _EVAL_33 & _EVAL_506;
  assign _EVAL_502 = _EVAL_33 & _EVAL_182;
  assign _EVAL_405 = _EVAL_285 | _EVAL_28;
  assign _EVAL_452 = _EVAL_405 == 1'h0;
  assign _EVAL_423 = _EVAL_33 & _EVAL_388;
  assign _EVAL_195 = _EVAL_559 ? _EVAL_416 : 1'h0;
  assign _EVAL_210 = _EVAL_195 | _EVAL_28;
  assign _EVAL_155 = _EVAL_488 + 32'h1;
  assign _EVAL_660 = _EVAL_210 == 1'h0;
  assign _EVAL_378 = _EVAL_247 == 1'h0;
  assign _EVAL_106 = _EVAL_26 & _EVAL_284;
  assign _EVAL_268 = _EVAL_635 == 1'h0;
  assign _EVAL_459 = _EVAL_22 & _EVAL_413;
  assign _EVAL_151 = _EVAL_103 == 1'h0;
  assign _EVAL_591 = _EVAL_9 == 3'h3;
  assign _EVAL_143 = _EVAL_11 == 3'h2;
  assign _EVAL_643 = _EVAL_670 == 1'h0;
  assign _EVAL_54 = _EVAL_498 == 1'h0;
  assign _EVAL_278 = _EVAL_26 & _EVAL_143;
  assign _EVAL_120 = _EVAL_107 == 1'h0;
  assign _EVAL_42 = _EVAL_605 | _EVAL_28;
  assign _EVAL_632 = _EVAL_42 == 1'h0;
  assign _EVAL_539 = _EVAL_404 | _EVAL_28;
  assign _EVAL_266 = _EVAL_539 == 1'h0;
  assign _EVAL_633 = _EVAL_458 == 1'h0;
  assign _EVAL_419 = _EVAL_599 == 1'h0;
  assign _EVAL_330 = _EVAL_33 & _EVAL_591;
  assign _EVAL_309 = _EVAL_174 == 1'h0;
  assign _EVAL_387 = _EVAL_197 | _EVAL_628;
  assign _EVAL_295 = _EVAL_387 & _EVAL_588;
  assign _EVAL_467 = _EVAL_518 == 1'h0;
  assign _EVAL_202 = _EVAL_187 == 1'h0;
  assign _EVAL_274 = _EVAL_528 == 1'h0;
  assign _EVAL_363 = _EVAL_32 >= 4'h3;
  assign _EVAL_289 = _EVAL_363 | _EVAL_28;
  assign _EVAL_219 = _EVAL_289 == 1'h0;
  assign _EVAL_470 = _EVAL_281 == 1'h0;
  assign _EVAL_221 = _EVAL_22 & _EVAL_460;
  assign _EVAL_513 = _EVAL_181 == 1'h0;
  assign _EVAL_94 = _EVAL_570 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_148 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_162 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_167 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_173 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_183 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_197 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_232 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_245 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_311 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_316 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_369 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_370 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_411 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_420 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_439 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_471 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_488 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_495 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_503 = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_512 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_530 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_551 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_567 = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_615 = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_631 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_641 = _RAND_25[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_651 = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_667 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_28) begin
      _EVAL_148 <= 5'h0;
    end else begin
      if (_EVAL_321) begin
        if (_EVAL_517) begin
          _EVAL_148 <= 5'h0;
        end else begin
          _EVAL_148 <= _EVAL_49;
        end
      end
    end
    if (_EVAL_541) begin
      _EVAL_162 <= _EVAL_27;
    end
    if (_EVAL_469) begin
      _EVAL_167 <= _EVAL_23;
    end
    if (_EVAL_541) begin
      _EVAL_173 <= _EVAL_6;
    end
    if (_EVAL_540) begin
      _EVAL_183 <= _EVAL_25;
    end
    if (_EVAL_28) begin
      _EVAL_197 <= 9'h0;
    end else begin
      _EVAL_197 <= _EVAL_295;
    end
    if (_EVAL_35) begin
      _EVAL_232 <= _EVAL_14;
    end
    if (_EVAL_35) begin
      _EVAL_245 <= _EVAL_32;
    end
    if (_EVAL_35) begin
      _EVAL_311 <= _EVAL_1;
    end
    if (_EVAL_469) begin
      _EVAL_316 <= _EVAL_15;
    end
    if (_EVAL_540) begin
      _EVAL_369 <= _EVAL_9;
    end
    if (_EVAL_541) begin
      _EVAL_370 <= _EVAL_31;
    end
    if (_EVAL_28) begin
      _EVAL_411 <= 5'h0;
    end else begin
      if (_EVAL_510) begin
        if (_EVAL_157) begin
          if (_EVAL_630) begin
            _EVAL_411 <= _EVAL_544;
          end else begin
            _EVAL_411 <= 5'h0;
          end
        end else begin
          _EVAL_411 <= _EVAL_401;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_420 <= 5'h0;
    end else begin
      if (_EVAL_510) begin
        if (_EVAL_69) begin
          if (_EVAL_630) begin
            _EVAL_420 <= _EVAL_544;
          end else begin
            _EVAL_420 <= 5'h0;
          end
        end else begin
          _EVAL_420 <= _EVAL_358;
        end
      end
    end
    if (_EVAL_540) begin
      _EVAL_439 <= _EVAL_12;
    end
    if (_EVAL_35) begin
      _EVAL_471 <= _EVAL_13;
    end
    if (_EVAL_28) begin
      _EVAL_488 <= 32'h0;
    end else begin
      if (_EVAL_664) begin
        _EVAL_488 <= 32'h0;
      end else begin
        _EVAL_488 <= _EVAL_155;
      end
    end
    if (_EVAL_28) begin
      _EVAL_495 <= 5'h0;
    end else begin
      if (_EVAL_58) begin
        if (_EVAL_634) begin
          if (_EVAL_63) begin
            _EVAL_495 <= _EVAL_141;
          end else begin
            _EVAL_495 <= 5'h0;
          end
        end else begin
          _EVAL_495 <= _EVAL_666;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_503 <= 5'h0;
    end else begin
      if (_EVAL_485) begin
        if (_EVAL_123) begin
          if (_EVAL_505) begin
            _EVAL_503 <= _EVAL_523;
          end else begin
            _EVAL_503 <= 5'h0;
          end
        end else begin
          _EVAL_503 <= _EVAL_140;
        end
      end
    end
    if (_EVAL_541) begin
      _EVAL_512 <= _EVAL_11;
    end
    if (_EVAL_35) begin
      _EVAL_530 <= _EVAL_8;
    end
    if (_EVAL_35) begin
      _EVAL_551 <= _EVAL_19;
    end
    if (_EVAL_28) begin
      _EVAL_567 <= 5'h0;
    end else begin
      if (_EVAL_510) begin
        if (_EVAL_352) begin
          if (_EVAL_630) begin
            _EVAL_567 <= _EVAL_544;
          end else begin
            _EVAL_567 <= 5'h0;
          end
        end else begin
          _EVAL_567 <= _EVAL_622;
        end
      end
    end
    if (_EVAL_540) begin
      _EVAL_615 <= _EVAL_21;
    end
    if (_EVAL_541) begin
      _EVAL_631 <= _EVAL;
    end
    if (_EVAL_540) begin
      _EVAL_641 <= _EVAL_5;
    end
    if (_EVAL_28) begin
      _EVAL_651 <= 5'h0;
    end else begin
      if (_EVAL_485) begin
        if (_EVAL_111) begin
          if (_EVAL_505) begin
            _EVAL_651 <= _EVAL_523;
          end else begin
            _EVAL_651 <= 5'h0;
          end
        end else begin
          _EVAL_651 <= _EVAL_196;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_667 <= 2'h0;
    end else begin
      _EVAL_667 <= _EVAL_341;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_356) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44e915c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce929b95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_576) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a81ffd56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d0a23c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_514) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(722e5464)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41ba611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fa7a3ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_660) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(364219ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5f08e64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78cd3ba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee945b64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_362) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84fbc5b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_397) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(378f2b26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(247f822a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_419) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c47810)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81f2149c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a3709fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(872f79e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e32377b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_627) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7646043)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1850202c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98b3cfcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_403) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87943366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_643) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d73671a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c14f8f53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0e7e83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_522 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4b66f9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_356) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f1505ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_643) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_633) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f82c34e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4e5f947)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3794b660)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_419) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_507) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_403) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_621) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a546718)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb532850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_593) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71fd6dc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf03057f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc0ae1b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a7f91a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4652f71a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb5dda70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb0f91b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6d514fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1c98597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_633) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(577b5262)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_514) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d6b0770)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d544cc71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_627) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_397) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_621) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c299dbe1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_467) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_397) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(604c2046)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52c2956a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(379c3099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee65ef8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b03327f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63f7444f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_419) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_419) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d93a6235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90863b78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8010ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f895c69e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea938a39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_507) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89f7ea59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e777f17c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f111eb23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2aa7d02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_673) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb959071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_574) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1e88d10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82bb839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_657) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c16fb6d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_400) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(248eab7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_514) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_362) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9c2da0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69c7ff71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_627) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_362) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e774ced9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c9de0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbedeb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_419) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b3990e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_657) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e94fb26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ceef36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_419) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df6d00bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7215ac50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_467) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_400) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf4cab53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91271924)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_652) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90355e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7b2e9a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d0d146e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb2f8920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(babe3fd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(670732e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e888049)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_419) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb0326)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_576) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_514) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8409446f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ad184f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816c0c09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be206040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7f0dd3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_633) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_507) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c775b00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0ae3af4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e68535c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1311be9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_362) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_419) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(220419a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9caee567)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9db0ca3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_660) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(755e5c4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_514) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d267084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac288431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_673) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a05dab4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_397) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e369831e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc9f0b8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e264d31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_507) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1456870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_501) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf573a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_467) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54a11a7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b71a7cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caa34fd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18c5b941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_574) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eecb581b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_445 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_513) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b163484)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55095b15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4d5e85d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_633) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af0dc422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(905b53f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c47f15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_514) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c44e2667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_627) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b842d402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(296caa3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_513) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97b2e6ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39ae29b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9600976)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2948e21f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22960075)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_593) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2a7dc9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_514) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b653f757)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(422d7c22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_604) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(789d0501)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7d90e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_467) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a710bd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16c6fe94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_522 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(143d4ca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_514) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81cb4396)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_604) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(235f3bcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35aa0f95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_502 & _EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9f1de86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
