//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_84_assert(
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_7,
  input         _EVAL_9,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_22,
  input  [2:0]  _EVAL_25,
  input  [5:0]  _EVAL_34,
  input  [31:0] _EVAL_36,
  input  [3:0]  _EVAL_37,
  input  [2:0]  Queue_1__EVAL_14,
  input         Queue_1__EVAL_9,
  input         Queue_1__EVAL_5,
  input         Queue_1__EVAL_4,
  input         Queue_1__EVAL_3,
  input  [5:0]  Queue_1__EVAL_15,
  input  [3:0]  Queue_1__EVAL_11,
  input  [1:0]  Queue_1__EVAL_17,
  input         Queue__EVAL_4
);
  wire [5:0] TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire [3:0] TLMonitor__EVAL_1;
  wire [1:0] TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire [5:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [2:0] TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire [3:0] TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire [3:0] TLMonitor__EVAL_11;
  wire  TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [2:0] TLMonitor__EVAL_14;
  wire  TLMonitor__EVAL_15;
  wire [31:0] TLMonitor__EVAL_16;
  wire [2:0] TLMonitor__EVAL_17;
  wire  TLMonitor__EVAL_18;
  SiFive__EVAL_81_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18)
  );
  assign TLMonitor__EVAL_7 = Queue_1__EVAL_14;
  assign TLMonitor__EVAL = _EVAL_34;
  assign TLMonitor__EVAL_17 = _EVAL_25;
  assign TLMonitor__EVAL_12 = Queue_1__EVAL_9;
  assign TLMonitor__EVAL_5 = Queue_1__EVAL_5;
  assign TLMonitor__EVAL_6 = Queue_1__EVAL_4;
  assign TLMonitor__EVAL_18 = _EVAL_11;
  assign TLMonitor__EVAL_0 = Queue_1__EVAL_3;
  assign TLMonitor__EVAL_4 = Queue_1__EVAL_15;
  assign TLMonitor__EVAL_16 = _EVAL_36;
  assign TLMonitor__EVAL_3 = _EVAL_7;
  assign TLMonitor__EVAL_15 = _EVAL_22;
  assign TLMonitor__EVAL_1 = Queue_1__EVAL_11;
  assign TLMonitor__EVAL_9 = _EVAL_12;
  assign TLMonitor__EVAL_10 = _EVAL_9;
  assign TLMonitor__EVAL_11 = _EVAL_37;
  assign TLMonitor__EVAL_14 = _EVAL_2;
  assign TLMonitor__EVAL_2 = Queue_1__EVAL_17;
  assign TLMonitor__EVAL_13 = _EVAL_3;
  assign TLMonitor__EVAL_8 = Queue__EVAL_4;

endmodule
