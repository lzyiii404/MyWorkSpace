//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_34_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [7:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [30:0] _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [6:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [6:0]  _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_35;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_47;
  reg [31:0] _RAND_1;
  reg [6:0] _EVAL_51;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_113;
  reg [31:0] _RAND_3;
  reg  _EVAL_115;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_132;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_170;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_227;
  reg [31:0] _RAND_7;
  reg [30:0] _EVAL_240;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_248;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_251;
  reg [31:0] _RAND_10;
  reg [72:0] _EVAL_260;
  reg [95:0] _RAND_11;
  reg [6:0] _EVAL_278;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_295;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_324;
  reg [31:0] _RAND_14;
  wire [7:0] _EVAL_123;
  wire  _EVAL_312;
  wire  _EVAL_274;
  wire  _EVAL_283;
  wire  _EVAL_310;
  wire  _EVAL_202;
  wire  _EVAL_66;
  wire  _EVAL_99;
  wire [2:0] _EVAL_74;
  wire  _EVAL_166;
  wire  _EVAL_65;
  wire  _EVAL_130;
  wire  _EVAL_294;
  wire  _EVAL_127;
  wire [127:0] _EVAL_231;
  wire  _EVAL_242;
  wire  _EVAL_302;
  wire  _EVAL_168;
  wire  _EVAL_280;
  wire  _EVAL_33;
  wire [1:0] _EVAL_31;
  wire [3:0] _EVAL_134;
  wire [2:0] _EVAL_270;
  wire [2:0] _EVAL_330;
  wire  _EVAL_321;
  wire  _EVAL_271;
  wire  _EVAL_18;
  wire  _EVAL_315;
  wire  _EVAL_304;
  wire  _EVAL_228;
  wire  _EVAL_20;
  wire  _EVAL_298;
  wire  _EVAL_322;
  wire  _EVAL_284;
  wire  _EVAL_84;
  wire  _EVAL_275;
  wire  _EVAL_241;
  wire  _EVAL_329;
  wire  _EVAL_128;
  wire  _EVAL_316;
  wire  _EVAL_38;
  wire  _EVAL_229;
  wire  _EVAL_208;
  wire  _EVAL_263;
  wire  _EVAL_44;
  wire  _EVAL_68;
  wire  _EVAL_210;
  wire  _EVAL_186;
  wire  _EVAL_61;
  wire  _EVAL_89;
  wire  _EVAL_225;
  wire  _EVAL_60;
  wire  _EVAL_303;
  wire  _EVAL_237;
  wire  _EVAL_101;
  wire  _EVAL_238;
  wire  _EVAL_296;
  wire  _EVAL_48;
  wire  _EVAL_78;
  wire  _EVAL_254;
  wire  _EVAL_159;
  wire  _EVAL_222;
  wire  _EVAL_175;
  wire  _EVAL_328;
  wire  _EVAL_24;
  wire  _EVAL_158;
  wire  _EVAL_189;
  wire  _EVAL_37;
  wire  _EVAL_146;
  wire  _EVAL_286;
  wire  _EVAL_323;
  wire  _EVAL_67;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_156;
  wire  _EVAL_211;
  wire [7:0] _EVAL_39;
  wire [7:0] _EVAL_73;
  wire [7:0] _EVAL_59;
  wire  _EVAL_182;
  wire  _EVAL_326;
  wire  _EVAL_221;
  wire [2:0] _EVAL_178;
  wire [12:0] _EVAL_252;
  wire [5:0] _EVAL_309;
  wire [5:0] _EVAL_224;
  wire  _EVAL_95;
  wire  _EVAL_90;
  wire  _EVAL_288;
  wire  _EVAL_285;
  wire [2:0] _EVAL_45;
  wire  _EVAL_150;
  wire [12:0] _EVAL_169;
  wire [5:0] _EVAL_261;
  wire [5:0] _EVAL_291;
  wire [2:0] _EVAL_58;
  wire  _EVAL_318;
  wire  _EVAL_107;
  wire [31:0] _EVAL_198;
  wire [3:0] _EVAL_267;
  wire  _EVAL_234;
  wire  _EVAL_163;
  wire  _EVAL_119;
  wire  _EVAL_56;
  wire [3:0] _EVAL_147;
  wire  _EVAL_257;
  wire [2:0] _EVAL_193;
  wire  _EVAL_218;
  wire  _EVAL_292;
  wire  _EVAL_171;
  wire  _EVAL_49;
  wire  _EVAL_75;
  wire  _EVAL_97;
  wire  _EVAL_64;
  wire  _EVAL_103;
  wire  _EVAL_319;
  wire  _EVAL_290;
  wire  _EVAL_181;
  wire [127:0] _EVAL_149;
  wire  _EVAL_276;
  wire  _EVAL_53;
  wire  _EVAL_161;
  wire  _EVAL_183;
  wire  _EVAL_214;
  wire  _EVAL_122;
  wire [127:0] _EVAL_282;
  wire [72:0] _EVAL_300;
  wire  _EVAL_105;
  wire  _EVAL_143;
  wire  _EVAL_138;
  wire  _EVAL_55;
  wire  _EVAL_141;
  wire [127:0] _EVAL_86;
  wire [72:0] _EVAL_69;
  wire  _EVAL_54;
  wire  _EVAL_287;
  wire  _EVAL_76;
  wire [2:0] _EVAL_77;
  wire [72:0] _EVAL_165;
  wire  _EVAL_129;
  wire  _EVAL_30;
  wire  _EVAL_92;
  wire  _EVAL_188;
  wire  _EVAL_177;
  wire  _EVAL_83;
  wire [2:0] _EVAL_230;
  wire  _EVAL_87;
  wire  _EVAL_157;
  wire  _EVAL_26;
  wire  _EVAL_206;
  wire  _EVAL_245;
  wire  _EVAL_293;
  wire  _EVAL_301;
  wire  _EVAL_41;
  wire  _EVAL_111;
  wire  _EVAL_43;
  wire  _EVAL_209;
  wire  _EVAL_162;
  wire  _EVAL_80;
  wire  _EVAL_137;
  wire  _EVAL_320;
  wire  _EVAL_88;
  wire [2:0] _EVAL_289;
  wire  _EVAL_307;
  wire  _EVAL_223;
  wire  _EVAL_255;
  wire  _EVAL_313;
  wire  _EVAL_144;
  wire  _EVAL_154;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_19;
  wire  _EVAL_139;
  wire  _EVAL_277;
  wire  _EVAL_314;
  wire  _EVAL_265;
  wire [30:0] _EVAL_174;
  wire [31:0] _EVAL_79;
  wire [31:0] _EVAL_195;
  wire [31:0] _EVAL_172;
  wire  _EVAL_199;
  wire  _EVAL_71;
  wire  _EVAL_308;
  wire  _EVAL_262;
  wire  _EVAL_212;
  wire  _EVAL_120;
  wire  _EVAL_116;
  wire  _EVAL_125;
  wire  _EVAL_269;
  wire  _EVAL_217;
  wire  _EVAL_190;
  wire  _EVAL_21;
  wire  _EVAL_164;
  wire [72:0] _EVAL_327;
  wire [72:0] _EVAL_331;
  wire  _EVAL_179;
  wire  _EVAL_133;
  wire  _EVAL_243;
  wire  _EVAL_63;
  wire  _EVAL_23;
  wire  _EVAL_299;
  wire  _EVAL_136;
  wire  _EVAL_94;
  wire  _EVAL_256;
  wire  _EVAL_215;
  wire  _EVAL_268;
  wire [30:0] _EVAL_259;
  wire [30:0] _EVAL_180;
  wire  _EVAL_197;
  wire  _EVAL_140;
  wire  _EVAL_100;
  wire  _EVAL_264;
  wire [72:0] _EVAL_42;
  wire [72:0] _EVAL_249;
  wire [72:0] _EVAL_233;
  wire  _EVAL_239;
  wire  _EVAL_118;
  wire  _EVAL_184;
  wire  _EVAL_213;
  wire  _EVAL_108;
  wire  _EVAL_226;
  wire  _EVAL_325;
  wire  _EVAL_273;
  wire  _EVAL_17;
  wire  _EVAL_176;
  wire  _EVAL_152;
  wire  _EVAL_194;
  wire  _EVAL_148;
  wire  _EVAL_279;
  wire  _EVAL_297;
  wire  _EVAL_98;
  wire  _EVAL_29;
  wire  _EVAL_85;
  wire  _EVAL_121;
  wire  _EVAL_185;
  wire  _EVAL_50;
  wire  _EVAL_81;
  wire  _EVAL_236;
  wire  _EVAL_205;
  wire  _EVAL_203;
  wire  _EVAL_96;
  wire  _EVAL_82;
  wire  _EVAL_216;
  wire  _EVAL_32;
  wire  _EVAL_109;
  wire  _EVAL_196;
  wire  _EVAL_253;
  wire  _EVAL_160;
  wire  _EVAL_52;
  wire  _EVAL_258;
  wire  _EVAL_167;
  wire  _EVAL_151;
  wire  _EVAL_306;
  wire  _EVAL_27;
  wire  _EVAL_246;
  wire  _EVAL_201;
  wire  _EVAL_187;
  wire  _EVAL_244;
  wire  _EVAL_207;
  wire  _EVAL_110;
  wire  _EVAL_70;
  wire  _EVAL_22;
  wire  _EVAL_155;
  wire  _EVAL_91;
  wire  _EVAL_235;
  wire  _EVAL_142;
  wire  _EVAL_153;
  wire  _EVAL_72;
  wire  _EVAL_106;
  wire  _EVAL_145;
  wire  _EVAL_131;
  wire  _EVAL_281;
  wire  _EVAL_25;
  wire  _EVAL_36;
  wire  _EVAL_40;
  wire  _EVAL_232;
  wire  _EVAL_28;
  wire  _EVAL_204;
  wire  _EVAL_220;
  wire  _EVAL_250;
  wire  _EVAL_135;
  wire  _EVAL_93;
  wire  _EVAL_247;
  wire  _EVAL_272;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_123 = ~ _EVAL_5;
  assign _EVAL_312 = _EVAL_123 == 8'h0;
  assign _EVAL_274 = _EVAL_312 | _EVAL_1;
  assign _EVAL_283 = _EVAL_35 == 3'h0;
  assign _EVAL_310 = _EVAL_283 == 1'h0;
  assign _EVAL_202 = _EVAL_0 == 3'h1;
  assign _EVAL_66 = _EVAL_8 & _EVAL_202;
  assign _EVAL_99 = _EVAL_11 != 3'h0;
  assign _EVAL_74 = _EVAL_35 - 3'h1;
  assign _EVAL_166 = _EVAL & _EVAL_8;
  assign _EVAL_65 = _EVAL_170 == 3'h0;
  assign _EVAL_130 = _EVAL_166 & _EVAL_65;
  assign _EVAL_294 = _EVAL_9[0];
  assign _EVAL_127 = _EVAL_294 == 1'h0;
  assign _EVAL_231 = 128'h1 << _EVAL_15;
  assign _EVAL_242 = _EVAL_260 != 73'h0;
  assign _EVAL_302 = _EVAL_242 == 1'h0;
  assign _EVAL_168 = plusarg_reader_out == 32'h0;
  assign _EVAL_280 = _EVAL_302 | _EVAL_168;
  assign _EVAL_33 = _EVAL_2 >= 3'h3;
  assign _EVAL_31 = _EVAL_2[1:0];
  assign _EVAL_134 = 4'h1 << _EVAL_31;
  assign _EVAL_270 = _EVAL_134[2:0];
  assign _EVAL_330 = _EVAL_270 | 3'h1;
  assign _EVAL_321 = _EVAL_330[2];
  assign _EVAL_271 = _EVAL_9[2];
  assign _EVAL_18 = _EVAL_321 & _EVAL_271;
  assign _EVAL_315 = _EVAL_33 | _EVAL_18;
  assign _EVAL_304 = _EVAL_330[1];
  assign _EVAL_228 = _EVAL_9[1];
  assign _EVAL_20 = _EVAL_271 & _EVAL_228;
  assign _EVAL_298 = _EVAL_304 & _EVAL_20;
  assign _EVAL_322 = _EVAL_315 | _EVAL_298;
  assign _EVAL_284 = _EVAL_330[0];
  assign _EVAL_84 = _EVAL_20 & _EVAL_127;
  assign _EVAL_275 = _EVAL_284 & _EVAL_84;
  assign _EVAL_241 = _EVAL_322 | _EVAL_275;
  assign _EVAL_329 = _EVAL_11 == 3'h0;
  assign _EVAL_128 = _EVAL_329 | _EVAL_1;
  assign _EVAL_316 = _EVAL_128 == 1'h0;
  assign _EVAL_38 = _EVAL_11 == _EVAL_47;
  assign _EVAL_229 = _EVAL_38 | _EVAL_1;
  assign _EVAL_208 = _EVAL_20 & _EVAL_294;
  assign _EVAL_263 = _EVAL_284 & _EVAL_208;
  assign _EVAL_44 = _EVAL_322 | _EVAL_263;
  assign _EVAL_68 = _EVAL_228 == 1'h0;
  assign _EVAL_210 = _EVAL_271 & _EVAL_68;
  assign _EVAL_186 = _EVAL_304 & _EVAL_210;
  assign _EVAL_61 = _EVAL_315 | _EVAL_186;
  assign _EVAL_89 = _EVAL_210 & _EVAL_294;
  assign _EVAL_225 = _EVAL_284 & _EVAL_89;
  assign _EVAL_60 = _EVAL_61 | _EVAL_225;
  assign _EVAL_303 = _EVAL_210 & _EVAL_127;
  assign _EVAL_237 = _EVAL_284 & _EVAL_303;
  assign _EVAL_101 = _EVAL_61 | _EVAL_237;
  assign _EVAL_238 = _EVAL_271 == 1'h0;
  assign _EVAL_296 = _EVAL_321 & _EVAL_238;
  assign _EVAL_48 = _EVAL_33 | _EVAL_296;
  assign _EVAL_78 = _EVAL_238 & _EVAL_228;
  assign _EVAL_254 = _EVAL_304 & _EVAL_78;
  assign _EVAL_159 = _EVAL_48 | _EVAL_254;
  assign _EVAL_222 = _EVAL_78 & _EVAL_294;
  assign _EVAL_175 = _EVAL_284 & _EVAL_222;
  assign _EVAL_328 = _EVAL_159 | _EVAL_175;
  assign _EVAL_24 = _EVAL_78 & _EVAL_127;
  assign _EVAL_158 = _EVAL_284 & _EVAL_24;
  assign _EVAL_189 = _EVAL_159 | _EVAL_158;
  assign _EVAL_37 = _EVAL_238 & _EVAL_68;
  assign _EVAL_146 = _EVAL_304 & _EVAL_37;
  assign _EVAL_286 = _EVAL_48 | _EVAL_146;
  assign _EVAL_323 = _EVAL_37 & _EVAL_294;
  assign _EVAL_67 = _EVAL_284 & _EVAL_323;
  assign _EVAL_112 = _EVAL_286 | _EVAL_67;
  assign _EVAL_114 = _EVAL_37 & _EVAL_127;
  assign _EVAL_156 = _EVAL_284 & _EVAL_114;
  assign _EVAL_211 = _EVAL_286 | _EVAL_156;
  assign _EVAL_39 = {_EVAL_44,_EVAL_241,_EVAL_60,_EVAL_101,_EVAL_328,_EVAL_189,_EVAL_112,_EVAL_211};
  assign _EVAL_73 = ~ _EVAL_39;
  assign _EVAL_59 = _EVAL_5 & _EVAL_73;
  assign _EVAL_182 = _EVAL_59 == 8'h0;
  assign _EVAL_326 = _EVAL_182 | _EVAL_1;
  assign _EVAL_221 = _EVAL_326 == 1'h0;
  assign _EVAL_178 = _EVAL_170 - 3'h1;
  assign _EVAL_252 = 13'h3f << _EVAL_2;
  assign _EVAL_309 = _EVAL_252[5:0];
  assign _EVAL_224 = ~ _EVAL_309;
  assign _EVAL_95 = _EVAL_12 == 1'h0;
  assign _EVAL_90 = _EVAL_2 <= 3'h6;
  assign _EVAL_288 = _EVAL_0[2];
  assign _EVAL_285 = _EVAL_288 == 1'h0;
  assign _EVAL_45 = _EVAL_224[5:3];
  assign _EVAL_150 = _EVAL_14[0];
  assign _EVAL_169 = 13'h3f << _EVAL_4;
  assign _EVAL_261 = _EVAL_169[5:0];
  assign _EVAL_291 = ~ _EVAL_261;
  assign _EVAL_58 = _EVAL_291[5:3];
  assign _EVAL_318 = _EVAL_6 & _EVAL_7;
  assign _EVAL_107 = _EVAL_166 | _EVAL_318;
  assign _EVAL_198 = _EVAL_227 + 32'h1;
  assign _EVAL_267 = _EVAL_13[6:3];
  assign _EVAL_234 = _EVAL_267 == 4'h8;
  assign _EVAL_163 = _EVAL_15 == 7'h48;
  assign _EVAL_119 = _EVAL_15 == 7'h40;
  assign _EVAL_56 = _EVAL_163 | _EVAL_119;
  assign _EVAL_147 = _EVAL_15[6:3];
  assign _EVAL_257 = _EVAL_147 == 4'h8;
  assign _EVAL_193 = _EVAL_15[2:0];
  assign _EVAL_218 = 3'h1 <= _EVAL_193;
  assign _EVAL_292 = _EVAL_257 & _EVAL_218;
  assign _EVAL_171 = _EVAL_56 | _EVAL_292;
  assign _EVAL_49 = _EVAL_15 == 7'h20;
  assign _EVAL_75 = _EVAL_171 | _EVAL_49;
  assign _EVAL_97 = _EVAL_11 <= 3'h4;
  assign _EVAL_64 = _EVAL_97 | _EVAL_1;
  assign _EVAL_103 = _EVAL_64 == 1'h0;
  assign _EVAL_319 = _EVAL_147 == 4'h1;
  assign _EVAL_290 = _EVAL_14 == 3'h1;
  assign _EVAL_181 = _EVAL_7 & _EVAL_290;
  assign _EVAL_149 = 128'h1 << _EVAL_13;
  assign _EVAL_276 = _EVAL_0 == 3'h0;
  assign _EVAL_53 = _EVAL_8 & _EVAL_276;
  assign _EVAL_161 = _EVAL_3 == 1'h0;
  assign _EVAL_183 = _EVAL_161 | _EVAL_16;
  assign _EVAL_214 = _EVAL_183 | _EVAL_1;
  assign _EVAL_122 = _EVAL_214 == 1'h0;
  assign _EVAL_282 = _EVAL_130 ? _EVAL_231 : 128'h0;
  assign _EVAL_300 = _EVAL_282[72:0];
  assign _EVAL_105 = _EVAL_132 == 3'h0;
  assign _EVAL_143 = _EVAL_318 & _EVAL_105;
  assign _EVAL_138 = _EVAL_14 == 3'h6;
  assign _EVAL_55 = _EVAL_138 == 1'h0;
  assign _EVAL_141 = _EVAL_143 & _EVAL_55;
  assign _EVAL_86 = _EVAL_141 ? _EVAL_149 : 128'h0;
  assign _EVAL_69 = _EVAL_86[72:0];
  assign _EVAL_54 = _EVAL_300 != _EVAL_69;
  assign _EVAL_287 = _EVAL_15 == _EVAL_51;
  assign _EVAL_76 = _EVAL_248 == 3'h0;
  assign _EVAL_77 = _EVAL_248 - 3'h1;
  assign _EVAL_165 = _EVAL_260 >> _EVAL_15;
  assign _EVAL_129 = _EVAL_165[0];
  assign _EVAL_30 = _EVAL_129 == 1'h0;
  assign _EVAL_92 = _EVAL_227 < plusarg_reader_out;
  assign _EVAL_188 = _EVAL_280 | _EVAL_92;
  assign _EVAL_177 = _EVAL_13 == 7'h20;
  assign _EVAL_83 = _EVAL_0 == 3'h2;
  assign _EVAL_230 = _EVAL_13[2:0];
  assign _EVAL_87 = _EVAL_13 == 7'h48;
  assign _EVAL_157 = _EVAL_13 == 7'h40;
  assign _EVAL_26 = _EVAL_87 | _EVAL_157;
  assign _EVAL_206 = 3'h1 <= _EVAL_230;
  assign _EVAL_245 = _EVAL_234 & _EVAL_206;
  assign _EVAL_293 = _EVAL_26 | _EVAL_245;
  assign _EVAL_301 = _EVAL_293 | _EVAL_177;
  assign _EVAL_41 = _EVAL_267 == 4'h0;
  assign _EVAL_111 = _EVAL_301 | _EVAL_41;
  assign _EVAL_43 = _EVAL_267 == 4'h1;
  assign _EVAL_209 = _EVAL_111 | _EVAL_43;
  assign _EVAL_162 = _EVAL_267 == 4'h2;
  assign _EVAL_80 = _EVAL_209 | _EVAL_162;
  assign _EVAL_137 = _EVAL_267 == 4'h3;
  assign _EVAL_320 = _EVAL_80 | _EVAL_137;
  assign _EVAL_88 = _EVAL_320 | _EVAL_1;
  assign _EVAL_289 = _EVAL_132 - 3'h1;
  assign _EVAL_307 = _EVAL_0 == _EVAL_324;
  assign _EVAL_223 = _EVAL_307 | _EVAL_1;
  assign _EVAL_255 = _EVAL_223 == 1'h0;
  assign _EVAL_313 = _EVAL_14 <= 3'h6;
  assign _EVAL_144 = _EVAL_300 != 73'h0;
  assign _EVAL_154 = _EVAL_144 == 1'h0;
  assign _EVAL_191 = _EVAL_54 | _EVAL_154;
  assign _EVAL_192 = _EVAL_191 | _EVAL_1;
  assign _EVAL_19 = _EVAL_192 == 1'h0;
  assign _EVAL_139 = _EVAL_7 & _EVAL_138;
  assign _EVAL_277 = _EVAL_161 | _EVAL_1;
  assign _EVAL_314 = _EVAL_11 <= 3'h2;
  assign _EVAL_265 = _EVAL_314 | _EVAL_1;
  assign _EVAL_174 = _EVAL_9 ^ 31'h40000000;
  assign _EVAL_79 = {1'b0,$signed(_EVAL_174)};
  assign _EVAL_195 = $signed(_EVAL_79) & $signed(-32'sh2000);
  assign _EVAL_172 = $signed(_EVAL_195);
  assign _EVAL_199 = $signed(_EVAL_172) == $signed(32'sh0);
  assign _EVAL_71 = _EVAL_90 & _EVAL_199;
  assign _EVAL_308 = _EVAL_71 | _EVAL_1;
  assign _EVAL_262 = _EVAL_147 == 4'h0;
  assign _EVAL_212 = _EVAL_75 | _EVAL_262;
  assign _EVAL_120 = _EVAL_212 | _EVAL_319;
  assign _EVAL_116 = _EVAL_147 == 4'h2;
  assign _EVAL_125 = _EVAL_120 | _EVAL_116;
  assign _EVAL_269 = _EVAL_147 == 4'h3;
  assign _EVAL_217 = _EVAL_125 | _EVAL_269;
  assign _EVAL_190 = _EVAL_11 <= 3'h3;
  assign _EVAL_21 = _EVAL_190 | _EVAL_1;
  assign _EVAL_164 = _EVAL_313 | _EVAL_1;
  assign _EVAL_327 = _EVAL_300 | _EVAL_260;
  assign _EVAL_331 = _EVAL_327 >> _EVAL_13;
  assign _EVAL_179 = _EVAL_331[0];
  assign _EVAL_133 = _EVAL_179 | _EVAL_1;
  assign _EVAL_243 = _EVAL_133 == 1'h0;
  assign _EVAL_63 = _EVAL_33 | _EVAL_1;
  assign _EVAL_23 = _EVAL_16 == 1'h0;
  assign _EVAL_299 = _EVAL_14 == _EVAL_251;
  assign _EVAL_136 = _EVAL_299 | _EVAL_1;
  assign _EVAL_94 = _EVAL_274 == 1'h0;
  assign _EVAL_256 = _EVAL_5 == _EVAL_39;
  assign _EVAL_215 = _EVAL_256 | _EVAL_1;
  assign _EVAL_268 = _EVAL_215 == 1'h0;
  assign _EVAL_259 = {{25'd0}, _EVAL_224};
  assign _EVAL_180 = _EVAL_9 & _EVAL_259;
  assign _EVAL_197 = _EVAL_180 == 31'h0;
  assign _EVAL_140 = _EVAL_3 == _EVAL_115;
  assign _EVAL_100 = _EVAL_140 | _EVAL_1;
  assign _EVAL_264 = _EVAL_100 == 1'h0;
  assign _EVAL_42 = _EVAL_260 | _EVAL_300;
  assign _EVAL_249 = ~ _EVAL_69;
  assign _EVAL_233 = _EVAL_42 & _EVAL_249;
  assign _EVAL_239 = _EVAL_287 | _EVAL_1;
  assign _EVAL_118 = _EVAL_0 == 3'h6;
  assign _EVAL_184 = _EVAL_8 & _EVAL_118;
  assign _EVAL_213 = _EVAL_14 == 3'h2;
  assign _EVAL_108 = _EVAL_7 & _EVAL_213;
  assign _EVAL_226 = _EVAL_229 == 1'h0;
  assign _EVAL_325 = _EVAL_95 | _EVAL_1;
  assign _EVAL_273 = _EVAL_325 == 1'h0;
  assign _EVAL_17 = _EVAL_2 == _EVAL_295;
  assign _EVAL_176 = _EVAL_17 | _EVAL_1;
  assign _EVAL_152 = _EVAL_176 == 1'h0;
  assign _EVAL_194 = _EVAL_14 == 3'h0;
  assign _EVAL_148 = _EVAL_7 & _EVAL_194;
  assign _EVAL_279 = _EVAL_9 == _EVAL_240;
  assign _EVAL_297 = _EVAL_279 | _EVAL_1;
  assign _EVAL_98 = _EVAL_318 & _EVAL_283;
  assign _EVAL_29 = _EVAL_13 == _EVAL_278;
  assign _EVAL_85 = _EVAL_29 | _EVAL_1;
  assign _EVAL_121 = _EVAL_85 == 1'h0;
  assign _EVAL_185 = _EVAL_30 | _EVAL_1;
  assign _EVAL_50 = _EVAL_0 == 3'h3;
  assign _EVAL_81 = _EVAL_8 & _EVAL_50;
  assign _EVAL_236 = _EVAL_99 | _EVAL_1;
  assign _EVAL_205 = _EVAL_236 == 1'h0;
  assign _EVAL_203 = _EVAL_308 == 1'h0;
  assign _EVAL_96 = _EVAL_14 == 3'h5;
  assign _EVAL_82 = _EVAL_0 == 3'h5;
  assign _EVAL_216 = _EVAL_8 & _EVAL_82;
  assign _EVAL_32 = _EVAL_0 == 3'h7;
  assign _EVAL_109 = _EVAL_88 == 1'h0;
  assign _EVAL_196 = _EVAL_166 & _EVAL_76;
  assign _EVAL_253 = _EVAL_185 == 1'h0;
  assign _EVAL_160 = _EVAL_4 == _EVAL_113;
  assign _EVAL_52 = _EVAL_160 | _EVAL_1;
  assign _EVAL_258 = 3'h6 == _EVAL_2;
  assign _EVAL_167 = _EVAL_119 ? _EVAL_258 : 1'h0;
  assign _EVAL_151 = _EVAL_167 | _EVAL_1;
  assign _EVAL_306 = _EVAL_151 == 1'h0;
  assign _EVAL_27 = _EVAL_239 == 1'h0;
  assign _EVAL_246 = _EVAL_8 & _EVAL_83;
  assign _EVAL_201 = _EVAL_136 == 1'h0;
  assign _EVAL_187 = _EVAL_197 | _EVAL_1;
  assign _EVAL_244 = _EVAL_187 == 1'h0;
  assign _EVAL_207 = _EVAL_76 == 1'h0;
  assign _EVAL_110 = _EVAL_8 & _EVAL_207;
  assign _EVAL_70 = _EVAL_0 == 3'h4;
  assign _EVAL_22 = _EVAL_188 | _EVAL_1;
  assign _EVAL_155 = _EVAL_1 == 1'h0;
  assign _EVAL_91 = _EVAL_23 | _EVAL_1;
  assign _EVAL_235 = _EVAL_91 == 1'h0;
  assign _EVAL_142 = _EVAL_164 == 1'h0;
  assign _EVAL_153 = _EVAL_8 & _EVAL_70;
  assign _EVAL_72 = _EVAL_14 == 3'h4;
  assign _EVAL_106 = _EVAL_277 == 1'h0;
  assign _EVAL_145 = _EVAL_217 | _EVAL_1;
  assign _EVAL_131 = _EVAL_4 >= 3'h3;
  assign _EVAL_281 = _EVAL_52 == 1'h0;
  assign _EVAL_25 = _EVAL_131 | _EVAL_1;
  assign _EVAL_36 = _EVAL_25 == 1'h0;
  assign _EVAL_40 = _EVAL_7 & _EVAL_310;
  assign _EVAL_232 = _EVAL_21 == 1'h0;
  assign _EVAL_28 = _EVAL_7 & _EVAL_72;
  assign _EVAL_204 = _EVAL_265 == 1'h0;
  assign _EVAL_220 = _EVAL_22 == 1'h0;
  assign _EVAL_250 = _EVAL_297 == 1'h0;
  assign _EVAL_135 = _EVAL_145 == 1'h0;
  assign _EVAL_93 = _EVAL_8 & _EVAL_32;
  assign _EVAL_247 = _EVAL_7 & _EVAL_96;
  assign _EVAL_272 = _EVAL_63 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_35 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_47 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_51 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_113 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_115 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_132 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_170 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_227 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_240 = _RAND_8[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_248 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_251 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {3{`RANDOM}};
  _EVAL_260 = _RAND_11[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_278 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_295 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_324 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_10) begin
    if (_EVAL_1) begin
      _EVAL_35 <= 3'h0;
    end else begin
      if (_EVAL_318) begin
        if (_EVAL_283) begin
          if (_EVAL_150) begin
            _EVAL_35 <= _EVAL_58;
          end else begin
            _EVAL_35 <= 3'h0;
          end
        end else begin
          _EVAL_35 <= _EVAL_74;
        end
      end
    end
    if (_EVAL_196) begin
      _EVAL_47 <= _EVAL_11;
    end
    if (_EVAL_196) begin
      _EVAL_51 <= _EVAL_15;
    end
    if (_EVAL_98) begin
      _EVAL_113 <= _EVAL_4;
    end
    if (_EVAL_98) begin
      _EVAL_115 <= _EVAL_3;
    end
    if (_EVAL_1) begin
      _EVAL_132 <= 3'h0;
    end else begin
      if (_EVAL_318) begin
        if (_EVAL_105) begin
          if (_EVAL_150) begin
            _EVAL_132 <= _EVAL_58;
          end else begin
            _EVAL_132 <= 3'h0;
          end
        end else begin
          _EVAL_132 <= _EVAL_289;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_170 <= 3'h0;
    end else begin
      if (_EVAL_166) begin
        if (_EVAL_65) begin
          if (_EVAL_285) begin
            _EVAL_170 <= _EVAL_45;
          end else begin
            _EVAL_170 <= 3'h0;
          end
        end else begin
          _EVAL_170 <= _EVAL_178;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_227 <= 32'h0;
    end else begin
      if (_EVAL_107) begin
        _EVAL_227 <= 32'h0;
      end else begin
        _EVAL_227 <= _EVAL_198;
      end
    end
    if (_EVAL_196) begin
      _EVAL_240 <= _EVAL_9;
    end
    if (_EVAL_1) begin
      _EVAL_248 <= 3'h0;
    end else begin
      if (_EVAL_166) begin
        if (_EVAL_76) begin
          if (_EVAL_285) begin
            _EVAL_248 <= _EVAL_45;
          end else begin
            _EVAL_248 <= 3'h0;
          end
        end else begin
          _EVAL_248 <= _EVAL_77;
        end
      end
    end
    if (_EVAL_98) begin
      _EVAL_251 <= _EVAL_14;
    end
    if (_EVAL_1) begin
      _EVAL_260 <= 73'h0;
    end else begin
      _EVAL_260 <= _EVAL_233;
    end
    if (_EVAL_98) begin
      _EVAL_278 <= _EVAL_13;
    end
    if (_EVAL_196) begin
      _EVAL_295 <= _EVAL_2;
    end
    if (_EVAL_196) begin
      _EVAL_324 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ef356c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4a75bd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f467d77a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f71a3ab6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f51584b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c16c105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4c241fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c1c8aa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(905e7e3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf5bf044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c290e3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b780fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(168ca410)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8835be42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b484f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d317a93b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4c3f0cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d317b874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35736f01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7f4d543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feaa085e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ce43c39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25e8d8da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0950ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(814c0bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be987ff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3815352f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5fc133d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(210d240b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2815b3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(899a0b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a4391e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb64fa40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e6d1acc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61e0214f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaba50a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb51a35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a425f59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c39d62f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3216d65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f66e62e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a5de2af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23370815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a58cce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5e56b62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57b385c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71939e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6632e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0fb2f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61a0bd46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(394bcd60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(271be4c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b84ce40c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb1501c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6002024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9ba313a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30a3441c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(822cbee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c00bc045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0fcedf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eb770b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b2703a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(808af58c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54063205)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5af380a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc0c798)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15f1993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad724b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb8c432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78dc8ed3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4a55021)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83c68e65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e746b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30da9593)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16a7cada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(802f1cc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c4445ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc32fb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a4d080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0aeaf90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
