//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_290(
  input  [9:0]  _EVAL,
  input         _EVAL_0,
  output [4:0]  _EVAL_1,
  output [32:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [26:0] _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9
);
  wire  _EVAL_111;
  wire [8:0] _EVAL_131;
  wire [8:0] _EVAL_148;
  wire  _EVAL_110;
  wire [7:0] _EVAL_122;
  wire  _EVAL_33;
  wire [6:0] _EVAL_167;
  wire  _EVAL_100;
  wire [5:0] _EVAL_128;
  wire [64:0] _EVAL_45;
  wire [21:0] _EVAL_27;
  wire [15:0] _EVAL_162;
  wire [7:0] _EVAL_120;
  wire [15:0] _EVAL_207;
  wire [7:0] _EVAL_105;
  wire [15:0] _EVAL_133;
  wire [15:0] _EVAL_12;
  wire [15:0] _EVAL_14;
  wire [11:0] _EVAL_141;
  wire [15:0] _EVAL_53;
  wire [15:0] _EVAL_177;
  wire [11:0] _EVAL_178;
  wire [15:0] _EVAL_37;
  wire [15:0] _EVAL_49;
  wire [15:0] _EVAL_140;
  wire [13:0] _EVAL_58;
  wire [15:0] _EVAL_156;
  wire [15:0] _EVAL_164;
  wire [13:0] _EVAL_41;
  wire [15:0] _EVAL_174;
  wire [15:0] _EVAL_59;
  wire [15:0] _EVAL_69;
  wire [14:0] _EVAL_206;
  wire [15:0] _EVAL_79;
  wire [15:0] _EVAL_127;
  wire [14:0] _EVAL_86;
  wire [15:0] _EVAL_106;
  wire [15:0] _EVAL_60;
  wire [15:0] _EVAL_47;
  wire [5:0] _EVAL_194;
  wire [3:0] _EVAL_43;
  wire [1:0] _EVAL_143;
  wire  _EVAL_138;
  wire  _EVAL_152;
  wire [1:0] _EVAL_129;
  wire  _EVAL_201;
  wire  _EVAL_65;
  wire [1:0] _EVAL_67;
  wire  _EVAL_17;
  wire  _EVAL_48;
  wire [21:0] _EVAL_132;
  wire [21:0] _EVAL_57;
  wire [21:0] _EVAL_118;
  wire [21:0] _EVAL_30;
  wire [24:0] _EVAL_189;
  wire [2:0] _EVAL_180;
  wire [1:0] _EVAL_179;
  wire  _EVAL_96;
  wire  _EVAL_63;
  wire  _EVAL_181;
  wire [2:0] _EVAL_169;
  wire [2:0] _EVAL_104;
  wire [24:0] _EVAL_154;
  wire [24:0] _EVAL_11;
  wire [24:0] _EVAL_190;
  wire [24:0] _EVAL_40;
  wire [26:0] _EVAL_16;
  wire  _EVAL_42;
  wire  _EVAL_117;
  wire  _EVAL_44;
  wire  _EVAL_72;
  wire  _EVAL_83;
  wire  _EVAL_66;
  wire  _EVAL_184;
  wire  _EVAL_87;
  wire  _EVAL_193;
  wire  _EVAL_25;
  wire  _EVAL_39;
  wire  _EVAL_191;
  wire  _EVAL_20;
  wire [25:0] _EVAL_52;
  wire [26:0] _EVAL_205;
  wire [26:0] _EVAL_26;
  wire [26:0] _EVAL_89;
  wire [26:0] _EVAL_204;
  wire  _EVAL_168;
  wire  _EVAL_70;
  wire  _EVAL_91;
  wire  _EVAL_123;
  wire  _EVAL_74;
  wire  _EVAL_173;
  wire  _EVAL_98;
  wire  _EVAL_81;
  wire [26:0] _EVAL_125;
  wire  _EVAL_88;
  wire  _EVAL_172;
  wire  _EVAL_90;
  wire  _EVAL_197;
  wire [26:0] _EVAL_166;
  wire [24:0] _EVAL_71;
  wire [25:0] _EVAL_61;
  wire  _EVAL_163;
  wire  _EVAL_115;
  wire  _EVAL_56;
  wire [25:0] _EVAL_85;
  wire [25:0] _EVAL_97;
  wire [25:0] _EVAL_198;
  wire [26:0] _EVAL_73;
  wire [26:0] _EVAL_203;
  wire [24:0] _EVAL_92;
  wire [25:0] _EVAL_158;
  wire  _EVAL_196;
  wire  _EVAL_54;
  wire [25:0] _EVAL_34;
  wire [25:0] _EVAL_13;
  wire [25:0] _EVAL_137;
  wire [25:0] _EVAL_84;
  wire [1:0] _EVAL_80;
  wire [2:0] _EVAL_121;
  wire [9:0] _EVAL_36;
  wire [10:0] _EVAL_82;
  wire [3:0] _EVAL_157;
  wire  _EVAL_22;
  wire  _EVAL_119;
  wire  _EVAL_202;
  wire  _EVAL_139;
  wire  _EVAL_31;
  wire [8:0] _EVAL_38;
  wire [1:0] _EVAL_29;
  wire  _EVAL_64;
  wire  _EVAL_68;
  wire  _EVAL_116;
  wire  _EVAL_113;
  wire  _EVAL_75;
  wire  _EVAL_183;
  wire  _EVAL_94;
  wire  _EVAL_112;
  wire  _EVAL_55;
  wire  _EVAL_146;
  wire  _EVAL_182;
  wire  _EVAL_185;
  wire  _EVAL_188;
  wire  _EVAL_195;
  wire  _EVAL_32;
  wire  _EVAL_95;
  wire [1:0] _EVAL_126;
  wire  _EVAL_103;
  wire  _EVAL_102;
  wire  _EVAL_130;
  wire  _EVAL_51;
  wire  _EVAL_171;
  wire  _EVAL_21;
  wire  _EVAL_76;
  wire  _EVAL_23;
  wire  _EVAL_107;
  wire [8:0] _EVAL_109;
  wire [8:0] _EVAL_176;
  wire  _EVAL_93;
  wire  _EVAL_62;
  wire  _EVAL_186;
  wire  _EVAL_155;
  wire  _EVAL_50;
  wire [8:0] _EVAL_10;
  wire [8:0] _EVAL_147;
  wire [22:0] _EVAL_114;
  wire [8:0] _EVAL_135;
  wire [8:0] _EVAL_134;
  wire  _EVAL_142;
  wire [8:0] _EVAL_124;
  wire [8:0] _EVAL_18;
  wire [8:0] _EVAL_28;
  wire [8:0] _EVAL_165;
  wire [8:0] _EVAL_15;
  wire [8:0] _EVAL_150;
  wire  _EVAL_200;
  wire  _EVAL_175;
  wire [8:0] _EVAL_77;
  wire [8:0] _EVAL_149;
  wire [8:0] _EVAL_187;
  wire [8:0] _EVAL_19;
  wire [8:0] _EVAL_136;
  wire [8:0] _EVAL_46;
  wire [8:0] _EVAL_151;
  wire [8:0] _EVAL_159;
  wire  _EVAL_78;
  wire [9:0] _EVAL_108;
  wire [2:0] _EVAL_199;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [22:0] _EVAL_145;
  wire [22:0] _EVAL_35;
  wire [22:0] _EVAL_99;
  wire [22:0] _EVAL_24;
  wire [22:0] _EVAL_192;
  wire [22:0] _EVAL_153;
  wire  _EVAL_170;
  wire  _EVAL_144;
  wire [1:0] _EVAL_101;
  assign _EVAL_111 = _EVAL_6[26];
  assign _EVAL_131 = _EVAL[8:0];
  assign _EVAL_148 = ~ _EVAL_131;
  assign _EVAL_110 = _EVAL_148[8];
  assign _EVAL_122 = _EVAL_148[7:0];
  assign _EVAL_33 = _EVAL_122[7];
  assign _EVAL_167 = _EVAL_122[6:0];
  assign _EVAL_100 = _EVAL_167[6];
  assign _EVAL_128 = _EVAL_167[5:0];
  assign _EVAL_45 = $signed(-65'sh10000000000000000) >>> _EVAL_128;
  assign _EVAL_27 = _EVAL_45[63:42];
  assign _EVAL_162 = _EVAL_27[15:0];
  assign _EVAL_120 = _EVAL_162[15:8];
  assign _EVAL_207 = {{8'd0}, _EVAL_120};
  assign _EVAL_105 = _EVAL_162[7:0];
  assign _EVAL_133 = {_EVAL_105, 8'h0};
  assign _EVAL_12 = _EVAL_133 & 16'hff00;
  assign _EVAL_14 = _EVAL_207 | _EVAL_12;
  assign _EVAL_141 = _EVAL_14[15:4];
  assign _EVAL_53 = {{4'd0}, _EVAL_141};
  assign _EVAL_177 = _EVAL_53 & 16'hf0f;
  assign _EVAL_178 = _EVAL_14[11:0];
  assign _EVAL_37 = {_EVAL_178, 4'h0};
  assign _EVAL_49 = _EVAL_37 & 16'hf0f0;
  assign _EVAL_140 = _EVAL_177 | _EVAL_49;
  assign _EVAL_58 = _EVAL_140[15:2];
  assign _EVAL_156 = {{2'd0}, _EVAL_58};
  assign _EVAL_164 = _EVAL_156 & 16'h3333;
  assign _EVAL_41 = _EVAL_140[13:0];
  assign _EVAL_174 = {_EVAL_41, 2'h0};
  assign _EVAL_59 = _EVAL_174 & 16'hcccc;
  assign _EVAL_69 = _EVAL_164 | _EVAL_59;
  assign _EVAL_206 = _EVAL_69[15:1];
  assign _EVAL_79 = {{1'd0}, _EVAL_206};
  assign _EVAL_127 = _EVAL_79 & 16'h5555;
  assign _EVAL_86 = _EVAL_69[14:0];
  assign _EVAL_106 = {_EVAL_86, 1'h0};
  assign _EVAL_60 = _EVAL_106 & 16'haaaa;
  assign _EVAL_47 = _EVAL_127 | _EVAL_60;
  assign _EVAL_194 = _EVAL_27[21:16];
  assign _EVAL_43 = _EVAL_194[3:0];
  assign _EVAL_143 = _EVAL_43[1:0];
  assign _EVAL_138 = _EVAL_143[0];
  assign _EVAL_152 = _EVAL_143[1];
  assign _EVAL_129 = _EVAL_43[3:2];
  assign _EVAL_201 = _EVAL_129[0];
  assign _EVAL_65 = _EVAL_129[1];
  assign _EVAL_67 = _EVAL_194[5:4];
  assign _EVAL_17 = _EVAL_67[0];
  assign _EVAL_48 = _EVAL_67[1];
  assign _EVAL_132 = {_EVAL_47,_EVAL_138,_EVAL_152,_EVAL_201,_EVAL_65,_EVAL_17,_EVAL_48};
  assign _EVAL_57 = ~ _EVAL_132;
  assign _EVAL_118 = _EVAL_100 ? 22'h0 : _EVAL_57;
  assign _EVAL_30 = ~ _EVAL_118;
  assign _EVAL_189 = {_EVAL_30,3'h7};
  assign _EVAL_180 = _EVAL_45[2:0];
  assign _EVAL_179 = _EVAL_180[1:0];
  assign _EVAL_96 = _EVAL_179[0];
  assign _EVAL_63 = _EVAL_179[1];
  assign _EVAL_181 = _EVAL_180[2];
  assign _EVAL_169 = {_EVAL_96,_EVAL_63,_EVAL_181};
  assign _EVAL_104 = _EVAL_100 ? _EVAL_169 : 3'h0;
  assign _EVAL_154 = _EVAL_33 ? _EVAL_189 : {{22'd0}, _EVAL_104};
  assign _EVAL_11 = _EVAL_110 ? _EVAL_154 : 25'h0;
  assign _EVAL_190 = {{24'd0}, _EVAL_111};
  assign _EVAL_40 = _EVAL_11 | _EVAL_190;
  assign _EVAL_16 = {_EVAL_40,2'h3};
  assign _EVAL_42 = _EVAL_16[3];
  assign _EVAL_117 = _EVAL_16[2];
  assign _EVAL_44 = _EVAL_111 ? _EVAL_42 : _EVAL_117;
  assign _EVAL_72 = _EVAL_5 | _EVAL_9;
  assign _EVAL_83 = _EVAL_0 | _EVAL_8;
  assign _EVAL_66 = _EVAL_83 == 1'h0;
  assign _EVAL_184 = _EVAL_72 == 1'h0;
  assign _EVAL_87 = _EVAL_66 & _EVAL_184;
  assign _EVAL_193 = _EVAL_3 == 1'h0;
  assign _EVAL_25 = _EVAL_87 & _EVAL_193;
  assign _EVAL_39 = _EVAL_7 == 3'h0;
  assign _EVAL_191 = _EVAL_7 == 3'h4;
  assign _EVAL_20 = _EVAL_39 | _EVAL_191;
  assign _EVAL_52 = _EVAL_16[26:1];
  assign _EVAL_205 = {1'h0,_EVAL_52};
  assign _EVAL_26 = ~ _EVAL_205;
  assign _EVAL_89 = _EVAL_26 & _EVAL_16;
  assign _EVAL_204 = _EVAL_6 & _EVAL_89;
  assign _EVAL_168 = _EVAL_204 != 27'h0;
  assign _EVAL_70 = _EVAL_20 & _EVAL_168;
  assign _EVAL_91 = _EVAL_7 == 3'h2;
  assign _EVAL_123 = _EVAL_91 & _EVAL_4;
  assign _EVAL_74 = _EVAL_7 == 3'h3;
  assign _EVAL_173 = _EVAL_4 == 1'h0;
  assign _EVAL_98 = _EVAL_74 & _EVAL_173;
  assign _EVAL_81 = _EVAL_123 | _EVAL_98;
  assign _EVAL_125 = _EVAL_6 & _EVAL_205;
  assign _EVAL_88 = _EVAL_125 != 27'h0;
  assign _EVAL_172 = _EVAL_168 | _EVAL_88;
  assign _EVAL_90 = _EVAL_81 & _EVAL_172;
  assign _EVAL_197 = _EVAL_70 | _EVAL_90;
  assign _EVAL_166 = _EVAL_6 | _EVAL_16;
  assign _EVAL_71 = _EVAL_166[26:2];
  assign _EVAL_61 = _EVAL_71 + 25'h1;
  assign _EVAL_163 = _EVAL_39 & _EVAL_168;
  assign _EVAL_115 = _EVAL_88 == 1'h0;
  assign _EVAL_56 = _EVAL_163 & _EVAL_115;
  assign _EVAL_85 = _EVAL_56 ? _EVAL_52 : 26'h0;
  assign _EVAL_97 = ~ _EVAL_85;
  assign _EVAL_198 = _EVAL_61 & _EVAL_97;
  assign _EVAL_73 = ~ _EVAL_16;
  assign _EVAL_203 = _EVAL_6 & _EVAL_73;
  assign _EVAL_92 = _EVAL_203[26:2];
  assign _EVAL_158 = {{1'd0}, _EVAL_92};
  assign _EVAL_196 = _EVAL_7 == 3'h6;
  assign _EVAL_54 = _EVAL_196 & _EVAL_172;
  assign _EVAL_34 = _EVAL_89[26:1];
  assign _EVAL_13 = _EVAL_54 ? _EVAL_34 : 26'h0;
  assign _EVAL_137 = _EVAL_158 | _EVAL_13;
  assign _EVAL_84 = _EVAL_197 ? _EVAL_198 : _EVAL_137;
  assign _EVAL_80 = _EVAL_84[25:24];
  assign _EVAL_121 = {1'b0,$signed(_EVAL_80)};
  assign _EVAL_36 = {{7{_EVAL_121[2]}},_EVAL_121};
  assign _EVAL_82 = $signed(_EVAL) + $signed(_EVAL_36);
  assign _EVAL_157 = _EVAL_82[10:7];
  assign _EVAL_22 = $signed(_EVAL_157) >= $signed(4'sh3);
  assign _EVAL_119 = _EVAL_25 & _EVAL_22;
  assign _EVAL_202 = _EVAL_20 | _EVAL_81;
  assign _EVAL_139 = _EVAL_119 & _EVAL_202;
  assign _EVAL_31 = _EVAL_72 | _EVAL_139;
  assign _EVAL_38 = _EVAL_31 ? 9'h180 : 9'h0;
  assign _EVAL_29 = _EVAL[9:8];
  assign _EVAL_64 = $signed(_EVAL_29) <= $signed(2'sh0);
  assign _EVAL_68 = _EVAL_172 & _EVAL_64;
  assign _EVAL_116 = _EVAL_68 & _EVAL_44;
  assign _EVAL_113 = _EVAL_16[4];
  assign _EVAL_75 = _EVAL_111 ? _EVAL_113 : _EVAL_42;
  assign _EVAL_183 = _EVAL_75 == 1'h0;
  assign _EVAL_94 = _EVAL_84[25];
  assign _EVAL_112 = _EVAL_84[24];
  assign _EVAL_55 = _EVAL_111 ? _EVAL_94 : _EVAL_112;
  assign _EVAL_146 = _EVAL_183 & _EVAL_55;
  assign _EVAL_182 = _EVAL_146 & _EVAL_168;
  assign _EVAL_185 = _EVAL_6[2];
  assign _EVAL_188 = _EVAL_6[1];
  assign _EVAL_195 = _EVAL_111 ? _EVAL_185 : _EVAL_188;
  assign _EVAL_32 = _EVAL_20 & _EVAL_195;
  assign _EVAL_95 = _EVAL_111 & _EVAL_185;
  assign _EVAL_126 = _EVAL_6[1:0];
  assign _EVAL_103 = _EVAL_126 != 2'h0;
  assign _EVAL_102 = _EVAL_95 | _EVAL_103;
  assign _EVAL_130 = _EVAL_81 & _EVAL_102;
  assign _EVAL_51 = _EVAL_32 | _EVAL_130;
  assign _EVAL_171 = _EVAL_182 & _EVAL_51;
  assign _EVAL_21 = _EVAL_171 == 1'h0;
  assign _EVAL_76 = _EVAL_116 & _EVAL_21;
  assign _EVAL_23 = _EVAL_202 == 1'h0;
  assign _EVAL_107 = _EVAL_119 & _EVAL_23;
  assign _EVAL_109 = _EVAL_107 ? 9'h17f : 9'h0;
  assign _EVAL_176 = _EVAL_107 ? 9'h80 : 9'h0;
  assign _EVAL_93 = _EVAL_83 | _EVAL_3;
  assign _EVAL_62 = $signed(_EVAL_82) < $signed(11'sh6b);
  assign _EVAL_186 = _EVAL_25 & _EVAL_62;
  assign _EVAL_155 = _EVAL_81 | _EVAL_196;
  assign _EVAL_50 = _EVAL_186 & _EVAL_155;
  assign _EVAL_10 = _EVAL_50 ? 9'h194 : 9'h0;
  assign _EVAL_147 = ~ _EVAL_10;
  assign _EVAL_114 = _EVAL_84[22:0];
  assign _EVAL_135 = _EVAL_50 ? 9'h6b : 9'h0;
  assign _EVAL_134 = _EVAL_82[8:0];
  assign _EVAL_142 = _EVAL_3 | _EVAL_62;
  assign _EVAL_124 = _EVAL_142 ? 9'h1c0 : 9'h0;
  assign _EVAL_18 = ~ _EVAL_124;
  assign _EVAL_28 = _EVAL_134 & _EVAL_18;
  assign _EVAL_165 = _EVAL_28 & _EVAL_147;
  assign _EVAL_15 = ~ _EVAL_176;
  assign _EVAL_150 = _EVAL_165 & _EVAL_15;
  assign _EVAL_200 = _EVAL_62 | _EVAL_172;
  assign _EVAL_175 = _EVAL_25 & _EVAL_200;
  assign _EVAL_77 = _EVAL_31 ? 9'h40 : 9'h0;
  assign _EVAL_149 = ~ _EVAL_77;
  assign _EVAL_187 = _EVAL_150 & _EVAL_149;
  assign _EVAL_19 = _EVAL_187 | _EVAL_135;
  assign _EVAL_136 = _EVAL_19 | _EVAL_109;
  assign _EVAL_46 = _EVAL_136 | _EVAL_38;
  assign _EVAL_151 = _EVAL_83 ? 9'h1c0 : 9'h0;
  assign _EVAL_159 = _EVAL_46 | _EVAL_151;
  assign _EVAL_78 = _EVAL_83 ? 1'h0 : _EVAL_4;
  assign _EVAL_108 = {_EVAL_78,_EVAL_159};
  assign _EVAL_199 = {_EVAL_0,_EVAL_5,_EVAL_119};
  assign _EVAL_160 = _EVAL_119 | _EVAL_175;
  assign _EVAL_161 = _EVAL_93 | _EVAL_62;
  assign _EVAL_145 = _EVAL_83 ? 23'h400000 : 23'h0;
  assign _EVAL_35 = _EVAL_84[23:1];
  assign _EVAL_99 = _EVAL_111 ? _EVAL_35 : _EVAL_114;
  assign _EVAL_24 = _EVAL_161 ? _EVAL_145 : _EVAL_99;
  assign _EVAL_192 = _EVAL_107 ? 23'h7fffff : 23'h0;
  assign _EVAL_153 = _EVAL_24 | _EVAL_192;
  assign _EVAL_170 = _EVAL_62 | _EVAL_76;
  assign _EVAL_144 = _EVAL_25 & _EVAL_170;
  assign _EVAL_101 = {_EVAL_144,_EVAL_160};
  assign _EVAL_2 = {_EVAL_108,_EVAL_153};
  assign _EVAL_1 = {_EVAL_199,_EVAL_101};
endmodule
