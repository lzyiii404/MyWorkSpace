//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_308(
  output         _EVAL,
  output [4:0]   _EVAL_0,
  input          _EVAL_1,
  output [127:0] _EVAL_2,
  output         _EVAL_3,
  output         _EVAL_4,
  output         _EVAL_5,
  input          _EVAL_6,
  output         _EVAL_7,
  input  [8:0]   _EVAL_8,
  input  [1:0]   _EVAL_9,
  output [2:0]   _EVAL_10,
  output         _EVAL_11,
  input          _EVAL_12,
  input          _EVAL_13,
  output         _EVAL_14,
  output [1:0]   _EVAL_15,
  output         _EVAL_16,
  output         _EVAL_17,
  output         _EVAL_18,
  input          _EVAL_19,
  output         _EVAL_20,
  output         _EVAL_21,
  output         _EVAL_22,
  output         _EVAL_23,
  input          _EVAL_24,
  input  [1:0]   _EVAL_25,
  input          _EVAL_26,
  input  [31:0]  _EVAL_27,
  output         _EVAL_28,
  input          _EVAL_29,
  output [1:0]   _EVAL_30,
  input          _EVAL_31,
  input          _EVAL_32,
  input  [63:0]  _EVAL_33,
  output         _EVAL_34,
  output         _EVAL_35,
  output         _EVAL_36,
  output         _EVAL_37,
  output [4:0]   _EVAL_38,
  input          _EVAL_39,
  output         _EVAL_40,
  output [4:0]   _EVAL_41,
  input          _EVAL_42,
  input  [2:0]   _EVAL_43,
  input  [31:0]  _EVAL_44,
  output         _EVAL_45,
  output         _EVAL_46,
  input          _EVAL_47,
  input          _EVAL_48,
  input          _EVAL_49,
  output         _EVAL_50,
  input          _EVAL_51,
  input          _EVAL_52,
  input          _EVAL_53,
  output         _EVAL_54,
  output         _EVAL_55,
  input  [1:0]   _EVAL_56,
  input          _EVAL_57,
  output         _EVAL_58,
  output [8:0]   _EVAL_59,
  input          _EVAL_60,
  input          _EVAL_61,
  output         _EVAL_62,
  output [4:0]   _EVAL_63,
  input          _EVAL_64,
  output         _EVAL_65,
  input          _EVAL_66,
  input          _EVAL_67,
  output         _EVAL_68,
  output         _EVAL_69,
  output         _EVAL_70,
  output         _EVAL_71,
  input          _EVAL_72,
  input          _EVAL_73,
  output         _EVAL_74,
  input          _EVAL_75,
  output         _EVAL_76,
  input          _EVAL_77,
  output         _EVAL_78,
  input          _EVAL_79,
  output [14:0]  _EVAL_80,
  output         _EVAL_81,
  output [2:0]   _EVAL_82,
  output         _EVAL_83,
  output         _EVAL_84,
  output         _EVAL_85,
  output         _EVAL_86,
  output         _EVAL_87,
  output [6:0]   _EVAL_88,
  input          _EVAL_89,
  input          _EVAL_90,
  input          _EVAL_91,
  input  [1:0]   _EVAL_92,
  output [14:0]  _EVAL_93,
  output [8:0]   _EVAL_94,
  input          _EVAL_95,
  output [4:0]   _EVAL_96,
  output         _EVAL_97,
  input  [1:0]   _EVAL_98,
  output         _EVAL_99,
  input  [2:0]   _EVAL_100,
  output         _EVAL_101,
  input  [31:0]  _EVAL_102,
  output         _EVAL_103,
  input          _EVAL_104,
  output         _EVAL_105,
  output         _EVAL_106,
  input          _EVAL_107,
  input  [14:0]  _EVAL_108,
  output         _EVAL_109,
  input          _EVAL_110,
  output [4:0]   _EVAL_111,
  output         _EVAL_112,
  output         _EVAL_113,
  output         _EVAL_114,
  output         _EVAL_115,
  output         _EVAL_116,
  input  [127:0] _EVAL_117,
  output         _EVAL_118,
  output [31:0]  _EVAL_119,
  output         _EVAL_120,
  output         _EVAL_121,
  input          _EVAL_122,
  output [4:0]   _EVAL_123,
  output         _EVAL_124,
  output [127:0] _EVAL_125,
  input  [31:0]  _EVAL_126,
  input          _EVAL_127,
  output         _EVAL_128,
  output         _EVAL_129,
  output [31:0]  _EVAL_130,
  output [2:0]   _EVAL_131,
  input          _EVAL_132,
  output         _EVAL_133,
  output         _EVAL_134,
  output         _EVAL_135,
  input  [31:0]  _EVAL_136,
  output [2:0]   _EVAL_137,
  output         _EVAL_138,
  input  [1:0]   _EVAL_139,
  output         _EVAL_140,
  output         _EVAL_141,
  input          _EVAL_142,
  input          _EVAL_143,
  input          _EVAL_144,
  input          _EVAL_145,
  output [2:0]   _EVAL_146,
  input          _EVAL_147,
  output [2:0]   _EVAL_148,
  output         _EVAL_149,
  output [6:0]   _EVAL_150,
  output         _EVAL_151,
  input  [2:0]   _EVAL_152,
  output         _EVAL_153,
  input          _EVAL_154,
  output         _EVAL_155,
  input          _EVAL_156,
  output         _EVAL_157,
  output [4:0]   _EVAL_158,
  output         _EVAL_159
);
  reg  _EVAL_372;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_701;
  reg [31:0] _RAND_1;
  reg  _EVAL_717;
  reg [31:0] _RAND_2;
  reg  _EVAL_718;
  reg [31:0] _RAND_3;
  reg  _EVAL_788;
  reg [31:0] _RAND_4;
  reg  _EVAL_815;
  reg [31:0] _RAND_5;
  reg  _EVAL_1171;
  reg [31:0] _RAND_6;
  reg  _EVAL_1563;
  reg [31:0] _RAND_7;
  reg  _EVAL_1726;
  reg [31:0] _RAND_8;
  reg  _EVAL_2135;
  reg [31:0] _RAND_9;
  reg  _EVAL_2202;
  reg [31:0] _RAND_10;
  reg  _EVAL_2241;
  reg [31:0] _RAND_11;
  reg [8:0] _EVAL_2281;
  reg [31:0] _RAND_12;
  reg [127:0] _EVAL_2740;
  reg [127:0] _RAND_13;
  reg [1:0] _EVAL_3403;
  reg [31:0] _RAND_14;
  reg  _EVAL_3526;
  reg [31:0] _RAND_15;
  reg  _EVAL_3907;
  reg [31:0] _RAND_16;
  reg  _EVAL_4123;
  reg [31:0] _RAND_17;
  reg  _EVAL_4261;
  reg [31:0] _RAND_18;
  reg [1:0] _EVAL_4273;
  reg [31:0] _RAND_19;
  reg [31:0] _EVAL_4664;
  reg [31:0] _RAND_20;
  reg  _EVAL_4774;
  reg [31:0] _RAND_21;
  reg  _EVAL_4793;
  reg [31:0] _RAND_22;
  reg [15:0] _EVAL_5094;
  reg [31:0] _RAND_23;
  reg  _EVAL_5165;
  reg [31:0] _RAND_24;
  reg [2:0] _EVAL_5225;
  reg [31:0] _RAND_25;
  reg  _EVAL_5335;
  reg [31:0] _RAND_26;
  reg  _EVAL_5437;
  reg [31:0] _RAND_27;
  reg  _EVAL_5648;
  reg [31:0] _RAND_28;
  reg  _EVAL_5701;
  reg [31:0] _RAND_29;
  reg  _EVAL_5994;
  reg [31:0] _RAND_30;
  reg [14:0] _EVAL_6019;
  reg [31:0] _RAND_31;
  wire [15:0] _EVAL_2666;
  wire [15:0] _EVAL_4292;
  wire [15:0] _EVAL_5159;
  wire [47:0] _EVAL_3455;
  wire [2:0] _EVAL_4071;
  wire  _EVAL_4669;
  wire  _EVAL_241;
  wire [2:0] _EVAL_4901;
  wire  _EVAL_2996;
  wire [6:0] _EVAL_1346;
  wire [1:0] _EVAL_1939;
  wire [2:0] _EVAL_3926;
  wire [2:0] _EVAL_4872;
  wire [4:0] _EVAL_5992;
  wire [26:0] _EVAL_1643;
  wire  _EVAL_2288;
  wire [26:0] _EVAL_4563;
  wire  _EVAL_453;
  wire [1:0] _EVAL_5278;
  wire [7:0] _EVAL_5928;
  wire [2:0] _EVAL_2821;
  wire [4:0] _EVAL_1749;
  wire [27:0] _EVAL_3859;
  wire  _EVAL_936;
  wire [26:0] _EVAL_3053;
  wire  _EVAL_1674;
  wire [26:0] _EVAL_3821;
  wire  _EVAL_597;
  wire [26:0] _EVAL_2991;
  wire  _EVAL_5755;
  wire [27:0] _EVAL_2246;
  wire [3:0] _EVAL_4532;
  wire [1:0] _EVAL_5956;
  wire [29:0] _EVAL_1848;
  wire [29:0] _EVAL_812;
  wire [29:0] _EVAL_173;
  wire [29:0] _EVAL_2725;
  wire [29:0] _EVAL_2541;
  wire [29:0] _EVAL_4645;
  wire [29:0] _EVAL_3736;
  wire [29:0] _EVAL_3595;
  wire [31:0] _EVAL_2164;
  wire [31:0] _EVAL_1690;
  wire  _EVAL_4293;
  wire [31:0] _EVAL_5077;
  wire  _EVAL_3471;
  wire  _EVAL_2314;
  wire [31:0] _EVAL_877;
  wire  _EVAL_4098;
  wire  _EVAL_1135;
  wire [31:0] _EVAL_1286;
  wire  _EVAL_4327;
  wire  _EVAL_2655;
  wire [31:0] _EVAL_1215;
  wire  _EVAL_5365;
  wire  _EVAL_2407;
  wire [31:0] _EVAL_5699;
  wire  _EVAL_3701;
  wire  _EVAL_4420;
  wire [31:0] _EVAL_3778;
  wire  _EVAL_1131;
  wire  _EVAL_5931;
  wire [31:0] _EVAL_764;
  wire  _EVAL_3234;
  wire  _EVAL_447;
  wire [31:0] _EVAL_6097;
  wire  _EVAL_4305;
  wire  _EVAL_5238;
  wire [31:0] _EVAL_645;
  wire  _EVAL_836;
  wire  _EVAL_4330;
  wire [31:0] _EVAL_4039;
  wire  _EVAL_367;
  wire  _EVAL_210;
  wire [31:0] _EVAL_3250;
  wire  _EVAL_1116;
  wire  _EVAL_2096;
  wire  _EVAL_4777;
  wire  _EVAL_2982;
  wire [31:0] _EVAL_3891;
  wire  _EVAL_687;
  wire  _EVAL_1570;
  wire  _EVAL_6053;
  wire  _EVAL_1771;
  wire [31:0] _EVAL_5477;
  wire  _EVAL_3235;
  wire  _EVAL_3436;
  wire [31:0] _EVAL_2614;
  wire  _EVAL_4022;
  wire  _EVAL_4755;
  wire [31:0] _EVAL_3440;
  wire  _EVAL_3096;
  wire  _EVAL_2790;
  wire [31:0] _EVAL_2778;
  wire  _EVAL_2477;
  wire  _EVAL_4155;
  wire [31:0] _EVAL_171;
  wire  _EVAL_262;
  wire  _EVAL_4260;
  wire [31:0] _EVAL_2457;
  wire  _EVAL_3049;
  wire  _EVAL_3000;
  wire [31:0] _EVAL_5743;
  wire  _EVAL_3229;
  wire  _EVAL_2362;
  wire  _EVAL_2629;
  wire  _EVAL_2143;
  wire [3:0] _EVAL_5731;
  wire [1:0] _EVAL_4188;
  wire [3:0] _EVAL_3997;
  wire [15:0] _EVAL_3588;
  wire [79:0] _EVAL_654;
  wire [31:0] _EVAL_4702;
  wire [31:0] _EVAL_4125;
  wire [1:0] _EVAL_2935;
  wire [10:0] _EVAL_2290;
  wire  _EVAL_3023;
  wire [31:0] _EVAL_2277;
  wire [2:0] _EVAL_808;
  wire  _EVAL_1088;
  wire [3:0] _EVAL_3841;
  wire [7:0] _EVAL_738;
  wire [2:0] _EVAL_3877;
  wire [4:0] _EVAL_1321;
  wire [4:0] _EVAL_694;
  wire [27:0] _EVAL_3043;
  wire  _EVAL_537;
  wire [27:0] _EVAL_5721;
  wire  _EVAL_1378;
  wire [2:0] _EVAL_4771;
  wire [2:0] _EVAL_2483;
  wire [8:0] _EVAL_5892;
  wire [3:0] _EVAL_4114;
  wire [4:0] _EVAL_4538;
  wire [28:0] _EVAL_3320;
  wire  _EVAL_4440;
  wire  _EVAL_3082;
  wire  _EVAL_2173;
  wire [4:0] _EVAL_4094;
  wire [24:0] _EVAL_759;
  wire  _EVAL_1360;
  wire [24:0] _EVAL_4100;
  wire [24:0] _EVAL_2188;
  wire [17:0] _EVAL_3216;
  wire [24:0] _EVAL_938;
  wire [24:0] _EVAL_448;
  wire [24:0] _EVAL_1277;
  wire [24:0] _EVAL_4791;
  wire [24:0] _EVAL_1610;
  wire [24:0] _EVAL_947;
  wire [24:0] _EVAL_1568;
  wire  _EVAL_761;
  wire [1:0] _EVAL_4347;
  wire [2:0] _EVAL_2114;
  wire [27:0] _EVAL_3139;
  wire  _EVAL_5989;
  wire [27:0] _EVAL_3138;
  wire  _EVAL_3016;
  wire [2:0] _EVAL_2231;
  wire [1:0] _EVAL_4575;
  wire [28:0] _EVAL_2397;
  wire [25:0] _EVAL_1481;
  wire [28:0] _EVAL_2014;
  wire [28:0] _EVAL_2350;
  wire [28:0] _EVAL_3048;
  wire [28:0] _EVAL_583;
  wire [28:0] _EVAL_327;
  wire [28:0] _EVAL_2482;
  wire [28:0] _EVAL_4396;
  wire [31:0] _EVAL_3078;
  wire [31:0] _EVAL_4897;
  wire  _EVAL_4008;
  wire [31:0] _EVAL_2032;
  wire  _EVAL_1754;
  wire  _EVAL_4659;
  wire [31:0] _EVAL_4518;
  wire  _EVAL_2788;
  wire  _EVAL_1008;
  wire [31:0] _EVAL_2628;
  wire  _EVAL_1860;
  wire  _EVAL_4503;
  wire [31:0] _EVAL_4163;
  wire  _EVAL_5214;
  wire  _EVAL_5228;
  wire [31:0] _EVAL_4951;
  wire  _EVAL_4400;
  wire  _EVAL_4544;
  wire [31:0] _EVAL_2517;
  wire  _EVAL_1021;
  wire  _EVAL_2838;
  wire [31:0] _EVAL_5223;
  wire  _EVAL_5145;
  wire  _EVAL_4103;
  wire [31:0] _EVAL_4594;
  wire  _EVAL_5654;
  wire  _EVAL_3674;
  wire [31:0] _EVAL_2087;
  wire  _EVAL_2442;
  wire  _EVAL_1507;
  wire [31:0] _EVAL_4591;
  wire  _EVAL_5913;
  wire  _EVAL_4603;
  wire [31:0] _EVAL_5143;
  wire  _EVAL_1641;
  wire  _EVAL_3239;
  wire [31:0] _EVAL_4268;
  wire [2:0] _EVAL_771;
  wire  _EVAL_5623;
  wire [1:0] _EVAL_263;
  wire [3:0] _EVAL_3602;
  wire [7:0] _EVAL_3330;
  wire [2:0] _EVAL_762;
  wire [4:0] _EVAL_3553;
  wire [4:0] _EVAL_871;
  wire [27:0] _EVAL_2908;
  wire  _EVAL_5053;
  wire [27:0] _EVAL_5618;
  wire  _EVAL_2321;
  wire [2:0] _EVAL_3871;
  wire [2:0] _EVAL_2808;
  wire [8:0] _EVAL_1025;
  wire [3:0] _EVAL_2831;
  wire [4:0] _EVAL_2613;
  wire [28:0] _EVAL_1479;
  wire  _EVAL_3712;
  wire  _EVAL_5439;
  wire  _EVAL_1657;
  wire [4:0] _EVAL_932;
  wire [24:0] _EVAL_2026;
  wire  _EVAL_3685;
  wire [24:0] _EVAL_4034;
  wire [24:0] _EVAL_3296;
  wire [17:0] _EVAL_1863;
  wire [24:0] _EVAL_4578;
  wire [24:0] _EVAL_4876;
  wire [24:0] _EVAL_3519;
  wire [24:0] _EVAL_4673;
  wire [24:0] _EVAL_5005;
  wire [24:0] _EVAL_282;
  wire [24:0] _EVAL_4515;
  wire  _EVAL_1743;
  wire [1:0] _EVAL_5411;
  wire [2:0] _EVAL_626;
  wire [27:0] _EVAL_2036;
  wire  _EVAL_4038;
  wire [27:0] _EVAL_1073;
  wire  _EVAL_5573;
  wire [2:0] _EVAL_763;
  wire [1:0] _EVAL_167;
  wire [28:0] _EVAL_3823;
  wire [25:0] _EVAL_341;
  wire [28:0] _EVAL_180;
  wire [28:0] _EVAL_1110;
  wire [28:0] _EVAL_4831;
  wire [28:0] _EVAL_1996;
  wire [28:0] _EVAL_227;
  wire [28:0] _EVAL_3987;
  wire [28:0] _EVAL_2410;
  wire [31:0] _EVAL_3006;
  wire [31:0] _EVAL_2462;
  wire  _EVAL_5041;
  wire [31:0] _EVAL_3952;
  wire  _EVAL_4113;
  wire  _EVAL_4830;
  wire [31:0] _EVAL_1111;
  wire  _EVAL_3150;
  wire  _EVAL_3757;
  wire [31:0] _EVAL_1137;
  wire  _EVAL_470;
  wire  _EVAL_5979;
  wire [63:0] _EVAL_5386;
  wire [2:0] _EVAL_1136;
  wire  _EVAL_4999;
  wire  _EVAL_287;
  wire [2:0] _EVAL_688;
  wire  _EVAL_2964;
  wire [6:0] _EVAL_3443;
  wire [1:0] _EVAL_746;
  wire [2:0] _EVAL_1418;
  wire [2:0] _EVAL_5546;
  wire [4:0] _EVAL_1050;
  wire [26:0] _EVAL_2013;
  wire  _EVAL_4185;
  wire [26:0] _EVAL_4065;
  wire  _EVAL_3493;
  wire [1:0] _EVAL_5289;
  wire [7:0] _EVAL_3643;
  wire [2:0] _EVAL_3861;
  wire [4:0] _EVAL_5112;
  wire [27:0] _EVAL_5044;
  wire  _EVAL_3261;
  wire [26:0] _EVAL_343;
  wire  _EVAL_268;
  wire [26:0] _EVAL_4834;
  wire  _EVAL_179;
  wire [26:0] _EVAL_5270;
  wire  _EVAL_2175;
  wire [27:0] _EVAL_3947;
  wire [3:0] _EVAL_4465;
  wire [1:0] _EVAL_3341;
  wire [29:0] _EVAL_2263;
  wire [29:0] _EVAL_3834;
  wire [29:0] _EVAL_997;
  wire [29:0] _EVAL_1859;
  wire [29:0] _EVAL_5281;
  wire [29:0] _EVAL_1799;
  wire [29:0] _EVAL_2373;
  wire [29:0] _EVAL_1455;
  wire [31:0] _EVAL_386;
  wire [31:0] _EVAL_2259;
  wire  _EVAL_2390;
  wire [31:0] _EVAL_1473;
  wire  _EVAL_706;
  wire  _EVAL_983;
  wire [1:0] _EVAL_476;
  wire [3:0] _EVAL_4927;
  wire [7:0] _EVAL_1900;
  wire [2:0] _EVAL_2067;
  wire [4:0] _EVAL_2075;
  wire [4:0] _EVAL_4281;
  wire [27:0] _EVAL_3343;
  wire [27:0] _EVAL_4648;
  wire [8:0] _EVAL_5823;
  wire [3:0] _EVAL_4096;
  wire [4:0] _EVAL_822;
  wire [28:0] _EVAL_6068;
  wire  _EVAL_735;
  wire  _EVAL_1516;
  wire [4:0] _EVAL_3655;
  wire [24:0] _EVAL_3062;
  wire  _EVAL_863;
  wire [24:0] _EVAL_1869;
  wire [24:0] _EVAL_5542;
  wire [17:0] _EVAL_3808;
  wire [24:0] _EVAL_5624;
  wire [24:0] _EVAL_3593;
  wire [24:0] _EVAL_3134;
  wire [24:0] _EVAL_1119;
  wire [24:0] _EVAL_5616;
  wire [24:0] _EVAL_543;
  wire [24:0] _EVAL_2595;
  wire [1:0] _EVAL_2351;
  wire [2:0] _EVAL_5138;
  wire [27:0] _EVAL_569;
  wire [27:0] _EVAL_578;
  wire [28:0] _EVAL_4655;
  wire [25:0] _EVAL_272;
  wire [28:0] _EVAL_5476;
  wire [28:0] _EVAL_1189;
  wire [28:0] _EVAL_3708;
  wire [28:0] _EVAL_3613;
  wire [28:0] _EVAL_785;
  wire [28:0] _EVAL_593;
  wire [28:0] _EVAL_1348;
  wire [31:0] _EVAL_2039;
  wire [31:0] _EVAL_957;
  wire  _EVAL_2132;
  wire [31:0] _EVAL_3434;
  wire  _EVAL_2712;
  wire  _EVAL_5529;
  wire [31:0] _EVAL_5802;
  wire  _EVAL_4128;
  wire  _EVAL_5560;
  wire [31:0] _EVAL_5355;
  wire  _EVAL_3991;
  wire  _EVAL_5696;
  wire [31:0] _EVAL_3844;
  wire  _EVAL_4210;
  wire  _EVAL_5945;
  wire [31:0] _EVAL_2398;
  wire  _EVAL_644;
  wire  _EVAL_4110;
  wire [31:0] _EVAL_5061;
  wire  _EVAL_4386;
  wire  _EVAL_3478;
  wire [31:0] _EVAL_5686;
  wire  _EVAL_6118;
  wire  _EVAL_1707;
  wire [31:0] _EVAL_1164;
  wire  _EVAL_255;
  wire  _EVAL_3880;
  wire [31:0] _EVAL_335;
  wire  _EVAL_2153;
  wire  _EVAL_568;
  wire [31:0] _EVAL_4841;
  wire  _EVAL_6112;
  wire  _EVAL_2897;
  wire [31:0] _EVAL_5329;
  wire  _EVAL_2769;
  wire  _EVAL_2848;
  wire  _EVAL_5113;
  wire  _EVAL_3410;
  wire [31:0] _EVAL_2663;
  wire  _EVAL_5344;
  wire  _EVAL_3795;
  wire  _EVAL_861;
  wire  _EVAL_5070;
  wire [31:0] _EVAL_5078;
  wire  _EVAL_2802;
  wire  _EVAL_5069;
  wire [31:0] _EVAL_3300;
  wire  _EVAL_2197;
  wire  _EVAL_3874;
  wire [31:0] _EVAL_4267;
  wire  _EVAL_4618;
  wire  _EVAL_203;
  wire [31:0] _EVAL_4796;
  wire  _EVAL_2412;
  wire  _EVAL_264;
  wire [31:0] _EVAL_5455;
  wire  _EVAL_801;
  wire  _EVAL_2360;
  wire [31:0] _EVAL_4191;
  wire  _EVAL_5897;
  wire  _EVAL_1134;
  wire [31:0] _EVAL_4944;
  wire  _EVAL_548;
  wire  _EVAL_3574;
  wire  _EVAL_2849;
  wire  _EVAL_892;
  wire [31:0] _EVAL_3840;
  wire  _EVAL_2742;
  wire  _EVAL_1290;
  wire  _EVAL_4399;
  wire  _EVAL_2736;
  wire [31:0] _EVAL_234;
  wire  _EVAL_2598;
  wire  _EVAL_1520;
  wire [31:0] _EVAL_2890;
  wire  _EVAL_4216;
  wire  _EVAL_1398;
  wire [2:0] _EVAL_4535;
  wire  _EVAL_418;
  wire  _EVAL_1583;
  wire [4:0] _EVAL_2657;
  wire [1:0] _EVAL_3105;
  wire  _EVAL_5775;
  wire [1:0] _EVAL_2671;
  wire [1:0] _EVAL_3182;
  wire [12:0] _EVAL_269;
  wire  _EVAL_6027;
  wire [5:0] _EVAL_4693;
  wire [2:0] _EVAL_1375;
  wire [3:0] _EVAL_3642;
  wire  _EVAL_3414;
  wire [31:0] _EVAL_4233;
  wire  _EVAL_5821;
  wire [31:0] _EVAL_4762;
  wire  _EVAL_2644;
  wire [9:0] _EVAL_2268;
  wire  _EVAL_5309;
  wire [1:0] _EVAL_4709;
  wire  _EVAL_5340;
  wire  _EVAL_882;
  wire  _EVAL_3287;
  wire [2:0] _EVAL_3748;
  wire [20:0] _EVAL_3811;
  wire  _EVAL_2989;
  wire [9:0] _EVAL_2920;
  wire  _EVAL_5236;
  wire [7:0] _EVAL_1128;
  wire [31:0] _EVAL_5753;
  wire  _EVAL_4202;
  wire  _EVAL_5825;
  wire [2:0] _EVAL_5741;
  wire [2:0] _EVAL_1612;
  wire  _EVAL_5920;
  wire  _EVAL_4348;
  wire  _EVAL_3827;
  wire  _EVAL_346;
  wire  _EVAL_2219;
  wire  _EVAL_2608;
  wire  _EVAL_1784;
  wire [2:0] _EVAL_1778;
  wire [2:0] _EVAL_5864;
  wire [2:0] _EVAL_4324;
  wire [2:0] _EVAL_937;
  wire [2:0] _EVAL_350;
  wire [2:0] _EVAL_5404;
  wire [2:0] _EVAL_2308;
  wire [6:0] _EVAL_4551;
  wire [24:0] _EVAL_1161;
  wire [30:0] _EVAL_2572;
  wire  _EVAL_3966;
  wire [30:0] _EVAL_1339;
  wire [30:0] _EVAL_620;
  wire  _EVAL_647;
  wire [6:0] _EVAL_2409;
  wire [4:0] _EVAL_4489;
  wire [31:0] _EVAL_2776;
  wire  _EVAL_1181;
  wire [25:0] _EVAL_4695;
  wire [30:0] _EVAL_4933;
  wire [30:0] _EVAL_2664;
  wire [30:0] _EVAL_1112;
  wire [31:0] _EVAL_3909;
  wire [31:0] _EVAL_1839;
  wire  _EVAL_4352;
  wire [4:0] _EVAL_5023;
  wire  _EVAL_3277;
  wire [2:0] _EVAL_2576;
  wire  _EVAL_1329;
  wire [31:0] _EVAL_477;
  wire [14:0] _EVAL_1713;
  wire [31:0] _EVAL_3263;
  wire [19:0] _EVAL_3826;
  wire [31:0] _EVAL_3311;
  wire [31:0] _EVAL_3412;
  wire  _EVAL_1014;
  wire [31:0] _EVAL_1003;
  wire  _EVAL_630;
  wire [31:0] _EVAL_1962;
  wire [31:0] _EVAL_1235;
  wire [31:0] _EVAL_1320;
  wire [31:0] _EVAL_4467;
  wire [31:0] _EVAL_1727;
  wire [31:0] _EVAL_1493;
  wire [31:0] _EVAL_3372;
  wire [31:0] _EVAL_3906;
  wire [31:0] _EVAL_1362;
  wire [31:0] _EVAL_1096;
  wire  _EVAL_5421;
  wire [2:0] _EVAL_2600;
  wire  _EVAL_5872;
  wire  _EVAL_5387;
  wire  _EVAL_5474;
  wire  _EVAL_392;
  wire  _EVAL_4750;
  wire  _EVAL_4809;
  wire  _EVAL_1551;
  wire [2:0] _EVAL_4531;
  wire [2:0] _EVAL_3094;
  wire [2:0] _EVAL_5638;
  wire [2:0] _EVAL_6071;
  wire [2:0] _EVAL_6140;
  wire [2:0] _EVAL_3910;
  wire [2:0] _EVAL_3630;
  wire [6:0] _EVAL_4250;
  wire [24:0] _EVAL_3408;
  wire [4:0] _EVAL_3385;
  wire  _EVAL_218;
  wire [1:0] _EVAL_948;
  wire [1:0] _EVAL_3864;
  wire [12:0] _EVAL_334;
  wire [5:0] _EVAL_5403;
  wire [1:0] _EVAL_4728;
  wire  _EVAL_5952;
  wire  _EVAL_4111;
  wire [4:0] _EVAL_2534;
  wire  _EVAL_3920;
  wire [1:0] _EVAL_3636;
  wire [1:0] _EVAL_5034;
  wire [12:0] _EVAL_502;
  wire  _EVAL_707;
  wire [5:0] _EVAL_876;
  wire [3:0] _EVAL_5766;
  wire  _EVAL_650;
  wire [31:0] _EVAL_5831;
  wire [31:0] _EVAL_2480;
  wire [9:0] _EVAL_2912;
  wire  _EVAL_3183;
  wire [1:0] _EVAL_745;
  wire  _EVAL_2546;
  wire  _EVAL_3106;
  wire [2:0] _EVAL_1759;
  wire [20:0] _EVAL_4715;
  wire  _EVAL_2592;
  wire [9:0] _EVAL_3210;
  wire  _EVAL_2251;
  wire [7:0] _EVAL_1182;
  wire [31:0] _EVAL_5304;
  wire  _EVAL_896;
  wire [2:0] _EVAL_4176;
  wire  _EVAL_4036;
  wire  _EVAL_4845;
  wire  _EVAL_4391;
  wire  _EVAL_5613;
  wire  _EVAL_6020;
  wire  _EVAL_5356;
  wire  _EVAL_2174;
  wire [2:0] _EVAL_2242;
  wire [2:0] _EVAL_3710;
  wire [2:0] _EVAL_5357;
  wire [2:0] _EVAL_3395;
  wire [2:0] _EVAL_2668;
  wire [2:0] _EVAL_2414;
  wire [2:0] _EVAL_1443;
  wire [6:0] _EVAL_3839;
  wire [24:0] _EVAL_1890;
  wire [30:0] _EVAL_3767;
  wire  _EVAL_3470;
  wire [30:0] _EVAL_3378;
  wire [30:0] _EVAL_553;
  wire  _EVAL_4751;
  wire [6:0] _EVAL_1746;
  wire [4:0] _EVAL_2272;
  wire [31:0] _EVAL_3621;
  wire  _EVAL_1824;
  wire [25:0] _EVAL_1970;
  wire [30:0] _EVAL_4916;
  wire [30:0] _EVAL_4429;
  wire [30:0] _EVAL_1678;
  wire [31:0] _EVAL_3761;
  wire [31:0] _EVAL_5015;
  wire [4:0] _EVAL_4374;
  wire  _EVAL_3004;
  wire [2:0] _EVAL_757;
  wire [31:0] _EVAL_3218;
  wire [14:0] _EVAL_2157;
  wire [31:0] _EVAL_5760;
  wire [19:0] _EVAL_5101;
  wire [31:0] _EVAL_837;
  wire [31:0] _EVAL_2568;
  wire [31:0] _EVAL_4390;
  wire [31:0] _EVAL_6047;
  wire [31:0] _EVAL_1954;
  wire [31:0] _EVAL_5009;
  wire [31:0] _EVAL_4338;
  wire [31:0] _EVAL_5428;
  wire [31:0] _EVAL_1416;
  wire [31:0] _EVAL_3129;
  wire [31:0] _EVAL_1160;
  wire [31:0] _EVAL_4743;
  wire [4:0] _EVAL_5510;
  wire [4:0] _EVAL_5456;
  wire [4:0] _EVAL_5074;
  wire [1:0] _EVAL_3200;
  wire [3:0] _EVAL_2739;
  wire [7:0] _EVAL_4277;
  wire [2:0] _EVAL_2466;
  wire [4:0] _EVAL_1636;
  wire [27:0] _EVAL_3405;
  wire [27:0] _EVAL_5944;
  wire [2:0] _EVAL_821;
  wire [8:0] _EVAL_1036;
  wire [3:0] _EVAL_5503;
  wire [4:0] _EVAL_5874;
  wire [28:0] _EVAL_5265;
  wire  _EVAL_2327;
  wire [24:0] _EVAL_1152;
  wire  _EVAL_5924;
  wire [24:0] _EVAL_5441;
  wire [24:0] _EVAL_3534;
  wire [17:0] _EVAL_1041;
  wire [24:0] _EVAL_5904;
  wire [24:0] _EVAL_4112;
  wire [24:0] _EVAL_5615;
  wire [24:0] _EVAL_4812;
  wire [24:0] _EVAL_4730;
  wire [24:0] _EVAL_1536;
  wire [24:0] _EVAL_212;
  wire [1:0] _EVAL_4012;
  wire [2:0] _EVAL_1124;
  wire [27:0] _EVAL_5736;
  wire [27:0] _EVAL_4560;
  wire [28:0] _EVAL_2417;
  wire [25:0] _EVAL_3883;
  wire [28:0] _EVAL_5416;
  wire [28:0] _EVAL_436;
  wire [28:0] _EVAL_2883;
  wire [28:0] _EVAL_5490;
  wire [28:0] _EVAL_5515;
  wire [28:0] _EVAL_1358;
  wire [28:0] _EVAL_1162;
  wire [31:0] _EVAL_1978;
  wire [31:0] _EVAL_4366;
  wire [4:0] _EVAL_1747;
  wire  _EVAL_3677;
  wire [1:0] _EVAL_4680;
  wire [1:0] _EVAL_1092;
  wire [12:0] _EVAL_5804;
  wire  _EVAL_4021;
  wire [5:0] _EVAL_3474;
  wire [3:0] _EVAL_3014;
  wire  _EVAL_2266;
  wire [31:0] _EVAL_2779;
  wire [31:0] _EVAL_3091;
  wire [9:0] _EVAL_4449;
  wire  _EVAL_1100;
  wire [1:0] _EVAL_3102;
  wire  _EVAL_2711;
  wire  _EVAL_2003;
  wire  _EVAL_2525;
  wire [2:0] _EVAL_3498;
  wire [20:0] _EVAL_5465;
  wire  _EVAL_3881;
  wire [9:0] _EVAL_5580;
  wire  _EVAL_3307;
  wire [7:0] _EVAL_5562;
  wire [31:0] _EVAL_5948;
  wire  _EVAL_695;
  wire [2:0] _EVAL_1803;
  wire  _EVAL_4620;
  wire  _EVAL_5493;
  wire  _EVAL_1121;
  wire  _EVAL_5602;
  wire  _EVAL_1210;
  wire  _EVAL_3051;
  wire  _EVAL_2984;
  wire [2:0] _EVAL_4547;
  wire [2:0] _EVAL_2877;
  wire [2:0] _EVAL_3126;
  wire [2:0] _EVAL_6094;
  wire [2:0] _EVAL_3820;
  wire [2:0] _EVAL_3209;
  wire [2:0] _EVAL_690;
  wire [6:0] _EVAL_3616;
  wire [24:0] _EVAL_464;
  wire [30:0] _EVAL_1675;
  wire  _EVAL_243;
  wire [30:0] _EVAL_2022;
  wire [30:0] _EVAL_1807;
  wire  _EVAL_380;
  wire [6:0] _EVAL_3620;
  wire [31:0] _EVAL_2934;
  wire  _EVAL_5259;
  wire [25:0] _EVAL_4447;
  wire [30:0] _EVAL_4905;
  wire [30:0] _EVAL_1056;
  wire [30:0] _EVAL_1194;
  wire [31:0] _EVAL_3148;
  wire [31:0] _EVAL_5991;
  wire  _EVAL_2176;
  wire [2:0] _EVAL_2235;
  wire  _EVAL_3591;
  wire [31:0] _EVAL_5679;
  wire [14:0] _EVAL_2444;
  wire [31:0] _EVAL_1199;
  wire [19:0] _EVAL_5415;
  wire [31:0] _EVAL_4247;
  wire [31:0] _EVAL_3013;
  wire [31:0] _EVAL_6042;
  wire [31:0] _EVAL_4319;
  wire [31:0] _EVAL_5271;
  wire [31:0] _EVAL_3598;
  wire [31:0] _EVAL_3467;
  wire [31:0] _EVAL_4394;
  wire [31:0] _EVAL_1565;
  wire [31:0] _EVAL_4372;
  wire [31:0] _EVAL_3213;
  wire [31:0] _EVAL_4882;
  wire [31:0] _EVAL_411;
  wire  _EVAL_3011;
  wire [31:0] _EVAL_3065;
  wire [6:0] _EVAL_185;
  wire [1:0] _EVAL_3946;
  wire [4:0] _EVAL_6089;
  wire [26:0] _EVAL_3100;
  wire [26:0] _EVAL_5832;
  wire [7:0] _EVAL_2494;
  wire [2:0] _EVAL_6126;
  wire [4:0] _EVAL_522;
  wire [27:0] _EVAL_1065;
  wire [26:0] _EVAL_5132;
  wire [26:0] _EVAL_5338;
  wire [26:0] _EVAL_4120;
  wire [27:0] _EVAL_2122;
  wire [3:0] _EVAL_5636;
  wire [1:0] _EVAL_5612;
  wire [29:0] _EVAL_193;
  wire [29:0] _EVAL_4936;
  wire [29:0] _EVAL_1314;
  wire [29:0] _EVAL_6108;
  wire [29:0] _EVAL_306;
  wire [29:0] _EVAL_2752;
  wire [29:0] _EVAL_1177;
  wire [29:0] _EVAL_3496;
  wire [31:0] _EVAL_5133;
  wire [31:0] _EVAL_5578;
  wire  _EVAL_5723;
  wire  _EVAL_6081;
  wire  _EVAL_2110;
  wire  _EVAL_5564;
  wire  _EVAL_5718;
  wire  _EVAL_2396;
  wire  _EVAL_1206;
  wire [3:0] _EVAL_5440;
  wire [3:0] _EVAL_4264;
  wire  _EVAL_5087;
  wire  _EVAL_3382;
  wire  _EVAL_2532;
  wire  _EVAL_5393;
  wire [1:0] _EVAL_5211;
  wire  _EVAL_4914;
  wire [31:0] _EVAL_1992;
  wire [28:0] _EVAL_1854;
  wire [31:0] _EVAL_5390;
  wire [28:0] _EVAL_3822;
  wire  _EVAL_4204;
  wire  _EVAL_2127;
  wire [2:0] _EVAL_3117;
  wire  _EVAL_5381;
  wire  _EVAL_5561;
  wire  _EVAL_3293;
  wire  _EVAL_379;
  wire  _EVAL_4444;
  wire  _EVAL_481;
  wire  _EVAL_2618;
  wire  _EVAL_439;
  wire  _EVAL_550;
  wire  _EVAL_1763;
  wire  _EVAL_4397;
  wire [3:0] _EVAL_5705;
  wire [3:0] _EVAL_431;
  wire [2:0] _EVAL_1858;
  wire [3:0] _EVAL_3483;
  wire [3:0] _EVAL_4626;
  wire  _EVAL_1689;
  wire  _EVAL_3326;
  wire  _EVAL_1283;
  wire  _EVAL_4867;
  wire  _EVAL_6128;
  wire  _EVAL_4732;
  wire  _EVAL_5875;
  wire  _EVAL_4630;
  wire  _EVAL_3345;
  wire  _EVAL_2781;
  wire  _EVAL_977;
  wire [1:0] _EVAL_3807;
  wire  _EVAL_5680;
  wire [31:0] _EVAL_3560;
  wire [28:0] _EVAL_2209;
  wire  _EVAL_5844;
  wire  _EVAL_5549;
  wire [2:0] _EVAL_5107;
  wire  _EVAL_719;
  wire  _EVAL_5702;
  wire  _EVAL_1914;
  wire  _EVAL_3257;
  wire  _EVAL_2111;
  wire  _EVAL_2107;
  wire  _EVAL_5426;
  wire  _EVAL_1831;
  wire  _EVAL_1408;
  wire  _EVAL_3705;
  wire  _EVAL_5459;
  wire [3:0] _EVAL_3251;
  wire [3:0] _EVAL_5435;
  wire [2:0] _EVAL_5809;
  wire [3:0] _EVAL_4935;
  wire [3:0] _EVAL_920;
  wire  _EVAL_2163;
  wire  _EVAL_4460;
  wire  _EVAL_5220;
  wire  _EVAL_1006;
  wire  _EVAL_2524;
  wire  _EVAL_6001;
  wire  _EVAL_3477;
  wire  _EVAL_4922;
  wire  _EVAL_5668;
  wire  _EVAL_1173;
  wire  _EVAL_4437;
  wire  _EVAL_5698;
  wire  _EVAL_5324;
  wire  _EVAL_2252;
  wire  _EVAL_2993;
  wire  _EVAL_2093;
  wire  _EVAL_3169;
  wire  _EVAL_1383;
  wire  _EVAL_4063;
  wire  _EVAL_2293;
  wire  _EVAL_5967;
  wire  _EVAL_3336;
  wire  _EVAL_169;
  wire  _EVAL_3206;
  wire  _EVAL_3962;
  wire  _EVAL_376;
  wire  _EVAL_165;
  wire  _EVAL_4359;
  wire  _EVAL_4985;
  wire  _EVAL_3923;
  wire  _EVAL_3524;
  wire  _EVAL_209;
  wire  _EVAL_2108;
  wire  _EVAL_2606;
  wire  _EVAL_6086;
  wire  _EVAL_4214;
  wire  _EVAL_3846;
  wire  _EVAL_868;
  wire  _EVAL_2469;
  wire  _EVAL_881;
  wire  _EVAL_2491;
  wire  _EVAL_5443;
  wire  _EVAL_1322;
  wire  _EVAL_4104;
  wire [3:0] _EVAL_1700;
  wire  _EVAL_3143;
  wire  _EVAL_1633;
  wire  _EVAL_2213;
  wire  _EVAL_3402;
  wire  _EVAL_1342;
  wire [1:0] _EVAL_2837;
  wire  _EVAL_1958;
  wire  _EVAL_3242;
  wire [3:0] _EVAL_1670;
  wire  _EVAL_5385;
  wire [31:0] _EVAL_2375;
  wire [31:0] _EVAL_4964;
  wire [9:0] _EVAL_4199;
  wire  _EVAL_2817;
  wire [1:0] _EVAL_1211;
  wire  _EVAL_581;
  wire  _EVAL_4521;
  wire  _EVAL_2557;
  wire [2:0] _EVAL_2977;
  wire [20:0] _EVAL_5750;
  wire  _EVAL_3334;
  wire [9:0] _EVAL_673;
  wire  _EVAL_3399;
  wire [7:0] _EVAL_2699;
  wire [31:0] _EVAL_2011;
  wire  _EVAL_3863;
  wire [2:0] _EVAL_4148;
  wire  _EVAL_5258;
  wire  _EVAL_923;
  wire  _EVAL_1428;
  wire  _EVAL_5313;
  wire  _EVAL_2860;
  wire  _EVAL_2913;
  wire  _EVAL_175;
  wire [2:0] _EVAL_356;
  wire [2:0] _EVAL_5286;
  wire [2:0] _EVAL_1393;
  wire [2:0] _EVAL_1627;
  wire [2:0] _EVAL_2624;
  wire [2:0] _EVAL_1575;
  wire [2:0] _EVAL_4092;
  wire [6:0] _EVAL_1453;
  wire [24:0] _EVAL_5141;
  wire [30:0] _EVAL_2240;
  wire  _EVAL_278;
  wire [30:0] _EVAL_3972;
  wire [30:0] _EVAL_4308;
  wire  _EVAL_3802;
  wire [6:0] _EVAL_1802;
  wire [31:0] _EVAL_4154;
  wire  _EVAL_2914;
  wire [25:0] _EVAL_5870;
  wire [30:0] _EVAL_2134;
  wire [30:0] _EVAL_4842;
  wire [30:0] _EVAL_415;
  wire [31:0] _EVAL_2437;
  wire [31:0] _EVAL_5781;
  wire  _EVAL_4230;
  wire [2:0] _EVAL_5609;
  wire  _EVAL_1095;
  wire [31:0] _EVAL_5429;
  wire [14:0] _EVAL_2178;
  wire [31:0] _EVAL_1528;
  wire [19:0] _EVAL_755;
  wire [31:0] _EVAL_1950;
  wire [31:0] _EVAL_371;
  wire [31:0] _EVAL_3507;
  wire [31:0] _EVAL_3518;
  wire [31:0] _EVAL_642;
  wire [31:0] _EVAL_2214;
  wire [31:0] _EVAL_2200;
  wire [31:0] _EVAL_2279;
  wire [31:0] _EVAL_5175;
  wire [31:0] _EVAL_4697;
  wire [31:0] _EVAL_1498;
  wire [31:0] _EVAL_5813;
  wire [4:0] _EVAL_3032;
  wire [6:0] _EVAL_4947;
  wire [1:0] _EVAL_780;
  wire [4:0] _EVAL_5149;
  wire [26:0] _EVAL_1587;
  wire [26:0] _EVAL_1934;
  wire [7:0] _EVAL_3815;
  wire [2:0] _EVAL_4593;
  wire [4:0] _EVAL_3988;
  wire [27:0] _EVAL_6113;
  wire [26:0] _EVAL_2933;
  wire [26:0] _EVAL_4194;
  wire [26:0] _EVAL_1940;
  wire [27:0] _EVAL_2805;
  wire [3:0] _EVAL_2047;
  wire [1:0] _EVAL_252;
  wire [29:0] _EVAL_894;
  wire [29:0] _EVAL_328;
  wire [29:0] _EVAL_5593;
  wire [29:0] _EVAL_3319;
  wire [29:0] _EVAL_5487;
  wire [29:0] _EVAL_2597;
  wire [29:0] _EVAL_5123;
  wire [29:0] _EVAL_1103;
  wire [31:0] _EVAL_1947;
  wire [4:0] _EVAL_2720;
  wire [4:0] _EVAL_3562;
  wire [4:0] _EVAL_3628;
  wire  _EVAL_5099;
  wire [1:0] _EVAL_5712;
  wire [1:0] _EVAL_1187;
  wire [12:0] _EVAL_5663;
  wire  _EVAL_554;
  wire [5:0] _EVAL_1316;
  wire [3:0] _EVAL_2050;
  wire  _EVAL_3015;
  wire [31:0] _EVAL_4903;
  wire [31:0] _EVAL_5375;
  wire [9:0] _EVAL_5334;
  wire  _EVAL_1491;
  wire [1:0] _EVAL_4013;
  wire  _EVAL_1170;
  wire  _EVAL_2315;
  wire [2:0] _EVAL_1140;
  wire [20:0] _EVAL_5342;
  wire  _EVAL_5903;
  wire [9:0] _EVAL_5716;
  wire  _EVAL_5891;
  wire [7:0] _EVAL_2926;
  wire [31:0] _EVAL_1686;
  wire  _EVAL_4224;
  wire [30:0] _EVAL_913;
  wire  _EVAL_4827;
  wire [30:0] _EVAL_1169;
  wire [30:0] _EVAL_5533;
  wire  _EVAL_4062;
  wire [6:0] _EVAL_2007;
  wire [31:0] _EVAL_3113;
  wire  _EVAL_2461;
  wire [25:0] _EVAL_2113;
  wire [30:0] _EVAL_512;
  wire [30:0] _EVAL_830;
  wire [30:0] _EVAL_4813;
  wire [31:0] _EVAL_2673;
  wire [31:0] _EVAL_2005;
  wire  _EVAL_1681;
  wire [2:0] _EVAL_4764;
  wire [31:0] _EVAL_705;
  wire [14:0] _EVAL_4362;
  wire [31:0] _EVAL_3453;
  wire [19:0] _EVAL_2749;
  wire [31:0] _EVAL_5689;
  wire [31:0] _EVAL_5672;
  wire [31:0] _EVAL_4561;
  wire [31:0] _EVAL_4799;
  wire [31:0] _EVAL_2503;
  wire [31:0] _EVAL_4894;
  wire [31:0] _EVAL_5759;
  wire [31:0] _EVAL_1927;
  wire [31:0] _EVAL_5964;
  wire [31:0] _EVAL_5076;
  wire [31:0] _EVAL_479;
  wire [31:0] _EVAL_1242;
  wire [31:0] _EVAL_5851;
  wire  _EVAL_1280;
  wire [31:0] _EVAL_2710;
  wire  _EVAL_4647;
  wire [31:0] _EVAL_5315;
  wire  _EVAL_4478;
  wire [31:0] _EVAL_2445;
  wire  _EVAL_1275;
  wire  _EVAL_5396;
  wire [31:0] _EVAL_5938;
  wire  _EVAL_449;
  wire  _EVAL_4286;
  wire [31:0] _EVAL_365;
  wire [31:0] _EVAL_4689;
  wire [28:0] _EVAL_5201;
  wire  _EVAL_4226;
  wire [1:0] _EVAL_4177;
  wire  _EVAL_383;
  wire  _EVAL_5369;
  wire  _EVAL_5505;
  wire  _EVAL_486;
  wire  _EVAL_4172;
  wire  _EVAL_4140;
  wire  _EVAL_5893;
  wire [3:0] _EVAL_3550;
  wire [3:0] _EVAL_3406;
  wire [2:0] _EVAL_1773;
  wire [2:0] _EVAL_2975;
  wire [3:0] _EVAL_4318;
  wire [3:0] _EVAL_4784;
  wire  _EVAL_5997;
  wire  _EVAL_2968;
  wire  _EVAL_3370;
  wire  _EVAL_1779;
  wire  _EVAL_3679;
  wire  _EVAL_1808;
  wire [3:0] _EVAL_4633;
  wire  _EVAL_1323;
  wire  _EVAL_646;
  wire  _EVAL_5187;
  wire  _EVAL_935;
  wire  _EVAL_2547;
  wire  _EVAL_2371;
  wire  _EVAL_5740;
  wire  _EVAL_4050;
  wire  _EVAL_4302;
  wire [3:0] _EVAL_1715;
  wire  _EVAL_2486;
  wire  _EVAL_2758;
  wire  _EVAL_952;
  wire  _EVAL_2194;
  wire  _EVAL_6065;
  wire  _EVAL_3460;
  wire [31:0] _EVAL_1882;
  wire  _EVAL_222;
  wire  _EVAL_574;
  wire  _EVAL_1649;
  wire  _EVAL_600;
  wire [3:0] _EVAL_284;
  wire [3:0] _EVAL_651;
  wire  _EVAL_4453;
  wire  _EVAL_4492;
  wire  _EVAL_2940;
  wire  _EVAL_5039;
  wire [1:0] _EVAL_1766;
  wire  _EVAL_4291;
  wire [31:0] _EVAL_2539;
  wire [28:0] _EVAL_2382;
  wire  _EVAL_1310;
  wire  _EVAL_584;
  wire [2:0] _EVAL_3401;
  wire  _EVAL_979;
  wire  _EVAL_1429;
  wire  _EVAL_505;
  wire  _EVAL_1969;
  wire  _EVAL_4193;
  wire  _EVAL_2372;
  wire  _EVAL_1905;
  wire  _EVAL_1336;
  wire  _EVAL_2585;
  wire  _EVAL_5867;
  wire  _EVAL_4513;
  wire [3:0] _EVAL_4534;
  wire [3:0] _EVAL_1289;
  wire [2:0] _EVAL_4221;
  wire [3:0] _EVAL_5530;
  wire [3:0] _EVAL_3975;
  wire  _EVAL_3373;
  wire  _EVAL_4200;
  wire  _EVAL_2651;
  wire  _EVAL_1558;
  wire  _EVAL_4719;
  wire  _EVAL_2646;
  wire  _EVAL_4220;
  wire  _EVAL_2255;
  wire  _EVAL_5826;
  wire [3:0] _EVAL_2642;
  wire  _EVAL_2874;
  wire  _EVAL_1084;
  wire  _EVAL_2430;
  wire  _EVAL_1928;
  wire  _EVAL_3392;
  wire  _EVAL_1365;
  wire [31:0] _EVAL_1395;
  wire  _EVAL_3570;
  wire [31:0] _EVAL_1184;
  wire  _EVAL_1302;
  wire [31:0] _EVAL_2555;
  wire  _EVAL_4333;
  wire  _EVAL_1477;
  wire [31:0] _EVAL_5093;
  wire  _EVAL_410;
  wire  _EVAL_4325;
  wire [31:0] _EVAL_4211;
  wire  _EVAL_1265;
  wire  _EVAL_5227;
  wire [31:0] _EVAL_4801;
  wire  _EVAL_2845;
  wire  _EVAL_3957;
  wire [31:0] _EVAL_2937;
  wire  _EVAL_1384;
  wire  _EVAL_2777;
  wire [31:0] _EVAL_2819;
  wire  _EVAL_2150;
  wire  _EVAL_5754;
  wire  _EVAL_4501;
  wire  _EVAL_1910;
  wire [31:0] _EVAL_1255;
  wire  _EVAL_2545;
  wire  _EVAL_841;
  wire [31:0] _EVAL_446;
  wire  _EVAL_4572;
  wire  _EVAL_5462;
  wire [31:0] _EVAL_3041;
  wire  _EVAL_662;
  wire  _EVAL_1244;
  wire [31:0] _EVAL_2505;
  wire  _EVAL_2782;
  wire  _EVAL_5570;
  wire  _EVAL_3538;
  wire  _EVAL_463;
  wire [31:0] _EVAL_322;
  wire  _EVAL_4892;
  wire  _EVAL_2559;
  wire  _EVAL_5359;
  wire  _EVAL_689;
  wire [31:0] _EVAL_5420;
  wire  _EVAL_1560;
  wire  _EVAL_377;
  wire [31:0] _EVAL_4808;
  wire  _EVAL_4208;
  wire  _EVAL_3157;
  wire [31:0] _EVAL_4482;
  wire  _EVAL_3054;
  wire  _EVAL_2785;
  wire [31:0] _EVAL_480;
  wire  _EVAL_3970;
  wire  _EVAL_1724;
  wire [31:0] _EVAL_3608;
  wire  _EVAL_5391;
  wire  _EVAL_4654;
  wire [31:0] _EVAL_2947;
  wire  _EVAL_162;
  wire  _EVAL_4817;
  wire [31:0] _EVAL_2714;
  wire [31:0] _EVAL_4361;
  wire  _EVAL_2672;
  wire  _EVAL_197;
  wire  _EVAL_1525;
  wire  _EVAL_5845;
  wire [1:0] _EVAL_3010;
  wire [1:0] _EVAL_3528;
  wire  _EVAL_1371;
  wire  _EVAL_5276;
  wire  _EVAL_5833;
  wire  _EVAL_4360;
  wire  _EVAL_2513;
  wire  _EVAL_1061;
  wire  _EVAL_3052;
  wire [1:0] _EVAL_3573;
  wire  _EVAL_2970;
  wire  _EVAL_4887;
  wire  _EVAL_2051;
  wire  _EVAL_3045;
  wire  _EVAL_2142;
  wire [1:0] _EVAL_2797;
  wire [1:0] _EVAL_4231;
  wire [6:0] _EVAL_1213;
  wire [1:0] _EVAL_5685;
  wire [4:0] _EVAL_2915;
  wire [26:0] _EVAL_5067;
  wire [26:0] _EVAL_2744;
  wire [7:0] _EVAL_4236;
  wire [2:0] _EVAL_1545;
  wire [4:0] _EVAL_747;
  wire [27:0] _EVAL_3951;
  wire [26:0] _EVAL_595;
  wire [26:0] _EVAL_4337;
  wire [26:0] _EVAL_2622;
  wire [27:0] _EVAL_4314;
  wire [3:0] _EVAL_667;
  wire [1:0] _EVAL_3835;
  wire [29:0] _EVAL_5603;
  wire [29:0] _EVAL_1544;
  wire [29:0] _EVAL_3752;
  wire [29:0] _EVAL_6003;
  wire [29:0] _EVAL_3614;
  wire [29:0] _EVAL_708;
  wire [29:0] _EVAL_5962;
  wire [29:0] _EVAL_2878;
  wire [31:0] _EVAL_3271;
  wire [31:0] _EVAL_3897;
  wire  _EVAL_2771;
  wire [31:0] _EVAL_2034;
  wire  _EVAL_1077;
  wire  _EVAL_1079;
  wire [31:0] _EVAL_6088;
  wire  _EVAL_2192;
  wire  _EVAL_3280;
  wire [31:0] _EVAL_205;
  wire  _EVAL_4368;
  wire  _EVAL_3650;
  wire [31:0] _EVAL_5535;
  wire  _EVAL_1855;
  wire  _EVAL_5970;
  wire [31:0] _EVAL_1413;
  wire  _EVAL_4228;
  wire  _EVAL_5969;
  wire [31:0] _EVAL_303;
  wire  _EVAL_4726;
  wire  _EVAL_571;
  wire [31:0] _EVAL_5115;
  wire  _EVAL_1531;
  wire  _EVAL_5675;
  wire [31:0] _EVAL_3380;
  wire  _EVAL_1328;
  wire  _EVAL_3867;
  wire [31:0] _EVAL_3678;
  wire  _EVAL_1542;
  wire  _EVAL_683;
  wire [31:0] _EVAL_3309;
  wire  _EVAL_2183;
  wire  _EVAL_427;
  wire [31:0] _EVAL_5836;
  wire  _EVAL_1971;
  wire  _EVAL_2520;
  wire  _EVAL_3684;
  wire  _EVAL_5190;
  wire [31:0] _EVAL_3112;
  wire  _EVAL_3118;
  wire  _EVAL_2792;
  wire  _EVAL_2156;
  wire  _EVAL_4474;
  wire [31:0] _EVAL_2391;
  wire  _EVAL_5695;
  wire  _EVAL_3506;
  wire [31:0] _EVAL_5860;
  wire  _EVAL_5543;
  wire  _EVAL_2892;
  wire [31:0] _EVAL_401;
  wire  _EVAL_1639;
  wire  _EVAL_1029;
  wire [31:0] _EVAL_4878;
  wire  _EVAL_1075;
  wire  _EVAL_652;
  wire [31:0] _EVAL_2078;
  wire  _EVAL_3407;
  wire  _EVAL_775;
  wire [31:0] _EVAL_5930;
  wire  _EVAL_4946;
  wire  _EVAL_2930;
  wire [31:0] _EVAL_4219;
  wire  _EVAL_5687;
  wire  _EVAL_3584;
  wire  _EVAL_1098;
  wire  _EVAL_3398;
  wire [31:0] _EVAL_1731;
  wire  _EVAL_3850;
  wire [31:0] _EVAL_2680;
  wire  _EVAL_4875;
  wire  _EVAL_4025;
  wire [31:0] _EVAL_1671;
  wire  _EVAL_955;
  wire  _EVAL_909;
  wire  _EVAL_4554;
  wire [4:0] _EVAL_4968;
  wire [4:0] _EVAL_1682;
  wire [4:0] _EVAL_374;
  wire [4:0] _EVAL_2057;
  wire [4:0] _EVAL_4536;
  wire  _EVAL_4681;
  wire  _EVAL_2723;
  wire [31:0] _EVAL_4164;
  wire  _EVAL_3297;
  wire  _EVAL_4256;
  wire [31:0] _EVAL_4183;
  wire  _EVAL_579;
  wire [31:0] _EVAL_5311;
  wire [31:0] _EVAL_5114;
  wire  _EVAL_607;
  wire [31:0] _EVAL_3979;
  wire  _EVAL_4530;
  wire  _EVAL_4748;
  wire [31:0] _EVAL_1733;
  wire  _EVAL_1483;
  wire  _EVAL_1650;
  wire [31:0] _EVAL_3166;
  wire  _EVAL_2422;
  wire  _EVAL_4571;
  wire [31:0] _EVAL_1805;
  wire  _EVAL_3361;
  wire  _EVAL_2304;
  wire [31:0] _EVAL_3292;
  wire  _EVAL_373;
  wire [31:0] _EVAL_614;
  wire  _EVAL_3423;
  wire  _EVAL_4345;
  wire  _EVAL_2681;
  wire  _EVAL_3641;
  wire [31:0] _EVAL_3956;
  wire  _EVAL_570;
  wire  _EVAL_4059;
  wire [31:0] _EVAL_2030;
  wire  _EVAL_5532;
  wire  _EVAL_1817;
  wire  _EVAL_5926;
  wire  _EVAL_1074;
  wire [31:0] _EVAL_4939;
  wire  _EVAL_4862;
  wire [31:0] _EVAL_777;
  wire  _EVAL_1961;
  wire  _EVAL_4493;
  wire [31:0] _EVAL_3076;
  wire  _EVAL_3260;
  wire  _EVAL_2902;
  wire [31:0] _EVAL_2648;
  wire  _EVAL_2589;
  wire  _EVAL_2835;
  wire [31:0] _EVAL_2190;
  wire  _EVAL_5292;
  wire  _EVAL_1367;
  wire [31:0] _EVAL_4718;
  wire  _EVAL_4869;
  wire [31:0] _EVAL_852;
  wire  _EVAL_5171;
  wire  _EVAL_5346;
  wire [31:0] _EVAL_2438;
  wire  _EVAL_2471;
  wire  _EVAL_2698;
  wire [31:0] _EVAL_2128;
  wire  _EVAL_577;
  wire  _EVAL_1157;
  wire [31:0] _EVAL_5674;
  wire  _EVAL_5127;
  wire  _EVAL_2025;
  wire  _EVAL_2187;
  wire  _EVAL_3973;
  wire  _EVAL_5811;
  wire  _EVAL_4448;
  wire [1:0] _EVAL_3558;
  wire [2:0] _EVAL_1720;
  wire [31:0] _EVAL_960;
  wire [31:0] _EVAL_2463;
  wire [31:0] _EVAL_3111;
  wire  _EVAL_1679;
  wire  _EVAL_4085;
  wire [31:0] _EVAL_2965;
  wire  _EVAL_2924;
  wire  _EVAL_3087;
  wire  _EVAL_2950;
  wire  _EVAL_6059;
  wire [31:0] _EVAL_5006;
  wire  _EVAL_259;
  wire  _EVAL_1880;
  wire [31:0] _EVAL_5151;
  wire  _EVAL_1745;
  wire  _EVAL_1051;
  wire [31:0] _EVAL_5320;
  wire  _EVAL_5043;
  wire  _EVAL_315;
  wire [31:0] _EVAL_3607;
  wire  _EVAL_3925;
  wire  _EVAL_2577;
  wire [31:0] _EVAL_3644;
  wire  _EVAL_2364;
  wire  _EVAL_1009;
  wire [31:0] _EVAL_2451;
  wire  _EVAL_192;
  wire  _EVAL_536;
  wire [31:0] _EVAL_3391;
  wire  _EVAL_4651;
  wire  _EVAL_4297;
  wire  _EVAL_1830;
  wire  _EVAL_348;
  wire [31:0] _EVAL_4430;
  wire  _EVAL_3744;
  wire  _EVAL_1034;
  wire  _EVAL_5088;
  wire  _EVAL_1130;
  wire [31:0] _EVAL_1201;
  wire  _EVAL_5066;
  wire  _EVAL_3669;
  wire [31:0] _EVAL_643;
  wire  _EVAL_4349;
  wire  _EVAL_2001;
  wire  _EVAL_2353;
  wire  _EVAL_1058;
  wire [31:0] _EVAL_2248;
  wire  _EVAL_5789;
  wire  _EVAL_3581;
  wire [31:0] _EVAL_1591;
  wire  _EVAL_1722;
  wire [31:0] _EVAL_3927;
  wire  _EVAL_4217;
  wire  _EVAL_2938;
  wire [31:0] _EVAL_2827;
  wire  _EVAL_5949;
  wire  _EVAL_1078;
  wire [31:0] _EVAL_4806;
  wire  _EVAL_6045;
  wire [1:0] _EVAL_1647;
  wire  _EVAL_5690;
  wire [31:0] _EVAL_1585;
  wire  _EVAL_2784;
  wire [31:0] _EVAL_878;
  wire  _EVAL_2221;
  wire  _EVAL_3692;
  wire [31:0] _EVAL_5004;
  wire  _EVAL_3390;
  wire  _EVAL_1908;
  wire  _EVAL_2378;
  wire  _EVAL_2901;
  wire [31:0] _EVAL_2367;
  wire  _EVAL_5771;
  wire [31:0] _EVAL_5020;
  wire  _EVAL_4213;
  wire  _EVAL_3922;
  wire [31:0] _EVAL_5539;
  wire  _EVAL_2101;
  wire  _EVAL_559;
  wire [31:0] _EVAL_3986;
  wire  _EVAL_4419;
  wire  _EVAL_172;
  wire  _EVAL_5327;
  wire  _EVAL_1270;
  wire  _EVAL_3232;
  wire  _EVAL_4190;
  wire  _EVAL_3473;
  wire  _EVAL_4923;
  wire [3:0] _EVAL_5322;
  wire [3:0] _EVAL_5959;
  wire  _EVAL_1644;
  wire  _EVAL_2801;
  wire  _EVAL_5244;
  wire  _EVAL_4115;
  wire  _EVAL_519;
  wire  _EVAL_5620;
  wire  _EVAL_1295;
  wire  _EVAL_1972;
  wire  _EVAL_2419;
  wire  _EVAL_5527;
  wire [3:0] _EVAL_5012;
  wire  _EVAL_5541;
  wire  _EVAL_2368;
  wire  _EVAL_4079;
  wire  _EVAL_3848;
  wire  _EVAL_6064;
  wire  _EVAL_3955;
  wire  _EVAL_2357;
  wire  _EVAL_527;
  wire  _EVAL_1086;
  wire  _EVAL_2198;
  wire  _EVAL_3829;
  wire  _EVAL_1595;
  wire  _EVAL_1566;
  wire [3:0] _EVAL_5606;
  wire  _EVAL_1022;
  wire  _EVAL_2021;
  wire  _EVAL_2256;
  wire  _EVAL_3123;
  wire  _EVAL_5174;
  wire  _EVAL_1660;
  wire  _EVAL_3758;
  wire  _EVAL_5472;
  wire  _EVAL_1048;
  wire  _EVAL_2053;
  wire  _EVAL_2348;
  wire  _EVAL_5853;
  wire  _EVAL_2383;
  wire  _EVAL_2374;
  wire  _EVAL_3377;
  wire  _EVAL_991;
  wire  _EVAL_5086;
  wire  _EVAL_1278;
  wire  _EVAL_3243;
  wire  _EVAL_1555;
  wire  _EVAL_606;
  wire  _EVAL_2713;
  wire  _EVAL_2615;
  wire [3:0] _EVAL_1602;
  wire  _EVAL_660;
  wire  _EVAL_3832;
  wire  _EVAL_5489;
  wire  _EVAL_5900;
  wire  _EVAL_4138;
  wire  _EVAL_2917;
  wire  _EVAL_704;
  wire  _EVAL_1777;
  wire  _EVAL_409;
  wire  _EVAL_5454;
  wire  _EVAL_4132;
  wire  _EVAL_4295;
  wire  _EVAL_4428;
  wire  _EVAL_4168;
  wire  _EVAL_2223;
  wire  _EVAL_2945;
  wire  _EVAL_1609;
  wire  _EVAL_5937;
  wire [3:0] _EVAL_3364;
  wire  _EVAL_378;
  wire  _EVAL_3437;
  wire  _EVAL_2707;
  wire  _EVAL_3887;
  wire  _EVAL_4484;
  wire  _EVAL_4389;
  wire  _EVAL_2062;
  wire  _EVAL_5332;
  wire [3:0] _EVAL_676;
  wire  _EVAL_5676;
  wire  _EVAL_3358;
  wire  _EVAL_1380;
  wire  _EVAL_202;
  wire  _EVAL_6029;
  wire  _EVAL_5373;
  wire  _EVAL_2418;
  wire  _EVAL_4959;
  wire  _EVAL_1523;
  wire  _EVAL_2498;
  wire  _EVAL_1629;
  wire  _EVAL_3001;
  wire  _EVAL_1628;
  wire  _EVAL_3658;
  wire  _EVAL_3870;
  wire  _EVAL_3444;
  wire  _EVAL_680;
  wire  _EVAL_2337;
  wire  _EVAL_859;
  wire  _EVAL_5943;
  wire  _EVAL_4043;
  wire  _EVAL_5976;
  wire  _EVAL_6052;
  wire  _EVAL_5135;
  wire  _EVAL_5024;
  wire  _EVAL_3967;
  wire  _EVAL_803;
  wire  _EVAL_2105;
  wire  _EVAL_4401;
  wire  _EVAL_1385;
  wire  _EVAL_5430;
  wire  _EVAL_5130;
  wire  _EVAL_357;
  wire [3:0] _EVAL_4731;
  wire  _EVAL_2939;
  wire  _EVAL_618;
  wire  _EVAL_2732;
  wire  _EVAL_2429;
  wire  _EVAL_3876;
  wire  _EVAL_5725;
  wire  _EVAL_5423;
  wire  _EVAL_4189;
  wire [3:0] _EVAL_1462;
  wire  _EVAL_3445;
  wire  _EVAL_2238;
  wire  _EVAL_4754;
  wire  _EVAL_3980;
  wire  _EVAL_2949;
  wire  _EVAL_4716;
  wire  _EVAL_4218;
  wire  _EVAL_1973;
  wire  _EVAL_2216;
  wire  _EVAL_3737;
  wire  _EVAL_3940;
  wire  _EVAL_1478;
  wire  _EVAL_1422;
  wire  _EVAL_4818;
  wire  _EVAL_3070;
  wire  _EVAL_2070;
  wire  _EVAL_4848;
  wire  _EVAL_3141;
  wire  _EVAL_3321;
  wire  _EVAL_6090;
  wire [3:0] _EVAL_5516;
  wire  _EVAL_2754;
  wire  _EVAL_1357;
  wire  _EVAL_4826;
  wire  _EVAL_3337;
  wire  _EVAL_5388;
  wire  _EVAL_1826;
  wire  _EVAL_726;
  wire  _EVAL_1597;
  wire  _EVAL_3272;
  wire  _EVAL_2706;
  wire  _EVAL_2225;
  wire [3:0] _EVAL_1183;
  wire [1:0] _EVAL_2389;
  wire  _EVAL_1069;
  wire  _EVAL_4441;
  wire  _EVAL_1010;
  wire  _EVAL_798;
  wire  _EVAL_3905;
  wire  _EVAL_5880;
  wire  _EVAL_5422;
  wire  _EVAL_4481;
  wire  _EVAL_867;
  wire  _EVAL_1505;
  wire  _EVAL_5579;
  wire  _EVAL_5985;
  wire  _EVAL_3676;
  wire  _EVAL_1613;
  wire  _EVAL_258;
  wire  _EVAL_5337;
  wire  _EVAL_5777;
  wire  _EVAL_4994;
  wire  _EVAL_3529;
  wire  _EVAL_1930;
  wire  _EVAL_3904;
  wire  _EVAL_4772;
  wire  _EVAL_6031;
  wire  _EVAL_1226;
  wire [3:0] _EVAL_3219;
  wire  _EVAL_1217;
  wire  _EVAL_2765;
  wire  _EVAL_1699;
  wire  _EVAL_2002;
  wire [3:0] _EVAL_5251;
  wire [3:0] _EVAL_907;
  wire [3:0] _EVAL_2058;
  wire [3:0] _EVAL_4445;
  wire [3:0] _EVAL_3266;
  wire [31:0] _EVAL_232;
  wire  _EVAL_3554;
  wire [31:0] _EVAL_1757;
  wire  _EVAL_360;
  wire  _EVAL_2867;
  wire [31:0] _EVAL_1291;
  wire [31:0] _EVAL_4961;
  wire [31:0] _EVAL_454;
  wire [31:0] _EVAL_532;
  wire [31:0] _EVAL_4856;
  wire [31:0] _EVAL_3893;
  wire  _EVAL_641;
  wire  _EVAL_2303;
  wire  _EVAL_3103;
  wire  _EVAL_3107;
  wire  _EVAL_914;
  wire  _EVAL_5770;
  wire  _EVAL_432;
  wire  _EVAL_5748;
  wire  _EVAL_3728;
  wire  _EVAL_6011;
  wire  _EVAL_391;
  wire [31:0] _EVAL_740;
  wire [31:0] _EVAL_4622;
  wire  _EVAL_6009;
  wire [31:0] _EVAL_3996;
  wire  _EVAL_1191;
  wire [31:0] _EVAL_5801;
  wire  _EVAL_4737;
  wire  _EVAL_3387;
  wire [31:0] _EVAL_3680;
  wire  _EVAL_4232;
  wire  _EVAL_1272;
  wire [31:0] _EVAL_3618;
  wire  _EVAL_1764;
  wire [31:0] _EVAL_4343;
  wire  _EVAL_1709;
  wire  _EVAL_3575;
  wire [31:0] _EVAL_4930;
  wire  _EVAL_4636;
  wire  _EVAL_467;
  wire [31:0] _EVAL_5820;
  wire [31:0] _EVAL_4227;
  wire [31:0] _EVAL_362;
  wire  _EVAL_4434;
  wire [31:0] _EVAL_2696;
  wire  _EVAL_426;
  wire  _EVAL_1845;
  wire [31:0] _EVAL_5778;
  wire  _EVAL_3899;
  wire  _EVAL_968;
  wire [4:0] _EVAL_4490;
  wire [4:0] _EVAL_1621;
  wire [4:0] _EVAL_3256;
  wire [4:0] _EVAL_5155;
  wire [4:0] _EVAL_329;
  wire [4:0] _EVAL_880;
  wire [31:0] _EVAL_2144;
  wire  _EVAL_1433;
  wire [31:0] _EVAL_4790;
  wire  _EVAL_4271;
  wire  _EVAL_4136;
  wire  _EVAL_1361;
  wire [31:0] _EVAL_3654;
  wire  _EVAL_2020;
  wire  _EVAL_3755;
  wire [31:0] _EVAL_5191;
  wire  _EVAL_1781;
  wire  _EVAL_1975;
  wire [1:0] _EVAL_2341;
  wire [3:0] _EVAL_2439;
  wire [7:0] _EVAL_1666;
  wire [2:0] _EVAL_462;
  wire [4:0] _EVAL_772;
  wire [27:0] _EVAL_4956;
  wire [27:0] _EVAL_3193;
  wire [8:0] _EVAL_1968;
  wire [3:0] _EVAL_5604;
  wire [4:0] _EVAL_3146;
  wire [28:0] _EVAL_1926;
  wire  _EVAL_3798;
  wire [24:0] _EVAL_2603;
  wire  _EVAL_5207;
  wire [24:0] _EVAL_4020;
  wire [24:0] _EVAL_3416;
  wire [17:0] _EVAL_1109;
  wire [24:0] _EVAL_2325;
  wire [24:0] _EVAL_4404;
  wire [24:0] _EVAL_3939;
  wire [24:0] _EVAL_5815;
  wire [24:0] _EVAL_455;
  wire [24:0] _EVAL_3329;
  wire [24:0] _EVAL_3768;
  wire [1:0] _EVAL_5183;
  wire [2:0] _EVAL_1842;
  wire [27:0] _EVAL_2215;
  wire [27:0] _EVAL_3291;
  wire [28:0] _EVAL_5363;
  wire [25:0] _EVAL_4807;
  wire [28:0] _EVAL_5785;
  wire [28:0] _EVAL_592;
  wire [28:0] _EVAL_5203;
  wire [28:0] _EVAL_1663;
  wire [28:0] _EVAL_430;
  wire [28:0] _EVAL_2497;
  wire [28:0] _EVAL_2440;
  wire [31:0] _EVAL_888;
  wire [31:0] _EVAL_2898;
  wire  _EVAL_6120;
  wire [11:0] _EVAL_5634;
  wire  _EVAL_4843;
  wire  _EVAL_5966;
  wire  _EVAL_526;
  wire  _EVAL_1986;
  wire [31:0] _EVAL_3164;
  wire  _EVAL_5713;
  wire  _EVAL_5504;
  wire  _EVAL_4711;
  wire [31:0] _EVAL_3160;
  wire [31:0] _EVAL_1618;
  wire  _EVAL_5724;
  wire [31:0] _EVAL_4982;
  wire  _EVAL_1355;
  wire [31:0] _EVAL_1368;
  wire  _EVAL_4987;
  wire  _EVAL_3046;
  wire [31:0] _EVAL_1832;
  wire  _EVAL_3545;
  wire  _EVAL_6105;
  wire [31:0] _EVAL_5364;
  wire  _EVAL_5715;
  wire  _EVAL_2709;
  wire [31:0] _EVAL_2690;
  wire  _EVAL_2063;
  wire  _EVAL_1638;
  wire [31:0] _EVAL_4864;
  wire  _EVAL_1646;
  wire  _EVAL_1944;
  wire [31:0] _EVAL_6022;
  wire  _EVAL_1864;
  wire  _EVAL_4810;
  wire [31:0] _EVAL_3794;
  wire  _EVAL_3645;
  wire  _EVAL_1651;
  wire [31:0] _EVAL_3869;
  wire  _EVAL_1853;
  wire  _EVAL_1937;
  wire [31:0] _EVAL_5219;
  wire  _EVAL_1407;
  wire  _EVAL_5119;
  wire [31:0] _EVAL_2029;
  wire  _EVAL_5661;
  wire  _EVAL_5089;
  wire [31:0] _EVAL_996;
  wire  _EVAL_2936;
  wire  _EVAL_2048;
  wire  _EVAL_5947;
  wire  _EVAL_4237;
  wire [31:0] _EVAL_5054;
  wire  _EVAL_5253;
  wire  _EVAL_2307;
  wire  _EVAL_4658;
  wire  _EVAL_1102;
  wire [31:0] _EVAL_2456;
  wire  _EVAL_3439;
  wire  _EVAL_2299;
  wire [31:0] _EVAL_3954;
  wire  _EVAL_2780;
  wire  _EVAL_4823;
  wire [31:0] _EVAL_5287;
  wire  _EVAL_5596;
  wire  _EVAL_887;
  wire [31:0] _EVAL_1604;
  wire  _EVAL_5095;
  wire  _EVAL_5483;
  wire [31:0] _EVAL_3180;
  wire  _EVAL_2016;
  wire  _EVAL_5231;
  wire [31:0] _EVAL_2322;
  wire  _EVAL_5398;
  wire  _EVAL_4351;
  wire [31:0] _EVAL_1956;
  wire  _EVAL_4665;
  wire  _EVAL_4663;
  wire  _EVAL_601;
  wire  _EVAL_3119;
  wire [31:0] _EVAL_2627;
  wire  _EVAL_3020;
  wire  _EVAL_987;
  wire  _EVAL_1045;
  wire  _EVAL_5519;
  wire [31:0] _EVAL_3278;
  wire  _EVAL_1510;
  wire  _EVAL_1239;
  wire [31:0] _EVAL_4496;
  wire  _EVAL_2208;
  wire [7:0] _EVAL_4931;
  wire  _EVAL_2558;
  wire  _EVAL_2979;
  wire  _EVAL_4388;
  wire  _EVAL_2179;
  wire  _EVAL_5305;
  wire  _EVAL_2770;
  wire [31:0] _EVAL_4950;
  wire  _EVAL_3379;
  wire [31:0] _EVAL_5665;
  wire  _EVAL_2866;
  wire [31:0] _EVAL_3255;
  wire [31:0] _EVAL_3985;
  wire [31:0] _EVAL_389;
  wire [31:0] _EVAL_3298;
  wire  _EVAL_1702;
  wire [31:0] _EVAL_4821;
  wire  _EVAL_1680;
  wire [31:0] _EVAL_6070;
  wire  _EVAL_942;
  wire  _EVAL_1013;
  wire  _EVAL_1578;
  wire [31:0] _EVAL_5323;
  wire  _EVAL_3447;
  wire  _EVAL_5575;
  wire [31:0] _EVAL_1458;
  wire [31:0] _EVAL_1974;
  wire  _EVAL_617;
  wire [31:0] _EVAL_621;
  wire  _EVAL_2449;
  wire [31:0] _EVAL_1550;
  wire  _EVAL_4779;
  wire  _EVAL_3713;
  wire [31:0] _EVAL_4301;
  wire  _EVAL_1015;
  wire  _EVAL_5787;
  wire  _EVAL_3843;
  wire  _EVAL_5164;
  wire [31:0] _EVAL_5854;
  wire [31:0] _EVAL_6084;
  wire  _EVAL_2941;
  wire [31:0] _EVAL_1642;
  wire  _EVAL_4567;
  wire  _EVAL_2052;
  wire [31:0] _EVAL_1804;
  wire  _EVAL_6080;
  wire  _EVAL_1829;
  wire [31:0] _EVAL_1259;
  wire  _EVAL_787;
  wire [31:0] _EVAL_2678;
  wire  _EVAL_3715;
  wire  _EVAL_609;
  wire [31:0] _EVAL_2090;
  wire  _EVAL_1197;
  wire  _EVAL_1203;
  wire [31:0] _EVAL_540;
  wire  _EVAL_4403;
  wire  _EVAL_3890;
  wire [31:0] _EVAL_5072;
  wire [31:0] _EVAL_5400;
  wire  _EVAL_5224;
  wire [31:0] _EVAL_2130;
  wire  _EVAL_1448;
  wire  _EVAL_5899;
  wire [4:0] _EVAL_3215;
  wire [1:0] _EVAL_736;
  wire  _EVAL_3722;
  wire  _EVAL_3659;
  wire [14:0] _EVAL_4425;
  wire  _EVAL_359;
  wire [31:0] _EVAL_4334;
  wire  _EVAL_4045;
  wire  _EVAL_4858;
  wire [31:0] _EVAL_4602;
  wire  _EVAL_1634;
  wire [31:0] _EVAL_516;
  wire  _EVAL_3286;
  wire  _EVAL_2154;
  wire [31:0] _EVAL_3417;
  wire [31:0] _EVAL_4466;
  wire [31:0] _EVAL_4660;
  wire  _EVAL_1936;
  wire [31:0] _EVAL_4031;
  wire  _EVAL_975;
  wire  _EVAL_2233;
  wire  _EVAL_604;
  wire [31:0] _EVAL_5325;
  wire  _EVAL_2334;
  wire  _EVAL_3836;
  wire [31:0] _EVAL_5999;
  wire  _EVAL_3098;
  wire [10:0] _EVAL_4355;
  wire  _EVAL_2795;
  wire  _EVAL_1236;
  wire  _EVAL_1598;
  wire  _EVAL_4920;
  wire  _EVAL_5008;
  wire  _EVAL_2116;
  wire  _EVAL_846;
  wire [31:0] _EVAL_4646;
  wire  _EVAL_2329;
  wire  _EVAL_1007;
  wire [31:0] _EVAL_6137;
  wire  _EVAL_4639;
  wire  _EVAL_3310;
  wire [31:0] _EVAL_5463;
  wire  _EVAL_5215;
  wire  _EVAL_3731;
  wire  _EVAL_4244;
  wire  _EVAL_4239;
  wire [31:0] _EVAL_4671;
  wire  _EVAL_293;
  wire  _EVAL_5268;
  wire [31:0] _EVAL_5622;
  wire  _EVAL_2147;
  wire  _EVAL_1652;
  wire  _EVAL_4829;
  wire  _EVAL_6006;
  wire  _EVAL_4282;
  wire  _EVAL_5384;
  wire  _EVAL_2669;
  wire  _EVAL_1669;
  wire  _EVAL_1537;
  wire [31:0] _EVAL_4583;
  wire  _EVAL_5738;
  wire  _EVAL_1856;
  wire [31:0] _EVAL_3133;
  wire  _EVAL_5912;
  wire  _EVAL_3451;
  wire [31:0] _EVAL_5582;
  wire  _EVAL_2741;
  wire  _EVAL_2296;
  wire [31:0] _EVAL_939;
  wire  _EVAL_4998;
  wire  _EVAL_1317;
  wire [31:0] _EVAL_3609;
  wire  _EVAL_2952;
  wire  _EVAL_2516;
  wire  _EVAL_5756;
  wire  _EVAL_4004;
  wire  _EVAL_5060;
  wire [31:0] _EVAL_1912;
  wire  _EVAL_1027;
  wire [31:0] _EVAL_1541;
  wire  _EVAL_3323;
  wire [31:0] _EVAL_3018;
  wire [31:0] _EVAL_246;
  wire  _EVAL_715;
  wire [4:0] _EVAL_5303;
  wire [4:0] _EVAL_1163;
  wire [4:0] _EVAL_1324;
  wire [4:0] _EVAL_4638;
  wire [4:0] _EVAL_5452;
  wire [4:0] _EVAL_3003;
  wire [4:0] _EVAL_2570;
  wire [31:0] _EVAL_2405;
  wire  _EVAL_4978;
  wire  _EVAL_4462;
  wire [31:0] _EVAL_2811;
  wire [31:0] _EVAL_2858;
  wire  _EVAL_624;
  wire [31:0] _EVAL_5670;
  wire  _EVAL_1868;
  wire  _EVAL_1356;
  wire [31:0] _EVAL_3194;
  wire  _EVAL_677;
  wire  _EVAL_213;
  wire [31:0] _EVAL_2500;
  wire  _EVAL_1846;
  wire  _EVAL_4206;
  wire [31:0] _EVAL_5908;
  wire  _EVAL_950;
  wire  _EVAL_5438;
  wire [31:0] _EVAL_3088;
  wire  _EVAL_4890;
  wire  _EVAL_6037;
  wire  _EVAL_2607;
  wire  _EVAL_1464;
  wire  _EVAL_2274;
  wire [31:0] _EVAL_1697;
  wire  _EVAL_1327;
  wire  _EVAL_397;
  wire [31:0] _EVAL_5222;
  wire  _EVAL_4354;
  wire  _EVAL_270;
  wire  _EVAL_3413;
  wire  _EVAL_5525;
  wire  _EVAL_5062;
  wire  _EVAL_1451;
  wire  _EVAL_4350;
  wire  _EVAL_3426;
  wire  _EVAL_2152;
  wire  _EVAL_4510;
  wire  _EVAL_351;
  wire  _EVAL_3787;
  wire  _EVAL_6131;
  wire [31:0] _EVAL_4373;
  wire  _EVAL_4084;
  wire  _EVAL_1985;
  wire  _EVAL_5521;
  wire  _EVAL_3318;
  wire [31:0] _EVAL_638;
  wire  _EVAL_2879;
  wire  _EVAL_4528;
  wire [31:0] _EVAL_6040;
  wire  _EVAL_1264;
  wire  _EVAL_5601;
  wire [31:0] _EVAL_5495;
  wire  _EVAL_1205;
  wire  _EVAL_300;
  wire [31:0] _EVAL_4504;
  wire  _EVAL_1399;
  wire  _EVAL_1219;
  wire  _EVAL_4055;
  wire  _EVAL_2692;
  wire [31:0] _EVAL_6125;
  wire  _EVAL_3435;
  wire  _EVAL_3600;
  wire [31:0] _EVAL_4596;
  wire  _EVAL_2806;
  wire  _EVAL_1005;
  wire [31:0] _EVAL_5822;
  wire  _EVAL_445;
  wire  _EVAL_3931;
  wire  _EVAL_5432;
  wire  _EVAL_3732;
  wire [31:0] _EVAL_1844;
  wire  _EVAL_4209;
  wire  _EVAL_2865;
  wire [31:0] _EVAL_2843;
  wire  _EVAL_6132;
  wire  _EVAL_5326;
  wire  _EVAL_5173;
  wire  _EVAL_2076;
  wire [31:0] _EVAL_2452;
  wire  _EVAL_5193;
  wire [31:0] _EVAL_4704;
  wire  _EVAL_1955;
  wire [31:0] _EVAL_1879;
  wire  _EVAL_3770;
  wire [31:0] _EVAL_3911;
  wire  _EVAL_5611;
  wire  _EVAL_752;
  wire [31:0] _EVAL_1515;
  wire  _EVAL_2895;
  wire  _EVAL_473;
  wire [31:0] _EVAL_1851;
  wire  _EVAL_988;
  wire  _EVAL_1893;
  wire [31:0] _EVAL_6075;
  wire  _EVAL_247;
  wire  _EVAL_2875;
  wire [31:0] _EVAL_4548;
  wire  _EVAL_1390;
  wire  _EVAL_3739;
  wire [31:0] _EVAL_260;
  wire  _EVAL_1819;
  wire  _EVAL_340;
  wire [31:0] _EVAL_4383;
  wire  _EVAL_3097;
  wire  _EVAL_1370;
  wire [31:0] _EVAL_1665;
  wire  _EVAL_4729;
  wire  _EVAL_5876;
  wire [31:0] _EVAL_2028;
  wire  _EVAL_3606;
  wire  _EVAL_1285;
  wire [31:0] _EVAL_4174;
  wire  _EVAL_4788;
  wire  _EVAL_3711;
  wire [31:0] _EVAL_518;
  wire  _EVAL_1511;
  wire  _EVAL_2229;
  wire  _EVAL_2393;
  wire  _EVAL_3214;
  wire [31:0] _EVAL_5709;
  wire  _EVAL_5855;
  wire  _EVAL_5745;
  wire  _EVAL_4541;
  wire  _EVAL_3211;
  wire [31:0] _EVAL_1708;
  wire  _EVAL_3784;
  wire  _EVAL_5014;
  wire [31:0] _EVAL_5058;
  wire  _EVAL_3961;
  wire  _EVAL_1230;
  wire [31:0] _EVAL_3605;
  wire  _EVAL_3419;
  wire  _EVAL_3792;
  wire [31:0] _EVAL_2338;
  wire  _EVAL_1540;
  wire  _EVAL_546;
  wire [31:0] _EVAL_4942;
  wire  _EVAL_2320;
  wire  _EVAL_710;
  wire [31:0] _EVAL_2587;
  wire  _EVAL_5792;
  wire  _EVAL_731;
  wire  _EVAL_2980;
  wire  _EVAL_3700;
  wire  _EVAL_4980;
  wire  _EVAL_5284;
  wire [31:0] _EVAL_1374;
  wire  _EVAL_1221;
  wire  _EVAL_3719;
  wire  _EVAL_2578;
  wire  _EVAL_5482;
  wire [31:0] _EVAL_5392;
  wire  _EVAL_2571;
  wire  _EVAL_3533;
  wire [31:0] _EVAL_5464;
  wire  _EVAL_4989;
  wire  _EVAL_5488;
  wire [31:0] _EVAL_5584;
  wire  _EVAL_5784;
  wire  _EVAL_5234;
  wire [31:0] _EVAL_503;
  wire  _EVAL_2783;
  wire [31:0] _EVAL_596;
  wire  _EVAL_929;
  wire  _EVAL_585;
  wire [31:0] _EVAL_6051;
  wire  _EVAL_848;
  wire  _EVAL_3063;
  wire [31:0] _EVAL_4835;
  wire  _EVAL_2854;
  wire  _EVAL_891;
  wire  _EVAL_5186;
  wire  _EVAL_1151;
  wire [31:0] _EVAL_3071;
  wire  _EVAL_5167;
  wire  _EVAL_1822;
  wire [31:0] _EVAL_4432;
  wire  _EVAL_4517;
  wire  _EVAL_5056;
  wire [31:0] _EVAL_238;
  wire  _EVAL_4657;
  wire  _EVAL_4016;
  wire [31:0] _EVAL_5664;
  wire  _EVAL_1257;
  wire  _EVAL_2239;
  wire [31:0] _EVAL_3074;
  wire  _EVAL_5028;
  wire  _EVAL_3056;
  wire [31:0] _EVAL_1590;
  wire  _EVAL_2493;
  wire  _EVAL_4052;
  wire [31:0] _EVAL_2244;
  wire  _EVAL_1420;
  wire  _EVAL_3515;
  wire [31:0] _EVAL_3741;
  wire  _EVAL_1018;
  wire  _EVAL_5898;
  wire [31:0] _EVAL_2976;
  wire  _EVAL_2961;
  wire  _EVAL_484;
  wire [31:0] _EVAL_1292;
  wire  _EVAL_679;
  wire  _EVAL_4151;
  wire [31:0] _EVAL_6111;
  wire  _EVAL_297;
  wire  _EVAL_2684;
  wire  _EVAL_564;
  wire  _EVAL_3369;
  wire [31:0] _EVAL_279;
  wire  _EVAL_5446;
  wire  _EVAL_5232;
  wire  _EVAL_4060;
  wire  _EVAL_4171;
  wire [31:0] _EVAL_4795;
  wire  _EVAL_4409;
  wire  _EVAL_5783;
  wire [31:0] _EVAL_895;
  wire  _EVAL_5491;
  wire  _EVAL_2905;
  wire [31:0] _EVAL_5776;
  wire [4:0] _EVAL_4076;
  wire [31:0] _EVAL_1224;
  wire  _EVAL_2759;
  wire [31:0] _EVAL_3693;
  wire  _EVAL_1685;
  wire  _EVAL_5621;
  wire [31:0] _EVAL_3729;
  wire  _EVAL_4415;
  wire  _EVAL_728;
  wire [31:0] _EVAL_4263;
  wire  _EVAL_3521;
  wire  _EVAL_344;
  wire [31:0] _EVAL_273;
  wire  _EVAL_5494;
  wire  _EVAL_5688;
  wire [31:0] _EVAL_3638;
  wire  _EVAL_5978;
  wire [31:0] _EVAL_1501;
  wire  _EVAL_4468;
  wire  _EVAL_3806;
  wire [31:0] _EVAL_337;
  wire  _EVAL_4269;
  wire  _EVAL_1315;
  wire [31:0] _EVAL_2148;
  wire  _EVAL_1559;
  wire  _EVAL_1835;
  wire [31:0] _EVAL_2685;
  wire  _EVAL_5581;
  wire [31:0] _EVAL_499;
  wire  _EVAL_497;
  wire  _EVAL_2161;
  wire  _EVAL_4913;
  wire [31:0] _EVAL_2530;
  wire  _EVAL_2697;
  wire  _EVAL_4142;
  wire [31:0] _EVAL_2881;
  wire  _EVAL_4863;
  wire  _EVAL_4509;
  wire [31:0] _EVAL_3208;
  wire  _EVAL_4512;
  wire  _EVAL_1126;
  wire [31:0] _EVAL_2910;
  wire  _EVAL_4129;
  wire  _EVAL_3660;
  wire [31:0] _EVAL_2574;
  wire  _EVAL_3724;
  wire  _EVAL_3322;
  wire [31:0] _EVAL_1068;
  wire  _EVAL_5524;
  wire  _EVAL_3264;
  wire [31:0] _EVAL_739;
  wire  _EVAL_3639;
  wire  _EVAL_4644;
  wire [31:0] _EVAL_2193;
  wire  _EVAL_5117;
  wire  _EVAL_5749;
  wire [31:0] _EVAL_5274;
  wire  _EVAL_4725;
  wire  _EVAL_5633;
  wire  _EVAL_1057;
  wire  _EVAL_5182;
  wire [31:0] _EVAL_5919;
  wire  _EVAL_5773;
  wire  _EVAL_3040;
  wire  _EVAL_3661;
  wire  _EVAL_3184;
  wire [31:0] _EVAL_3135;
  wire  _EVAL_1546;
  wire  _EVAL_3734;
  wire [31:0] _EVAL_3374;
  wire  _EVAL_1241;
  wire  _EVAL_2882;
  wire [31:0] _EVAL_5646;
  wire  _EVAL_495;
  wire  _EVAL_1790;
  wire [31:0] _EVAL_2829;
  wire  _EVAL_5752;
  wire  _EVAL_4971;
  wire [31:0] _EVAL_5240;
  wire  _EVAL_1933;
  wire  _EVAL_2459;
  wire [31:0] _EVAL_3522;
  wire  _EVAL_332;
  wire  _EVAL_354;
  wire [31:0] _EVAL_4973;
  wire  _EVAL_666;
  wire  _EVAL_4724;
  wire  _EVAL_4668;
  wire  _EVAL_629;
  wire [31:0] _EVAL_2074;
  wire  _EVAL_5479;
  wire  _EVAL_4859;
  wire  _EVAL_5105;
  wire  _EVAL_5808;
  wire [31:0] _EVAL_3686;
  wire  _EVAL_2196;
  wire  _EVAL_5907;
  wire [31:0] _EVAL_3696;
  wire  _EVAL_6077;
  wire  _EVAL_4977;
  wire [31:0] _EVAL_1620;
  wire  _EVAL_2386;
  wire  _EVAL_954;
  wire [31:0] _EVAL_5029;
  wire  _EVAL_2185;
  wire  _EVAL_3036;
  wire  _EVAL_962;
  wire  _EVAL_504;
  wire [31:0] _EVAL_1300;
  wire  _EVAL_3577;
  wire [31:0] _EVAL_4069;
  wire  _EVAL_4074;
  wire [31:0] _EVAL_5170;
  wire  _EVAL_3788;
  wire  _EVAL_4451;
  wire [31:0] _EVAL_2863;
  wire  _EVAL_4965;
  wire  _EVAL_741;
  wire [31:0] _EVAL_5883;
  wire  _EVAL_4495;
  wire  _EVAL_450;
  wire [31:0] _EVAL_4604;
  wire  _EVAL_3222;
  wire  _EVAL_321;
  wire [31:0] _EVAL_1673;
  wire  _EVAL_3115;
  wire  _EVAL_4235;
  wire [31:0] _EVAL_4692;
  wire  _EVAL_4439;
  wire  _EVAL_460;
  wire [31:0] _EVAL_3121;
  wire  _EVAL_4255;
  wire  _EVAL_911;
  wire [31:0] _EVAL_4708;
  wire  _EVAL_5176;
  wire  _EVAL_4511;
  wire [31:0] _EVAL_2519;
  wire  _EVAL_2612;
  wire  _EVAL_1392;
  wire [31:0] _EVAL_533;
  wire  _EVAL_6117;
  wire  _EVAL_5586;
  wire [31:0] _EVAL_5990;
  wire  _EVAL_5637;
  wire  _EVAL_5189;
  wire [31:0] _EVAL_4739;
  wire  _EVAL_3290;
  wire  _EVAL_353;
  wire  _EVAL_2868;
  wire  _EVAL_4545;
  wire [31:0] _EVAL_4048;
  wire  _EVAL_5585;
  wire  _EVAL_1877;
  wire  _EVAL_3851;
  wire  _EVAL_1435;
  wire [31:0] _EVAL_1732;
  wire  _EVAL_1417;
  wire  _EVAL_404;
  wire [31:0] _EVAL_4011;
  wire  _EVAL_985;
  wire  _EVAL_5590;
  wire [31:0] _EVAL_6014;
  wire  _EVAL_2431;
  wire  _EVAL_5097;
  wire [31:0] _EVAL_1989;
  wire  _EVAL_714;
  wire  _EVAL_2809;
  wire [31:0] _EVAL_368;
  wire  _EVAL_3484;
  wire  _EVAL_5316;
  wire [31:0] _EVAL_1311;
  wire  _EVAL_857;
  wire  _EVAL_2623;
  wire  _EVAL_1099;
  wire  _EVAL_2473;
  wire  _EVAL_3915;
  wire  _EVAL_2097;
  wire [31:0] _EVAL_364;
  wire  _EVAL_615;
  wire  _EVAL_5694;
  wire  _EVAL_5458;
  wire  _EVAL_978;
  wire [31:0] _EVAL_3549;
  wire  _EVAL_4857;
  wire  _EVAL_1167;
  wire  _EVAL_1144;
  wire [31:0] _EVAL_637;
  wire  _EVAL_993;
  wire  _EVAL_236;
  wire [31:0] _EVAL_2694;
  wire [31:0] _EVAL_4589;
  wire [31:0] _EVAL_4064;
  wire  _EVAL_4598;
  wire  _EVAL_3487;
  wire  _EVAL_2851;
  wire [31:0] _EVAL_3415;
  wire [31:0] _EVAL_2344;
  wire  _EVAL_6074;
  wire  _EVAL_5772;
  wire [31:0] _EVAL_1960;
  wire  _EVAL_1484;
  wire  _EVAL_2703;
  wire [31:0] _EVAL_2460;
  wire [31:0] _EVAL_4159;
  wire  _EVAL_5558;
  wire  _EVAL_3785;
  wire  _EVAL_394;
  wire [31:0] _EVAL_5739;
  wire  _EVAL_4413;
  wire  _EVAL_2944;
  wire [31:0] _EVAL_3022;
  wire [31:0] _EVAL_4606;
  wire  _EVAL_2069;
  wire [10:0] _EVAL_730;
  wire [31:0] _EVAL_2844;
  wire  _EVAL_974;
  wire [31:0] _EVAL_5691;
  wire  _EVAL_2772;
  wire  _EVAL_767;
  wire [31:0] _EVAL_471;
  wire  _EVAL_567;
  wire  _EVAL_5569;
  wire [31:0] _EVAL_5350;
  wire  _EVAL_628;
  wire  _EVAL_3509;
  wire  _EVAL_4953;
  wire  _EVAL_889;
  wire [31:0] _EVAL_6026;
  wire  _EVAL_2064;
  wire [31:0] _EVAL_4941;
  wire  _EVAL_697;
  wire  _EVAL_2853;
  wire  _EVAL_4395;
  wire [31:0] _EVAL_927;
  wire  _EVAL_1460;
  wire [4:0] _EVAL_5297;
  wire  _EVAL_4371;
  wire [31:0] _EVAL_5657;
  wire [31:0] _EVAL_5124;
  wire  _EVAL_3635;
  wire  _EVAL_3029;
  wire [31:0] _EVAL_1318;
  wire  _EVAL_4749;
  wire  _EVAL_2509;
  wire [31:0] _EVAL_4106;
  wire  _EVAL_1667;
  wire  _EVAL_653;
  wire [31:0] _EVAL_267;
  wire  _EVAL_1693;
  wire  _EVAL_3332;
  wire [31:0] _EVAL_4412;
  wire  _EVAL_3192;
  wire  _EVAL_4804;
  wire [31:0] _EVAL_565;
  wire  _EVAL_5360;
  wire  _EVAL_3790;
  wire [31:0] _EVAL_5389;
  wire  _EVAL_4187;
  wire  _EVAL_5194;
  wire [31:0] _EVAL_3262;
  wire  _EVAL_3963;
  wire  _EVAL_2359;
  wire [31:0] _EVAL_2825;
  wire  _EVAL_5496;
  wire  _EVAL_2054;
  wire [31:0] _EVAL_5531;
  wire  _EVAL_1866;
  wire  _EVAL_634;
  wire [31:0] _EVAL_2465;
  wire  _EVAL_3428;
  wire  _EVAL_5932;
  wire  _EVAL_4167;
  wire  _EVAL_4450;
  wire [31:0] _EVAL_2012;
  wire  _EVAL_5896;
  wire  _EVAL_5210;
  wire  _EVAL_2476;
  wire  _EVAL_3632;
  wire [31:0] _EVAL_2191;
  wire [4:0] _EVAL_1635;
  wire [4:0] _EVAL_1662;
  wire [4:0] _EVAL_5293;
  wire [4:0] _EVAL_2862;
  wire [4:0] _EVAL_1332;
  wire [10:0] _EVAL_3514;
  wire  _EVAL_769;
  wire  _EVAL_1364;
  wire  _EVAL_5923;
  wire  _EVAL_5104;
  wire  _EVAL_2464;
  wire [31:0] _EVAL_1198;
  wire [31:0] _EVAL_1935;
  wire [11:0] _EVAL_1573;
  wire  _EVAL_5245;
  wire  _EVAL_4002;
  wire  _EVAL_3675;
  wire  _EVAL_922;
  wire  _EVAL_1350;
  wire  _EVAL_5243;
  wire  _EVAL_1405;
  wire [31:0] _EVAL_1263;
  wire  _EVAL_2411;
  wire  _EVAL_6083;
  wire  _EVAL_5925;
  wire  _EVAL_2550;
  wire [31:0] _EVAL_2434;
  wire  _EVAL_524;
  wire  _EVAL_1800;
  wire  _EVAL_5300;
  wire  _EVAL_5589;
  wire [31:0] _EVAL_2234;
  wire  _EVAL_542;
  wire  _EVAL_1820;
  wire [31:0] _EVAL_280;
  wire  _EVAL_3976;
  wire  _EVAL_307;
  wire [3:0] _EVAL_304;
  wire [31:0] _EVAL_4463;
  wire  _EVAL_1495;
  wire [31:0] _EVAL_1995;
  wire  _EVAL_5658;
  wire [31:0] _EVAL_3348;
  wire  _EVAL_1728;
  wire [31:0] _EVAL_5528;
  wire  _EVAL_610;
  wire  _EVAL_2687;
  wire  _EVAL_4421;
  wire [31:0] _EVAL_3499;
  wire  _EVAL_850;
  wire [31:0] _EVAL_4118;
  wire  _EVAL_1186;
  wire  _EVAL_345;
  wire [31:0] _EVAL_2287;
  wire  _EVAL_528;
  wire  _EVAL_5202;
  wire [31:0] _EVAL_2146;
  wire  _EVAL_5818;
  wire  _EVAL_1059;
  wire [31:0] _EVAL_1083;
  wire  _EVAL_582;
  wire  _EVAL_758;
  wire [31:0] _EVAL_1942;
  wire  _EVAL_849;
  wire  _EVAL_4473;
  wire [31:0] _EVAL_3424;
  wire  _EVAL_4197;
  wire  _EVAL_813;
  wire [31:0] _EVAL_5348;
  wire  _EVAL_4649;
  wire  _EVAL_4505;
  wire [31:0] _EVAL_2757;
  wire  _EVAL_4860;
  wire  _EVAL_1783;
  wire [31:0] _EVAL_5501;
  wire  _EVAL_2872;
  wire  _EVAL_5862;
  wire [31:0] _EVAL_5877;
  wire  _EVAL_5280;
  wire  _EVAL_2269;
  wire [31:0] _EVAL_3796;
  wire  _EVAL_2502;
  wire  _EVAL_5233;
  wire  _EVAL_177;
  wire  _EVAL_3394;
  wire [31:0] _EVAL_2072;
  wire  _EVAL_1261;
  wire  _EVAL_2527;
  wire  _EVAL_2748;
  wire  _EVAL_2746;
  wire [31:0] _EVAL_5144;
  wire  _EVAL_1104;
  wire  _EVAL_5110;
  wire [31:0] _EVAL_2083;
  wire  _EVAL_3599;
  wire  _EVAL_1442;
  wire  _EVAL_623;
  wire  _EVAL_2123;
  wire [31:0] _EVAL_3067;
  wire  _EVAL_2859;
  wire  _EVAL_4086;
  wire [31:0] _EVAL_2581;
  wire  _EVAL_2201;
  wire  _EVAL_2507;
  wire  _EVAL_1064;
  wire  _EVAL_915;
  wire  _EVAL_4192;
  wire  _EVAL_2485;
  wire [31:0] _EVAL_240;
  wire  _EVAL_6082;
  wire [31:0] _EVAL_5449;
  wire  _EVAL_5033;
  wire [31:0] _EVAL_294;
  wire  _EVAL_5037;
  wire  _EVAL_5905;
  wire [31:0] _EVAL_5206;
  wire [31:0] _EVAL_333;
  wire [31:0] _EVAL_6032;
  wire [31:0] _EVAL_3769;
  wire [31:0] _EVAL_5641;
  wire  _EVAL_3130;
  wire  _EVAL_3892;
  wire [31:0] _EVAL_3057;
  wire  _EVAL_5733;
  wire  _EVAL_1668;
  wire [31:0] _EVAL_3172;
  wire  _EVAL_5002;
  wire [31:0] _EVAL_1755;
  wire  _EVAL_4133;
  wire  _EVAL_1761;
  wire [31:0] _EVAL_4562;
  wire  _EVAL_5786;
  wire  _EVAL_4141;
  wire [31:0] _EVAL_4353;
  wire  _EVAL_4745;
  wire  _EVAL_4928;
  wire [31:0] _EVAL_530;
  wire [31:0] _EVAL_3637;
  wire [31:0] _EVAL_1506;
  wire  _EVAL_5719;
  wire  _EVAL_493;
  wire [31:0] _EVAL_2640;
  wire  _EVAL_4398;
  wire  _EVAL_375;
  wire [31:0] _EVAL_3458;
  wire  _EVAL_4685;
  wire [31:0] _EVAL_3706;
  wire [31:0] _EVAL_5720;
  wire  _EVAL_5790;
  wire [31:0] _EVAL_5283;
  wire  _EVAL_4382;
  wire [31:0] _EVAL_4601;
  wire  _EVAL_1250;
  wire  _EVAL_4696;
  wire [31:0] _EVAL_2392;
  wire  _EVAL_6054;
  wire  _EVAL_5000;
  wire [31:0] _EVAL_3984;
  wire  _EVAL_1576;
  wire  _EVAL_1840;
  wire [31:0] _EVAL_1200;
  wire  _EVAL_1607;
  wire  _EVAL_2639;
  wire [31:0] _EVAL_6129;
  wire  _EVAL_5834;
  wire  _EVAL_2900;
  wire  _EVAL_5863;
  wire  _EVAL_4089;
  wire  _EVAL_4558;
  wire  _EVAL_1437;
  wire  _EVAL_1696;
  wire  _EVAL_5885;
  wire  _EVAL_352;
  wire [31:0] _EVAL_5302;
  wire  _EVAL_827;
  wire [7:0] _EVAL_1269;
  wire  _EVAL_3854;
  wire  _EVAL_1920;
  wire  _EVAL_2129;
  wire  _EVAL_5993;
  wire [31:0] _EVAL_806;
  wire  _EVAL_1705;
  wire  _EVAL_781;
  wire  _EVAL_870;
  wire  _EVAL_2563;
  wire  _EVAL_3610;
  wire  _EVAL_3253;
  wire  _EVAL_1334;
  wire  _EVAL_3328;
  wire  _EVAL_1471;
  wire  _EVAL_2841;
  wire  _EVAL_2521;
  wire  _EVAL_4686;
  wire  _EVAL_3050;
  wire  _EVAL_668;
  wire  _EVAL_3937;
  wire  _EVAL_4570;
  wire  _EVAL_969;
  wire  _EVAL_4461;
  wire  _EVAL_5328;
  wire [31:0] _EVAL_1262;
  wire  _EVAL_4909;
  wire  _EVAL_1388;
  wire [31:0] _EVAL_3845;
  wire  _EVAL_4047;
  wire  _EVAL_2611;
  wire [31:0] _EVAL_3690;
  wire  _EVAL_2305;
  wire  _EVAL_1605;
  wire [31:0] _EVAL_2919;
  wire  _EVAL_2258;
  wire [31:0] _EVAL_4017;
  wire  _EVAL_2384;
  wire [31:0] _EVAL_3448;
  wire  _EVAL_1414;
  wire  _EVAL_1499;
  wire  _EVAL_295;
  wire  _EVAL_4816;
  wire [31:0] _EVAL_5469;
  wire  _EVAL_602;
  wire  _EVAL_905;
  wire [31:0] _EVAL_2102;
  wire  _EVAL_2346;
  wire  _EVAL_2625;
  wire [31:0] _EVAL_823;
  wire  _EVAL_1768;
  wire  _EVAL_2552;
  wire [31:0] _EVAL_1672;
  wire  _EVAL_4229;
  wire  _EVAL_1243;
  wire [31:0] _EVAL_3099;
  wire  _EVAL_1843;
  wire  _EVAL_4580;
  wire [31:0] _EVAL_4627;
  wire  _EVAL_5001;
  wire  _EVAL_999;
  wire [31:0] _EVAL_3472;
  wire  _EVAL_274;
  wire  _EVAL_2923;
  wire [31:0] _EVAL_5828;
  wire  _EVAL_4054;
  wire  _EVAL_4752;
  wire [31:0] _EVAL_924;
  wire  _EVAL_253;
  wire  _EVAL_2885;
  wire  _EVAL_1209;
  wire  _EVAL_5003;
  wire [31:0] _EVAL_4487;
  wire  _EVAL_466;
  wire  _EVAL_5649;
  wire  _EVAL_725;
  wire  _EVAL_2855;
  wire [31:0] _EVAL_4364;
  wire  _EVAL_879;
  wire  _EVAL_3245;
  wire [31:0] _EVAL_2719;
  wire  _EVAL_4769;
  wire  _EVAL_4529;
  wire [31:0] _EVAL_4744;
  wire  _EVAL_2181;
  wire  _EVAL_3885;
  wire [31:0] _EVAL_2328;
  wire  _EVAL_2762;
  wire  _EVAL_4893;
  wire [31:0] _EVAL_1653;
  wire  _EVAL_1988;
  wire  _EVAL_5981;
  wire [31:0] _EVAL_3386;
  wire  _EVAL_3136;
  wire [2:0] _EVAL_1984;
  wire [2:0] _EVAL_4908;
  wire [2:0] _EVAL_3849;
  wire [2:0] _EVAL_2514;
  wire [2:0] _EVAL_3125;
  wire [2:0] _EVAL_4634;
  wire [2:0] _EVAL_4698;
  wire [2:0] _EVAL_3351;
  wire [2:0] _EVAL_2112;
  wire [2:0] _EVAL_5617;
  wire [2:0] _EVAL_5842;
  wire [2:0] _EVAL_1622;
  wire [2:0] _EVAL_3513;
  wire [2:0] _EVAL_5806;
  wire [2:0] _EVAL_2151;
  wire [2:0] _EVAL_4798;
  wire [2:0] _EVAL_4608;
  wire [2:0] _EVAL_5935;
  wire [2:0] _EVAL_1977;
  wire [2:0] _EVAL_5858;
  wire [2:0] _EVAL_4722;
  wire [2:0] _EVAL_1486;
  wire [2:0] _EVAL_2656;
  wire [2:0] _EVAL_1363;
  wire [31:0] _EVAL_4262;
  wire  _EVAL_4309;
  wire [31:0] _EVAL_1179;
  wire  _EVAL_1475;
  wire  _EVAL_1297;
  wire [31:0] _EVAL_4126;
  wire  _EVAL_4329;
  wire  _EVAL_1040;
  wire [31:0] _EVAL_4932;
  wire  _EVAL_5331;
  wire [31:0] _EVAL_2427;
  wire  _EVAL_1450;
  wire  _EVAL_2566;
  wire [31:0] _EVAL_3468;
  wire  _EVAL_4770;
  wire  _EVAL_2120;
  wire [31:0] _EVAL_1921;
  wire  _EVAL_4617;
  wire [31:0] _EVAL_1703;
  wire  _EVAL_2433;
  wire  _EVAL_782;
  wire [31:0] _EVAL_456;
  wire  _EVAL_1739;
  wire  _EVAL_3207;
  wire  _EVAL_4266;
  wire  _EVAL_3224;
  wire  _EVAL_4733;
  wire [31:0] _EVAL_2027;
  wire [31:0] _EVAL_206;
  wire  _EVAL_2475;
  wire [31:0] _EVAL_4027;
  wire [31:0] _EVAL_2166;
  wire  _EVAL_2833;
  wire [31:0] _EVAL_4945;
  wire  _EVAL_6063;
  wire  _EVAL_4524;
  wire  _EVAL_407;
  wire [31:0] _EVAL_3344;
  wire  _EVAL_1698;
  wire [31:0] _EVAL_3432;
  wire  _EVAL_3308;
  wire  _EVAL_3932;
  wire  _EVAL_5168;
  wire [31:0] _EVAL_3203;
  wire  _EVAL_2247;
  wire  _EVAL_5597;
  wire  _EVAL_1337;
  wire  _EVAL_1333;
  wire  _EVAL_3198;
  wire  _EVAL_3170;
  wire [31:0] _EVAL_4370;
  wire  _EVAL_1412;
  wire [31:0] _EVAL_3179;
  wire  _EVAL_4546;
  wire  _EVAL_2282;
  wire [31:0] _EVAL_1874;
  wire  _EVAL_5204;
  wire  _EVAL_2261;
  wire [31:0] _EVAL_1496;
  wire  _EVAL_4507;
  wire [31:0] _EVAL_3204;
  wire  _EVAL_3640;
  wire  _EVAL_1857;
  wire [31:0] _EVAL_3301;
  wire  _EVAL_2428;
  wire  _EVAL_3541;
  wire  _EVAL_6133;
  wire [31:0] _EVAL_2626;
  wire  _EVAL_4061;
  wire [31:0] _EVAL_4023;
  wire  _EVAL_3212;
  wire  _EVAL_1146;
  wire  _EVAL_2649;
  wire  _EVAL_3727;
  wire [31:0] _EVAL_5902;
  wire  _EVAL_3517;
  wire  _EVAL_1172;
  wire [31:0] _EVAL_1000;
  wire  _EVAL_3896;
  wire  _EVAL_5779;
  wire [31:0] _EVAL_3824;
  wire  _EVAL_3305;
  wire  _EVAL_3879;
  wire [31:0] _EVAL_4181;
  wire  _EVAL_311;
  wire  _EVAL_1603;
  wire [31:0] _EVAL_4363;
  wire  _EVAL_3902;
  wire  _EVAL_2302;
  wire [31:0] _EVAL_5881;
  wire  _EVAL_5677;
  wire  _EVAL_561;
  wire [31:0] _EVAL_1149;
  wire  _EVAL_4838;
  wire [31:0] _EVAL_5796;
  wire  _EVAL_1287;
  wire  _EVAL_5758;
  wire [31:0] _EVAL_4344;
  wire  _EVAL_2301;
  wire  _EVAL_4760;
  wire [31:0] _EVAL_3446;
  wire  _EVAL_831;
  wire  _EVAL_3730;
  wire [31:0] _EVAL_2876;
  wire  _EVAL_3617;
  wire  _EVAL_2284;
  wire [31:0] _EVAL_2583;
  wire  _EVAL_3557;
  wire [31:0] _EVAL_1719;
  wire  _EVAL_4839;
  wire  _EVAL_2091;
  wire [31:0] _EVAL_2794;
  wire  _EVAL_4166;
  wire  _EVAL_509;
  wire [31:0] _EVAL_2297;
  wire  _EVAL_2932;
  wire  _EVAL_2312;
  wire [31:0] _EVAL_1153;
  wire  _EVAL_3895;
  wire  _EVAL_5082;
  wire  _EVAL_5252;
  wire  _EVAL_1922;
  wire  _EVAL_4632;
  wire  _EVAL_4356;
  wire [31:0] _EVAL_188;
  wire  _EVAL_4822;
  wire [31:0] _EVAL_4387;
  wire  _EVAL_3764;
  wire  _EVAL_3465;
  wire  _EVAL_2104;
  wire  _EVAL_3847;
  wire  _EVAL_3726;
  wire [31:0] _EVAL_1212;
  wire  _EVAL_3027;
  wire  _EVAL_2326;
  wire [4:0] _EVAL_5057;
  wire  _EVAL_4574;
  wire  _EVAL_842;
  wire  _EVAL_1120;
  wire  _EVAL_2370;
  wire  _EVAL_2115;
  wire [31:0] _EVAL_1567;
  wire  _EVAL_1504;
  wire  _EVAL_5500;
  wire [31:0] _EVAL_1282;
  wire  _EVAL_4550;
  wire  _EVAL_4026;
  wire [31:0] _EVAL_5732;
  wire  _EVAL_2441;
  wire  _EVAL_807;
  wire [31:0] _EVAL_3520;
  wire  _EVAL_754;
  wire  _EVAL_1915;
  wire [31:0] _EVAL_1925;
  wire  _EVAL_1729;
  wire  _EVAL_2056;
  wire [31:0] _EVAL_5354;
  wire  _EVAL_3559;
  wire  _EVAL_6005;
  wire  _EVAL_3978;
  wire  _EVAL_4041;
  wire  _EVAL_1899;
  wire [7:0] _EVAL_632;
  wire  _EVAL_5213;
  wire  _EVAL_1684;
  wire  _EVAL_250;
  wire  _EVAL_4242;
  wire  _EVAL_5693;
  wire  _EVAL_5178;
  wire  _EVAL_1564;
  wire  _EVAL_1825;
  wire  _EVAL_1601;
  wire [31:0] _EVAL_1571;
  wire  _EVAL_4458;
  wire  _EVAL_5402;
  wire  _EVAL_3142;
  wire [31:0] _EVAL_457;
  wire  _EVAL_2487;
  wire  _EVAL_972;
  wire [31:0] _EVAL_4553;
  wire  _EVAL_1997;
  wire  _EVAL_898;
  wire [31:0] _EVAL_5196;
  wire  _EVAL_5448;
  wire  _EVAL_5075;
  wire [31:0] _EVAL_2084;
  wire  _EVAL_1979;
  wire  _EVAL_2467;
  wire [31:0] _EVAL_2904;
  wire  _EVAL_6021;
  wire  _EVAL_4436;
  wire [31:0] _EVAL_2347;
  wire  _EVAL_1894;
  wire  _EVAL_1411;
  wire [31:0] _EVAL_2232;
  wire  _EVAL_1439;
  wire  _EVAL_1423;
  wire [31:0] _EVAL_5071;
  wire  _EVAL_875;
  wire  _EVAL_1849;
  wire [31:0] _EVAL_3580;
  wire  _EVAL_6038;
  wire  _EVAL_5625;
  wire [31:0] _EVAL_3101;
  wire  _EVAL_3578;
  wire  _EVAL_3702;
  wire  _EVAL_1549;
  wire  _EVAL_2554;
  wire [31:0] _EVAL_3360;
  wire  _EVAL_3750;
  wire  _EVAL_2846;
  wire  _EVAL_1016;
  wire  _EVAL_4537;
  wire [31:0] _EVAL_5632;
  wire  _EVAL_6139;
  wire  _EVAL_4081;
  wire [31:0] _EVAL_2332;
  wire  _EVAL_3903;
  wire  _EVAL_5017;
  wire [31:0] _EVAL_1788;
  wire  _EVAL_4014;
  wire  _EVAL_1581;
  wire [31:0] _EVAL_3999;
  wire  _EVAL_4717;
  wire  _EVAL_820;
  wire [31:0] _EVAL_874;
  wire  _EVAL_4763;
  wire  _EVAL_1798;
  wire [31:0] _EVAL_494;
  wire  _EVAL_1929;
  wire  _EVAL_4153;
  wire [31:0] _EVAL_1331;
  wire  _EVAL_1249;
  wire  _EVAL_4037;
  wire  _EVAL_4418;
  wire  _EVAL_5064;
  wire [31:0] _EVAL_4119;
  wire  _EVAL_1721;
  wire  _EVAL_903;
  wire  _EVAL_1394;
  wire  _EVAL_3233;
  wire [31:0] _EVAL_3749;
  wire  _EVAL_3965;
  wire  _EVAL_3622;
  wire [31:0] _EVAL_1557;
  wire  _EVAL_3662;
  wire  _EVAL_3275;
  wire [31:0] _EVAL_5555;
  wire  _EVAL_5692;
  wire  _EVAL_5163;
  wire  _EVAL_1953;
  wire  _EVAL_2009;
  wire  _EVAL_560;
  wire  _EVAL_5816;
  wire [31:0] _EVAL_2579;
  wire  _EVAL_2222;
  wire  _EVAL_3543;
  wire [31:0] _EVAL_5401;
  wire  _EVAL_5958;
  wire  _EVAL_4911;
  wire  _EVAL_3090;
  wire  _EVAL_1751;
  wire  _EVAL_5894;
  wire [31:0] _EVAL_520;
  wire  _EVAL_1990;
  wire  _EVAL_320;
  wire  _EVAL_4289;
  wire  _EVAL_1881;
  wire  _EVAL_1175;
  wire  _EVAL_6050;
  wire [31:0] _EVAL_5729;
  wire  _EVAL_656;
  wire [11:0] _EVAL_805;
  wire  _EVAL_6046;
  wire  _EVAL_2609;
  wire  _EVAL_1142;
  wire  _EVAL_640;
  wire  _EVAL_3355;
  wire  _EVAL_800;
  wire  _EVAL_5563;
  wire [31:0] _EVAL_4687;
  wire  _EVAL_576;
  wire [31:0] _EVAL_4937;
  wire  _EVAL_5812;
  wire  _EVAL_1532;
  wire  _EVAL_4592;
  wire  _EVAL_4641;
  wire [31:0] _EVAL_1718;
  wire  _EVAL_4001;
  wire  _EVAL_5697;
  wire [31:0] _EVAL_2654;
  wire  _EVAL_776;
  wire  _EVAL_562;
  wire  _EVAL_2017;
  wire  _EVAL_1366;
  wire [31:0] _EVAL_3418;
  wire  _EVAL_5568;
  wire  _EVAL_5453;
  wire  _EVAL_4306;
  wire [31:0] _EVAL_865;
  wire  _EVAL_3781;
  wire  _EVAL_164;
  wire  _EVAL_5548;
  wire [31:0] _EVAL_4427;
  wire  _EVAL_5478;
  wire  _EVAL_963;
  wire [31:0] _EVAL_1035;
  wire  _EVAL_4661;
  wire  _EVAL_2880;
  wire [31:0] _EVAL_5857;
  wire  _EVAL_2106;
  wire [31:0] _EVAL_3338;
  wire  _EVAL_5829;
  wire  _EVAL_2170;
  wire  _EVAL_1789;
  wire [31:0] _EVAL_1614;
  wire  _EVAL_4070;
  wire  _EVAL_1994;
  wire [31:0] _EVAL_1113;
  wire  _EVAL_1967;
  wire  _EVAL_810;
  wire  _EVAL_5208;
  wire  _EVAL_5909;
  wire  _EVAL_1982;
  wire  _EVAL_1325;
  wire  _EVAL_3623;
  wire [31:0] _EVAL_4542;
  wire  _EVAL_1876;
  wire [31:0] _EVAL_5109;
  wire  _EVAL_1816;
  wire  _EVAL_3285;
  wire [31:0] _EVAL_544;
  wire  _EVAL_1811;
  wire  _EVAL_4480;
  wire [31:0] _EVAL_6096;
  wire  _EVAL_1382;
  wire  _EVAL_1381;
  wire [31:0] _EVAL_5314;
  wire  _EVAL_3149;
  wire  _EVAL_2289;
  wire [31:0] _EVAL_5195;
  wire  _EVAL_5794;
  wire  _EVAL_3315;
  wire [31:0] _EVAL_4740;
  wire  _EVAL_3579;
  wire  _EVAL_1780;
  wire [31:0] _EVAL_1600;
  wire  _EVAL_214;
  wire  _EVAL_1026;
  wire [31:0] _EVAL_501;
  wire  _EVAL_5817;
  wire  _EVAL_3908;
  wire [31:0] _EVAL_1951;
  wire  _EVAL_1795;
  wire  _EVAL_3228;
  wire [31:0] _EVAL_5065;
  wire  _EVAL_703;
  wire  _EVAL_1535;
  wire [31:0] _EVAL_3306;
  wire  _EVAL_5007;
  wire  _EVAL_3187;
  wire  _EVAL_1123;
  wire  _EVAL_2262;
  wire [31:0] _EVAL_4078;
  wire  _EVAL_1812;
  wire  _EVAL_4926;
  wire  _EVAL_5511;
  wire  _EVAL_3837;
  wire [31:0] _EVAL_4042;
  wire  _EVAL_2665;
  wire  _EVAL_2182;
  wire [31:0] _EVAL_4385;
  wire  _EVAL_2292;
  wire  _EVAL_3738;
  wire [31:0] _EVAL_4080;
  wire  _EVAL_1246;
  wire  _EVAL_1892;
  wire [31:0] _EVAL_2987;
  wire  _EVAL_2006;
  wire  _EVAL_1980;
  wire [3:0] _EVAL_2250;
  wire [2:0] _EVAL_3461;
  wire [1:0] _EVAL_919;
  wire [1:0] _EVAL_4832;
  wire [1:0] _EVAL_2822;
  wire [2:0] _EVAL_858;
  wire [31:0] _EVAL_3083;
  wire  _EVAL_4088;
  wire [3:0] _EVAL_2260;
  wire  _EVAL_4577;
  wire  _EVAL_5600;
  wire  _EVAL_2086;
  wire  _EVAL_5417;
  wire  _EVAL_1904;
  wire  _EVAL_1114;
  wire  _EVAL_5217;
  wire  _EVAL_4758;
  wire  _EVAL_964;
  wire  _EVAL_5918;
  wire  _EVAL_2526;
  wire  _EVAL_3544;
  wire  _EVAL_5298;
  wire  _EVAL_2245;
  wire  _EVAL_965;
  wire  _EVAL_3376;
  wire  _EVAL_2645;
  wire  _EVAL_4879;
  wire [3:0] _EVAL_1330;
  wire  _EVAL_5788;
  wire  _EVAL_1299;
  wire  _EVAL_2956;
  wire  _EVAL_3196;
  wire [3:0] _EVAL_1809;
  wire [3:0] _EVAL_2031;
  wire [3:0] _EVAL_4375;
  wire [3:0] _EVAL_4170;
  wire [3:0] _EVAL_4984;
  wire [3:0] _EVAL_5671;
  wire  _EVAL_5588;
  wire  _EVAL_4426;
  wire [31:0] _EVAL_4087;
  wire [6:0] _EVAL_5282;
  wire [31:0] _EVAL_515;
  wire  _EVAL_5631;
  wire [31:0] _EVAL_4741;
  wire  _EVAL_6023;
  wire  _EVAL_2602;
  wire  _EVAL_6016;
  wire  _EVAL_590;
  wire [31:0] _EVAL_292;
  wire [31:0] _EVAL_2387;
  wire  _EVAL_5882;
  wire [31:0] _EVAL_3186;
  wire  _EVAL_161;
  wire [31:0] _EVAL_4066;
  wire  _EVAL_989;
  wire  _EVAL_4175;
  wire [31:0] _EVAL_3247;
  wire  _EVAL_2693;
  wire  _EVAL_1129;
  wire [31:0] _EVAL_5166;
  wire  _EVAL_310;
  wire  _EVAL_961;
  wire [31:0] _EVAL_2206;
  wire  _EVAL_2264;
  wire  _EVAL_223;
  wire [31:0] _EVAL_3612;
  wire  _EVAL_2584;
  wire  _EVAL_3327;
  wire [31:0] _EVAL_5376;
  wire  _EVAL_1409;
  wire  _EVAL_5512;
  wire [31:0] _EVAL_2773;
  wire  _EVAL_1888;
  wire  _EVAL_1617;
  wire [31:0] _EVAL_678;
  wire  _EVAL_3281;
  wire  _EVAL_3284;
  wire [31:0] _EVAL_6010;
  wire  _EVAL_1837;
  wire  _EVAL_5835;
  wire  _EVAL_2249;
  wire  _EVAL_3333;
  wire [31:0] _EVAL_5197;
  wire  _EVAL_3147;
  wire  _EVAL_1734;
  wire  _EVAL_1611;
  wire  _EVAL_3393;
  wire [31:0] _EVAL_408;
  wire  _EVAL_3695;
  wire  _EVAL_783;
  wire  _EVAL_1474;
  wire  _EVAL_1949;
  wire  _EVAL_5717;
  wire [31:0] _EVAL_6121;
  wire  _EVAL_2542;
  wire  _EVAL_2948;
  wire [31:0] _EVAL_3930;
  wire  _EVAL_3995;
  wire  _EVAL_750;
  wire [31:0] _EVAL_5209;
  wire  _EVAL_420;
  wire  _EVAL_1082;
  wire [31:0] _EVAL_1993;
  wire  _EVAL_3454;
  wire  _EVAL_1216;
  wire  _EVAL_2401;
  wire  _EVAL_1245;
  wire [31:0] _EVAL_1502;
  wire  _EVAL_2077;
  wire  _EVAL_2750;
  wire  _EVAL_5351;
  wire  _EVAL_2972;
  wire [31:0] _EVAL_981;
  wire  _EVAL_3667;
  wire  _EVAL_6008;
  wire  _EVAL_1030;
  wire  _EVAL_4201;
  wire [31:0] _EVAL_2891;
  wire  _EVAL_3673;
  wire [31:0] _EVAL_4581;
  wire  _EVAL_2999;
  wire  _EVAL_5063;
  wire [31:0] _EVAL_1656;
  wire  _EVAL_3707;
  wire  _EVAL_3363;
  wire [31:0] _EVAL_3202;
  wire  _EVAL_670;
  wire  _EVAL_3459;
  wire [31:0] _EVAL_3168;
  wire [31:0] _EVAL_219;
  wire [31:0] _EVAL_1023;
  wire  _EVAL_2008;
  wire [31:0] _EVAL_3682;
  wire  _EVAL_5567;
  wire [31:0] _EVAL_1645;
  wire  _EVAL_1688;
  wire  _EVAL_4483;
  wire [31:0] _EVAL_3163;
  wire [31:0] _EVAL_4642;
  wire  _EVAL_1284;
  wire  _EVAL_5667;
  wire [31:0] _EVAL_5847;
  wire [31:0] _EVAL_6123;
  wire  _EVAL_1917;
  wire [31:0] _EVAL_587;
  wire  _EVAL_4640;
  wire  _EVAL_3691;
  wire [31:0] _EVAL_2909;
  wire  _EVAL_4525;
  wire  _EVAL_4670;
  wire [31:0] _EVAL_3759;
  wire  _EVAL_1032;
  wire [31:0] _EVAL_3068;
  wire  _EVAL_5339;
  wire  _EVAL_3037;
  wire [31:0] _EVAL_1440;
  wire  _EVAL_4457;
  wire  _EVAL_4072;
  wire  _EVAL_3611;
  wire  _EVAL_4161;
  wire  _EVAL_2856;
  wire [31:0] _EVAL_5795;
  wire [31:0] _EVAL_2253;
  wire  _EVAL_1716;
  wire [31:0] _EVAL_4825;
  wire  _EVAL_2973;
  wire [31:0] _EVAL_2647;
  wire  _EVAL_4316;
  wire  _EVAL_5285;
  wire [31:0] _EVAL_2955;
  wire  _EVAL_5011;
  wire  _EVAL_4974;
  wire [31:0] _EVAL_3480;
  wire  _EVAL_4853;
  wire [31:0] _EVAL_4963;
  wire  _EVAL_3131;
  wire  _EVAL_2816;
  wire [31:0] _EVAL_2610;
  wire [31:0] _EVAL_3875;
  wire  _EVAL_5102;
  wire  _EVAL_5318;
  wire [31:0] _EVAL_2079;
  wire  _EVAL_4500;
  wire  _EVAL_4499;
  wire [31:0] _EVAL_845;
  wire  _EVAL_580;
  wire  _EVAL_2404;
  wire [31:0] _EVAL_5565;
  wire  _EVAL_2335;
  wire [31:0] _EVAL_608;
  wire  _EVAL_682;
  wire [4:0] _EVAL_2786;
  wire [4:0] _EVAL_2745;
  wire [4:0] _EVAL_3449;
  wire [4:0] _EVAL_897;
  wire [4:0] _EVAL_2511;
  wire [4:0] _EVAL_5080;
  wire [4:0] _EVAL_3929;
  wire [4:0] _EVAL_5607;
  wire [4:0] _EVAL_3882;
  wire [4:0] _EVAL_5734;
  wire [4:0] _EVAL_4781;
  wire [4:0] _EVAL_2958;
  wire [4:0] _EVAL_5295;
  wire [4:0] _EVAL_1093;
  wire [4:0] _EVAL_4800;
  wire [4:0] _EVAL_4753;
  wire [4:0] _EVAL_3340;
  wire [4:0] _EVAL_1907;
  wire [4:0] _EVAL_1296;
  wire [4:0] _EVAL_5577;
  wire [4:0] _EVAL_1431;
  wire [4:0] _EVAL_627;
  wire [4:0] _EVAL_308;
  wire [4:0] _EVAL_531;
  wire [4:0] _EVAL_945;
  wire [4:0] _EVAL_3026;
  wire [4:0] _EVAL_3857;
  wire [4:0] _EVAL_285;
  wire [4:0] _EVAL_458;
  wire [4:0] _EVAL_5797;
  wire [4:0] _EVAL_5226;
  wire [4:0] _EVAL_4180;
  wire [4:0] _EVAL_3983;
  wire [31:0] _EVAL_1465;
  wire  _EVAL_5442;
  wire [31:0] _EVAL_1723;
  wire  _EVAL_3656;
  wire  _EVAL_5255;
  wire  _EVAL_1004;
  wire  _EVAL_6055;
  wire  _EVAL_1081;
  wire  _EVAL_1630;
  wire  _EVAL_2510;
  wire  _EVAL_3508;
  wire  _EVAL_3950;
  wire  _EVAL_183;
  wire  _EVAL_5841;
  wire  _EVAL_5136;
  wire  _EVAL_4573;
  wire  _EVAL_4294;
  wire  _EVAL_1903;
  wire  _EVAL_2594;
  wire  _EVAL_5140;
  wire  _EVAL_283;
  wire  _EVAL_239;
  wire  _EVAL_4880;
  wire  _EVAL_5583;
  wire  _EVAL_5473;
  wire [3:0] _EVAL_2385;
  wire [3:0] _EVAL_3012;
  wire [31:0] _EVAL_2394;
  wire [31:0] _EVAL_4044;
  wire  _EVAL_5480;
  wire [31:0] _EVAL_1897;
  wire  _EVAL_5933;
  wire  _EVAL_4734;
  wire [31:0] _EVAL_224;
  wire  _EVAL_2596;
  wire  _EVAL_4836;
  wire [4:0] _EVAL_2839;
  wire [31:0] _EVAL_3396;
  wire  _EVAL_1267;
  wire [31:0] _EVAL_2470;
  wire  _EVAL_1606;
  wire [31:0] _EVAL_4677;
  wire  _EVAL_675;
  wire  _EVAL_2911;
  wire [31:0] _EVAL_1582;
  wire  _EVAL_290;
  wire  _EVAL_4625;
  wire [31:0] _EVAL_5158;
  wire  _EVAL_1553;
  wire  _EVAL_3137;
  wire  _EVAL_1415;
  wire [31:0] _EVAL_388;
  wire  _EVAL_5540;
  wire [31:0] _EVAL_3295;
  wire  _EVAL_5188;
  wire [31:0] _EVAL_4402;
  wire [31:0] _EVAL_2653;
  wire  _EVAL_4225;
  wire [31:0] _EVAL_4662;
  wire  _EVAL_4868;
  wire  _EVAL_598;
  wire [31:0] _EVAL_498;
  wire  _EVAL_4134;
  wire  _EVAL_3583;
  wire  _EVAL_959;
  wire [31:0] _EVAL_2228;
  wire  _EVAL_2540;
  wire  _EVAL_5156;
  wire [31:0] _EVAL_5408;
  wire  _EVAL_2323;
  wire  _EVAL_3081;
  wire [4:0] _EVAL_1592;
  wire [4:0] _EVAL_181;
  wire [31:0] _EVAL_2311;
  wire [31:0] _EVAL_2479;
  wire [31:0] _EVAL_286;
  wire [31:0] _EVAL_3942;
  wire  _EVAL_3482;
  wire [31:0] _EVAL_3898;
  wire  _EVAL_2455;
  wire  _EVAL_884;
  wire  _EVAL_4248;
  wire [31:0] _EVAL_2702;
  wire  _EVAL_3564;
  wire [31:0] _EVAL_3842;
  wire  _EVAL_2236;
  wire  _EVAL_1661;
  wire  _EVAL_2798;
  wire  _EVAL_4969;
  wire [31:0] _EVAL_4290;
  wire  _EVAL_778;
  wire  _EVAL_4332;
  wire [31:0] _EVAL_1446;
  wire  _EVAL_5229;
  wire [31:0] _EVAL_4960;
  wire  _EVAL_1524;
  wire [31:0] _EVAL_4674;
  wire  _EVAL_1891;
  wire  _EVAL_4278;
  wire [31:0] _EVAL_451;
  wire  _EVAL_5988;
  wire  _EVAL_3009;
  wire [31:0] _EVAL_2088;
  wire  _EVAL_4683;
  wire  _EVAL_1071;
  wire [31:0] _EVAL_2708;
  wire  _EVAL_2033;
  wire  _EVAL_3809;
  wire [31:0] _EVAL_4910;
  wire  _EVAL_3486;
  wire  _EVAL_2907;
  wire [31:0] _EVAL_1312;
  wire  _EVAL_5946;
  wire  _EVAL_789;
  wire  _EVAL_3886;
  wire  _EVAL_5382;
  wire [31:0] _EVAL_429;
  wire  _EVAL_2888;
  wire  _EVAL_5260;
  wire [31:0] _EVAL_6101;
  wire  _EVAL_3060;
  wire  _EVAL_3586;
  wire [31:0] _EVAL_2316;
  wire  _EVAL_5116;
  wire  _EVAL_2533;
  wire  _EVAL_4628;
  wire  _EVAL_2489;
  wire  _EVAL_5544;
  wire  _EVAL_6110;
  wire  _EVAL_1053;
  wire [31:0] _EVAL_3034;
  wire  _EVAL_1814;
  wire  _EVAL_4018;
  wire [31:0] _EVAL_6130;
  wire  _EVAL_2421;
  wire  _EVAL_4559;
  wire [31:0] _EVAL_2138;
  wire  _EVAL_5470;
  wire  _EVAL_5895;
  wire [31:0] _EVAL_1938;
  wire  _EVAL_2118;
  wire  _EVAL_1214;
  wire [31:0] _EVAL_437;
  wire  _EVAL_3346;
  wire  _EVAL_1202;
  wire [31:0] _EVAL_5879;
  wire  _EVAL_1400;
  wire  _EVAL_5929;
  wire [31:0] _EVAL_1218;
  wire  _EVAL_3777;
  wire  _EVAL_5643;
  wire  _EVAL_3152;
  wire  _EVAL_1463;
  wire  _EVAL_5049;
  wire  _EVAL_3924;
  wire  _EVAL_2580;
  wire  _EVAL_657;
  wire  _EVAL_4108;
  wire [31:0] _EVAL_1543;
  wire  _EVAL_1107;
  wire [31:0] _EVAL_5380;
  wire  _EVAL_4288;
  wire [31:0] _EVAL_4471;
  wire  _EVAL_5272;
  wire  _EVAL_3008;
  wire [31:0] _EVAL_3086;
  wire  _EVAL_5419;
  wire  _EVAL_1577;
  wire [31:0] _EVAL_1793;
  wire  _EVAL_4367;
  wire  _EVAL_2538;
  wire [31:0] _EVAL_3231;
  wire  _EVAL_4714;
  wire [31:0] _EVAL_4925;
  wire  _EVAL_1072;
  wire  _EVAL_838;
  wire  _EVAL_3238;
  wire [31:0] _EVAL_591;
  wire [31:0] _EVAL_5466;
  wire  _EVAL_2309;
  wire  _EVAL_3783;
  wire [31:0] _EVAL_549;
  wire  _EVAL_5262;
  wire  _EVAL_4712;
  wire [31:0] _EVAL_1631;
  wire  _EVAL_2061;
  wire  _EVAL_4783;
  wire [31:0] _EVAL_5814;
  wire  _EVAL_5451;
  wire  _EVAL_182;
  wire  _EVAL_946;
  wire  _EVAL_393;
  wire  _EVAL_4109;
  wire  _EVAL_1063;
  wire  _EVAL_1810;
  wire  _EVAL_3069;
  wire  _EVAL_4410;
  wire  _EVAL_3077;
  wire [31:0] _EVAL_4701;
  wire  _EVAL_4756;
  wire  _EVAL_2667;
  wire  _EVAL_3268;
  wire  _EVAL_1019;
  wire [31:0] _EVAL_2582;
  wire  _EVAL_1717;
  wire  _EVAL_2735;
  wire [31:0] _EVAL_2826;
  wire  _EVAL_4948;
  wire  _EVAL_558;
  wire [31:0] _EVAL_5538;
  wire  _EVAL_299;
  wire  _EVAL_2400;
  wire  _EVAL_4506;
  wire  _EVAL_4918;
  wire  _EVAL_2349;
  wire [31:0] _EVAL_1875;
  wire  _EVAL_1273;
  wire  _EVAL_2857;
  wire  _EVAL_2899;
  wire  _EVAL_3457;
  wire [31:0] _EVAL_2055;
  wire  _EVAL_3516;
  wire  _EVAL_5727;
  wire [31:0] _EVAL_3024;
  wire  _EVAL_3775;
  wire  _EVAL_2840;
  wire [31:0] _EVAL_5405;
  wire  _EVAL_2512;
  wire  _EVAL_2099;
  wire  _EVAL_3948;
  wire  _EVAL_3279;
  wire [31:0] _EVAL_1736;
  wire  _EVAL_1534;
  wire  _EVAL_3943;
  wire  _EVAL_3017;
  wire  _EVAL_438;
  wire [31:0] _EVAL_1469;
  wire  _EVAL_4526;
  wire  _EVAL_163;
  wire  _EVAL_3760;
  wire  _EVAL_4854;
  wire [31:0] _EVAL_5608;
  wire  _EVAL_331;
  wire  _EVAL_6092;
  wire [31:0] _EVAL_5277;
  wire  _EVAL_3576;
  wire  _EVAL_2023;
  wire  _EVAL_5347;
  wire  _EVAL_1775;
  wire [31:0] _EVAL_474;
  wire  _EVAL_2066;
  wire  _EVAL_3028;
  wire [31:0] _EVAL_4392;
  wire  _EVAL_4891;
  wire  _EVAL_2501;
  wire  _EVAL_3831;
  wire  _EVAL_4303;
  wire [31:0] _EVAL_3596;
  wire  _EVAL_5556;
  wire  _EVAL_3803;
  wire  _EVAL_4117;
  wire  _EVAL_366;
  wire [31:0] _EVAL_2522;
  wire  _EVAL_795;
  wire  _EVAL_2960;
  wire  _EVAL_2189;
  wire  _EVAL_4678;
  wire [31:0] _EVAL_1467;
  wire  _EVAL_2599;
  wire  _EVAL_6044;
  wire [31:0] _EVAL_1792;
  wire  _EVAL_3425;
  wire  _EVAL_251;
  wire [31:0] _EVAL_6043;
  wire  _EVAL_3165;
  wire  _EVAL_4995;
  wire [31:0] _EVAL_1452;
  wire  _EVAL_5036;
  wire  _EVAL_6073;
  wire  _EVAL_944;
  wire [31:0] _EVAL_2544;
  wire  _EVAL_5934;
  wire  _EVAL_2481;
  wire  _EVAL_665;
  wire  _EVAL_3627;
  wire  _EVAL_2454;
  wire  _EVAL_5296;
  wire [7:0] _EVAL_3830;
  wire  _EVAL_2092;
  wire  _EVAL_2635;
  wire  _EVAL_2408;
  wire  _EVAL_3371;
  wire  _EVAL_5100;
  wire  _EVAL_1193;
  wire  _EVAL_3671;
  wire  _EVAL_2453;
  wire  _EVAL_2425;
  wire [31:0] _EVAL_6056;
  wire  _EVAL_4003;
  wire  _EVAL_4082;
  wire [31:0] _EVAL_2149;
  wire  _EVAL_696;
  wire  _EVAL_1039;
  wire  _EVAL_658;
  wire  _EVAL_2171;
  wire [31:0] _EVAL_5762;
  wire  _EVAL_6124;
  wire  _EVAL_3058;
  wire  _EVAL_825;
  wire  _EVAL_5508;
  wire  _EVAL_4780;
  wire  _EVAL_4446;
  wire  _EVAL_4284;
  wire  _EVAL_4147;
  wire  _EVAL_4296;
  wire [31:0] _EVAL_2971;
  wire  _EVAL_5083;
  wire  _EVAL_1494;
  wire [31:0] _EVAL_2137;
  wire  _EVAL_3582;
  wire  _EVAL_3365;
  wire  _EVAL_1125;
  wire  _EVAL_2432;
  wire [31:0] _EVAL_5799;
  wire  _EVAL_4814;
  wire [31:0] _EVAL_4747;
  wire  _EVAL_6013;
  wire  _EVAL_753;
  wire  _EVAL_1821;
  wire  _EVAL_2180;
  wire  _EVAL_276;
  wire [31:0] _EVAL_4212;
  wire  _EVAL_1834;
  wire  _EVAL_2492;
  wire [31:0] _EVAL_1569;
  wire  _EVAL_733;
  wire  _EVAL_1676;
  wire [31:0] _EVAL_4405;
  wire  _EVAL_720;
  wire  _EVAL_4502;
  wire [31:0] _EVAL_433;
  wire  _EVAL_3162;
  wire  _EVAL_4962;
  wire [31:0] _EVAL_1787;
  wire  _EVAL_3765;
  wire  _EVAL_1389;
  wire [31:0] _EVAL_5866;
  wire  _EVAL_3120;
  wire  _EVAL_3109;
  wire [31:0] _EVAL_2306;
  wire  _EVAL_1987;
  wire  _EVAL_1379;
  wire  _EVAL_5246;
  wire  _EVAL_1155;
  wire  _EVAL_5139;
  wire [31:0] _EVAL_2098;
  wire  _EVAL_5185;
  wire  _EVAL_5662;
  wire  _EVAL_5499;
  wire  _EVAL_4207;
  wire  _EVAL_4746;
  wire  _EVAL_2643;
  wire [31:0] _EVAL_2082;
  wire  _EVAL_1227;
  wire  _EVAL_3005;
  wire [31:0] _EVAL_2992;
  wire  _EVAL_3779;
  wire  _EVAL_734;
  wire [31:0] _EVAL_3776;
  wire  _EVAL_1251;
  wire  _EVAL_1207;
  wire [31:0] _EVAL_1108;
  wire  _EVAL_1965;
  wire  _EVAL_1293;
  wire [31:0] _EVAL_934;
  wire  _EVAL_3497;
  wire  _EVAL_1432;
  wire [31:0] _EVAL_4285;
  wire  _EVAL_3634;
  wire  _EVAL_1744;
  wire  _EVAL_6066;
  wire  _EVAL_900;
  wire  _EVAL_5160;
  wire  _EVAL_4954;
  wire  _EVAL_1305;
  wire [31:0] _EVAL_2659;
  wire  _EVAL_4336;
  wire  _EVAL_4160;
  wire  _EVAL_5181;
  wire  _EVAL_3354;
  wire  _EVAL_3504;
  wire  _EVAL_4637;
  wire [31:0] _EVAL_1060;
  wire  _EVAL_5522;
  wire  _EVAL_3888;
  wire  _EVAL_3933;
  wire  _EVAL_1067;
  wire [31:0] _EVAL_2733;
  wire  _EVAL_5502;
  wire  _EVAL_3225;
  wire  _EVAL_2842;
  wire  _EVAL_3381;
  wire  _EVAL_5050;
  wire  _EVAL_2100;
  wire  _EVAL_3699;
  wire  _EVAL_3747;
  wire  _EVAL_5264;
  wire  _EVAL_5523;
  wire  _EVAL_3397;
  wire [31:0] _EVAL_5172;
  wire  _EVAL_215;
  wire  _EVAL_2046;
  wire [31:0] _EVAL_3709;
  wire  _EVAL_5887;
  wire  _EVAL_1192;
  wire [31:0] _EVAL_4699;
  wire  _EVAL_5610;
  wire  _EVAL_4767;
  wire [31:0] _EVAL_1485;
  wire  _EVAL_2734;
  wire  _EVAL_4030;
  wire  _EVAL_5653;
  wire [31:0] _EVAL_3797;
  wire  _EVAL_5301;
  wire  _EVAL_5868;
  wire [31:0] _EVAL_4631;
  wire  _EVAL_2675;
  wire  _EVAL_5137;
  wire  _EVAL_338;
  wire  _EVAL_766;
  wire  _EVAL_756;
  wire  _EVAL_5294;
  wire  _EVAL_5319;
  wire  _EVAL_2403;
  wire  _EVAL_6030;
  wire [31:0] _EVAL_228;
  wire  _EVAL_2616;
  wire  _EVAL_2807;
  wire [31:0] _EVAL_1640;
  wire  _EVAL_4317;
  wire  _EVAL_3267;
  wire [31:0] _EVAL_2068;
  wire  _EVAL_2701;
  wire  _EVAL_2285;
  wire [31:0] _EVAL_2270;
  wire  _EVAL_1141;
  wire  _EVAL_4803;
  wire [31:0] _EVAL_1349;
  wire  _EVAL_557;
  wire  _EVAL_4417;
  wire [31:0] _EVAL_4833;
  wire  _EVAL_4040;
  wire  _EVAL_1911;
  wire [31:0] _EVAL_2237;
  wire  _EVAL_296;
  wire  _EVAL_2804;
  wire  _EVAL_2676;
  wire  _EVAL_3921;
  wire [10:0] _EVAL_4924;
  wire  _EVAL_4075;
  wire  _EVAL_3766;
  wire  _EVAL_288;
  wire  _EVAL_1369;
  wire  _EVAL_563;
  wire  _EVAL_3774;
  wire  _EVAL_1122;
  wire  _EVAL_843;
  wire [31:0] _EVAL_2870;
  wire  _EVAL_1677;
  wire  _EVAL_5595;
  wire  _EVAL_4988;
  wire [31:0] _EVAL_613;
  wire  _EVAL_4590;
  wire  _EVAL_3089;
  wire [31:0] _EVAL_1225;
  wire  _EVAL_1352;
  wire  _EVAL_413;
  wire [31:0] _EVAL_3462;
  wire  _EVAL_839;
  wire  _EVAL_3772;
  wire [31:0] _EVAL_3075;
  wire  _EVAL_3501;
  wire  _EVAL_1090;
  wire [31:0] _EVAL_403;
  wire  _EVAL_906;
  wire  _EVAL_5026;
  wire  _EVAL_5254;
  wire  _EVAL_3721;
  wire  _EVAL_1089;
  wire  _EVAL_2674;
  wire [31:0] _EVAL_4993;
  wire  _EVAL_211;
  wire  _EVAL_1461;
  wire [31:0] _EVAL_770;
  wire  _EVAL_4871;
  wire  _EVAL_1948;
  wire [31:0] _EVAL_3441;
  wire  _EVAL_2379;
  wire  _EVAL_2921;
  wire [31:0] _EVAL_5514;
  wire  _EVAL_406;
  wire  _EVAL_6072;
  wire  _EVAL_2109;
  wire  _EVAL_5048;
  wire [31:0] _EVAL_4929;
  wire  _EVAL_4101;
  wire  _EVAL_2045;
  wire [31:0] _EVAL_885;
  wire  _EVAL_3254;
  wire  _EVAL_231;
  wire  _EVAL_4552;
  wire  _EVAL_4393;
  wire  _EVAL_3916;
  wire  _EVAL_1916;
  wire  _EVAL_3108;
  wire  _EVAL_545;
  wire  _EVAL_6004;
  wire  _EVAL_1459;
  wire [31:0] _EVAL_699;
  wire  _EVAL_817;
  wire  _EVAL_3567;
  wire [31:0] _EVAL_1031;
  wire  _EVAL_3236;
  wire  _EVAL_5509;
  wire  _EVAL_3490;
  wire  _EVAL_2217;
  wire [31:0] _EVAL_2019;
  wire  _EVAL_5142;
  wire  _EVAL_4904;
  wire  _EVAL_4607;
  wire [31:0] _EVAL_2420;
  wire  _EVAL_539;
  wire  _EVAL_3154;
  wire [31:0] _EVAL_1335;
  wire  _EVAL_2738;
  wire  _EVAL_3532;
  wire [31:0] _EVAL_2435;
  wire  _EVAL_5551;
  wire  _EVAL_700;
  wire [31:0] _EVAL_3657;
  wire  _EVAL_2342;
  wire  _EVAL_4313;
  wire [31:0] _EVAL_1281;
  wire  _EVAL_4073;
  wire  _EVAL_4776;
  wire [31:0] _EVAL_1196;
  wire  _EVAL_1204;
  wire  _EVAL_2499;
  wire [31:0] _EVAL_1776;
  wire  _EVAL_2633;
  wire  _EVAL_3649;
  wire  _EVAL_4497;
  wire  _EVAL_424;
  wire  _EVAL_4886;
  wire [11:0] _EVAL_4407;
  wire  _EVAL_4539;
  wire  _EVAL_6091;
  wire  _EVAL_774;
  wire  _EVAL_2774;
  wire  _EVAL_5444;
  wire  _EVAL_3571;
  wire  _EVAL_6039;
  wire [31:0] _EVAL_5343;
  wire  _EVAL_1132;
  wire  _EVAL_5890;
  wire [31:0] _EVAL_940;
  wire  _EVAL_4408;
  wire  _EVAL_3325;
  wire [31:0] _EVAL_1712;
  wire  _EVAL_3409;
  wire  _EVAL_5371;
  wire [31:0] _EVAL_5288;
  wire  _EVAL_4149;
  wire  _EVAL_1256;
  wire [31:0] _EVAL_4881;
  wire  _EVAL_5635;
  wire  _EVAL_809;
  wire [31:0] _EVAL_1785;
  wire  _EVAL_5940;
  wire  _EVAL_5200;
  wire [31:0] _EVAL_4609;
  wire  _EVAL_4707;
  wire  _EVAL_3025;
  wire  _EVAL_4785;
  wire  _EVAL_4238;
  wire  _EVAL_4990;
  wire [7:0] _EVAL_500;
  wire  _EVAL_5914;
  wire  _EVAL_1909;
  wire  _EVAL_2632;
  wire  _EVAL_2474;
  wire  _EVAL_5256;
  wire  _EVAL_326;
  wire  _EVAL_902;
  wire  _EVAL_3055;
  wire  _EVAL_1833;
  wire [31:0] _EVAL_5134;
  wire  _EVAL_5682;
  wire  _EVAL_4477;
  wire  _EVAL_4705;
  wire  _EVAL_847;
  wire [31:0] _EVAL_4527;
  wire  _EVAL_5921;
  wire  _EVAL_1354;
  wire [31:0] _EVAL_547;
  wire  _EVAL_4102;
  wire  _EVAL_3663;
  wire  _EVAL_1741;
  wire [31:0] _EVAL_5757;
  wire  _EVAL_3725;
  wire  _EVAL_2136;
  wire  _EVAL_5782;
  wire [31:0] _EVAL_2426;
  wire  _EVAL_5791;
  wire  _EVAL_4253;
  wire  _EVAL_1873;
  wire  _EVAL_2085;
  wire  _EVAL_2871;
  wire  _EVAL_6127;
  wire  _EVAL_1952;
  wire  _EVAL_5619;
  wire  _EVAL_178;
  wire  _EVAL_2300;
  wire  _EVAL_1750;
  wire [31:0] _EVAL_2508;
  wire [31:0] _EVAL_4865;
  wire  _EVAL_2126;
  wire [31:0] _EVAL_5131;
  wire  _EVAL_1037;
  wire [31:0] _EVAL_3527;
  wire  _EVAL_1608;
  wire  _EVAL_4438;
  wire  _EVAL_1704;
  wire  _EVAL_1304;
  wire  _EVAL_3936;
  wire  _EVAL_4222;
  wire  _EVAL_5052;
  wire [31:0] _EVAL_1850;
  wire [11:0] _EVAL_792;
  wire [4:0] _EVAL_4765;
  wire [4:0] _EVAL_3551;
  wire [4:0] _EVAL_1847;
  wire [4:0] _EVAL_421;
  wire [4:0] _EVAL_3913;
  wire [4:0] _EVAL_1710;
  wire [4:0] _EVAL_698;
  wire  _EVAL_1434;
  wire  _EVAL_5378;
  wire  _EVAL_4579;
  wire  _EVAL_612;
  wire  _EVAL_198;
  wire  _EVAL_6078;
  wire [31:0] _EVAL_1945;
  wire  _EVAL_2119;
  wire  _EVAL_1782;
  wire [31:0] _EVAL_6109;
  wire  _EVAL_4610;
  wire  _EVAL_729;
  wire [31:0] _EVAL_4870;
  wire  _EVAL_4735;
  wire  _EVAL_4019;
  wire  _EVAL_1174;
  wire  _EVAL_1492;
  wire [4:0] _EVAL_5878;
  wire  _EVAL_1797;
  wire  _EVAL_1340;
  wire [31:0] _EVAL_1248;
  wire  _EVAL_425;
  wire  _EVAL_1828;
  wire [4:0] _EVAL_6087;
  wire  _EVAL_4955;
  wire  _EVAL_541;
  wire  _EVAL_3563;
  wire  _EVAL_1827;
  wire  _EVAL_4454;
  wire  _EVAL_4416;
  wire  _EVAL_1105;
  wire  _EVAL_465;
  wire  _EVAL_1185;
  wire [1:0] _EVAL_4381;
  wire [1:0] _EVAL_5481;
  wire [2:0] _EVAL_3299;
  wire [1:0] _EVAL_2638;
  wire [2:0] _EVAL_298;
  wire [3:0] _EVAL_184;
  wire [3:0] _EVAL_3061;
  wire [3:0] _EVAL_1472;
  wire [1:0] _EVAL_722;
  wire [3:0] _EVAL_2791;
  wire [3:0] _EVAL_712;
  wire [3:0] _EVAL_6085;
  wire [3:0] _EVAL_2943;
  wire [3:0] _EVAL_693;
  wire  _EVAL_358;
  wire  _EVAL_5859;
  wire  _EVAL_3810;
  wire [31:0] _EVAL_5126;
  wire  _EVAL_1616;
  wire  _EVAL_2543;
  wire [31:0] _EVAL_511;
  wire  _EVAL_1449;
  wire [31:0] _EVAL_2588;
  wire  _EVAL_4051;
  wire  _EVAL_2230;
  wire  _EVAL_2767;
  wire [31:0] _EVAL_2931;
  wire  _EVAL_2704;
  wire  _EVAL_3258;
  wire [31:0] _EVAL_5486;
  wire  _EVAL_4251;
  wire  _EVAL_417;
  wire  _EVAL_4058;
  wire  _EVAL_2376;
  wire  _EVAL_3626;
  wire  _EVAL_1487;
  wire  _EVAL_5650;
  wire  _EVAL_4508;
  wire  _EVAL_3716;
  wire  _EVAL_3878;
  wire  _EVAL_2345;
  wire  _EVAL_5027;
  wire [31:0] _EVAL_3934;
  wire  _EVAL_4249;
  wire  _EVAL_325;
  wire [31:0] _EVAL_2689;
  wire  _EVAL_5290;
  wire [31:0] _EVAL_3540;
  wire  _EVAL_3384;
  wire  _EVAL_1180;
  wire [31:0] _EVAL_1659;
  wire  _EVAL_2747;
  wire  _EVAL_4736;
  wire  _EVAL_2569;
  wire  _EVAL_3566;
  wire  _EVAL_5333;
  wire  _EVAL_5518;
  wire  _EVAL_811;
  wire  _EVAL_4682;
  wire [31:0] _EVAL_3740;
  wire  _EVAL_3167;
  wire [31:0] _EVAL_318;
  wire  _EVAL_2049;
  wire  _EVAL_1529;
  wire [31:0] _EVAL_339;
  wire  _EVAL_1156;
  wire  _EVAL_2823;
  wire [31:0] _EVAL_5735;
  wire  _EVAL_4792;
  wire  _EVAL_1148;
  wire  _EVAL_4898;
  wire [31:0] _EVAL_4384;
  wire  _EVAL_5838;
  wire  _EVAL_669;
  wire [31:0] _EVAL_1426;
  wire  _EVAL_1964;
  wire  _EVAL_4376;
  wire [31:0] _EVAL_1143;
  wire  _EVAL_2661;
  wire  _EVAL_4778;
  wire  _EVAL_2812;
  wire [31:0] _EVAL_835;
  wire  _EVAL_5954;
  wire  _EVAL_5161;
  wire [31:0] _EVAL_2226;
  wire  _EVAL_4690;
  wire [31:0] _EVAL_323;
  wire  _EVAL_1998;
  wire  _EVAL_4797;
  wire  _EVAL_4196;
  wire  _EVAL_1271;
  wire [31:0] _EVAL_6093;
  wire  _EVAL_1806;
  wire  _EVAL_1232;
  wire [31:0] _EVAL_4957;
  wire  _EVAL_4091;
  wire  _EVAL_3763;
  wire  _EVAL_4245;
  wire  _EVAL_3274;
  wire  _EVAL_4029;
  wire  _EVAL_3912;
  wire  _EVAL_5599;
  wire  _EVAL_3542;
  wire  _EVAL_1396;
  wire  _EVAL_992;
  wire  _EVAL_1238;
  wire  _EVAL_1234;
  wire  _EVAL_953;
  wire [31:0] _EVAL_1976;
  wire  _EVAL_4028;
  wire [31:0] _EVAL_2537;
  wire  _EVAL_395;
  wire  _EVAL_6067;
  wire  _EVAL_5798;
  wire  _EVAL_671;
  wire [31:0] _EVAL_6079;
  wire  _EVAL_5025;
  wire  _EVAL_5425;
  wire  _EVAL_195;
  wire [31:0] _EVAL_982;
  wire  _EVAL_3201;
  wire [31:0] _EVAL_916;
  wire  _EVAL_5407;
  wire  _EVAL_2549;
  wire [31:0] _EVAL_3813;
  wire  _EVAL_5263;
  wire  _EVAL_3536;
  wire  _EVAL_3084;
  wire  _EVAL_5683;
  wire [31:0] _EVAL_4819;
  wire  _EVAL_3317;
  wire  _EVAL_4272;
  wire [31:0] _EVAL_5513;
  wire  _EVAL_5856;
  wire [31:0] _EVAL_552;
  wire  _EVAL_2753;
  wire  _EVAL_5108;
  wire  _EVAL_2165;
  wire  _EVAL_5587;
  wire  _EVAL_3687;
  wire  _EVAL_6061;
  wire [31:0] _EVAL_5963;
  wire  _EVAL_2729;
  wire  _EVAL_1738;
  wire  _EVAL_4949;
  wire  _EVAL_5764;
  wire  _EVAL_5129;
  wire  _EVAL_5299;
  wire [31:0] _EVAL_4861;
  wire  _EVAL_3085;
  wire [31:0] _EVAL_5819;
  wire  _EVAL_2953;
  wire  _EVAL_2682;
  wire [31:0] _EVAL_2828;
  wire  _EVAL_3007;
  wire  _EVAL_655;
  wire  _EVAL_6099;
  wire [31:0] _EVAL_4519;
  wire  _EVAL_2158;
  wire [31:0] _EVAL_4274;
  wire  _EVAL_3191;
  wire  _EVAL_4156;
  wire  _EVAL_226;
  wire  _EVAL_5850;
  wire  _EVAL_5460;
  wire  _EVAL_3368;
  wire  _EVAL_5955;
  wire [31:0] _EVAL_853;
  wire  _EVAL_2679;
  wire  _EVAL_4566;
  wire  _EVAL_6100;
  wire [31:0] _EVAL_3714;
  wire  _EVAL_5728;
  wire  _EVAL_1596;
  wire [31:0] _EVAL_3977;
  wire  _EVAL_3476;
  wire [31:0] _EVAL_5526;
  wire  _EVAL_5598;
  wire  _EVAL_434;
  wire [31:0] _EVAL_3825;
  wire  _EVAL_3653;
  wire  _EVAL_3555;
  wire  _EVAL_3316;
  wire  _EVAL_4520;
  wire  _EVAL_220;
  wire  _EVAL_2094;
  wire  _EVAL_4672;
  wire  _EVAL_1943;
  wire  _EVAL_3181;
  wire  _EVAL_2565;
  wire [31:0] _EVAL_4757;
  wire  _EVAL_2065;
  wire  _EVAL_385;
  wire [31:0] _EVAL_1872;
  wire  _EVAL_4912;
  wire  _EVAL_3185;
  wire  _EVAL_1561;
  wire  _EVAL_4549;
  wire  _EVAL_3773;
  wire  _EVAL_1932;
  wire  _EVAL_5177;
  wire  _EVAL_2395;
  wire  _EVAL_235;
  wire  _EVAL_3601;
  wire  _EVAL_4378;
  wire  _EVAL_3161;
  wire [31:0] _EVAL_5436;
  wire  _EVAL_5751;
  wire  _EVAL_2227;
  wire  _EVAL_4981;
  wire  _EVAL_3664;
  wire  _EVAL_984;
  wire  _EVAL_5018;
  wire  _EVAL_5169;
  wire  _EVAL_5148;
  wire  _EVAL_2562;
  wire  _EVAL_3176;
  wire  _EVAL_1626;
  wire  _EVAL_727;
  wire [3:0] _EVAL_3900;
  wire [3:0] _EVAL_5125;
  wire  _EVAL_1020;
  wire  _EVAL_3804;
  wire  _EVAL_773;
  wire  _EVAL_917;
  wire  _EVAL_275;
  wire  _EVAL_1427;
  wire  _EVAL_4095;
  wire  _EVAL_4794;
  wire  _EVAL_631;
  wire [31:0] _EVAL_5911;
  wire  _EVAL_1562;
  wire  _EVAL_1774;
  wire  _EVAL_556;
  wire  _EVAL_910;
  wire [31:0] _EVAL_5865;
  wire  _EVAL_444;
  wire [31:0] _EVAL_3647;
  wire  _EVAL_507;
  wire  _EVAL_217;
  wire [31:0] _EVAL_2472;
  wire  _EVAL_1509;
  wire  _EVAL_5307;
  wire  _EVAL_5073;
  wire  _EVAL_3805;
  wire  _EVAL_3269;
  wire  _EVAL_5704;
  wire  _EVAL_799;
  wire [31:0] _EVAL_225;
  wire  _EVAL_4479;
  wire [31:0] _EVAL_4975;
  wire  _EVAL_1344;
  wire  _EVAL_793;
  wire [31:0] _EVAL_3227;
  wire  _EVAL_2504;
  wire [31:0] _EVAL_1404;
  wire  _EVAL_4907;
  wire  _EVAL_3220;
  wire  _EVAL_5091;
  wire  _EVAL_2787;
  wire  _EVAL_1410;
  wire  _EVAL_1139;
  wire [31:0] _EVAL_5974;
  wire  _EVAL_956;
  wire  _EVAL_5098;
  wire [31:0] _EVAL_1796;
  wire  _EVAL_5571;
  wire  _EVAL_3603;
  wire [31:0] _EVAL_967;
  wire [31:0] _EVAL_6115;
  wire  _EVAL_3289;
  wire  _EVAL_5399;
  wire  _EVAL_1373;
  wire  _EVAL_2705;
  wire  _EVAL_3353;
  wire  _EVAL_3938;
  wire  _EVAL_2124;
  wire  _EVAL_3283;
  wire [31:0] _EVAL_5090;
  wire  _EVAL_1258;
  wire  _EVAL_4270;
  wire [31:0] _EVAL_851;
  wire  _EVAL_4331;
  wire  _EVAL_4850;
  wire [31:0] _EVAL_2861;
  wire  _EVAL_3110;
  wire  _EVAL_4165;
  wire  _EVAL_2041;
  wire [31:0] _EVAL_5471;
  wire  _EVAL_4124;
  wire  _EVAL_3683;
  wire  _EVAL_5267;
  wire  _EVAL_3633;
  wire [31:0] _EVAL_4684;
  wire  _EVAL_2133;
  wire [31:0] _EVAL_1253;
  wire  _EVAL_1359;
  wire [31:0] _EVAL_4341;
  wire  _EVAL_4121;
  wire  _EVAL_4287;
  wire  _EVAL_3512;
  wire  _EVAL_4921;
  wire [31:0] _EVAL_3145;
  wire  _EVAL_6057;
  wire [31:0] _EVAL_2024;
  wire  _EVAL_1220;
  wire  _EVAL_6062;
  wire [31:0] _EVAL_1223;
  wire  _EVAL_2310;
  wire  _EVAL_616;
  wire  _EVAL_2103;
  wire [31:0] _EVAL_1457;
  wire  _EVAL_242;
  wire  _EVAL_361;
  wire  _EVAL_469;
  wire [31:0] _EVAL_370;
  wire  _EVAL_2756;
  wire [31:0] _EVAL_1042;
  wire  _EVAL_2636;
  wire  _EVAL_369;
  wire [31:0] _EVAL_2212;
  wire  _EVAL_160;
  wire  _EVAL_2836;
  wire  _EVAL_4614;
  wire  _EVAL_3651;
  wire  _EVAL_4258;
  wire [31:0] _EVAL_1919;
  wire  _EVAL_648;
  wire [31:0] _EVAL_4369;
  wire  _EVAL_1735;
  wire  _EVAL_1878;
  wire [31:0] _EVAL_1228;
  wire  _EVAL_4811;
  wire  _EVAL_302;
  wire  _EVAL_3589;
  wire [31:0] _EVAL_5341;
  wire [31:0] _EVAL_2276;
  wire  _EVAL_768;
  wire  _EVAL_1222;
  wire  _EVAL_2590;
  wire  _EVAL_5361;
  wire  _EVAL_2951;
  wire  _EVAL_2963;
  wire  _EVAL_254;
  wire  _EVAL_2211;
  wire [31:0] _EVAL_5410;
  wire  _EVAL_1730;
  wire  _EVAL_4906;
  wire [31:0] _EVAL_872;
  wire  _EVAL_3958;
  wire [31:0] _EVAL_2224;
  wire  _EVAL_2339;
  wire  _EVAL_6135;
  wire [31:0] _EVAL_1981;
  wire  _EVAL_4406;
  wire  _EVAL_1772;
  wire [6:0] _EVAL_4469;
  wire [6:0] _EVAL_3817;
  wire [6:0] _EVAL_2894;
  wire [6:0] _EVAL_5628;
  wire [6:0] _EVAL_3488;
  wire [31:0] _EVAL_2929;
  wire [31:0] _EVAL_3994;
  wire  _EVAL_3866;
  wire  _EVAL_5630;
  wire [31:0] _EVAL_1654;
  wire  _EVAL_1931;
  wire  _EVAL_864;
  wire [6:0] _EVAL_490;
  wire [31:0] _EVAL_3042;
  wire  _EVAL_4787;
  wire  _EVAL_4057;
  wire [31:0] _EVAL_1313;
  wire  _EVAL_330;
  wire  _EVAL_2000;
  wire [31:0] _EVAL_1133;
  wire  _EVAL_5927;
  wire  _EVAL_5269;
  wire  _EVAL_2662;
  wire  _EVAL_3666;
  wire  _EVAL_4056;
  wire  _EVAL_3745;
  wire [31:0] _EVAL_3800;
  wire  _EVAL_6076;
  wire  _EVAL_5431;
  wire [31:0] _EVAL_2365;
  wire  _EVAL_4157;
  wire  _EVAL_4688;
  wire [31:0] _EVAL_1260;
  wire  _EVAL_3964;
  wire  _EVAL_1648;
  wire [31:0] _EVAL_760;
  wire  _EVAL_4629;
  wire  _EVAL_3537;
  wire [31:0] _EVAL_2406;
  wire  _EVAL_1655;
  wire  _EVAL_4934;
  wire  _EVAL_826;
  wire  _EVAL_2071;
  wire  _EVAL_3047;
  wire  _EVAL_2641;
  wire  _EVAL_201;
  wire [31:0] _EVAL_1070;
  wire  _EVAL_4653;
  wire  _EVAL_4322;
  wire [31:0] _EVAL_5406;
  wire  _EVAL_3031;
  wire  _EVAL_6136;
  wire  _EVAL_4340;
  wire  _EVAL_1538;
  wire  _EVAL_3173;
  wire  _EVAL_4773;
  wire [31:0] _EVAL_1168;
  wire  _EVAL_2884;
  wire  _EVAL_2766;
  wire [1:0] _EVAL_3992;
  wire [1:0] _EVAL_5574;
  wire  _EVAL_3080;
  wire  _EVAL_2458;
  wire [31:0] _EVAL_5418;
  wire [4:0] _EVAL_4470;
  wire [4:0] _EVAL_5153;
  wire [4:0] _EVAL_5261;
  wire [4:0] _EVAL_4919;
  wire [4:0] _EVAL_2141;
  wire [4:0] _EVAL_3703;
  wire [4:0] _EVAL_2336;
  wire [4:0] _EVAL_4223;
  wire [4:0] _EVAL_2388;
  wire [4:0] _EVAL_1276;
  wire [4:0] _EVAL_1593;
  wire [4:0] _EVAL_5377;
  wire [4:0] _EVAL_3104;
  wire [4:0] _EVAL_4491;
  wire [4:0] _EVAL_794;
  wire [4:0] _EVAL_4846;
  wire [4:0] _EVAL_3594;
  wire [4:0] _EVAL_261;
  wire [4:0] _EVAL_166;
  wire [4:0] _EVAL_5965;
  wire [4:0] _EVAL_5128;
  wire [4:0] _EVAL_3548;
  wire [4:0] _EVAL_5492;
  wire [4:0] _EVAL_1028;
  wire [4:0] _EVAL_2343;
  wire [4:0] _EVAL_639;
  wire [31:0] _EVAL_4486;
  wire  _EVAL_317;
  wire  _EVAL_3969;
  wire  _EVAL_4339;
  wire  _EVAL_5572;
  wire [31:0] _EVAL_4585;
  wire  _EVAL_5247;
  wire [4:0] _EVAL_3259;
  wire [4:0] _EVAL_2496;
  wire [4:0] _EVAL_5520;
  wire [4:0] _EVAL_3059;
  wire [31:0] _EVAL_3828;
  wire [31:0] _EVAL_1887;
  wire  _EVAL_400;
  wire [31:0] _EVAL_3140;
  wire  _EVAL_2139;
  wire  _EVAL_229;
  wire [31:0] _EVAL_1338;
  wire  _EVAL_381;
  wire  _EVAL_4320;
  wire  _EVAL_928;
  wire  _EVAL_2717;
  wire [31:0] _EVAL_3404;
  wire  _EVAL_2986;
  wire  _EVAL_534;
  wire [31:0] _EVAL_5397;
  wire  _EVAL_1424;
  wire  _EVAL_4476;
  wire [31:0] _EVAL_5016;
  wire  _EVAL_2906;
  wire  _EVAL_2631;
  wire [31:0] _EVAL_3629;
  wire  _EVAL_832;
  wire  _EVAL_489;
  wire  _EVAL_4254;
  wire  _EVAL_5986;
  wire  _EVAL_3248;
  wire  _EVAL_5445;
  wire [31:0] _EVAL_514;
  wire  _EVAL_5157;
  wire  _EVAL_2355;
  wire [31:0] _EVAL_5906;
  wire  _EVAL_2763;
  wire  _EVAL_1518;
  wire [31:0] _EVAL_4144;
  wire  _EVAL_749;
  wire  _EVAL_4346;
  wire [31:0] _EVAL_1017;
  wire  _EVAL_5306;
  wire  _EVAL_4840;
  wire  _EVAL_893;
  wire  _EVAL_5150;
  wire  _EVAL_3450;
  wire [31:0] _EVAL_194;
  wire  _EVAL_2220;
  wire  _EVAL_5374;
  wire  _EVAL_3155;
  wire  _EVAL_5022;
  wire  _EVAL_1043;
  wire  _EVAL_4877;
  wire [31:0] _EVAL_174;
  wire  _EVAL_412;
  wire  _EVAL_4766;
  wire [31:0] _EVAL_5032;
  wire  _EVAL_2591;
  wire [31:0] _EVAL_441;
  wire [31:0] _EVAL_4328;
  wire  _EVAL_2317;
  wire [31:0] _EVAL_4252;
  wire  _EVAL_3799;
  wire [31:0] _EVAL_196;
  wire  _EVAL_2038;
  wire  _EVAL_3282;
  wire  _EVAL_4365;
  wire  _EVAL_1691;
  wire  _EVAL_384;
  wire [31:0] _EVAL_5678;
  wire  _EVAL_5230;
  wire  _EVAL_566;
  wire [31:0] _EVAL_4623;
  wire  _EVAL_4243;
  wire [31:0] _EVAL_4442;
  wire  _EVAL_6106;
  wire  _EVAL_204;
  wire  _EVAL_5980;
  wire [31:0] _EVAL_1658;
  wire  _EVAL_1923;
  wire [31:0] _EVAL_2488;
  wire  _EVAL_281;
  wire  _EVAL_2415;
  wire  _EVAL_3273;
  wire [31:0] _EVAL_3244;
  wire  _EVAL_2620;
  wire  _EVAL_2815;
  wire [31:0] _EVAL_3856;
  wire  _EVAL_1445;
  wire  _EVAL_5059;
  wire [31:0] _EVAL_3865;
  wire  _EVAL_2803;
  wire  _EVAL_5968;
  wire  _EVAL_5972;
  wire  _EVAL_521;
  wire  _EVAL_1343;
  wire  _EVAL_4315;
  wire [31:0] _EVAL_3313;
  wire  _EVAL_5310;
  wire  _EVAL_6122;
  wire  _EVAL_4032;
  wire  _EVAL_4090;
  wire [31:0] _EVAL_1901;
  wire  _EVAL_4035;
  wire  _EVAL_5871;
  wire [31:0] _EVAL_5146;
  wire  _EVAL_737;
  wire  _EVAL_5235;
  wire [31:0] _EVAL_1625;
  wire  _EVAL_1714;
  wire  _EVAL_248;
  wire  _EVAL_2366;
  wire  _EVAL_1548;
  wire  _EVAL_1966;
  wire  _EVAL_1401;
  wire [31:0] _EVAL_6024;
  wire  _EVAL_2450;
  wire  _EVAL_4498;
  wire [31:0] _EVAL_5827;
  wire  _EVAL_535;
  wire  _EVAL_5805;
  wire [31:0] _EVAL_3092;
  wire  _EVAL_1288;
  wire  _EVAL_599;
  wire  _EVAL_4298;
  wire  _EVAL_4158;
  wire [4:0] _EVAL_5447;
  wire  _EVAL_5767;
  wire [31:0] _EVAL_2995;
  wire  _EVAL_573;
  wire  _EVAL_2650;
  wire  _EVAL_5726;
  wire [31:0] _EVAL_995;
  wire  _EVAL_3511;
  wire  _EVAL_1397;
  wire  _EVAL_305;
  wire  _EVAL_2331;
  wire  _EVAL_1999;
  wire [31:0] _EVAL_5803;
  wire  _EVAL_4900;
  wire  _EVAL_5742;
  wire [4:0] _EVAL_190;
  wire  _EVAL_266;
  wire  _EVAL_4377;
  wire  _EVAL_4706;
  wire  _EVAL_3197;
  wire  _EVAL_572;
  wire  _EVAL_6114;
  wire [31:0] _EVAL_2402;
  wire  _EVAL_4307;
  wire  _EVAL_5873;
  wire [31:0] _EVAL_2155;
  wire  _EVAL_5084;
  wire  _EVAL_5468;
  wire  _EVAL_1237;
  wire  _EVAL_4555;
  wire  _EVAL_3205;
  wire [31:0] _EVAL_5507;
  wire  _EVAL_4130;
  wire [31:0] _EVAL_2832;
  wire  _EVAL_1786;
  wire  _EVAL_4195;
  wire [31:0] _EVAL_5035;
  wire  _EVAL_4616;
  wire  _EVAL_3427;
  wire [31:0] _EVAL_3688;
  wire  _EVAL_5910;
  wire  _EVAL_1584;
  wire  _EVAL_216;
  wire  _EVAL_1055;
  wire  _EVAL_2716;
  wire [31:0] _EVAL_4205;
  wire  _EVAL_3442;
  wire  _EVAL_428;
  wire [31:0] _EVAL_4005;
  wire  _EVAL_5545;
  wire  _EVAL_3171;
  wire [31:0] _EVAL_5950;
  wire  _EVAL_1480;
  wire  _EVAL_2978;
  wire [31:0] _EVAL_3652;
  wire  _EVAL_3565;
  wire  _EVAL_784;
  wire  _EVAL_589;
  wire  _EVAL_1308;
  wire [31:0] _EVAL_625;
  wire  _EVAL_4721;
  wire  _EVAL_4010;
  wire [31:0] _EVAL_3252;
  wire  _EVAL_819;
  wire  _EVAL_4851;
  wire  _EVAL_4007;
  wire  _EVAL_3159;
  wire  _EVAL_3858;
  wire  _EVAL_1517;
  wire  _EVAL_3568;
  wire  _EVAL_485;
  wire  _EVAL_5180;
  wire [4:0] _EVAL_4150;
  wire  _EVAL_844;
  wire  _EVAL_862;
  wire [4:0] _EVAL_488;
  wire  _EVAL_3791;
  wire  _EVAL_4611;
  wire  _EVAL_5103;
  wire  _EVAL_4424;
  wire  _EVAL_4015;
  wire  _EVAL_4259;
  wire [31:0] _EVAL_958;
  wire [31:0] _EVAL_5370;
  wire  _EVAL_2446;
  wire  _EVAL_5279;
  wire [31:0] _EVAL_4599;
  wire  _EVAL_5085;
  wire  _EVAL_1913;
  wire [31:0] _EVAL_5747;
  wire  _EVAL_189;
  wire  _EVAL_523;
  wire  _EVAL_2695;
  wire [31:0] _EVAL_5241;
  wire  _EVAL_931;
  wire  _EVAL_4943;
  wire  _EVAL_2700;
  wire  _EVAL_3304;
  wire [31:0] _EVAL_319;
  wire  _EVAL_1298;
  wire [31:0] _EVAL_4423;
  wire  _EVAL_1946;
  wire  _EVAL_419;
  wire  _EVAL_4516;
  wire [31:0] _EVAL_4899;
  wire  _EVAL_840;
  wire  _EVAL_3122;
  wire  _EVAL_3422;
  wire [31:0] _EVAL_5626;
  wire  _EVAL_3230;
  wire  _EVAL_3375;
  wire  _EVAL_3981;
  wire  _EVAL_3044;
  wire  _EVAL_221;
  wire  _EVAL_1615;
  wire  _EVAL_314;
  wire  _EVAL_2760;
  wire  _EVAL_475;
  wire  _EVAL_2593;
  wire  _EVAL_5852;
  wire  _EVAL_4240;
  wire [31:0] _EVAL_5450;
  wire  _EVAL_4844;
  wire  _EVAL_3697;
  wire [31:0] _EVAL_4414;
  wire  _EVAL_4569;
  wire  _EVAL_6036;
  wire [31:0] _EVAL_786;
  wire  _EVAL_2793;
  wire  _EVAL_1632;
  wire [31:0] _EVAL_899;
  wire  _EVAL_686;
  wire  _EVAL_5218;
  wire  _EVAL_1522;
  wire  _EVAL_5353;
  wire  _EVAL_4983;
  wire  _EVAL_743;
  wire  _EVAL_2824;
  wire  _EVAL_2927;
  wire  _EVAL_4837;
  wire  _EVAL_4323;
  wire  _EVAL_4300;
  wire  _EVAL_2730;
  wire  _EVAL_3668;
  wire  _EVAL_2495;
  wire  _EVAL_5257;
  wire  _EVAL_6025;
  wire  _EVAL_2162;
  wire  _EVAL_5996;
  wire  _EVAL_2637;
  wire  _EVAL_3151;
  wire  _EVAL_663;
  wire  _EVAL_186;
  wire  _EVAL_3742;
  wire  _EVAL_2160;
  wire  _EVAL_1094;
  wire  _EVAL_1619;
  wire  _EVAL_5824;
  wire  _EVAL_4676;
  wire  _EVAL_1038;
  wire  _EVAL_4068;
  wire  _EVAL_399;
  wire  _EVAL_4472;
  wire  _EVAL_2728;
  wire  _EVAL_2966;
  wire  _EVAL_716;
  wire  _EVAL_2169;
  wire  _EVAL_2413;
  wire  _EVAL_2925;
  wire [3:0] _EVAL_1889;
  wire [3:0] _EVAL_4595;
  wire  _EVAL_4006;
  wire  _EVAL_2447;
  wire [31:0] _EVAL_2218;
  wire  _EVAL_2942;
  wire  _EVAL_2990;
  wire  _EVAL_692;
  wire  _EVAL_816;
  wire  _EVAL_4849;
  wire  _EVAL_1178;
  wire [31:0] _EVAL_1240;
  wire  _EVAL_2095;
  wire  _EVAL_5536;
  wire [31:0] _EVAL_5358;
  wire  _EVAL_4169;
  wire  _EVAL_1818;
  wire [31:0] _EVAL_5730;
  wire  _EVAL_866;
  wire  _EVAL_4162;
  wire  _EVAL_349;
  wire [31:0] _EVAL_2254;
  wire  _EVAL_1683;
  wire  _EVAL_3464;
  wire [31:0] _EVAL_1046;
  wire  _EVAL_3226;
  wire  _EVAL_4464;
  wire [31:0] _EVAL_5485;
  wire  _EVAL_2688;
  wire  _EVAL_2893;
  wire  _EVAL_5412;
  wire  _EVAL_5647;
  wire  _EVAL_4279;
  wire  _EVAL_5554;
  wire [31:0] _EVAL_5917;
  wire  _EVAL_2356;
  wire  _EVAL_4523;
  wire [31:0] _EVAL_3556;
  wire  _EVAL_5936;
  wire  _EVAL_3127;
  wire  _EVAL_2536;
  wire  _EVAL_1252;
  wire  _EVAL_5592;
  wire  _EVAL_176;
  wire  _EVAL_2601;
  wire [31:0] _EVAL_4312;
  wire  _EVAL_1533;
  wire  _EVAL_869;
  wire [31:0] _EVAL_5467;
  wire  _EVAL_5922;
  wire  _EVAL_1229;
  wire  _EVAL_2518;
  wire  _EVAL_6142;
  wire  _EVAL_5266;
  wire  _EVAL_3132;
  wire  _EVAL_5763;
  wire  _EVAL_5040;
  wire  _EVAL_5395;
  wire [31:0] _EVAL_529;
  wire  _EVAL_5106;
  wire  _EVAL_2686;
  wire [31:0] _EVAL_5627;
  wire  _EVAL_3429;
  wire  _EVAL_4761;
  wire  _EVAL_1767;
  wire  _EVAL_5457;
  wire [31:0] _EVAL_3095;
  wire  _EVAL_5184;
  wire  _EVAL_873;
  wire  _EVAL_5349;
  wire  _EVAL_3237;
  wire  _EVAL_1147;
  wire  _EVAL_3569;
  wire  _EVAL_4600;
  wire  _EVAL_2634;
  wire  _EVAL_2630;
  wire  _EVAL_5984;
  wire [31:0] _EVAL_5706;
  wire  _EVAL_3743;
  wire [31:0] _EVAL_5681;
  wire  _EVAL_199;
  wire  _EVAL_2852;
  wire  _EVAL_2764;
  wire  _EVAL_4053;
  wire  _EVAL_5684;
  wire  _EVAL_1497;
  wire [31:0] _EVAL_1012;
  wire  _EVAL_711;
  wire  _EVAL_990;
  wire  _EVAL_1011;
  wire  _EVAL_170;
  wire  _EVAL_3019;
  wire [31:0] _EVAL_2286;
  wire  _EVAL_5031;
  wire  _EVAL_933;
  wire [31:0] _EVAL_765;
  wire  _EVAL_713;
  wire  _EVAL_4650;
  wire [31:0] _EVAL_1301;
  wire  _EVAL_4459;
  wire  _EVAL_5998;
  wire  _EVAL_4380;
  wire [31:0] _EVAL_3505;
  wire  _EVAL_3195;
  wire  _EVAL_3547;
  wire  _EVAL_622;
  wire  _EVAL_2553;
  wire  _EVAL_2974;
  wire [31:0] _EVAL_5710;
  wire  _EVAL_912;
  wire  _EVAL_4958;
  wire [3:0] _EVAL_3771;
  wire  _EVAL_4675;
  wire [31:0] _EVAL_4411;
  wire  _EVAL_5111;
  wire  _EVAL_1637;
  wire  _EVAL_5030;
  wire  _EVAL_1841;
  wire [31:0] _EVAL_2298;
  wire  _EVAL_723;
  wire  _EVAL_4093;
  wire [31:0] _EVAL_2922;
  wire  _EVAL_1024;
  wire  _EVAL_208;
  wire [31:0] _EVAL_3615;
  wire  _EVAL_4938;
  wire  _EVAL_3889;
  wire  _EVAL_3572;
  wire  _EVAL_2478;
  wire [31:0] _EVAL_802;
  wire  _EVAL_4046;
  wire  _EVAL_5982;
  wire [31:0] _EVAL_5639;
  wire  _EVAL_2560;
  wire  _EVAL_1838;
  wire [31:0] _EVAL_5983;
  wire  _EVAL_1503;
  wire  _EVAL_2369;
  wire [31:0] _EVAL_3523;
  wire  _EVAL_2354;
  wire  _EVAL_2810;
  wire [31:0] _EVAL_508;
  wire  _EVAL_1815;
  wire  _EVAL_1195;
  wire  _EVAL_1347;
  wire  _EVAL_1885;
  wire [31:0] _EVAL_2775;
  wire  _EVAL_949;
  wire  _EVAL_482;
  wire  _EVAL_3539;
  wire  _EVAL_1001;
  wire [31:0] _EVAL_2660;
  wire  _EVAL_6095;
  wire  _EVAL_1664;
  wire [31:0] _EVAL_4433;
  wire  _EVAL_4107;
  wire  _EVAL_3362;
  wire [31:0] _EVAL_664;
  wire  _EVAL_3124;
  wire  _EVAL_244;
  wire [31:0] _EVAL_6060;
  wire  _EVAL_4215;
  wire  _EVAL_5152;
  wire  _EVAL_2361;
  wire  _EVAL_2283;
  wire  _EVAL_5839;
  wire [31:0] _EVAL_6058;
  wire  _EVAL_930;
  wire  _EVAL_5046;
  wire  _EVAL_313;
  wire  _EVAL_3158;
  wire  _EVAL_230;
  wire  _EVAL_442;
  wire  _EVAL_4310;
  wire  _EVAL_2015;
  wire [31:0] _EVAL_387;
  wire  _EVAL_1049;
  wire  _EVAL_4357;
  wire  _EVAL_1725;
  wire [31:0] _EVAL_3592;
  wire  _EVAL_2363;
  wire  _EVAL_1514;
  wire [31:0] _EVAL_3357;
  wire  _EVAL_4299;
  wire  _EVAL_925;
  wire  _EVAL_1895;
  wire  _EVAL_1770;
  wire [31:0] _EVAL_4582;
  wire  _EVAL_5205;
  wire  _EVAL_1154;
  wire [31:0] _EVAL_3342;
  wire  _EVAL_2813;
  wire [6:0] _EVAL_4824;
  wire [4:0] _EVAL_5192;
  wire [4:0] _EVAL_4605;
  wire [4:0] _EVAL_2873;
  wire [4:0] _EVAL_5849;
  wire [4:0] _EVAL_3754;
  wire  _EVAL_1188;
  wire [31:0] _EVAL_791;
  wire  _EVAL_5317;
  wire [31:0] _EVAL_2864;
  wire  _EVAL_271;
  wire  _EVAL_6134;
  wire [4:0] _EVAL_1294;
  wire [3:0] _EVAL_4624;
  wire [3:0] _EVAL_586;
  wire [4:0] _EVAL_5793;
  wire [4:0] _EVAL_3033;
  wire [4:0] _EVAL_3689;
  wire [4:0] _EVAL_3456;
  wire [4:0] _EVAL_2294;
  wire [4:0] _EVAL_1692;
  wire [4:0] _EVAL_4612;
  wire [4:0] _EVAL_1091;
  wire [4:0] _EVAL_390;
  wire [4:0] _EVAL_5248;
  wire [4:0] _EVAL_5312;
  wire [4:0] _EVAL_2291;
  wire  _EVAL_2273;
  wire  _EVAL_1002;
  wire [31:0] _EVAL_3389;
  wire  _EVAL_191;
  wire  _EVAL_1438;
  wire [31:0] _EVAL_3335;
  wire  _EVAL_1345;
  wire  _EVAL_3388;
  wire [31:0] _EVAL_5154;
  wire  _EVAL_1247;
  wire  _EVAL_2333;
  wire [31:0] _EVAL_3093;
  wire  _EVAL_4564;
  wire  _EVAL_1902;
  wire  _EVAL_4888;
  wire  _EVAL_3868;
  wire  _EVAL_5830;
  wire  _EVAL_1403;
  wire  _EVAL_3998;
  wire [31:0] _EVAL_3665;
  wire  _EVAL_398;
  wire  _EVAL_487;
  wire  _EVAL_4379;
  wire [31:0] _EVAL_1306;
  wire  _EVAL_363;
  wire  _EVAL_3993;
  wire  _EVAL_1801;
  wire  _EVAL_555;
  wire [31:0] _EVAL_3156;
  wire  _EVAL_941;
  wire  _EVAL_3175;
  wire [31:0] _EVAL_5055;
  wire  _EVAL_5366;
  wire  _EVAL_2768;
  wire  _EVAL_2195;
  wire [31:0] _EVAL_2985;
  wire  _EVAL_3552;
  wire  _EVAL_1512;
  wire  _EVAL_2448;
  wire  _EVAL_5092;
  wire [31:0] _EVAL_3350;
  wire  _EVAL_3919;
  wire  _EVAL_443;
  wire  _EVAL_1117;
  wire  _EVAL_1521;
  wire  _EVAL_459;
  wire  _EVAL_2946;
  wire [31:0] _EVAL_5199;
  wire  _EVAL_3753;
  wire  _EVAL_4666;
  wire  _EVAL_980;
  wire  _EVAL_2726;
  wire  _EVAL_828;
  wire  _EVAL_472;
  wire  _EVAL_3894;
  wire [31:0] _EVAL_3780;
  wire  _EVAL_5068;
  wire  _EVAL_5901;
  wire  _EVAL_3174;
  wire [31:0] _EVAL_4246;
  wire  _EVAL_1963;
  wire  _EVAL_4456;
  wire [31:0] _EVAL_2243;
  wire  _EVAL_2424;
  wire  _EVAL_4565;
  wire  _EVAL_5861;
  wire  _EVAL_342;
  wire  _EVAL_901;
  wire  _EVAL_1861;
  wire  _EVAL_3188;
  wire [31:0] _EVAL_681;
  wire  _EVAL_833;
  wire  _EVAL_5121;
  wire  _EVAL_4619;
  wire  _EVAL_3366;
  wire  _EVAL_3217;
  wire  _EVAL_2988;
  wire  _EVAL_3270;
  wire  _EVAL_661;
  wire  _EVAL_233;
  wire  _EVAL_2436;
  wire  _EVAL_4700;
  wire  _EVAL_1870;
  wire  _EVAL_5846;
  wire  _EVAL_890;
  wire  _EVAL_4889;
  wire  _EVAL_3367;
  wire  _EVAL_3604;
  wire  _EVAL_5221;
  wire  _EVAL_3597;
  wire  _EVAL_478;
  wire  _EVAL_4723;
  wire  _EVAL_2168;
  wire  _EVAL_742;
  wire  _EVAL_1886;
  wire  _EVAL_6069;
  wire  _EVAL_5566;
  wire  _EVAL_2340;
  wire  _EVAL_603;
  wire  _EVAL_4241;
  wire  _EVAL_2918;
  wire  _EVAL_1436;
  wire  _EVAL_1087;
  wire  _EVAL_814;
  wire [3:0] _EVAL_2089;
  wire  _EVAL_1554;
  wire  _EVAL_1165;
  wire  _EVAL_973;
  wire [31:0] _EVAL_525;
  wire  _EVAL_918;
  wire [4:0] _EVAL_2652;
  wire  _EVAL_5414;
  wire [31:0] _EVAL_4615;
  wire  _EVAL_994;
  wire  _EVAL_4587;
  wire  _EVAL_883;
  wire  _EVAL_3199;
  wire  _EVAL_3625;
  wire  _EVAL_4710;
  wire  _EVAL_2381;
  wire  _EVAL_1145;
  wire [31:0] _EVAL_3153;
  wire  _EVAL_4105;
  wire  _EVAL_4679;
  wire  _EVAL_2586;
  wire  _EVAL_5506;
  wire  _EVAL_5655;
  wire  _EVAL_3525;
  wire [31:0] _EVAL_1386;
  wire  _EVAL_1756;
  wire  _EVAL_4873;
  wire [31:0] _EVAL_1468;
  wire  _EVAL_2998;
  wire  _EVAL_3144;
  wire [31:0] _EVAL_1574;
  wire  _EVAL_2267;
  wire [4:0] _EVAL_5237;
  wire  _EVAL_5250;
  wire [31:0] _EVAL_249;
  wire  _EVAL_4621;
  wire  _EVAL_336;
  wire  _EVAL_619;
  wire  _EVAL_2619;
  wire  _EVAL_2319;
  wire  _EVAL_2677;
  wire [31:0] _EVAL_4915;
  wire  _EVAL_517;
  wire [31:0] _EVAL_4597;
  wire  _EVAL_4275;
  wire  _EVAL_4000;
  wire [31:0] _EVAL_1794;
  wire  _EVAL_5120;
  wire  _EVAL_1865;
  wire [31:0] _EVAL_2172;
  wire  _EVAL_2928;
  wire  _EVAL_4514;
  wire [31:0] _EVAL_1159;
  wire  _EVAL_4986;
  wire  _EVAL_1883;
  wire [31:0] _EVAL_2265;
  wire  _EVAL_2416;
  wire  _EVAL_2814;
  wire  _EVAL_6141;
  wire [31:0] _EVAL_1303;
  wire  _EVAL_649;
  wire  _EVAL_1599;
  wire [31:0] _EVAL_2969;
  wire  _EVAL_414;
  wire  _EVAL_3717;
  wire [31:0] _EVAL_3704;
  wire  _EVAL_2983;
  wire  _EVAL_1372;
  wire [31:0] _EVAL_3038;
  wire  _EVAL_492;
  wire  _EVAL_2755;
  wire  _EVAL_3982;
  wire  _EVAL_4568;
  wire  _EVAL_5198;
  wire [31:0] _EVAL_207;
  wire  _EVAL_1941;
  wire  _EVAL_4952;
  wire  _EVAL_3303;
  wire [31:0] _EVAL_790;
  wire  _EVAL_5550;
  wire  _EVAL_4137;
  wire [31:0] _EVAL_4789;
  wire  _EVAL_5021;
  wire  _EVAL_4805;
  wire [31:0] _EVAL_2731;
  wire  _EVAL_5216;
  wire  _EVAL_886;
  wire  _EVAL_5321;
  wire [31:0] _EVAL_3968;
  wire  _EVAL_2159;
  wire [31:0] _EVAL_3114;
  wire  _EVAL_2954;
  wire  _EVAL_2573;
  wire [31:0] _EVAL_3221;
  wire  _EVAL_3530;
  wire  _EVAL_1508;
  wire  _EVAL_5433;
  wire  _EVAL_3276;
  wire  _EVAL_1274;
  wire  _EVAL_1547;
  wire  _EVAL_2081;
  wire  _EVAL_5703;
  wire  _EVAL_3718;
  wire  _EVAL_1898;
  wire  _EVAL_636;
  wire  _EVAL_5987;
  wire  _EVAL_2605;
  wire [31:0] _EVAL_5118;
  wire  _EVAL_5673;
  wire  _EVAL_3510;
  wire [31:0] _EVAL_1231;
  wire  _EVAL_2556;
  wire  _EVAL_2275;
  wire [31:0] _EVAL_5939;
  wire  _EVAL_1580;
  wire  _EVAL_491;
  wire [31:0] _EVAL_1309;
  wire  _EVAL_4768;
  wire  _EVAL_5576;
  wire  _EVAL_5973;
  wire  _EVAL_4556;
  wire [31:0] _EVAL_2121;
  wire  _EVAL_423;
  wire  _EVAL_5345;
  wire  _EVAL_237;
  wire  _EVAL_3479;
  wire  _EVAL_5557;
  wire  _EVAL_3066;
  wire  _EVAL_3989;
  wire  _EVAL_6035;
  wire  _EVAL_5746;
  wire [31:0] _EVAL_2059;
  wire  _EVAL_5614;
  wire  _EVAL_5645;
  wire  _EVAL_5889;
  wire  _EVAL_1454;
  wire  _EVAL_4452;
  wire  _EVAL_5840;
  wire [31:0] _EVAL_3331;
  wire  _EVAL_6107;
  wire  _EVAL_6103;
  wire  _EVAL_1760;
  wire [31:0] _EVAL_2018;
  wire  _EVAL_1441;
  wire  _EVAL_5424;
  wire [31:0] _EVAL_2604;
  wire  _EVAL_751;
  wire  _EVAL_3485;
  wire [31:0] _EVAL_2184;
  wire  _EVAL_5659;
  wire  _EVAL_2523;
  wire  _EVAL_3723;
  wire  _EVAL_2278;
  wire [31:0] _EVAL_4422;
  wire  _EVAL_4143;
  wire  _EVAL_2352;
  wire  _EVAL_1482;
  wire  _EVAL_5942;
  wire  _EVAL_5737;
  wire  _EVAL_684;
  wire  _EVAL_452;
  wire  _EVAL_4883;
  wire  _EVAL_3433;
  wire [31:0] _EVAL_5916;
  wire  _EVAL_1589;
  wire [31:0] _EVAL_1623;
  wire  _EVAL_496;
  wire  _EVAL_2850;
  wire [31:0] _EVAL_2761;
  wire [31:0] _EVAL_5038;
  wire  _EVAL_3782;
  wire  _EVAL_3974;
  wire [31:0] _EVAL_904;
  wire  _EVAL_2670;
  wire  _EVAL_3039;
  wire  _EVAL_1624;
  wire  _EVAL_1737;
  wire  _EVAL_5475;
  wire [31:0] _EVAL_1791;
  wire [4:0] _EVAL_4304;
  wire [4:0] _EVAL_3720;
  wire [4:0] _EVAL_6138;
  wire [4:0] _EVAL_5843;
  wire [4:0] _EVAL_2561;
  wire [31:0] _EVAL_2313;
  wire  _EVAL_4852;
  wire [31:0] _EVAL_1489;
  wire  _EVAL_2737;
  wire  _EVAL_3735;
  wire [31:0] _EVAL_1588;
  wire  _EVAL_324;
  wire  _EVAL_4435;
  wire [31:0] _EVAL_3481;
  wire  _EVAL_3535;
  wire [31:0] _EVAL_6049;
  wire  _EVAL_3349;
  wire  _EVAL_5019;
  wire  _EVAL_5042;
  wire  _EVAL_4976;
  wire  _EVAL_986;
  wire  _EVAL_402;
  wire  _EVAL_2683;
  wire  _EVAL_4135;
  wire [31:0] _EVAL_5147;
  wire  _EVAL_4198;
  wire  _EVAL_1594;
  wire [31:0] _EVAL_3178;
  wire  _EVAL_5081;
  wire  _EVAL_4557;
  wire  _EVAL_5888;
  wire  _EVAL_5652;
  wire [31:0] _EVAL_1208;
  wire  _EVAL_5768;
  wire  _EVAL_5975;
  wire  _EVAL_4184;
  wire  _EVAL_3420;
  wire  _EVAL_5394;
  wire  _EVAL_3624;
  wire  _EVAL_4902;
  wire [31:0] _EVAL_3002;
  wire [31:0] _EVAL_5336;
  wire [31:0] _EVAL_5497;
  wire  _EVAL_2916;
  wire  _EVAL_4970;
  wire [31:0] _EVAL_1047;
  wire  _EVAL_4828;
  wire  _EVAL_1319;
  wire  _EVAL_4485;
  wire  _EVAL_3079;
  wire  _EVAL_4667;
  wire [31:0] _EVAL_721;
  wire  _EVAL_1762;
  wire [31:0] _EVAL_4802;
  wire  _EVAL_1513;
  wire  _EVAL_5807;
  wire [31:0] _EVAL_3694;
  wire  _EVAL_1490;
  wire  _EVAL_4173;
  wire [31:0] _EVAL_1097;
  wire  _EVAL_824;
  wire  _EVAL_3495;
  wire [31:0] _EVAL_4691;
  wire  _EVAL_3751;
  wire  _EVAL_5413;
  wire  _EVAL_277;
  wire  _EVAL_2722;
  wire  _EVAL_4145;
  wire [31:0] _EVAL_860;
  wire  _EVAL_4049;
  wire [31:0] _EVAL_5884;
  wire  _EVAL_5239;
  wire  _EVAL_3917;
  wire  _EVAL_2131;
  wire  _EVAL_289;
  wire  _EVAL_854;
  wire [31:0] _EVAL_5660;
  wire  _EVAL_659;
  wire  _EVAL_5957;
  wire  _EVAL_5537;
  wire  _EVAL_5605;
  wire [31:0] _EVAL_2271;
  wire  _EVAL_1991;
  wire  _EVAL_5162;
  wire  _EVAL_4024;
  wire  _EVAL_2257;
  wire  _EVAL_3438;
  wire  _EVAL_4656;
  wire [31:0] _EVAL_2280;
  wire  _EVAL_513;
  wire  _EVAL_5362;
  wire  _EVAL_1519;
  wire  _EVAL_2789;
  wire  _EVAL_2042;
  wire  _EVAL_2834;
  wire  _EVAL_5461;
  wire [6:0] _EVAL_1527;
  wire [6:0] _EVAL_2295;
  wire [6:0] _EVAL_4576;
  wire [6:0] _EVAL_1419;
  wire [6:0] _EVAL_5848;
  wire [6:0] _EVAL_5915;
  wire [6:0] _EVAL_4759;
  wire [6:0] _EVAL_2967;
  wire [6:0] _EVAL_594;
  wire [6:0] _EVAL_4694;
  wire [6:0] _EVAL_3762;
  wire [6:0] _EVAL_1836;
  wire [6:0] _EVAL_5800;
  wire [6:0] _EVAL_3430;
  wire [6:0] _EVAL_2324;
  wire [6:0] _EVAL_1918;
  wire [6:0] _EVAL_4009;
  wire [6:0] _EVAL_4152;
  wire [6:0] _EVAL_1552;
  wire [6:0] _EVAL_1066;
  wire [6:0] _EVAL_1353;
  wire [6:0] _EVAL_468;
  wire  _EVAL_797;
  wire [31:0] _EVAL_575;
  wire  _EVAL_4643;
  wire  _EVAL_1753;
  wire  _EVAL_2715;
  wire  _EVAL_3812;
  wire  _EVAL_5941;
  wire  _EVAL_926;
  wire  _EVAL_6000;
  wire [31:0] _EVAL_3953;
  wire  _EVAL_461;
  wire  _EVAL_4855;
  wire  _EVAL_2818;
  wire  _EVAL_3681;
  wire  _EVAL_4083;
  wire [31:0] _EVAL_779;
  wire  _EVAL_3746;
  wire  _EVAL_4885;
  wire [31:0] _EVAL_3860;
  wire  _EVAL_4540;
  wire  _EVAL_3347;
  wire  _EVAL_5547;
  wire  _EVAL_3814;
  wire  _EVAL_5995;
  wire  _EVAL_6007;
  wire  _EVAL_2567;
  wire  _EVAL_4182;
  wire  _EVAL_316;
  wire  _EVAL_5122;
  wire  _EVAL_5273;
  wire  _EVAL_2035;
  wire  _EVAL_5951;
  wire [31:0] _EVAL_1402;
  wire  _EVAL_2529;
  wire [31:0] _EVAL_5517;
  wire [4:0] _EVAL_5352;
  wire  _EVAL_2330;
  wire  _EVAL_1556;
  wire [4:0] _EVAL_3990;
  wire [4:0] _EVAL_748;
  wire  _EVAL_6017;
  wire  _EVAL_3352;
  wire [31:0] _EVAL_2443;
  wire  _EVAL_2468;
  wire  _EVAL_3491;
  wire  _EVAL_855;
  wire  _EVAL_1326;
  wire  _EVAL_5711;
  wire  _EVAL_1268;
  wire [31:0] _EVAL_2490;
  wire  _EVAL_3502;
  wire  _EVAL_1769;
  wire  _EVAL_1586;
  wire  _EVAL_3030;
  wire  _EVAL_3189;
  wire [31:0] _EVAL_3855;
  wire  _EVAL_5249;
  wire  _EVAL_3670;
  wire  _EVAL_2800;
  wire  _EVAL_2060;
  wire [31:0] _EVAL_3631;
  wire  _EVAL_5096;
  wire  _EVAL_5640;
  wire [31:0] _EVAL_2658;
  wire  _EVAL_2043;
  wire  _EVAL_291;
  wire  _EVAL_2318;
  wire  _EVAL_3288;
  wire  _EVAL_4443;
  wire [31:0] _EVAL_6002;
  wire  _EVAL_2177;
  wire  _EVAL_856;
  wire  _EVAL_3265;
  wire  _EVAL_971;
  wire  _EVAL_2718;
  wire  _EVAL_5275;
  wire  _EVAL_2621;
  wire  _EVAL_2358;
  wire  _EVAL_6028;
  wire [31:0] _EVAL_1377;
  wire  _EVAL_3816;
  wire  _EVAL_1421;
  wire  _EVAL_5179;
  wire  _EVAL_265;
  wire  _EVAL_2140;
  wire  _EVAL_3872;
  wire  _EVAL_3884;
  wire  _EVAL_2886;
  wire  _EVAL_3619;
  wire [4:0] _EVAL_633;
  wire [4:0] _EVAL_5368;
  wire  _EVAL_976;
  wire  _EVAL_3503;
  wire  _EVAL_1062;
  wire  _EVAL_5434;
  wire  _EVAL_5498;
  wire  _EVAL_3819;
  wire  _EVAL_5594;
  wire  _EVAL_2820;
  wire  _EVAL_5651;
  wire  _EVAL_2117;
  wire  _EVAL_1470;
  wire  _EVAL_4635;
  wire  _EVAL_5047;
  wire  _EVAL_672;
  wire  _EVAL_4997;
  wire  _EVAL_2203;
  wire  _EVAL_4326;
  wire [4:0] _EVAL_5291;
  wire [4:0] _EVAL_1054;
  wire [4:0] _EVAL_4067;
  wire [4:0] _EVAL_1852;
  wire [4:0] _EVAL_5484;
  wire [4:0] _EVAL_3945;
  wire [2:0] _EVAL_3314;
  wire [31:0] _EVAL_4116;
  wire  _EVAL_3294;
  wire [31:0] _EVAL_4896;
  wire  _EVAL_4727;
  wire  _EVAL_3672;
  wire  _EVAL_1871;
  wire  _EVAL_1957;
  wire  _EVAL_1341;
  wire  _EVAL_2145;
  wire  _EVAL_1085;
  wire  _EVAL_2186;
  wire  _EVAL_1033;
  wire  _EVAL_2531;
  wire  _EVAL_3944;
  wire  _EVAL_3648;
  wire  _EVAL_1959;
  wire  _EVAL_1106;
  wire  _EVAL_2799;
  wire  _EVAL_691;
  wire  _EVAL_6015;
  wire  _EVAL_2205;
  wire  _EVAL_1080;
  wire [31:0] _EVAL_1579;
  wire  _EVAL_3585;
  wire  _EVAL_6018;
  wire [31:0] _EVAL_3463;
  wire  _EVAL_1695;
  wire  _EVAL_5708;
  wire  _EVAL_4992;
  wire  _EVAL_4652;
  wire  _EVAL_5559;
  wire  _EVAL_1176;
  wire  _EVAL_1150;
  wire  _EVAL_4895;
  wire  _EVAL_5886;
  wire [31:0] _EVAL_1488;
  wire  _EVAL_1376;
  wire  _EVAL_187;
  wire  _EVAL_5013;
  wire  _EVAL_1044;
  wire  _EVAL_6048;
  wire  _EVAL_1539;
  wire [2:0] _EVAL_2044;
  wire [2:0] _EVAL_3021;
  wire [2:0] _EVAL_3546;
  wire [2:0] _EVAL_4234;
  wire [2:0] _EVAL_1266;
  wire [2:0] _EVAL_5656;
  wire [2:0] _EVAL_1391;
  wire [2:0] _EVAL_3249;
  wire  _EVAL_347;
  wire [31:0] _EVAL_2484;
  wire  _EVAL_2207;
  wire  _EVAL_3411;
  wire  _EVAL_483;
  wire  _EVAL_4775;
  wire  _EVAL_5330;
  wire [31:0] _EVAL_3901;
  wire  _EVAL_3116;
  wire  _EVAL_4146;
  wire  _EVAL_1476;
  wire  _EVAL_4283;
  wire  _EVAL_2617;
  wire  _EVAL_5553;
  wire  _EVAL_2377;
  wire [31:0] _EVAL_168;
  wire  _EVAL_3475;
  wire [2:0] _EVAL_3852;
  wire [4:0] _EVAL_1983;
  wire  _EVAL_551;
  wire  _EVAL_3646;
  wire [2:0] _EVAL_2751;
  wire [2:0] _EVAL_382;
  wire [2:0] _EVAL_3246;
  wire [2:0] _EVAL_5960;
  wire [2:0] _EVAL_3064;
  wire [2:0] _EVAL_538;
  wire [2:0] _EVAL_4455;
  wire  _EVAL_245;
  wire  _EVAL_908;
  wire  _EVAL_2896;
  wire  _EVAL_4131;
  wire  _EVAL_4543;
  wire  _EVAL_301;
  wire  _EVAL_3452;
  wire  _EVAL_3421;
  wire  _EVAL_3789;
  wire  _EVAL_3928;
  wire  _EVAL_5010;
  wire  _EVAL_5051;
  wire  _EVAL_3949;
  wire  _EVAL_256;
  wire  _EVAL_1279;
  wire  _EVAL_4820;
  wire  _EVAL_2399;
  wire  _EVAL_5642;
  wire [31:0] _EVAL_4972;
  wire  _EVAL_3190;
  wire  _EVAL_405;
  wire  _EVAL_1307;
  wire  _EVAL_674;
  wire [31:0] _EVAL_5700;
  wire  _EVAL_2994;
  wire  _EVAL_1823;
  wire  _EVAL_2551;
  wire  _EVAL_3431;
  wire  _EVAL_3971;
  wire  _EVAL_1115;
  wire  _EVAL_4358;
  wire  _EVAL_4342;
  wire  _EVAL_1752;
  wire  _EVAL_4588;
  wire  _EVAL_3531;
  wire  _EVAL_4139;
  wire  _EVAL_1351;
  wire  _EVAL_2727;
  wire  _EVAL_1166;
  wire [31:0] _EVAL_3914;
  wire [31:0] _EVAL_4311;
  wire  _EVAL_1867;
  wire  _EVAL_5427;
  wire  _EVAL_1254;
  wire  _EVAL_2080;
  wire  _EVAL_5780;
  wire  _EVAL_1500;
  wire  _EVAL_605;
  wire  _EVAL_416;
  wire [31:0] _EVAL_2981;
  wire  _EVAL_6041;
  wire  _EVAL_5774;
  wire  _EVAL_732;
  wire  _EVAL_3587;
  wire  _EVAL_5367;
  wire [31:0] _EVAL_4979;
  wire  _EVAL_435;
  wire  _EVAL_312;
  wire  _EVAL_804;
  wire [31:0] _EVAL_3838;
  wire  _EVAL_396;
  wire  _EVAL_4586;
  wire  _EVAL_355;
  wire [31:0] _EVAL_4782;
  wire  _EVAL_3302;
  wire  _EVAL_921;
  wire  _EVAL_3489;
  wire  _EVAL_4203;
  wire  _EVAL_1466;
  wire  _EVAL_4488;
  wire [31:0] _EVAL_1862;
  wire  _EVAL_3786;
  wire  _EVAL_2125;
  wire  _EVAL_4786;
  wire  _EVAL_2548;
  wire  _EVAL_3356;
  wire  _EVAL_4713;
  wire  _EVAL_1687;
  wire  _EVAL_2515;
  wire  _EVAL_3177;
  wire  _EVAL_834;
  wire  _EVAL_4127;
  wire  _EVAL_2535;
  wire  _EVAL_5761;
  wire  _EVAL_3873;
  wire  _EVAL_4276;
  wire  _EVAL_5644;
  wire  _EVAL_2073;
  wire  _EVAL_3833;
  wire  _EVAL_4874;
  wire  _EVAL_1233;
  wire  _EVAL_3494;
  wire  _EVAL_3941;
  wire  _EVAL_3561;
  wire  _EVAL_3492;
  wire  _EVAL_3400;
  wire  _EVAL_3818;
  wire [1:0] _EVAL_1118;
  wire  _EVAL_2889;
  wire  _EVAL_5242;
  wire [31:0] _EVAL_3853;
  wire  _EVAL_3312;
  wire  _EVAL_702;
  wire  _EVAL_4940;
  wire [4:0] _EVAL_4742;
  wire [4:0] _EVAL_2037;
  wire  _EVAL_2830;
  wire  _EVAL_6104;
  wire [31:0] _EVAL_2957;
  wire  _EVAL_2847;
  wire  _EVAL_2903;
  wire  _EVAL_5837;
  wire  _EVAL_2691;
  wire  _EVAL_2423;
  wire  _EVAL_309;
  wire  _EVAL_1138;
  wire  _EVAL_1425;
  wire  _EVAL_1444;
  wire  _EVAL_1706;
  wire  _EVAL_3935;
  wire  _EVAL_1387;
  wire  _EVAL_4494;
  wire [31:0] _EVAL_943;
  wire  _EVAL_4866;
  wire  _EVAL_3756;
  wire  _EVAL_506;
  wire [2:0] _EVAL_5552;
  wire  _EVAL_4720;
  wire  _EVAL_5669;
  wire  _EVAL_3733;
  wire  _EVAL_5769;
  wire  _EVAL_5534;
  wire  _EVAL_5409;
  wire  _EVAL_966;
  wire [4:0] _EVAL_6033;
  wire [4:0] _EVAL_4847;
  wire [4:0] _EVAL_3223;
  wire [3:0] _EVAL_2167;
  wire [31:0] _EVAL_5722;
  wire [6:0] _EVAL_3793;
  wire [6:0] _EVAL_5869;
  wire [6:0] _EVAL_829;
  wire [6:0] _EVAL_1906;
  wire  _EVAL_796;
  wire  _EVAL_2199;
  wire  _EVAL_2564;
  wire  _EVAL_1572;
  wire  _EVAL_5372;
  wire [2:0] _EVAL_3960;
  wire [2:0] _EVAL_4321;
  wire [4:0] _EVAL_4703;
  wire [4:0] _EVAL_5953;
  wire  _EVAL_4738;
  wire  _EVAL_3035;
  wire [4:0] _EVAL_4917;
  wire  _EVAL_4884;
  wire  _EVAL_4584;
  wire  _EVAL_4178;
  wire  _EVAL_2040;
  wire  _EVAL_3469;
  wire  _EVAL_1711;
  wire  _EVAL_4475;
  wire  _EVAL_3698;
  wire [4:0] _EVAL_2959;
  wire [4:0] _EVAL_685;
  wire  _EVAL_1884;
  wire  _EVAL_4099;
  wire [6:0] _EVAL_3072;
  wire [6:0] _EVAL_588;
  wire [6:0] _EVAL_3500;
  wire [6:0] _EVAL_3240;
  wire [3:0] _EVAL_2796;
  wire  _EVAL_1406;
  wire  _EVAL_4097;
  wire  _EVAL_2010;
  wire  _EVAL_3339;
  wire  _EVAL_1052;
  wire [2:0] _EVAL_200;
  wire  _EVAL_4179;
  wire  _EVAL_257;
  wire [6:0] _EVAL_709;
  wire [6:0] _EVAL_1456;
  wire [6:0] _EVAL_5765;
  wire  _EVAL_6116;
  wire [6:0] _EVAL_2887;
  wire [6:0] _EVAL_2575;
  wire  _EVAL_5079;
  wire  _EVAL_3128;
  wire  _EVAL_611;
  wire  _EVAL_4996;
  wire  _EVAL_4522;
  wire  _EVAL_4280;
  wire  _EVAL_422;
  wire  _EVAL_5707;
  wire [127:0] _EVAL_1530;
  wire [4:0] _EVAL_3383;
  wire  _EVAL_2004;
  wire  _EVAL_818;
  wire  _EVAL_4967;
  wire  _EVAL_1740;
  wire [3:0] _EVAL_4265;
  wire  _EVAL_2997;
  wire  _EVAL_4335;
  wire  _EVAL_4033;
  wire  _EVAL_4431;
  wire  _EVAL_5379;
  wire  _EVAL_4077;
  wire  _EVAL_2380;
  wire  _EVAL_3862;
  wire  _EVAL_1127;
  wire [4:0] _EVAL_5308;
  wire [4:0] _EVAL_1190;
  wire  _EVAL_3073;
  wire  _EVAL_1813;
  wire  _EVAL_1447;
  wire  _EVAL_1748;
  wire  _EVAL_3324;
  wire  _EVAL_4122;
  wire  _EVAL_5666;
  wire [4:0] _EVAL_970;
  wire [8:0] _EVAL_6102;
  wire [4:0] _EVAL_3959;
  wire  _EVAL_4966;
  wire  _EVAL_1765;
  wire  _EVAL_2721;
  wire  _EVAL_1758;
  wire  _EVAL_5591;
  wire  _EVAL_5045;
  wire  _EVAL_724;
  wire  _EVAL_1158;
  wire  _EVAL_3801;
  wire  _EVAL_440;
  wire [31:0] _EVAL_4533;
  wire  _EVAL_6098;
  wire  _EVAL_2743;
  wire  _EVAL_3918;
  wire  _EVAL_1694;
  wire  _EVAL_1896;
  wire  _EVAL_3359;
  wire [3:0] _EVAL_5212;
  wire [3:0] _EVAL_2869;
  wire  _EVAL_2724;
  wire  _EVAL_2962;
  assign _EVAL_2666 = _EVAL_33[63:48];
  assign _EVAL_4292 = _EVAL_33[47:32];
  assign _EVAL_5159 = _EVAL_33[31:16];
  assign _EVAL_3455 = {_EVAL_2666,_EVAL_4292,_EVAL_5159};
  assign _EVAL_4071 = _EVAL_3455[15:13];
  assign _EVAL_4669 = _EVAL_4071 == 3'h7;
  assign _EVAL_241 = _EVAL_3455[5];
  assign _EVAL_4901 = _EVAL_3455[12:10];
  assign _EVAL_2996 = _EVAL_3455[6];
  assign _EVAL_1346 = {_EVAL_241,_EVAL_4901,_EVAL_2996,2'h0};
  assign _EVAL_1939 = _EVAL_1346[6:5];
  assign _EVAL_3926 = _EVAL_3455[4:2];
  assign _EVAL_4872 = _EVAL_3455[9:7];
  assign _EVAL_5992 = _EVAL_1346[4:0];
  assign _EVAL_1643 = {_EVAL_1939,2'h1,_EVAL_3926,2'h1,_EVAL_4872,3'h2,_EVAL_5992,7'h27};
  assign _EVAL_2288 = _EVAL_4071 == 3'h6;
  assign _EVAL_4563 = {_EVAL_1939,2'h1,_EVAL_3926,2'h1,_EVAL_4872,3'h2,_EVAL_5992,7'h23};
  assign _EVAL_453 = _EVAL_4071 == 3'h5;
  assign _EVAL_5278 = _EVAL_3455[6:5];
  assign _EVAL_5928 = {_EVAL_5278,_EVAL_4901,3'h0};
  assign _EVAL_2821 = _EVAL_5928[7:5];
  assign _EVAL_1749 = _EVAL_5928[4:0];
  assign _EVAL_3859 = {_EVAL_2821,2'h1,_EVAL_3926,2'h1,_EVAL_4872,3'h3,_EVAL_1749,7'h27};
  assign _EVAL_936 = _EVAL_4071 == 3'h4;
  assign _EVAL_3053 = {_EVAL_1939,2'h1,_EVAL_3926,2'h1,_EVAL_4872,3'h0,_EVAL_5992,7'h27};
  assign _EVAL_1674 = _EVAL_4071 == 3'h3;
  assign _EVAL_3821 = {_EVAL_241,_EVAL_4901,_EVAL_2996,2'h0,2'h1,_EVAL_4872,3'h2,2'h1,_EVAL_3926,7'h7};
  assign _EVAL_597 = _EVAL_4071 == 3'h2;
  assign _EVAL_2991 = {_EVAL_241,_EVAL_4901,_EVAL_2996,2'h0,2'h1,_EVAL_4872,3'h2,2'h1,_EVAL_3926,7'h3};
  assign _EVAL_5755 = _EVAL_4071 == 3'h1;
  assign _EVAL_2246 = {_EVAL_5278,_EVAL_4901,3'h0,2'h1,_EVAL_4872,3'h3,2'h1,_EVAL_3926,7'h7};
  assign _EVAL_4532 = _EVAL_3455[10:7];
  assign _EVAL_5956 = _EVAL_3455[12:11];
  assign _EVAL_1848 = {_EVAL_4532,_EVAL_5956,_EVAL_241,_EVAL_2996,2'h0,5'h2,3'h0,2'h1,_EVAL_3926,7'h13};
  assign _EVAL_812 = _EVAL_5755 ? {{2'd0}, _EVAL_2246} : _EVAL_1848;
  assign _EVAL_173 = _EVAL_597 ? {{3'd0}, _EVAL_2991} : _EVAL_812;
  assign _EVAL_2725 = _EVAL_1674 ? {{3'd0}, _EVAL_3821} : _EVAL_173;
  assign _EVAL_2541 = _EVAL_936 ? {{3'd0}, _EVAL_3053} : _EVAL_2725;
  assign _EVAL_4645 = _EVAL_453 ? {{2'd0}, _EVAL_3859} : _EVAL_2541;
  assign _EVAL_3736 = _EVAL_2288 ? {{3'd0}, _EVAL_4563} : _EVAL_4645;
  assign _EVAL_3595 = _EVAL_4669 ? {{3'd0}, _EVAL_1643} : _EVAL_3736;
  assign _EVAL_2164 = {2'h0,_EVAL_3595};
  assign _EVAL_1690 = _EVAL_2164 & 32'h207f;
  assign _EVAL_4293 = _EVAL_1690 == 32'h3;
  assign _EVAL_5077 = _EVAL_2164 & 32'h607f;
  assign _EVAL_3471 = _EVAL_5077 == 32'hf;
  assign _EVAL_2314 = _EVAL_4293 | _EVAL_3471;
  assign _EVAL_877 = _EVAL_2164 & 32'h5f;
  assign _EVAL_4098 = _EVAL_877 == 32'h17;
  assign _EVAL_1135 = _EVAL_2314 | _EVAL_4098;
  assign _EVAL_1286 = _EVAL_2164 & 32'hfc00007f;
  assign _EVAL_4327 = _EVAL_1286 == 32'h33;
  assign _EVAL_2655 = _EVAL_1135 | _EVAL_4327;
  assign _EVAL_1215 = _EVAL_2164 & 32'hbe00707f;
  assign _EVAL_5365 = _EVAL_1215 == 32'h33;
  assign _EVAL_2407 = _EVAL_2655 | _EVAL_5365;
  assign _EVAL_5699 = _EVAL_2164 & 32'h6000073;
  assign _EVAL_3701 = _EVAL_5699 == 32'h43;
  assign _EVAL_4420 = _EVAL_2407 | _EVAL_3701;
  assign _EVAL_3778 = _EVAL_2164 & 32'he600007f;
  assign _EVAL_1131 = _EVAL_3778 == 32'h53;
  assign _EVAL_5931 = _EVAL_4420 | _EVAL_1131;
  assign _EVAL_764 = _EVAL_2164 & 32'h707b;
  assign _EVAL_3234 = _EVAL_764 == 32'h63;
  assign _EVAL_447 = _EVAL_5931 | _EVAL_3234;
  assign _EVAL_6097 = _EVAL_2164 & 32'h7f;
  assign _EVAL_4305 = _EVAL_6097 == 32'h6f;
  assign _EVAL_5238 = _EVAL_447 | _EVAL_4305;
  assign _EVAL_645 = _EVAL_2164 & 32'hffefffff;
  assign _EVAL_836 = _EVAL_645 == 32'h73;
  assign _EVAL_4330 = _EVAL_5238 | _EVAL_836;
  assign _EVAL_4039 = _EVAL_2164 & 32'hfe00305f;
  assign _EVAL_367 = _EVAL_4039 == 32'h1013;
  assign _EVAL_210 = _EVAL_4330 | _EVAL_367;
  assign _EVAL_3250 = _EVAL_2164 & 32'h705b;
  assign _EVAL_1116 = _EVAL_3250 == 32'h2003;
  assign _EVAL_2096 = _EVAL_210 | _EVAL_1116;
  assign _EVAL_4777 = _EVAL_1690 == 32'h2013;
  assign _EVAL_2982 = _EVAL_2096 | _EVAL_4777;
  assign _EVAL_3891 = _EVAL_2164 & 32'h1800707f;
  assign _EVAL_687 = _EVAL_3891 == 32'h202f;
  assign _EVAL_1570 = _EVAL_2982 | _EVAL_687;
  assign _EVAL_6053 = _EVAL_1690 == 32'h2073;
  assign _EVAL_1771 = _EVAL_1570 | _EVAL_6053;
  assign _EVAL_5477 = _EVAL_2164 & 32'hbe00705f;
  assign _EVAL_3235 = _EVAL_5477 == 32'h5013;
  assign _EVAL_3436 = _EVAL_1771 | _EVAL_3235;
  assign _EVAL_2614 = _EVAL_2164 & 32'he800707f;
  assign _EVAL_4022 = _EVAL_2614 == 32'h800202f;
  assign _EVAL_4755 = _EVAL_3436 | _EVAL_4022;
  assign _EVAL_3440 = _EVAL_2164 & 32'hf9f0707f;
  assign _EVAL_3096 = _EVAL_3440 == 32'h1000202f;
  assign _EVAL_2790 = _EVAL_4755 | _EVAL_3096;
  assign _EVAL_2778 = _EVAL_2164 & 32'hdfffffff;
  assign _EVAL_2477 = _EVAL_2778 == 32'h10500073;
  assign _EVAL_4155 = _EVAL_2790 | _EVAL_2477;
  assign _EVAL_171 = _EVAL_2164 & 32'hf600607f;
  assign _EVAL_262 = _EVAL_171 == 32'h20000053;
  assign _EVAL_4260 = _EVAL_4155 | _EVAL_262;
  assign _EVAL_2457 = _EVAL_2164 & 32'h7e00607f;
  assign _EVAL_3049 = _EVAL_2457 == 32'h20000053;
  assign _EVAL_3000 = _EVAL_4260 | _EVAL_3049;
  assign _EVAL_5743 = _EVAL_2164 & 32'h7e00507f;
  assign _EVAL_3229 = _EVAL_5743 == 32'h20000053;
  assign _EVAL_2362 = _EVAL_3000 | _EVAL_3229;
  assign _EVAL_2629 = _EVAL_91;
  assign _EVAL_2143 = _EVAL_19;
  assign _EVAL_5731 = {_EVAL_2629,1'h0,1'h0,_EVAL_2143};
  assign _EVAL_4188 = _EVAL_9;
  assign _EVAL_3997 = _EVAL_5731 >> _EVAL_4188;
  assign _EVAL_3588 = _EVAL_33[15:0];
  assign _EVAL_654 = {_EVAL_2666,_EVAL_4292,_EVAL_5159,_EVAL_3588,_EVAL_5094};
  assign _EVAL_4702 = _EVAL_654[31:0];
  assign _EVAL_4125 = _EVAL_4702 & 32'h7e00607f;
  assign _EVAL_2935 = _EVAL_654[8:7];
  assign _EVAL_2290 = _EVAL_3455[12:2];
  assign _EVAL_3023 = _EVAL_2290 != 11'h0;
  assign _EVAL_2277 = _EVAL_4702 & 32'h2000040;
  assign _EVAL_808 = _EVAL_654[15:13];
  assign _EVAL_1088 = _EVAL_808 == 3'h7;
  assign _EVAL_3841 = _EVAL_654[12:9];
  assign _EVAL_738 = {_EVAL_2935,_EVAL_3841,2'h0};
  assign _EVAL_3877 = _EVAL_738[7:5];
  assign _EVAL_1321 = _EVAL_654[6:2];
  assign _EVAL_694 = _EVAL_738[4:0];
  assign _EVAL_3043 = {_EVAL_3877,_EVAL_1321,5'h2,3'h2,_EVAL_694,7'h27};
  assign _EVAL_537 = _EVAL_808 == 3'h6;
  assign _EVAL_5721 = {_EVAL_3877,_EVAL_1321,5'h2,3'h2,_EVAL_694,7'h23};
  assign _EVAL_1378 = _EVAL_808 == 3'h5;
  assign _EVAL_4771 = _EVAL_654[9:7];
  assign _EVAL_2483 = _EVAL_654[12:10];
  assign _EVAL_5892 = {_EVAL_4771,_EVAL_2483,3'h0};
  assign _EVAL_4114 = _EVAL_5892[8:5];
  assign _EVAL_4538 = _EVAL_5892[4:0];
  assign _EVAL_3320 = {_EVAL_4114,_EVAL_1321,5'h2,3'h3,_EVAL_4538,7'h27};
  assign _EVAL_4440 = _EVAL_808 == 3'h4;
  assign _EVAL_3082 = _EVAL_654[12];
  assign _EVAL_2173 = _EVAL_1321 != 5'h0;
  assign _EVAL_4094 = _EVAL_654[11:7];
  assign _EVAL_759 = {_EVAL_1321,_EVAL_4094,3'h0,_EVAL_4094,7'h33};
  assign _EVAL_1360 = _EVAL_4094 != 5'h0;
  assign _EVAL_4100 = {_EVAL_1321,_EVAL_4094,3'h0,12'he7};
  assign _EVAL_2188 = {_EVAL_1321,_EVAL_4094,3'h0,12'h67};
  assign _EVAL_3216 = _EVAL_2188[24:7];
  assign _EVAL_938 = {_EVAL_3216,7'h73};
  assign _EVAL_448 = _EVAL_938 | 25'h100000;
  assign _EVAL_1277 = _EVAL_1360 ? _EVAL_4100 : _EVAL_448;
  assign _EVAL_4791 = _EVAL_2173 ? _EVAL_759 : _EVAL_1277;
  assign _EVAL_1610 = {_EVAL_1321,5'h0,3'h4,_EVAL_4094,7'h33};
  assign _EVAL_947 = _EVAL_2173 ? _EVAL_1610 : _EVAL_2188;
  assign _EVAL_1568 = _EVAL_3082 ? _EVAL_4791 : _EVAL_947;
  assign _EVAL_761 = _EVAL_808 == 3'h3;
  assign _EVAL_4347 = _EVAL_654[3:2];
  assign _EVAL_2114 = _EVAL_654[6:4];
  assign _EVAL_3139 = {_EVAL_4347,_EVAL_3082,_EVAL_2114,2'h0,5'h2,3'h2,_EVAL_4094,7'h7};
  assign _EVAL_5989 = _EVAL_808 == 3'h2;
  assign _EVAL_3138 = {_EVAL_4347,_EVAL_3082,_EVAL_2114,2'h0,5'h2,3'h2,_EVAL_4094,7'h3};
  assign _EVAL_3016 = _EVAL_808 == 3'h1;
  assign _EVAL_2231 = _EVAL_654[4:2];
  assign _EVAL_4575 = _EVAL_654[6:5];
  assign _EVAL_2397 = {_EVAL_2231,_EVAL_3082,_EVAL_4575,3'h0,5'h2,3'h3,_EVAL_4094,7'h7};
  assign _EVAL_1481 = {_EVAL_3082,_EVAL_1321,_EVAL_4094,3'h1,_EVAL_4094,7'h13};
  assign _EVAL_2014 = _EVAL_3016 ? _EVAL_2397 : {{3'd0}, _EVAL_1481};
  assign _EVAL_2350 = _EVAL_5989 ? {{1'd0}, _EVAL_3138} : _EVAL_2014;
  assign _EVAL_3048 = _EVAL_761 ? {{1'd0}, _EVAL_3139} : _EVAL_2350;
  assign _EVAL_583 = _EVAL_4440 ? {{4'd0}, _EVAL_1568} : _EVAL_3048;
  assign _EVAL_327 = _EVAL_1378 ? _EVAL_3320 : _EVAL_583;
  assign _EVAL_2482 = _EVAL_537 ? {{1'd0}, _EVAL_5721} : _EVAL_327;
  assign _EVAL_4396 = _EVAL_1088 ? {{1'd0}, _EVAL_3043} : _EVAL_2482;
  assign _EVAL_3078 = {3'h0,_EVAL_4396};
  assign _EVAL_4897 = _EVAL_3078 & 32'h207f;
  assign _EVAL_4008 = _EVAL_4897 == 32'h3;
  assign _EVAL_2032 = _EVAL_3078 & 32'h607f;
  assign _EVAL_1754 = _EVAL_2032 == 32'hf;
  assign _EVAL_4659 = _EVAL_4008 | _EVAL_1754;
  assign _EVAL_4518 = _EVAL_3078 & 32'h5f;
  assign _EVAL_2788 = _EVAL_4518 == 32'h17;
  assign _EVAL_1008 = _EVAL_4659 | _EVAL_2788;
  assign _EVAL_2628 = _EVAL_3078 & 32'hfc00007f;
  assign _EVAL_1860 = _EVAL_2628 == 32'h33;
  assign _EVAL_4503 = _EVAL_1008 | _EVAL_1860;
  assign _EVAL_4163 = _EVAL_3078 & 32'hbe00707f;
  assign _EVAL_5214 = _EVAL_4163 == 32'h33;
  assign _EVAL_5228 = _EVAL_4503 | _EVAL_5214;
  assign _EVAL_4951 = _EVAL_3078 & 32'h6000073;
  assign _EVAL_4400 = _EVAL_4951 == 32'h43;
  assign _EVAL_4544 = _EVAL_5228 | _EVAL_4400;
  assign _EVAL_2517 = _EVAL_3078 & 32'he600007f;
  assign _EVAL_1021 = _EVAL_2517 == 32'h53;
  assign _EVAL_2838 = _EVAL_4544 | _EVAL_1021;
  assign _EVAL_5223 = _EVAL_3078 & 32'h707b;
  assign _EVAL_5145 = _EVAL_5223 == 32'h63;
  assign _EVAL_4103 = _EVAL_2838 | _EVAL_5145;
  assign _EVAL_4594 = _EVAL_3078 & 32'h7f;
  assign _EVAL_5654 = _EVAL_4594 == 32'h6f;
  assign _EVAL_3674 = _EVAL_4103 | _EVAL_5654;
  assign _EVAL_2087 = _EVAL_3078 & 32'hffefffff;
  assign _EVAL_2442 = _EVAL_2087 == 32'h73;
  assign _EVAL_1507 = _EVAL_3674 | _EVAL_2442;
  assign _EVAL_4591 = _EVAL_3078 & 32'hfe00305f;
  assign _EVAL_5913 = _EVAL_4591 == 32'h1013;
  assign _EVAL_4603 = _EVAL_1507 | _EVAL_5913;
  assign _EVAL_5143 = _EVAL_3078 & 32'h705b;
  assign _EVAL_1641 = _EVAL_5143 == 32'h2003;
  assign _EVAL_3239 = _EVAL_4603 | _EVAL_1641;
  assign _EVAL_4268 = {_EVAL_2666,_EVAL_4292};
  assign _EVAL_771 = _EVAL_4268[15:13];
  assign _EVAL_5623 = _EVAL_771 == 3'h7;
  assign _EVAL_263 = _EVAL_4268[8:7];
  assign _EVAL_3602 = _EVAL_4268[12:9];
  assign _EVAL_3330 = {_EVAL_263,_EVAL_3602,2'h0};
  assign _EVAL_762 = _EVAL_3330[7:5];
  assign _EVAL_3553 = _EVAL_4268[6:2];
  assign _EVAL_871 = _EVAL_3330[4:0];
  assign _EVAL_2908 = {_EVAL_762,_EVAL_3553,5'h2,3'h2,_EVAL_871,7'h27};
  assign _EVAL_5053 = _EVAL_771 == 3'h6;
  assign _EVAL_5618 = {_EVAL_762,_EVAL_3553,5'h2,3'h2,_EVAL_871,7'h23};
  assign _EVAL_2321 = _EVAL_771 == 3'h5;
  assign _EVAL_3871 = _EVAL_4268[9:7];
  assign _EVAL_2808 = _EVAL_4268[12:10];
  assign _EVAL_1025 = {_EVAL_3871,_EVAL_2808,3'h0};
  assign _EVAL_2831 = _EVAL_1025[8:5];
  assign _EVAL_2613 = _EVAL_1025[4:0];
  assign _EVAL_1479 = {_EVAL_2831,_EVAL_3553,5'h2,3'h3,_EVAL_2613,7'h27};
  assign _EVAL_3712 = _EVAL_771 == 3'h4;
  assign _EVAL_5439 = _EVAL_4268[12];
  assign _EVAL_1657 = _EVAL_3553 != 5'h0;
  assign _EVAL_932 = _EVAL_4268[11:7];
  assign _EVAL_2026 = {_EVAL_3553,_EVAL_932,3'h0,_EVAL_932,7'h33};
  assign _EVAL_3685 = _EVAL_932 != 5'h0;
  assign _EVAL_4034 = {_EVAL_3553,_EVAL_932,3'h0,12'he7};
  assign _EVAL_3296 = {_EVAL_3553,_EVAL_932,3'h0,12'h67};
  assign _EVAL_1863 = _EVAL_3296[24:7];
  assign _EVAL_4578 = {_EVAL_1863,7'h73};
  assign _EVAL_4876 = _EVAL_4578 | 25'h100000;
  assign _EVAL_3519 = _EVAL_3685 ? _EVAL_4034 : _EVAL_4876;
  assign _EVAL_4673 = _EVAL_1657 ? _EVAL_2026 : _EVAL_3519;
  assign _EVAL_5005 = {_EVAL_3553,5'h0,3'h4,_EVAL_932,7'h33};
  assign _EVAL_282 = _EVAL_1657 ? _EVAL_5005 : _EVAL_3296;
  assign _EVAL_4515 = _EVAL_5439 ? _EVAL_4673 : _EVAL_282;
  assign _EVAL_1743 = _EVAL_771 == 3'h3;
  assign _EVAL_5411 = _EVAL_4268[3:2];
  assign _EVAL_626 = _EVAL_4268[6:4];
  assign _EVAL_2036 = {_EVAL_5411,_EVAL_5439,_EVAL_626,2'h0,5'h2,3'h2,_EVAL_932,7'h7};
  assign _EVAL_4038 = _EVAL_771 == 3'h2;
  assign _EVAL_1073 = {_EVAL_5411,_EVAL_5439,_EVAL_626,2'h0,5'h2,3'h2,_EVAL_932,7'h3};
  assign _EVAL_5573 = _EVAL_771 == 3'h1;
  assign _EVAL_763 = _EVAL_4268[4:2];
  assign _EVAL_167 = _EVAL_4268[6:5];
  assign _EVAL_3823 = {_EVAL_763,_EVAL_5439,_EVAL_167,3'h0,5'h2,3'h3,_EVAL_932,7'h7};
  assign _EVAL_341 = {_EVAL_5439,_EVAL_3553,_EVAL_932,3'h1,_EVAL_932,7'h13};
  assign _EVAL_180 = _EVAL_5573 ? _EVAL_3823 : {{3'd0}, _EVAL_341};
  assign _EVAL_1110 = _EVAL_4038 ? {{1'd0}, _EVAL_1073} : _EVAL_180;
  assign _EVAL_4831 = _EVAL_1743 ? {{1'd0}, _EVAL_2036} : _EVAL_1110;
  assign _EVAL_1996 = _EVAL_3712 ? {{4'd0}, _EVAL_4515} : _EVAL_4831;
  assign _EVAL_227 = _EVAL_2321 ? _EVAL_1479 : _EVAL_1996;
  assign _EVAL_3987 = _EVAL_5053 ? {{1'd0}, _EVAL_5618} : _EVAL_227;
  assign _EVAL_2410 = _EVAL_5623 ? {{1'd0}, _EVAL_2908} : _EVAL_3987;
  assign _EVAL_3006 = {3'h0,_EVAL_2410};
  assign _EVAL_2462 = _EVAL_3006 & 32'h80000010;
  assign _EVAL_5041 = _EVAL_2462 == 32'h10;
  assign _EVAL_3952 = _EVAL_3006 & 32'h50;
  assign _EVAL_4113 = _EVAL_3952 == 32'h10;
  assign _EVAL_4830 = _EVAL_5041 | _EVAL_4113;
  assign _EVAL_1111 = _EVAL_3006 & 32'h40000040;
  assign _EVAL_3150 = _EVAL_1111 == 32'h40;
  assign _EVAL_3757 = _EVAL_4830 | _EVAL_3150;
  assign _EVAL_1137 = _EVAL_3006 & 32'h20000040;
  assign _EVAL_470 = _EVAL_1137 == 32'h40;
  assign _EVAL_5979 = _EVAL_3757 | _EVAL_470;
  assign _EVAL_5386 = {_EVAL_2666,_EVAL_4292,_EVAL_5159,_EVAL_3588};
  assign _EVAL_1136 = _EVAL_5386[15:13];
  assign _EVAL_4999 = _EVAL_1136 == 3'h7;
  assign _EVAL_287 = _EVAL_5386[5];
  assign _EVAL_688 = _EVAL_5386[12:10];
  assign _EVAL_2964 = _EVAL_5386[6];
  assign _EVAL_3443 = {_EVAL_287,_EVAL_688,_EVAL_2964,2'h0};
  assign _EVAL_746 = _EVAL_3443[6:5];
  assign _EVAL_1418 = _EVAL_5386[4:2];
  assign _EVAL_5546 = _EVAL_5386[9:7];
  assign _EVAL_1050 = _EVAL_3443[4:0];
  assign _EVAL_2013 = {_EVAL_746,2'h1,_EVAL_1418,2'h1,_EVAL_5546,3'h2,_EVAL_1050,7'h27};
  assign _EVAL_4185 = _EVAL_1136 == 3'h6;
  assign _EVAL_4065 = {_EVAL_746,2'h1,_EVAL_1418,2'h1,_EVAL_5546,3'h2,_EVAL_1050,7'h23};
  assign _EVAL_3493 = _EVAL_1136 == 3'h5;
  assign _EVAL_5289 = _EVAL_5386[6:5];
  assign _EVAL_3643 = {_EVAL_5289,_EVAL_688,3'h0};
  assign _EVAL_3861 = _EVAL_3643[7:5];
  assign _EVAL_5112 = _EVAL_3643[4:0];
  assign _EVAL_5044 = {_EVAL_3861,2'h1,_EVAL_1418,2'h1,_EVAL_5546,3'h3,_EVAL_5112,7'h27};
  assign _EVAL_3261 = _EVAL_1136 == 3'h4;
  assign _EVAL_343 = {_EVAL_746,2'h1,_EVAL_1418,2'h1,_EVAL_5546,3'h0,_EVAL_1050,7'h27};
  assign _EVAL_268 = _EVAL_1136 == 3'h3;
  assign _EVAL_4834 = {_EVAL_287,_EVAL_688,_EVAL_2964,2'h0,2'h1,_EVAL_5546,3'h2,2'h1,_EVAL_1418,7'h7};
  assign _EVAL_179 = _EVAL_1136 == 3'h2;
  assign _EVAL_5270 = {_EVAL_287,_EVAL_688,_EVAL_2964,2'h0,2'h1,_EVAL_5546,3'h2,2'h1,_EVAL_1418,7'h3};
  assign _EVAL_2175 = _EVAL_1136 == 3'h1;
  assign _EVAL_3947 = {_EVAL_5289,_EVAL_688,3'h0,2'h1,_EVAL_5546,3'h3,2'h1,_EVAL_1418,7'h7};
  assign _EVAL_4465 = _EVAL_5386[10:7];
  assign _EVAL_3341 = _EVAL_5386[12:11];
  assign _EVAL_2263 = {_EVAL_4465,_EVAL_3341,_EVAL_287,_EVAL_2964,2'h0,5'h2,3'h0,2'h1,_EVAL_1418,7'h13};
  assign _EVAL_3834 = _EVAL_2175 ? {{2'd0}, _EVAL_3947} : _EVAL_2263;
  assign _EVAL_997 = _EVAL_179 ? {{3'd0}, _EVAL_5270} : _EVAL_3834;
  assign _EVAL_1859 = _EVAL_268 ? {{3'd0}, _EVAL_4834} : _EVAL_997;
  assign _EVAL_5281 = _EVAL_3261 ? {{3'd0}, _EVAL_343} : _EVAL_1859;
  assign _EVAL_1799 = _EVAL_3493 ? {{2'd0}, _EVAL_5044} : _EVAL_5281;
  assign _EVAL_2373 = _EVAL_4185 ? {{3'd0}, _EVAL_4065} : _EVAL_1799;
  assign _EVAL_1455 = _EVAL_4999 ? {{3'd0}, _EVAL_2013} : _EVAL_2373;
  assign _EVAL_386 = {2'h0,_EVAL_1455};
  assign _EVAL_2259 = _EVAL_386 & 32'h64;
  assign _EVAL_2390 = _EVAL_2259 == 32'h0;
  assign _EVAL_1473 = _EVAL_386 & 32'h50;
  assign _EVAL_706 = _EVAL_1473 == 32'h10;
  assign _EVAL_983 = _EVAL_2390 | _EVAL_706;
  assign _EVAL_476 = _EVAL_3455[8:7];
  assign _EVAL_4927 = _EVAL_3455[12:9];
  assign _EVAL_1900 = {_EVAL_476,_EVAL_4927,2'h0};
  assign _EVAL_2067 = _EVAL_1900[7:5];
  assign _EVAL_2075 = _EVAL_3455[6:2];
  assign _EVAL_4281 = _EVAL_1900[4:0];
  assign _EVAL_3343 = {_EVAL_2067,_EVAL_2075,5'h2,3'h2,_EVAL_4281,7'h27};
  assign _EVAL_4648 = {_EVAL_2067,_EVAL_2075,5'h2,3'h2,_EVAL_4281,7'h23};
  assign _EVAL_5823 = {_EVAL_4872,_EVAL_4901,3'h0};
  assign _EVAL_4096 = _EVAL_5823[8:5];
  assign _EVAL_822 = _EVAL_5823[4:0];
  assign _EVAL_6068 = {_EVAL_4096,_EVAL_2075,5'h2,3'h3,_EVAL_822,7'h27};
  assign _EVAL_735 = _EVAL_3455[12];
  assign _EVAL_1516 = _EVAL_2075 != 5'h0;
  assign _EVAL_3655 = _EVAL_3455[11:7];
  assign _EVAL_3062 = {_EVAL_2075,_EVAL_3655,3'h0,_EVAL_3655,7'h33};
  assign _EVAL_863 = _EVAL_3655 != 5'h0;
  assign _EVAL_1869 = {_EVAL_2075,_EVAL_3655,3'h0,12'he7};
  assign _EVAL_5542 = {_EVAL_2075,_EVAL_3655,3'h0,12'h67};
  assign _EVAL_3808 = _EVAL_5542[24:7];
  assign _EVAL_5624 = {_EVAL_3808,7'h73};
  assign _EVAL_3593 = _EVAL_5624 | 25'h100000;
  assign _EVAL_3134 = _EVAL_863 ? _EVAL_1869 : _EVAL_3593;
  assign _EVAL_1119 = _EVAL_1516 ? _EVAL_3062 : _EVAL_3134;
  assign _EVAL_5616 = {_EVAL_2075,5'h0,3'h4,_EVAL_3655,7'h33};
  assign _EVAL_543 = _EVAL_1516 ? _EVAL_5616 : _EVAL_5542;
  assign _EVAL_2595 = _EVAL_735 ? _EVAL_1119 : _EVAL_543;
  assign _EVAL_2351 = _EVAL_3455[3:2];
  assign _EVAL_5138 = _EVAL_3455[6:4];
  assign _EVAL_569 = {_EVAL_2351,_EVAL_735,_EVAL_5138,2'h0,5'h2,3'h2,_EVAL_3655,7'h7};
  assign _EVAL_578 = {_EVAL_2351,_EVAL_735,_EVAL_5138,2'h0,5'h2,3'h2,_EVAL_3655,7'h3};
  assign _EVAL_4655 = {_EVAL_3926,_EVAL_735,_EVAL_5278,3'h0,5'h2,3'h3,_EVAL_3655,7'h7};
  assign _EVAL_272 = {_EVAL_735,_EVAL_2075,_EVAL_3655,3'h1,_EVAL_3655,7'h13};
  assign _EVAL_5476 = _EVAL_5755 ? _EVAL_4655 : {{3'd0}, _EVAL_272};
  assign _EVAL_1189 = _EVAL_597 ? {{1'd0}, _EVAL_578} : _EVAL_5476;
  assign _EVAL_3708 = _EVAL_1674 ? {{1'd0}, _EVAL_569} : _EVAL_1189;
  assign _EVAL_3613 = _EVAL_936 ? {{4'd0}, _EVAL_2595} : _EVAL_3708;
  assign _EVAL_785 = _EVAL_453 ? _EVAL_6068 : _EVAL_3613;
  assign _EVAL_593 = _EVAL_2288 ? {{1'd0}, _EVAL_4648} : _EVAL_785;
  assign _EVAL_1348 = _EVAL_4669 ? {{1'd0}, _EVAL_3343} : _EVAL_593;
  assign _EVAL_2039 = {3'h0,_EVAL_1348};
  assign _EVAL_957 = _EVAL_2039 & 32'h207f;
  assign _EVAL_2132 = _EVAL_957 == 32'h3;
  assign _EVAL_3434 = _EVAL_2039 & 32'h607f;
  assign _EVAL_2712 = _EVAL_3434 == 32'hf;
  assign _EVAL_5529 = _EVAL_2132 | _EVAL_2712;
  assign _EVAL_5802 = _EVAL_2039 & 32'h5f;
  assign _EVAL_4128 = _EVAL_5802 == 32'h17;
  assign _EVAL_5560 = _EVAL_5529 | _EVAL_4128;
  assign _EVAL_5355 = _EVAL_2039 & 32'hfc00007f;
  assign _EVAL_3991 = _EVAL_5355 == 32'h33;
  assign _EVAL_5696 = _EVAL_5560 | _EVAL_3991;
  assign _EVAL_3844 = _EVAL_2039 & 32'hbe00707f;
  assign _EVAL_4210 = _EVAL_3844 == 32'h33;
  assign _EVAL_5945 = _EVAL_5696 | _EVAL_4210;
  assign _EVAL_2398 = _EVAL_2039 & 32'h6000073;
  assign _EVAL_644 = _EVAL_2398 == 32'h43;
  assign _EVAL_4110 = _EVAL_5945 | _EVAL_644;
  assign _EVAL_5061 = _EVAL_2039 & 32'he600007f;
  assign _EVAL_4386 = _EVAL_5061 == 32'h53;
  assign _EVAL_3478 = _EVAL_4110 | _EVAL_4386;
  assign _EVAL_5686 = _EVAL_2039 & 32'h707b;
  assign _EVAL_6118 = _EVAL_5686 == 32'h63;
  assign _EVAL_1707 = _EVAL_3478 | _EVAL_6118;
  assign _EVAL_1164 = _EVAL_2039 & 32'h7f;
  assign _EVAL_255 = _EVAL_1164 == 32'h6f;
  assign _EVAL_3880 = _EVAL_1707 | _EVAL_255;
  assign _EVAL_335 = _EVAL_2039 & 32'hffefffff;
  assign _EVAL_2153 = _EVAL_335 == 32'h73;
  assign _EVAL_568 = _EVAL_3880 | _EVAL_2153;
  assign _EVAL_4841 = _EVAL_2039 & 32'hfe00305f;
  assign _EVAL_6112 = _EVAL_4841 == 32'h1013;
  assign _EVAL_2897 = _EVAL_568 | _EVAL_6112;
  assign _EVAL_5329 = _EVAL_2039 & 32'h705b;
  assign _EVAL_2769 = _EVAL_5329 == 32'h2003;
  assign _EVAL_2848 = _EVAL_2897 | _EVAL_2769;
  assign _EVAL_5113 = _EVAL_957 == 32'h2013;
  assign _EVAL_3410 = _EVAL_2848 | _EVAL_5113;
  assign _EVAL_2663 = _EVAL_2039 & 32'h1800707f;
  assign _EVAL_5344 = _EVAL_2663 == 32'h202f;
  assign _EVAL_3795 = _EVAL_3410 | _EVAL_5344;
  assign _EVAL_861 = _EVAL_957 == 32'h2073;
  assign _EVAL_5070 = _EVAL_3795 | _EVAL_861;
  assign _EVAL_5078 = _EVAL_2039 & 32'hbe00705f;
  assign _EVAL_2802 = _EVAL_5078 == 32'h5013;
  assign _EVAL_5069 = _EVAL_5070 | _EVAL_2802;
  assign _EVAL_3300 = _EVAL_2039 & 32'he800707f;
  assign _EVAL_2197 = _EVAL_3300 == 32'h800202f;
  assign _EVAL_3874 = _EVAL_5069 | _EVAL_2197;
  assign _EVAL_4267 = _EVAL_2039 & 32'hf9f0707f;
  assign _EVAL_4618 = _EVAL_4267 == 32'h1000202f;
  assign _EVAL_203 = _EVAL_3874 | _EVAL_4618;
  assign _EVAL_4796 = _EVAL_2039 & 32'hdfffffff;
  assign _EVAL_2412 = _EVAL_4796 == 32'h10500073;
  assign _EVAL_264 = _EVAL_203 | _EVAL_2412;
  assign _EVAL_5455 = _EVAL_2039 & 32'hf600607f;
  assign _EVAL_801 = _EVAL_5455 == 32'h20000053;
  assign _EVAL_2360 = _EVAL_264 | _EVAL_801;
  assign _EVAL_4191 = _EVAL_2039 & 32'h7e00607f;
  assign _EVAL_5897 = _EVAL_4191 == 32'h20000053;
  assign _EVAL_1134 = _EVAL_2360 | _EVAL_5897;
  assign _EVAL_4944 = _EVAL_2039 & 32'h7e00507f;
  assign _EVAL_548 = _EVAL_4944 == 32'h20000053;
  assign _EVAL_3574 = _EVAL_1134 | _EVAL_548;
  assign _EVAL_2849 = _EVAL_2039 == 32'h30200073;
  assign _EVAL_892 = _EVAL_3574 | _EVAL_2849;
  assign _EVAL_3840 = _EVAL_2039 & 32'hfff0007f;
  assign _EVAL_2742 = _EVAL_3840 == 32'h58000053;
  assign _EVAL_1290 = _EVAL_892 | _EVAL_2742;
  assign _EVAL_4399 = _EVAL_2039 == 32'h7b200073;
  assign _EVAL_2736 = _EVAL_1290 | _EVAL_4399;
  assign _EVAL_234 = _EVAL_2039 & 32'hefe0007f;
  assign _EVAL_2598 = _EVAL_234 == 32'hc0000053;
  assign _EVAL_1520 = _EVAL_2736 | _EVAL_2598;
  assign _EVAL_2890 = _EVAL_2039 & 32'hfff0607f;
  assign _EVAL_4216 = _EVAL_2890 == 32'he0000053;
  assign _EVAL_1398 = _EVAL_1520 | _EVAL_4216;
  assign _EVAL_4535 = _EVAL_2666[15:13];
  assign _EVAL_418 = _EVAL_4535 == 3'h7;
  assign _EVAL_1583 = _EVAL_2666[12];
  assign _EVAL_2657 = _EVAL_1583 ? 5'h1f : 5'h0;
  assign _EVAL_3105 = _EVAL_2666[6:5];
  assign _EVAL_5775 = _EVAL_2666[2];
  assign _EVAL_2671 = _EVAL_2666[11:10];
  assign _EVAL_3182 = _EVAL_2666[4:3];
  assign _EVAL_269 = {_EVAL_2657,_EVAL_3105,_EVAL_5775,_EVAL_2671,_EVAL_3182,1'h0};
  assign _EVAL_6027 = _EVAL_269[12];
  assign _EVAL_4693 = _EVAL_269[10:5];
  assign _EVAL_1375 = _EVAL_2666[9:7];
  assign _EVAL_3642 = _EVAL_269[4:1];
  assign _EVAL_3414 = _EVAL_269[11];
  assign _EVAL_4233 = {_EVAL_6027,_EVAL_4693,5'h0,2'h1,_EVAL_1375,3'h1,_EVAL_3642,_EVAL_3414,7'h63};
  assign _EVAL_5821 = _EVAL_4535 == 3'h6;
  assign _EVAL_4762 = {_EVAL_6027,_EVAL_4693,5'h0,2'h1,_EVAL_1375,3'h0,_EVAL_3642,_EVAL_3414,7'h63};
  assign _EVAL_2644 = _EVAL_4535 == 3'h5;
  assign _EVAL_2268 = _EVAL_1583 ? 10'h3ff : 10'h0;
  assign _EVAL_5309 = _EVAL_2666[8];
  assign _EVAL_4709 = _EVAL_2666[10:9];
  assign _EVAL_5340 = _EVAL_2666[6];
  assign _EVAL_882 = _EVAL_2666[7];
  assign _EVAL_3287 = _EVAL_2666[11];
  assign _EVAL_3748 = _EVAL_2666[5:3];
  assign _EVAL_3811 = {_EVAL_2268,_EVAL_5309,_EVAL_4709,_EVAL_5340,_EVAL_882,_EVAL_5775,_EVAL_3287,_EVAL_3748,1'h0};
  assign _EVAL_2989 = _EVAL_3811[20];
  assign _EVAL_2920 = _EVAL_3811[10:1];
  assign _EVAL_5236 = _EVAL_3811[11];
  assign _EVAL_1128 = _EVAL_3811[19:12];
  assign _EVAL_5753 = {_EVAL_2989,_EVAL_2920,_EVAL_5236,_EVAL_1128,5'h0,7'h6f};
  assign _EVAL_4202 = _EVAL_4535 == 3'h4;
  assign _EVAL_5825 = _EVAL_2671 == 2'h3;
  assign _EVAL_5741 = _EVAL_2666[4:2];
  assign _EVAL_1612 = {_EVAL_1583,_EVAL_3105};
  assign _EVAL_5920 = _EVAL_1612 == 3'h7;
  assign _EVAL_4348 = _EVAL_1612 == 3'h6;
  assign _EVAL_3827 = _EVAL_1612 == 3'h5;
  assign _EVAL_346 = _EVAL_1612 == 3'h4;
  assign _EVAL_2219 = _EVAL_1612 == 3'h3;
  assign _EVAL_2608 = _EVAL_1612 == 3'h2;
  assign _EVAL_1784 = _EVAL_1612 == 3'h1;
  assign _EVAL_1778 = _EVAL_1784 ? 3'h4 : 3'h0;
  assign _EVAL_5864 = _EVAL_2608 ? 3'h6 : _EVAL_1778;
  assign _EVAL_4324 = _EVAL_2219 ? 3'h7 : _EVAL_5864;
  assign _EVAL_937 = _EVAL_346 ? 3'h0 : _EVAL_4324;
  assign _EVAL_350 = _EVAL_3827 ? 3'h0 : _EVAL_937;
  assign _EVAL_5404 = _EVAL_4348 ? 3'h2 : _EVAL_350;
  assign _EVAL_2308 = _EVAL_5920 ? 3'h3 : _EVAL_5404;
  assign _EVAL_4551 = _EVAL_1583 ? 7'h3b : 7'h33;
  assign _EVAL_1161 = {2'h1,_EVAL_5741,2'h1,_EVAL_1375,_EVAL_2308,2'h1,_EVAL_1375,_EVAL_4551};
  assign _EVAL_2572 = {{6'd0}, _EVAL_1161};
  assign _EVAL_3966 = _EVAL_3105 == 2'h0;
  assign _EVAL_1339 = {_EVAL_3966, 30'h0};
  assign _EVAL_620 = _EVAL_2572 | _EVAL_1339;
  assign _EVAL_647 = _EVAL_2671 == 2'h2;
  assign _EVAL_2409 = _EVAL_1583 ? 7'h7f : 7'h0;
  assign _EVAL_4489 = _EVAL_2666[6:2];
  assign _EVAL_2776 = {_EVAL_2409,_EVAL_4489,2'h1,_EVAL_1375,3'h7,2'h1,_EVAL_1375,7'h13};
  assign _EVAL_1181 = _EVAL_2671 == 2'h1;
  assign _EVAL_4695 = {_EVAL_1583,_EVAL_4489,2'h1,_EVAL_1375,3'h5,2'h1,_EVAL_1375,7'h13};
  assign _EVAL_4933 = {{5'd0}, _EVAL_4695};
  assign _EVAL_2664 = _EVAL_4933 | 31'h40000000;
  assign _EVAL_1112 = _EVAL_1181 ? _EVAL_2664 : {{5'd0}, _EVAL_4695};
  assign _EVAL_3909 = _EVAL_647 ? _EVAL_2776 : {{1'd0}, _EVAL_1112};
  assign _EVAL_1839 = _EVAL_5825 ? {{1'd0}, _EVAL_620} : _EVAL_3909;
  assign _EVAL_4352 = _EVAL_4535 == 3'h3;
  assign _EVAL_5023 = _EVAL_2666[11:7];
  assign _EVAL_3277 = _EVAL_5023 == 5'h2;
  assign _EVAL_2576 = _EVAL_1583 ? 3'h7 : 3'h0;
  assign _EVAL_1329 = _EVAL_2666[5];
  assign _EVAL_477 = {_EVAL_2576,_EVAL_3182,_EVAL_1329,_EVAL_5775,_EVAL_5340,4'h0,_EVAL_5023,3'h0,_EVAL_5023,7'h13};
  assign _EVAL_1713 = _EVAL_1583 ? 15'h7fff : 15'h0;
  assign _EVAL_3263 = {_EVAL_1713,_EVAL_4489,12'h0};
  assign _EVAL_3826 = _EVAL_3263[31:12];
  assign _EVAL_3311 = {_EVAL_3826,_EVAL_5023,7'h37};
  assign _EVAL_3412 = _EVAL_3277 ? _EVAL_477 : _EVAL_3311;
  assign _EVAL_1014 = _EVAL_4535 == 3'h2;
  assign _EVAL_1003 = {_EVAL_2409,_EVAL_4489,5'h0,3'h0,_EVAL_5023,7'h13};
  assign _EVAL_630 = _EVAL_4535 == 3'h1;
  assign _EVAL_1962 = {_EVAL_2989,_EVAL_2920,_EVAL_5236,_EVAL_1128,5'h1,7'h6f};
  assign _EVAL_1235 = {_EVAL_2409,_EVAL_4489,_EVAL_5023,3'h0,_EVAL_5023,7'h13};
  assign _EVAL_1320 = _EVAL_630 ? _EVAL_1962 : _EVAL_1235;
  assign _EVAL_4467 = _EVAL_1014 ? _EVAL_1003 : _EVAL_1320;
  assign _EVAL_1727 = _EVAL_4352 ? _EVAL_3412 : _EVAL_4467;
  assign _EVAL_1493 = _EVAL_4202 ? _EVAL_1839 : _EVAL_1727;
  assign _EVAL_3372 = _EVAL_2644 ? _EVAL_5753 : _EVAL_1493;
  assign _EVAL_3906 = _EVAL_5821 ? _EVAL_4762 : _EVAL_3372;
  assign _EVAL_1362 = _EVAL_418 ? _EVAL_4233 : _EVAL_3906;
  assign _EVAL_1096 = _EVAL_1362 & 32'h44;
  assign _EVAL_5421 = _EVAL_1096 == 32'h0;
  assign _EVAL_2600 = {_EVAL_735,_EVAL_5278};
  assign _EVAL_5872 = _EVAL_2600 == 3'h7;
  assign _EVAL_5387 = _EVAL_2600 == 3'h6;
  assign _EVAL_5474 = _EVAL_2600 == 3'h5;
  assign _EVAL_392 = _EVAL_2600 == 3'h4;
  assign _EVAL_4750 = _EVAL_2600 == 3'h3;
  assign _EVAL_4809 = _EVAL_2600 == 3'h2;
  assign _EVAL_1551 = _EVAL_2600 == 3'h1;
  assign _EVAL_4531 = _EVAL_1551 ? 3'h4 : 3'h0;
  assign _EVAL_3094 = _EVAL_4809 ? 3'h6 : _EVAL_4531;
  assign _EVAL_5638 = _EVAL_4750 ? 3'h7 : _EVAL_3094;
  assign _EVAL_6071 = _EVAL_392 ? 3'h0 : _EVAL_5638;
  assign _EVAL_6140 = _EVAL_5474 ? 3'h0 : _EVAL_6071;
  assign _EVAL_3910 = _EVAL_5387 ? 3'h2 : _EVAL_6140;
  assign _EVAL_3630 = _EVAL_5872 ? 3'h3 : _EVAL_3910;
  assign _EVAL_4250 = _EVAL_735 ? 7'h3b : 7'h33;
  assign _EVAL_3408 = {2'h1,_EVAL_3926,2'h1,_EVAL_4872,_EVAL_3630,2'h1,_EVAL_4872,_EVAL_4250};
  assign _EVAL_3385 = _EVAL_3082 ? 5'h1f : 5'h0;
  assign _EVAL_218 = _EVAL_654[2];
  assign _EVAL_948 = _EVAL_654[11:10];
  assign _EVAL_3864 = _EVAL_654[4:3];
  assign _EVAL_334 = {_EVAL_3385,_EVAL_4575,_EVAL_218,_EVAL_948,_EVAL_3864,1'h0};
  assign _EVAL_5403 = _EVAL_334[10:5];
  assign _EVAL_4728 = _EVAL_5386[1:0];
  assign _EVAL_5952 = _EVAL_4728 == 2'h1;
  assign _EVAL_4111 = _EVAL_5386[12];
  assign _EVAL_2534 = _EVAL_4111 ? 5'h1f : 5'h0;
  assign _EVAL_3920 = _EVAL_5386[2];
  assign _EVAL_3636 = _EVAL_5386[11:10];
  assign _EVAL_5034 = _EVAL_5386[4:3];
  assign _EVAL_502 = {_EVAL_2534,_EVAL_5289,_EVAL_3920,_EVAL_3636,_EVAL_5034,1'h0};
  assign _EVAL_707 = _EVAL_502[12];
  assign _EVAL_876 = _EVAL_502[10:5];
  assign _EVAL_5766 = _EVAL_502[4:1];
  assign _EVAL_650 = _EVAL_502[11];
  assign _EVAL_5831 = {_EVAL_707,_EVAL_876,5'h0,2'h1,_EVAL_5546,3'h1,_EVAL_5766,_EVAL_650,7'h63};
  assign _EVAL_2480 = {_EVAL_707,_EVAL_876,5'h0,2'h1,_EVAL_5546,3'h0,_EVAL_5766,_EVAL_650,7'h63};
  assign _EVAL_2912 = _EVAL_4111 ? 10'h3ff : 10'h0;
  assign _EVAL_3183 = _EVAL_5386[8];
  assign _EVAL_745 = _EVAL_5386[10:9];
  assign _EVAL_2546 = _EVAL_5386[7];
  assign _EVAL_3106 = _EVAL_5386[11];
  assign _EVAL_1759 = _EVAL_5386[5:3];
  assign _EVAL_4715 = {_EVAL_2912,_EVAL_3183,_EVAL_745,_EVAL_2964,_EVAL_2546,_EVAL_3920,_EVAL_3106,_EVAL_1759,1'h0};
  assign _EVAL_2592 = _EVAL_4715[20];
  assign _EVAL_3210 = _EVAL_4715[10:1];
  assign _EVAL_2251 = _EVAL_4715[11];
  assign _EVAL_1182 = _EVAL_4715[19:12];
  assign _EVAL_5304 = {_EVAL_2592,_EVAL_3210,_EVAL_2251,_EVAL_1182,5'h0,7'h6f};
  assign _EVAL_896 = _EVAL_3636 == 2'h3;
  assign _EVAL_4176 = {_EVAL_4111,_EVAL_5289};
  assign _EVAL_4036 = _EVAL_4176 == 3'h7;
  assign _EVAL_4845 = _EVAL_4176 == 3'h6;
  assign _EVAL_4391 = _EVAL_4176 == 3'h5;
  assign _EVAL_5613 = _EVAL_4176 == 3'h4;
  assign _EVAL_6020 = _EVAL_4176 == 3'h3;
  assign _EVAL_5356 = _EVAL_4176 == 3'h2;
  assign _EVAL_2174 = _EVAL_4176 == 3'h1;
  assign _EVAL_2242 = _EVAL_2174 ? 3'h4 : 3'h0;
  assign _EVAL_3710 = _EVAL_5356 ? 3'h6 : _EVAL_2242;
  assign _EVAL_5357 = _EVAL_6020 ? 3'h7 : _EVAL_3710;
  assign _EVAL_3395 = _EVAL_5613 ? 3'h0 : _EVAL_5357;
  assign _EVAL_2668 = _EVAL_4391 ? 3'h0 : _EVAL_3395;
  assign _EVAL_2414 = _EVAL_4845 ? 3'h2 : _EVAL_2668;
  assign _EVAL_1443 = _EVAL_4036 ? 3'h3 : _EVAL_2414;
  assign _EVAL_3839 = _EVAL_4111 ? 7'h3b : 7'h33;
  assign _EVAL_1890 = {2'h1,_EVAL_1418,2'h1,_EVAL_5546,_EVAL_1443,2'h1,_EVAL_5546,_EVAL_3839};
  assign _EVAL_3767 = {{6'd0}, _EVAL_1890};
  assign _EVAL_3470 = _EVAL_5289 == 2'h0;
  assign _EVAL_3378 = {_EVAL_3470, 30'h0};
  assign _EVAL_553 = _EVAL_3767 | _EVAL_3378;
  assign _EVAL_4751 = _EVAL_3636 == 2'h2;
  assign _EVAL_1746 = _EVAL_4111 ? 7'h7f : 7'h0;
  assign _EVAL_2272 = _EVAL_5386[6:2];
  assign _EVAL_3621 = {_EVAL_1746,_EVAL_2272,2'h1,_EVAL_5546,3'h7,2'h1,_EVAL_5546,7'h13};
  assign _EVAL_1824 = _EVAL_3636 == 2'h1;
  assign _EVAL_1970 = {_EVAL_4111,_EVAL_2272,2'h1,_EVAL_5546,3'h5,2'h1,_EVAL_5546,7'h13};
  assign _EVAL_4916 = {{5'd0}, _EVAL_1970};
  assign _EVAL_4429 = _EVAL_4916 | 31'h40000000;
  assign _EVAL_1678 = _EVAL_1824 ? _EVAL_4429 : {{5'd0}, _EVAL_1970};
  assign _EVAL_3761 = _EVAL_4751 ? _EVAL_3621 : {{1'd0}, _EVAL_1678};
  assign _EVAL_5015 = _EVAL_896 ? {{1'd0}, _EVAL_553} : _EVAL_3761;
  assign _EVAL_4374 = _EVAL_5386[11:7];
  assign _EVAL_3004 = _EVAL_4374 == 5'h2;
  assign _EVAL_757 = _EVAL_4111 ? 3'h7 : 3'h0;
  assign _EVAL_3218 = {_EVAL_757,_EVAL_5034,_EVAL_287,_EVAL_3920,_EVAL_2964,4'h0,_EVAL_4374,3'h0,_EVAL_4374,7'h13};
  assign _EVAL_2157 = _EVAL_4111 ? 15'h7fff : 15'h0;
  assign _EVAL_5760 = {_EVAL_2157,_EVAL_2272,12'h0};
  assign _EVAL_5101 = _EVAL_5760[31:12];
  assign _EVAL_837 = {_EVAL_5101,_EVAL_4374,7'h37};
  assign _EVAL_2568 = _EVAL_3004 ? _EVAL_3218 : _EVAL_837;
  assign _EVAL_4390 = {_EVAL_1746,_EVAL_2272,5'h0,3'h0,_EVAL_4374,7'h13};
  assign _EVAL_6047 = {_EVAL_2592,_EVAL_3210,_EVAL_2251,_EVAL_1182,5'h1,7'h6f};
  assign _EVAL_1954 = {_EVAL_1746,_EVAL_2272,_EVAL_4374,3'h0,_EVAL_4374,7'h13};
  assign _EVAL_5009 = _EVAL_2175 ? _EVAL_6047 : _EVAL_1954;
  assign _EVAL_4338 = _EVAL_179 ? _EVAL_4390 : _EVAL_5009;
  assign _EVAL_5428 = _EVAL_268 ? _EVAL_2568 : _EVAL_4338;
  assign _EVAL_1416 = _EVAL_3261 ? _EVAL_5015 : _EVAL_5428;
  assign _EVAL_3129 = _EVAL_3493 ? _EVAL_5304 : _EVAL_1416;
  assign _EVAL_1160 = _EVAL_4185 ? _EVAL_2480 : _EVAL_3129;
  assign _EVAL_4743 = _EVAL_4999 ? _EVAL_5831 : _EVAL_1160;
  assign _EVAL_5510 = _EVAL_4743[24:20];
  assign _EVAL_5456 = _EVAL_386[24:20];
  assign _EVAL_5074 = _EVAL_5952 ? _EVAL_5510 : _EVAL_5456;
  assign _EVAL_3200 = _EVAL_2666[8:7];
  assign _EVAL_2739 = _EVAL_2666[12:9];
  assign _EVAL_4277 = {_EVAL_3200,_EVAL_2739,2'h0};
  assign _EVAL_2466 = _EVAL_4277[7:5];
  assign _EVAL_1636 = _EVAL_4277[4:0];
  assign _EVAL_3405 = {_EVAL_2466,_EVAL_4489,5'h2,3'h2,_EVAL_1636,7'h27};
  assign _EVAL_5944 = {_EVAL_2466,_EVAL_4489,5'h2,3'h2,_EVAL_1636,7'h23};
  assign _EVAL_821 = _EVAL_2666[12:10];
  assign _EVAL_1036 = {_EVAL_1375,_EVAL_821,3'h0};
  assign _EVAL_5503 = _EVAL_1036[8:5];
  assign _EVAL_5874 = _EVAL_1036[4:0];
  assign _EVAL_5265 = {_EVAL_5503,_EVAL_4489,5'h2,3'h3,_EVAL_5874,7'h27};
  assign _EVAL_2327 = _EVAL_4489 != 5'h0;
  assign _EVAL_1152 = {_EVAL_4489,_EVAL_5023,3'h0,_EVAL_5023,7'h33};
  assign _EVAL_5924 = _EVAL_5023 != 5'h0;
  assign _EVAL_5441 = {_EVAL_4489,_EVAL_5023,3'h0,12'he7};
  assign _EVAL_3534 = {_EVAL_4489,_EVAL_5023,3'h0,12'h67};
  assign _EVAL_1041 = _EVAL_3534[24:7];
  assign _EVAL_5904 = {_EVAL_1041,7'h73};
  assign _EVAL_4112 = _EVAL_5904 | 25'h100000;
  assign _EVAL_5615 = _EVAL_5924 ? _EVAL_5441 : _EVAL_4112;
  assign _EVAL_4812 = _EVAL_2327 ? _EVAL_1152 : _EVAL_5615;
  assign _EVAL_4730 = {_EVAL_4489,5'h0,3'h4,_EVAL_5023,7'h33};
  assign _EVAL_1536 = _EVAL_2327 ? _EVAL_4730 : _EVAL_3534;
  assign _EVAL_212 = _EVAL_1583 ? _EVAL_4812 : _EVAL_1536;
  assign _EVAL_4012 = _EVAL_2666[3:2];
  assign _EVAL_1124 = _EVAL_2666[6:4];
  assign _EVAL_5736 = {_EVAL_4012,_EVAL_1583,_EVAL_1124,2'h0,5'h2,3'h2,_EVAL_5023,7'h7};
  assign _EVAL_4560 = {_EVAL_4012,_EVAL_1583,_EVAL_1124,2'h0,5'h2,3'h2,_EVAL_5023,7'h3};
  assign _EVAL_2417 = {_EVAL_5741,_EVAL_1583,_EVAL_3105,3'h0,5'h2,3'h3,_EVAL_5023,7'h7};
  assign _EVAL_3883 = {_EVAL_1583,_EVAL_4489,_EVAL_5023,3'h1,_EVAL_5023,7'h13};
  assign _EVAL_5416 = _EVAL_630 ? _EVAL_2417 : {{3'd0}, _EVAL_3883};
  assign _EVAL_436 = _EVAL_1014 ? {{1'd0}, _EVAL_4560} : _EVAL_5416;
  assign _EVAL_2883 = _EVAL_4352 ? {{1'd0}, _EVAL_5736} : _EVAL_436;
  assign _EVAL_5490 = _EVAL_4202 ? {{4'd0}, _EVAL_212} : _EVAL_2883;
  assign _EVAL_5515 = _EVAL_2644 ? _EVAL_5265 : _EVAL_5490;
  assign _EVAL_1358 = _EVAL_5821 ? {{1'd0}, _EVAL_5944} : _EVAL_5515;
  assign _EVAL_1162 = _EVAL_418 ? {{1'd0}, _EVAL_3405} : _EVAL_1358;
  assign _EVAL_1978 = {3'h0,_EVAL_1162};
  assign _EVAL_4366 = _EVAL_1978 & 32'h5f;
  assign _EVAL_1747 = _EVAL_5439 ? 5'h1f : 5'h0;
  assign _EVAL_3677 = _EVAL_4268[2];
  assign _EVAL_4680 = _EVAL_4268[11:10];
  assign _EVAL_1092 = _EVAL_4268[4:3];
  assign _EVAL_5804 = {_EVAL_1747,_EVAL_167,_EVAL_3677,_EVAL_4680,_EVAL_1092,1'h0};
  assign _EVAL_4021 = _EVAL_5804[12];
  assign _EVAL_3474 = _EVAL_5804[10:5];
  assign _EVAL_3014 = _EVAL_5804[4:1];
  assign _EVAL_2266 = _EVAL_5804[11];
  assign _EVAL_2779 = {_EVAL_4021,_EVAL_3474,5'h0,2'h1,_EVAL_3871,3'h1,_EVAL_3014,_EVAL_2266,7'h63};
  assign _EVAL_3091 = {_EVAL_4021,_EVAL_3474,5'h0,2'h1,_EVAL_3871,3'h0,_EVAL_3014,_EVAL_2266,7'h63};
  assign _EVAL_4449 = _EVAL_5439 ? 10'h3ff : 10'h0;
  assign _EVAL_1100 = _EVAL_4268[8];
  assign _EVAL_3102 = _EVAL_4268[10:9];
  assign _EVAL_2711 = _EVAL_4268[6];
  assign _EVAL_2003 = _EVAL_4268[7];
  assign _EVAL_2525 = _EVAL_4268[11];
  assign _EVAL_3498 = _EVAL_4268[5:3];
  assign _EVAL_5465 = {_EVAL_4449,_EVAL_1100,_EVAL_3102,_EVAL_2711,_EVAL_2003,_EVAL_3677,_EVAL_2525,_EVAL_3498,1'h0};
  assign _EVAL_3881 = _EVAL_5465[20];
  assign _EVAL_5580 = _EVAL_5465[10:1];
  assign _EVAL_3307 = _EVAL_5465[11];
  assign _EVAL_5562 = _EVAL_5465[19:12];
  assign _EVAL_5948 = {_EVAL_3881,_EVAL_5580,_EVAL_3307,_EVAL_5562,5'h0,7'h6f};
  assign _EVAL_695 = _EVAL_4680 == 2'h3;
  assign _EVAL_1803 = {_EVAL_5439,_EVAL_167};
  assign _EVAL_4620 = _EVAL_1803 == 3'h7;
  assign _EVAL_5493 = _EVAL_1803 == 3'h6;
  assign _EVAL_1121 = _EVAL_1803 == 3'h5;
  assign _EVAL_5602 = _EVAL_1803 == 3'h4;
  assign _EVAL_1210 = _EVAL_1803 == 3'h3;
  assign _EVAL_3051 = _EVAL_1803 == 3'h2;
  assign _EVAL_2984 = _EVAL_1803 == 3'h1;
  assign _EVAL_4547 = _EVAL_2984 ? 3'h4 : 3'h0;
  assign _EVAL_2877 = _EVAL_3051 ? 3'h6 : _EVAL_4547;
  assign _EVAL_3126 = _EVAL_1210 ? 3'h7 : _EVAL_2877;
  assign _EVAL_6094 = _EVAL_5602 ? 3'h0 : _EVAL_3126;
  assign _EVAL_3820 = _EVAL_1121 ? 3'h0 : _EVAL_6094;
  assign _EVAL_3209 = _EVAL_5493 ? 3'h2 : _EVAL_3820;
  assign _EVAL_690 = _EVAL_4620 ? 3'h3 : _EVAL_3209;
  assign _EVAL_3616 = _EVAL_5439 ? 7'h3b : 7'h33;
  assign _EVAL_464 = {2'h1,_EVAL_763,2'h1,_EVAL_3871,_EVAL_690,2'h1,_EVAL_3871,_EVAL_3616};
  assign _EVAL_1675 = {{6'd0}, _EVAL_464};
  assign _EVAL_243 = _EVAL_167 == 2'h0;
  assign _EVAL_2022 = {_EVAL_243, 30'h0};
  assign _EVAL_1807 = _EVAL_1675 | _EVAL_2022;
  assign _EVAL_380 = _EVAL_4680 == 2'h2;
  assign _EVAL_3620 = _EVAL_5439 ? 7'h7f : 7'h0;
  assign _EVAL_2934 = {_EVAL_3620,_EVAL_3553,2'h1,_EVAL_3871,3'h7,2'h1,_EVAL_3871,7'h13};
  assign _EVAL_5259 = _EVAL_4680 == 2'h1;
  assign _EVAL_4447 = {_EVAL_5439,_EVAL_3553,2'h1,_EVAL_3871,3'h5,2'h1,_EVAL_3871,7'h13};
  assign _EVAL_4905 = {{5'd0}, _EVAL_4447};
  assign _EVAL_1056 = _EVAL_4905 | 31'h40000000;
  assign _EVAL_1194 = _EVAL_5259 ? _EVAL_1056 : {{5'd0}, _EVAL_4447};
  assign _EVAL_3148 = _EVAL_380 ? _EVAL_2934 : {{1'd0}, _EVAL_1194};
  assign _EVAL_5991 = _EVAL_695 ? {{1'd0}, _EVAL_1807} : _EVAL_3148;
  assign _EVAL_2176 = _EVAL_932 == 5'h2;
  assign _EVAL_2235 = _EVAL_5439 ? 3'h7 : 3'h0;
  assign _EVAL_3591 = _EVAL_4268[5];
  assign _EVAL_5679 = {_EVAL_2235,_EVAL_1092,_EVAL_3591,_EVAL_3677,_EVAL_2711,4'h0,_EVAL_932,3'h0,_EVAL_932,7'h13};
  assign _EVAL_2444 = _EVAL_5439 ? 15'h7fff : 15'h0;
  assign _EVAL_1199 = {_EVAL_2444,_EVAL_3553,12'h0};
  assign _EVAL_5415 = _EVAL_1199[31:12];
  assign _EVAL_4247 = {_EVAL_5415,_EVAL_932,7'h37};
  assign _EVAL_3013 = _EVAL_2176 ? _EVAL_5679 : _EVAL_4247;
  assign _EVAL_6042 = {_EVAL_3620,_EVAL_3553,5'h0,3'h0,_EVAL_932,7'h13};
  assign _EVAL_4319 = {_EVAL_3881,_EVAL_5580,_EVAL_3307,_EVAL_5562,5'h1,7'h6f};
  assign _EVAL_5271 = {_EVAL_3620,_EVAL_3553,_EVAL_932,3'h0,_EVAL_932,7'h13};
  assign _EVAL_3598 = _EVAL_5573 ? _EVAL_4319 : _EVAL_5271;
  assign _EVAL_3467 = _EVAL_4038 ? _EVAL_6042 : _EVAL_3598;
  assign _EVAL_4394 = _EVAL_1743 ? _EVAL_3013 : _EVAL_3467;
  assign _EVAL_1565 = _EVAL_3712 ? _EVAL_5991 : _EVAL_4394;
  assign _EVAL_4372 = _EVAL_2321 ? _EVAL_5948 : _EVAL_1565;
  assign _EVAL_3213 = _EVAL_5053 ? _EVAL_3091 : _EVAL_4372;
  assign _EVAL_4882 = _EVAL_5623 ? _EVAL_2779 : _EVAL_3213;
  assign _EVAL_411 = _EVAL_4882 & 32'h44;
  assign _EVAL_3011 = _EVAL_411 == 32'h4;
  assign _EVAL_3065 = _EVAL_3006 & 32'h64;
  assign _EVAL_185 = {_EVAL_3591,_EVAL_2808,_EVAL_2711,2'h0};
  assign _EVAL_3946 = _EVAL_185[6:5];
  assign _EVAL_6089 = _EVAL_185[4:0];
  assign _EVAL_3100 = {_EVAL_3946,2'h1,_EVAL_763,2'h1,_EVAL_3871,3'h2,_EVAL_6089,7'h27};
  assign _EVAL_5832 = {_EVAL_3946,2'h1,_EVAL_763,2'h1,_EVAL_3871,3'h2,_EVAL_6089,7'h23};
  assign _EVAL_2494 = {_EVAL_167,_EVAL_2808,3'h0};
  assign _EVAL_6126 = _EVAL_2494[7:5];
  assign _EVAL_522 = _EVAL_2494[4:0];
  assign _EVAL_1065 = {_EVAL_6126,2'h1,_EVAL_763,2'h1,_EVAL_3871,3'h3,_EVAL_522,7'h27};
  assign _EVAL_5132 = {_EVAL_3946,2'h1,_EVAL_763,2'h1,_EVAL_3871,3'h0,_EVAL_6089,7'h27};
  assign _EVAL_5338 = {_EVAL_3591,_EVAL_2808,_EVAL_2711,2'h0,2'h1,_EVAL_3871,3'h2,2'h1,_EVAL_763,7'h7};
  assign _EVAL_4120 = {_EVAL_3591,_EVAL_2808,_EVAL_2711,2'h0,2'h1,_EVAL_3871,3'h2,2'h1,_EVAL_763,7'h3};
  assign _EVAL_2122 = {_EVAL_167,_EVAL_2808,3'h0,2'h1,_EVAL_3871,3'h3,2'h1,_EVAL_763,7'h7};
  assign _EVAL_5636 = _EVAL_4268[10:7];
  assign _EVAL_5612 = _EVAL_4268[12:11];
  assign _EVAL_193 = {_EVAL_5636,_EVAL_5612,_EVAL_3591,_EVAL_2711,2'h0,5'h2,3'h0,2'h1,_EVAL_763,7'h13};
  assign _EVAL_4936 = _EVAL_5573 ? {{2'd0}, _EVAL_2122} : _EVAL_193;
  assign _EVAL_1314 = _EVAL_4038 ? {{3'd0}, _EVAL_4120} : _EVAL_4936;
  assign _EVAL_6108 = _EVAL_1743 ? {{3'd0}, _EVAL_5338} : _EVAL_1314;
  assign _EVAL_306 = _EVAL_3712 ? {{3'd0}, _EVAL_5132} : _EVAL_6108;
  assign _EVAL_2752 = _EVAL_2321 ? {{2'd0}, _EVAL_1065} : _EVAL_306;
  assign _EVAL_1177 = _EVAL_5053 ? {{3'd0}, _EVAL_5832} : _EVAL_2752;
  assign _EVAL_3496 = _EVAL_5623 ? {{3'd0}, _EVAL_3100} : _EVAL_1177;
  assign _EVAL_5133 = {2'h0,_EVAL_3496};
  assign _EVAL_5578 = _EVAL_5133 & 32'h4024;
  assign _EVAL_5723 = _EVAL_5578 == 32'h20;
  assign _EVAL_6081 = _EVAL_53;
  assign _EVAL_2110 = _EVAL_6081 == 1'h0;
  assign _EVAL_5564 = _EVAL_142;
  assign _EVAL_5718 = _EVAL_5564 == 1'h0;
  assign _EVAL_2396 = _EVAL_107;
  assign _EVAL_1206 = _EVAL_145;
  assign _EVAL_5440 = {_EVAL_2396,1'h0,1'h0,_EVAL_1206};
  assign _EVAL_4264 = _EVAL_5440 >> _EVAL_4188;
  assign _EVAL_5087 = _EVAL_4264[0];
  assign _EVAL_3382 = _EVAL_5718 & _EVAL_5087;
  assign _EVAL_2532 = _EVAL_32;
  assign _EVAL_5393 = _EVAL_3382 & _EVAL_2532;
  assign _EVAL_5211 = _EVAL_98;
  assign _EVAL_4914 = _EVAL_5211[1];
  assign _EVAL_1992 = _EVAL_136;
  assign _EVAL_1854 = _EVAL_1992[31:3];
  assign _EVAL_5390 = _EVAL_44;
  assign _EVAL_3822 = _EVAL_5390[31:3];
  assign _EVAL_4204 = _EVAL_1854 < _EVAL_3822;
  assign _EVAL_2127 = _EVAL_1854 == _EVAL_3822;
  assign _EVAL_3117 = _EVAL_5390[2:0];
  assign _EVAL_5381 = 3'h4 < _EVAL_3117;
  assign _EVAL_5561 = _EVAL_2127 & _EVAL_5381;
  assign _EVAL_3293 = _EVAL_4204 | _EVAL_5561;
  assign _EVAL_379 = _EVAL_5211[0];
  assign _EVAL_4444 = _EVAL_3293 == _EVAL_379;
  assign _EVAL_481 = _EVAL_5390[0];
  assign _EVAL_2618 = _EVAL_379 & _EVAL_481;
  assign _EVAL_439 = _EVAL_5390[1];
  assign _EVAL_550 = _EVAL_2618 & _EVAL_439;
  assign _EVAL_1763 = _EVAL_5390[2];
  assign _EVAL_4397 = _EVAL_550 & _EVAL_1763;
  assign _EVAL_5705 = {_EVAL_4397,_EVAL_550,_EVAL_2618,_EVAL_379};
  assign _EVAL_431 = 4'h3 | _EVAL_5705;
  assign _EVAL_1858 = ~ _EVAL_3117;
  assign _EVAL_3483 = {{1'd0}, _EVAL_1858};
  assign _EVAL_4626 = _EVAL_3483 | _EVAL_5705;
  assign _EVAL_1689 = _EVAL_431 == _EVAL_4626;
  assign _EVAL_3326 = _EVAL_2127 & _EVAL_1689;
  assign _EVAL_1283 = _EVAL_4914 ? _EVAL_4444 : _EVAL_3326;
  assign _EVAL_4867 = _EVAL_5393 & _EVAL_1283;
  assign _EVAL_6128 = _EVAL_2110 & _EVAL_4867;
  assign _EVAL_4732 = _EVAL_57;
  assign _EVAL_5875 = _EVAL_4732 == 1'h0;
  assign _EVAL_4630 = _EVAL_3997[0];
  assign _EVAL_3345 = _EVAL_5718 & _EVAL_4630;
  assign _EVAL_2781 = _EVAL_64;
  assign _EVAL_977 = _EVAL_3345 & _EVAL_2781;
  assign _EVAL_3807 = _EVAL_25;
  assign _EVAL_5680 = _EVAL_3807[1];
  assign _EVAL_3560 = _EVAL_102;
  assign _EVAL_2209 = _EVAL_3560[31:3];
  assign _EVAL_5844 = _EVAL_1854 < _EVAL_2209;
  assign _EVAL_5549 = _EVAL_1854 == _EVAL_2209;
  assign _EVAL_5107 = _EVAL_3560[2:0];
  assign _EVAL_719 = 3'h4 < _EVAL_5107;
  assign _EVAL_5702 = _EVAL_5549 & _EVAL_719;
  assign _EVAL_1914 = _EVAL_5844 | _EVAL_5702;
  assign _EVAL_3257 = _EVAL_3807[0];
  assign _EVAL_2111 = _EVAL_1914 == _EVAL_3257;
  assign _EVAL_2107 = _EVAL_3560[0];
  assign _EVAL_5426 = _EVAL_3257 & _EVAL_2107;
  assign _EVAL_1831 = _EVAL_3560[1];
  assign _EVAL_1408 = _EVAL_5426 & _EVAL_1831;
  assign _EVAL_3705 = _EVAL_3560[2];
  assign _EVAL_5459 = _EVAL_1408 & _EVAL_3705;
  assign _EVAL_3251 = {_EVAL_5459,_EVAL_1408,_EVAL_5426,_EVAL_3257};
  assign _EVAL_5435 = 4'h3 | _EVAL_3251;
  assign _EVAL_5809 = ~ _EVAL_5107;
  assign _EVAL_4935 = {{1'd0}, _EVAL_5809};
  assign _EVAL_920 = _EVAL_4935 | _EVAL_3251;
  assign _EVAL_2163 = _EVAL_5435 == _EVAL_920;
  assign _EVAL_4460 = _EVAL_5549 & _EVAL_2163;
  assign _EVAL_5220 = _EVAL_5680 ? _EVAL_2111 : _EVAL_4460;
  assign _EVAL_1006 = _EVAL_977 & _EVAL_5220;
  assign _EVAL_2524 = _EVAL_5875 | _EVAL_1006;
  assign _EVAL_6001 = _EVAL_6128 & _EVAL_2524;
  assign _EVAL_3477 = _EVAL_31;
  assign _EVAL_4922 = _EVAL_3382 & _EVAL_3477;
  assign _EVAL_5668 = 29'h0 < _EVAL_3822;
  assign _EVAL_1173 = 29'h0 == _EVAL_3822;
  assign _EVAL_4437 = _EVAL_1173 & _EVAL_5381;
  assign _EVAL_5698 = _EVAL_5668 | _EVAL_4437;
  assign _EVAL_5324 = _EVAL_5698 == _EVAL_379;
  assign _EVAL_2252 = _EVAL_1173 & _EVAL_1689;
  assign _EVAL_2993 = _EVAL_4914 ? _EVAL_5324 : _EVAL_2252;
  assign _EVAL_2093 = _EVAL_4922 & _EVAL_2993;
  assign _EVAL_3169 = _EVAL_2110 & _EVAL_2093;
  assign _EVAL_1383 = _EVAL_89;
  assign _EVAL_4063 = _EVAL_3345 & _EVAL_1383;
  assign _EVAL_2293 = 29'h0 < _EVAL_2209;
  assign _EVAL_5967 = 29'h0 == _EVAL_2209;
  assign _EVAL_3336 = _EVAL_5967 & _EVAL_719;
  assign _EVAL_169 = _EVAL_2293 | _EVAL_3336;
  assign _EVAL_3206 = _EVAL_169 == _EVAL_3257;
  assign _EVAL_3962 = _EVAL_5967 & _EVAL_2163;
  assign _EVAL_376 = _EVAL_5680 ? _EVAL_3206 : _EVAL_3962;
  assign _EVAL_165 = _EVAL_4063 & _EVAL_376;
  assign _EVAL_4359 = _EVAL_5875 | _EVAL_165;
  assign _EVAL_4985 = _EVAL_3169 & _EVAL_4359;
  assign _EVAL_3923 = _EVAL_72;
  assign _EVAL_3524 = _EVAL_3382 & _EVAL_3923;
  assign _EVAL_209 = _EVAL_3524 & _EVAL_2993;
  assign _EVAL_2108 = _EVAL_2110 & _EVAL_209;
  assign _EVAL_2606 = _EVAL_6;
  assign _EVAL_6086 = _EVAL_3345 & _EVAL_2606;
  assign _EVAL_4214 = _EVAL_6086 & _EVAL_376;
  assign _EVAL_3846 = _EVAL_5875 | _EVAL_4214;
  assign _EVAL_868 = _EVAL_2108 & _EVAL_3846;
  assign _EVAL_2469 = _EVAL_4985 ? 1'h1 : _EVAL_868;
  assign _EVAL_881 = _EVAL_6001 ? 1'h1 : _EVAL_2469;
  assign _EVAL_2491 = 3'h0 < _EVAL_3117;
  assign _EVAL_5443 = _EVAL_1173 & _EVAL_2491;
  assign _EVAL_1322 = _EVAL_5668 | _EVAL_5443;
  assign _EVAL_4104 = _EVAL_1322 == _EVAL_379;
  assign _EVAL_1700 = 4'h7 | _EVAL_5705;
  assign _EVAL_3143 = _EVAL_1700 == _EVAL_4626;
  assign _EVAL_1633 = _EVAL_1173 & _EVAL_3143;
  assign _EVAL_2213 = _EVAL_4914 ? _EVAL_4104 : _EVAL_1633;
  assign _EVAL_3402 = _EVAL_3524 & _EVAL_2213;
  assign _EVAL_1342 = _EVAL_2110 & _EVAL_3402;
  assign _EVAL_2837 = _EVAL_654[1:0];
  assign _EVAL_1958 = _EVAL_2837 == 2'h1;
  assign _EVAL_3242 = _EVAL_334[12];
  assign _EVAL_1670 = _EVAL_334[4:1];
  assign _EVAL_5385 = _EVAL_334[11];
  assign _EVAL_2375 = {_EVAL_3242,_EVAL_5403,5'h0,2'h1,_EVAL_4771,3'h1,_EVAL_1670,_EVAL_5385,7'h63};
  assign _EVAL_4964 = {_EVAL_3242,_EVAL_5403,5'h0,2'h1,_EVAL_4771,3'h0,_EVAL_1670,_EVAL_5385,7'h63};
  assign _EVAL_4199 = _EVAL_3082 ? 10'h3ff : 10'h0;
  assign _EVAL_2817 = _EVAL_654[8];
  assign _EVAL_1211 = _EVAL_654[10:9];
  assign _EVAL_581 = _EVAL_654[6];
  assign _EVAL_4521 = _EVAL_654[7];
  assign _EVAL_2557 = _EVAL_654[11];
  assign _EVAL_2977 = _EVAL_654[5:3];
  assign _EVAL_5750 = {_EVAL_4199,_EVAL_2817,_EVAL_1211,_EVAL_581,_EVAL_4521,_EVAL_218,_EVAL_2557,_EVAL_2977,1'h0};
  assign _EVAL_3334 = _EVAL_5750[20];
  assign _EVAL_673 = _EVAL_5750[10:1];
  assign _EVAL_3399 = _EVAL_5750[11];
  assign _EVAL_2699 = _EVAL_5750[19:12];
  assign _EVAL_2011 = {_EVAL_3334,_EVAL_673,_EVAL_3399,_EVAL_2699,5'h0,7'h6f};
  assign _EVAL_3863 = _EVAL_948 == 2'h3;
  assign _EVAL_4148 = {_EVAL_3082,_EVAL_4575};
  assign _EVAL_5258 = _EVAL_4148 == 3'h7;
  assign _EVAL_923 = _EVAL_4148 == 3'h6;
  assign _EVAL_1428 = _EVAL_4148 == 3'h5;
  assign _EVAL_5313 = _EVAL_4148 == 3'h4;
  assign _EVAL_2860 = _EVAL_4148 == 3'h3;
  assign _EVAL_2913 = _EVAL_4148 == 3'h2;
  assign _EVAL_175 = _EVAL_4148 == 3'h1;
  assign _EVAL_356 = _EVAL_175 ? 3'h4 : 3'h0;
  assign _EVAL_5286 = _EVAL_2913 ? 3'h6 : _EVAL_356;
  assign _EVAL_1393 = _EVAL_2860 ? 3'h7 : _EVAL_5286;
  assign _EVAL_1627 = _EVAL_5313 ? 3'h0 : _EVAL_1393;
  assign _EVAL_2624 = _EVAL_1428 ? 3'h0 : _EVAL_1627;
  assign _EVAL_1575 = _EVAL_923 ? 3'h2 : _EVAL_2624;
  assign _EVAL_4092 = _EVAL_5258 ? 3'h3 : _EVAL_1575;
  assign _EVAL_1453 = _EVAL_3082 ? 7'h3b : 7'h33;
  assign _EVAL_5141 = {2'h1,_EVAL_2231,2'h1,_EVAL_4771,_EVAL_4092,2'h1,_EVAL_4771,_EVAL_1453};
  assign _EVAL_2240 = {{6'd0}, _EVAL_5141};
  assign _EVAL_278 = _EVAL_4575 == 2'h0;
  assign _EVAL_3972 = {_EVAL_278, 30'h0};
  assign _EVAL_4308 = _EVAL_2240 | _EVAL_3972;
  assign _EVAL_3802 = _EVAL_948 == 2'h2;
  assign _EVAL_1802 = _EVAL_3082 ? 7'h7f : 7'h0;
  assign _EVAL_4154 = {_EVAL_1802,_EVAL_1321,2'h1,_EVAL_4771,3'h7,2'h1,_EVAL_4771,7'h13};
  assign _EVAL_2914 = _EVAL_948 == 2'h1;
  assign _EVAL_5870 = {_EVAL_3082,_EVAL_1321,2'h1,_EVAL_4771,3'h5,2'h1,_EVAL_4771,7'h13};
  assign _EVAL_2134 = {{5'd0}, _EVAL_5870};
  assign _EVAL_4842 = _EVAL_2134 | 31'h40000000;
  assign _EVAL_415 = _EVAL_2914 ? _EVAL_4842 : {{5'd0}, _EVAL_5870};
  assign _EVAL_2437 = _EVAL_3802 ? _EVAL_4154 : {{1'd0}, _EVAL_415};
  assign _EVAL_5781 = _EVAL_3863 ? {{1'd0}, _EVAL_4308} : _EVAL_2437;
  assign _EVAL_4230 = _EVAL_4094 == 5'h2;
  assign _EVAL_5609 = _EVAL_3082 ? 3'h7 : 3'h0;
  assign _EVAL_1095 = _EVAL_654[5];
  assign _EVAL_5429 = {_EVAL_5609,_EVAL_3864,_EVAL_1095,_EVAL_218,_EVAL_581,4'h0,_EVAL_4094,3'h0,_EVAL_4094,7'h13};
  assign _EVAL_2178 = _EVAL_3082 ? 15'h7fff : 15'h0;
  assign _EVAL_1528 = {_EVAL_2178,_EVAL_1321,12'h0};
  assign _EVAL_755 = _EVAL_1528[31:12];
  assign _EVAL_1950 = {_EVAL_755,_EVAL_4094,7'h37};
  assign _EVAL_371 = _EVAL_4230 ? _EVAL_5429 : _EVAL_1950;
  assign _EVAL_3507 = {_EVAL_1802,_EVAL_1321,5'h0,3'h0,_EVAL_4094,7'h13};
  assign _EVAL_3518 = {_EVAL_3334,_EVAL_673,_EVAL_3399,_EVAL_2699,5'h1,7'h6f};
  assign _EVAL_642 = {_EVAL_1802,_EVAL_1321,_EVAL_4094,3'h0,_EVAL_4094,7'h13};
  assign _EVAL_2214 = _EVAL_3016 ? _EVAL_3518 : _EVAL_642;
  assign _EVAL_2200 = _EVAL_5989 ? _EVAL_3507 : _EVAL_2214;
  assign _EVAL_2279 = _EVAL_761 ? _EVAL_371 : _EVAL_2200;
  assign _EVAL_5175 = _EVAL_4440 ? _EVAL_5781 : _EVAL_2279;
  assign _EVAL_4697 = _EVAL_1378 ? _EVAL_2011 : _EVAL_5175;
  assign _EVAL_1498 = _EVAL_537 ? _EVAL_4964 : _EVAL_4697;
  assign _EVAL_5813 = _EVAL_1088 ? _EVAL_2375 : _EVAL_1498;
  assign _EVAL_3032 = _EVAL_5813[6:2];
  assign _EVAL_4947 = {_EVAL_1095,_EVAL_2483,_EVAL_581,2'h0};
  assign _EVAL_780 = _EVAL_4947[6:5];
  assign _EVAL_5149 = _EVAL_4947[4:0];
  assign _EVAL_1587 = {_EVAL_780,2'h1,_EVAL_2231,2'h1,_EVAL_4771,3'h2,_EVAL_5149,7'h27};
  assign _EVAL_1934 = {_EVAL_780,2'h1,_EVAL_2231,2'h1,_EVAL_4771,3'h2,_EVAL_5149,7'h23};
  assign _EVAL_3815 = {_EVAL_4575,_EVAL_2483,3'h0};
  assign _EVAL_4593 = _EVAL_3815[7:5];
  assign _EVAL_3988 = _EVAL_3815[4:0];
  assign _EVAL_6113 = {_EVAL_4593,2'h1,_EVAL_2231,2'h1,_EVAL_4771,3'h3,_EVAL_3988,7'h27};
  assign _EVAL_2933 = {_EVAL_780,2'h1,_EVAL_2231,2'h1,_EVAL_4771,3'h0,_EVAL_5149,7'h27};
  assign _EVAL_4194 = {_EVAL_1095,_EVAL_2483,_EVAL_581,2'h0,2'h1,_EVAL_4771,3'h2,2'h1,_EVAL_2231,7'h7};
  assign _EVAL_1940 = {_EVAL_1095,_EVAL_2483,_EVAL_581,2'h0,2'h1,_EVAL_4771,3'h2,2'h1,_EVAL_2231,7'h3};
  assign _EVAL_2805 = {_EVAL_4575,_EVAL_2483,3'h0,2'h1,_EVAL_4771,3'h3,2'h1,_EVAL_2231,7'h7};
  assign _EVAL_2047 = _EVAL_654[10:7];
  assign _EVAL_252 = _EVAL_654[12:11];
  assign _EVAL_894 = {_EVAL_2047,_EVAL_252,_EVAL_1095,_EVAL_581,2'h0,5'h2,3'h0,2'h1,_EVAL_2231,7'h13};
  assign _EVAL_328 = _EVAL_3016 ? {{2'd0}, _EVAL_2805} : _EVAL_894;
  assign _EVAL_5593 = _EVAL_5989 ? {{3'd0}, _EVAL_1940} : _EVAL_328;
  assign _EVAL_3319 = _EVAL_761 ? {{3'd0}, _EVAL_4194} : _EVAL_5593;
  assign _EVAL_5487 = _EVAL_4440 ? {{3'd0}, _EVAL_2933} : _EVAL_3319;
  assign _EVAL_2597 = _EVAL_1378 ? {{2'd0}, _EVAL_6113} : _EVAL_5487;
  assign _EVAL_5123 = _EVAL_537 ? {{3'd0}, _EVAL_1934} : _EVAL_2597;
  assign _EVAL_1103 = _EVAL_1088 ? {{3'd0}, _EVAL_1587} : _EVAL_5123;
  assign _EVAL_1947 = {2'h0,_EVAL_1103};
  assign _EVAL_2720 = _EVAL_1947[6:2];
  assign _EVAL_3562 = _EVAL_1958 ? _EVAL_3032 : _EVAL_2720;
  assign _EVAL_3628 = _EVAL_735 ? 5'h1f : 5'h0;
  assign _EVAL_5099 = _EVAL_3455[2];
  assign _EVAL_5712 = _EVAL_3455[11:10];
  assign _EVAL_1187 = _EVAL_3455[4:3];
  assign _EVAL_5663 = {_EVAL_3628,_EVAL_5278,_EVAL_5099,_EVAL_5712,_EVAL_1187,1'h0};
  assign _EVAL_554 = _EVAL_5663[12];
  assign _EVAL_1316 = _EVAL_5663[10:5];
  assign _EVAL_2050 = _EVAL_5663[4:1];
  assign _EVAL_3015 = _EVAL_5663[11];
  assign _EVAL_4903 = {_EVAL_554,_EVAL_1316,5'h0,2'h1,_EVAL_4872,3'h1,_EVAL_2050,_EVAL_3015,7'h63};
  assign _EVAL_5375 = {_EVAL_554,_EVAL_1316,5'h0,2'h1,_EVAL_4872,3'h0,_EVAL_2050,_EVAL_3015,7'h63};
  assign _EVAL_5334 = _EVAL_735 ? 10'h3ff : 10'h0;
  assign _EVAL_1491 = _EVAL_3455[8];
  assign _EVAL_4013 = _EVAL_3455[10:9];
  assign _EVAL_1170 = _EVAL_3455[7];
  assign _EVAL_2315 = _EVAL_3455[11];
  assign _EVAL_1140 = _EVAL_3455[5:3];
  assign _EVAL_5342 = {_EVAL_5334,_EVAL_1491,_EVAL_4013,_EVAL_2996,_EVAL_1170,_EVAL_5099,_EVAL_2315,_EVAL_1140,1'h0};
  assign _EVAL_5903 = _EVAL_5342[20];
  assign _EVAL_5716 = _EVAL_5342[10:1];
  assign _EVAL_5891 = _EVAL_5342[11];
  assign _EVAL_2926 = _EVAL_5342[19:12];
  assign _EVAL_1686 = {_EVAL_5903,_EVAL_5716,_EVAL_5891,_EVAL_2926,5'h0,7'h6f};
  assign _EVAL_4224 = _EVAL_5712 == 2'h3;
  assign _EVAL_913 = {{6'd0}, _EVAL_3408};
  assign _EVAL_4827 = _EVAL_5278 == 2'h0;
  assign _EVAL_1169 = {_EVAL_4827, 30'h0};
  assign _EVAL_5533 = _EVAL_913 | _EVAL_1169;
  assign _EVAL_4062 = _EVAL_5712 == 2'h2;
  assign _EVAL_2007 = _EVAL_735 ? 7'h7f : 7'h0;
  assign _EVAL_3113 = {_EVAL_2007,_EVAL_2075,2'h1,_EVAL_4872,3'h7,2'h1,_EVAL_4872,7'h13};
  assign _EVAL_2461 = _EVAL_5712 == 2'h1;
  assign _EVAL_2113 = {_EVAL_735,_EVAL_2075,2'h1,_EVAL_4872,3'h5,2'h1,_EVAL_4872,7'h13};
  assign _EVAL_512 = {{5'd0}, _EVAL_2113};
  assign _EVAL_830 = _EVAL_512 | 31'h40000000;
  assign _EVAL_4813 = _EVAL_2461 ? _EVAL_830 : {{5'd0}, _EVAL_2113};
  assign _EVAL_2673 = _EVAL_4062 ? _EVAL_3113 : {{1'd0}, _EVAL_4813};
  assign _EVAL_2005 = _EVAL_4224 ? {{1'd0}, _EVAL_5533} : _EVAL_2673;
  assign _EVAL_1681 = _EVAL_3655 == 5'h2;
  assign _EVAL_4764 = _EVAL_735 ? 3'h7 : 3'h0;
  assign _EVAL_705 = {_EVAL_4764,_EVAL_1187,_EVAL_241,_EVAL_5099,_EVAL_2996,4'h0,_EVAL_3655,3'h0,_EVAL_3655,7'h13};
  assign _EVAL_4362 = _EVAL_735 ? 15'h7fff : 15'h0;
  assign _EVAL_3453 = {_EVAL_4362,_EVAL_2075,12'h0};
  assign _EVAL_2749 = _EVAL_3453[31:12];
  assign _EVAL_5689 = {_EVAL_2749,_EVAL_3655,7'h37};
  assign _EVAL_5672 = _EVAL_1681 ? _EVAL_705 : _EVAL_5689;
  assign _EVAL_4561 = {_EVAL_2007,_EVAL_2075,5'h0,3'h0,_EVAL_3655,7'h13};
  assign _EVAL_4799 = {_EVAL_5903,_EVAL_5716,_EVAL_5891,_EVAL_2926,5'h1,7'h6f};
  assign _EVAL_2503 = {_EVAL_2007,_EVAL_2075,_EVAL_3655,3'h0,_EVAL_3655,7'h13};
  assign _EVAL_4894 = _EVAL_5755 ? _EVAL_4799 : _EVAL_2503;
  assign _EVAL_5759 = _EVAL_597 ? _EVAL_4561 : _EVAL_4894;
  assign _EVAL_1927 = _EVAL_1674 ? _EVAL_5672 : _EVAL_5759;
  assign _EVAL_5964 = _EVAL_936 ? _EVAL_2005 : _EVAL_1927;
  assign _EVAL_5076 = _EVAL_453 ? _EVAL_1686 : _EVAL_5964;
  assign _EVAL_479 = _EVAL_2288 ? _EVAL_5375 : _EVAL_5076;
  assign _EVAL_1242 = _EVAL_4669 ? _EVAL_4903 : _EVAL_479;
  assign _EVAL_5851 = _EVAL_1242 & 32'h705b;
  assign _EVAL_1280 = _EVAL_5851 == 32'h2003;
  assign _EVAL_2710 = _EVAL_1362 & 32'h207f;
  assign _EVAL_4647 = _EVAL_2710 == 32'h2073;
  assign _EVAL_5315 = _EVAL_2039 & 32'h80000010;
  assign _EVAL_4478 = _EVAL_5315 == 32'h10;
  assign _EVAL_2445 = _EVAL_2039 & 32'h50;
  assign _EVAL_1275 = _EVAL_2445 == 32'h10;
  assign _EVAL_5396 = _EVAL_4478 | _EVAL_1275;
  assign _EVAL_5938 = _EVAL_2039 & 32'h40000040;
  assign _EVAL_449 = _EVAL_5938 == 32'h40;
  assign _EVAL_4286 = _EVAL_5396 | _EVAL_449;
  assign _EVAL_365 = _EVAL_4882 & 32'h2048;
  assign _EVAL_4689 = _EVAL_27;
  assign _EVAL_5201 = _EVAL_4689[31:3];
  assign _EVAL_4226 = _EVAL_1854 == _EVAL_5201;
  assign _EVAL_4177 = _EVAL_139;
  assign _EVAL_383 = _EVAL_4177[0];
  assign _EVAL_5369 = _EVAL_4689[0];
  assign _EVAL_5505 = _EVAL_383 & _EVAL_5369;
  assign _EVAL_486 = _EVAL_4689[1];
  assign _EVAL_4172 = _EVAL_5505 & _EVAL_486;
  assign _EVAL_4140 = _EVAL_4689[2];
  assign _EVAL_5893 = _EVAL_4172 & _EVAL_4140;
  assign _EVAL_3550 = {_EVAL_5893,_EVAL_4172,_EVAL_5505,_EVAL_383};
  assign _EVAL_3406 = 4'h3 | _EVAL_3550;
  assign _EVAL_1773 = _EVAL_4689[2:0];
  assign _EVAL_2975 = ~ _EVAL_1773;
  assign _EVAL_4318 = {{1'd0}, _EVAL_2975};
  assign _EVAL_4784 = _EVAL_4318 | _EVAL_3550;
  assign _EVAL_5997 = _EVAL_3406 == _EVAL_4784;
  assign _EVAL_2968 = _EVAL_4226 & _EVAL_5997;
  assign _EVAL_3370 = 3'h2 < _EVAL_3117;
  assign _EVAL_1779 = _EVAL_1173 & _EVAL_3370;
  assign _EVAL_3679 = _EVAL_5668 | _EVAL_1779;
  assign _EVAL_1808 = _EVAL_3679 == _EVAL_379;
  assign _EVAL_4633 = 4'h5 | _EVAL_5705;
  assign _EVAL_1323 = _EVAL_4633 == _EVAL_4626;
  assign _EVAL_646 = _EVAL_1173 & _EVAL_1323;
  assign _EVAL_5187 = _EVAL_4914 ? _EVAL_1808 : _EVAL_646;
  assign _EVAL_935 = _EVAL_4922 & _EVAL_5187;
  assign _EVAL_2547 = _EVAL_2110 & _EVAL_935;
  assign _EVAL_2371 = 3'h2 < _EVAL_5107;
  assign _EVAL_5740 = _EVAL_5967 & _EVAL_2371;
  assign _EVAL_4050 = _EVAL_2293 | _EVAL_5740;
  assign _EVAL_4302 = _EVAL_4050 == _EVAL_3257;
  assign _EVAL_1715 = 4'h5 | _EVAL_3251;
  assign _EVAL_2486 = _EVAL_1715 == _EVAL_920;
  assign _EVAL_2758 = _EVAL_5967 & _EVAL_2486;
  assign _EVAL_952 = _EVAL_5680 ? _EVAL_4302 : _EVAL_2758;
  assign _EVAL_2194 = _EVAL_4063 & _EVAL_952;
  assign _EVAL_6065 = _EVAL_5875 | _EVAL_2194;
  assign _EVAL_3460 = _EVAL_2547 & _EVAL_6065;
  assign _EVAL_1882 = _EVAL_4743 & 32'h707b;
  assign _EVAL_222 = _EVAL_67;
  assign _EVAL_574 = _EVAL_222 == 1'h0;
  assign _EVAL_1649 = _EVAL_24;
  assign _EVAL_600 = _EVAL_156;
  assign _EVAL_284 = {_EVAL_1649,1'h0,1'h0,_EVAL_600};
  assign _EVAL_651 = _EVAL_284 >> _EVAL_4188;
  assign _EVAL_4453 = _EVAL_651[0];
  assign _EVAL_4492 = _EVAL_5718 & _EVAL_4453;
  assign _EVAL_2940 = _EVAL_147;
  assign _EVAL_5039 = _EVAL_4492 & _EVAL_2940;
  assign _EVAL_1766 = _EVAL_56;
  assign _EVAL_4291 = _EVAL_1766[1];
  assign _EVAL_2539 = _EVAL_126;
  assign _EVAL_2382 = _EVAL_2539[31:3];
  assign _EVAL_1310 = _EVAL_1854 < _EVAL_2382;
  assign _EVAL_584 = _EVAL_1854 == _EVAL_2382;
  assign _EVAL_3401 = _EVAL_2539[2:0];
  assign _EVAL_979 = 3'h6 < _EVAL_3401;
  assign _EVAL_1429 = _EVAL_584 & _EVAL_979;
  assign _EVAL_505 = _EVAL_1310 | _EVAL_1429;
  assign _EVAL_1969 = _EVAL_1766[0];
  assign _EVAL_4193 = _EVAL_505 == _EVAL_1969;
  assign _EVAL_2372 = _EVAL_2539[0];
  assign _EVAL_1905 = _EVAL_1969 & _EVAL_2372;
  assign _EVAL_1336 = _EVAL_2539[1];
  assign _EVAL_2585 = _EVAL_1905 & _EVAL_1336;
  assign _EVAL_5867 = _EVAL_2539[2];
  assign _EVAL_4513 = _EVAL_2585 & _EVAL_5867;
  assign _EVAL_4534 = {_EVAL_4513,_EVAL_2585,_EVAL_1905,_EVAL_1969};
  assign _EVAL_1289 = 4'h1 | _EVAL_4534;
  assign _EVAL_4221 = ~ _EVAL_3401;
  assign _EVAL_5530 = {{1'd0}, _EVAL_4221};
  assign _EVAL_3975 = _EVAL_5530 | _EVAL_4534;
  assign _EVAL_3373 = _EVAL_1289 == _EVAL_3975;
  assign _EVAL_4200 = _EVAL_584 & _EVAL_3373;
  assign _EVAL_2651 = _EVAL_4291 ? _EVAL_4193 : _EVAL_4200;
  assign _EVAL_1558 = _EVAL_5039 & _EVAL_2651;
  assign _EVAL_4719 = _EVAL_574 & _EVAL_1558;
  assign _EVAL_2646 = 3'h6 < _EVAL_3117;
  assign _EVAL_4220 = _EVAL_2127 & _EVAL_2646;
  assign _EVAL_2255 = _EVAL_4204 | _EVAL_4220;
  assign _EVAL_5826 = _EVAL_2255 == _EVAL_379;
  assign _EVAL_2642 = 4'h1 | _EVAL_5705;
  assign _EVAL_2874 = _EVAL_2642 == _EVAL_4626;
  assign _EVAL_1084 = _EVAL_2127 & _EVAL_2874;
  assign _EVAL_2430 = _EVAL_4914 ? _EVAL_5826 : _EVAL_1084;
  assign _EVAL_1928 = _EVAL_5393 & _EVAL_2430;
  assign _EVAL_3392 = _EVAL_2110 | _EVAL_1928;
  assign _EVAL_1365 = _EVAL_4719 & _EVAL_3392;
  assign _EVAL_1395 = _EVAL_5813 & 32'h10000060;
  assign _EVAL_3570 = _EVAL_4728 == 2'h2;
  assign _EVAL_1184 = _EVAL_4743 & 32'h207f;
  assign _EVAL_1302 = _EVAL_1184 == 32'h3;
  assign _EVAL_2555 = _EVAL_4743 & 32'h607f;
  assign _EVAL_4333 = _EVAL_2555 == 32'hf;
  assign _EVAL_1477 = _EVAL_1302 | _EVAL_4333;
  assign _EVAL_5093 = _EVAL_4743 & 32'h5f;
  assign _EVAL_410 = _EVAL_5093 == 32'h17;
  assign _EVAL_4325 = _EVAL_1477 | _EVAL_410;
  assign _EVAL_4211 = _EVAL_4743 & 32'hfc00007f;
  assign _EVAL_1265 = _EVAL_4211 == 32'h33;
  assign _EVAL_5227 = _EVAL_4325 | _EVAL_1265;
  assign _EVAL_4801 = _EVAL_4743 & 32'hbe00707f;
  assign _EVAL_2845 = _EVAL_4801 == 32'h33;
  assign _EVAL_3957 = _EVAL_5227 | _EVAL_2845;
  assign _EVAL_2937 = _EVAL_4743 & 32'h6000073;
  assign _EVAL_1384 = _EVAL_2937 == 32'h43;
  assign _EVAL_2777 = _EVAL_3957 | _EVAL_1384;
  assign _EVAL_2819 = _EVAL_4743 & 32'he600007f;
  assign _EVAL_2150 = _EVAL_2819 == 32'h53;
  assign _EVAL_5754 = _EVAL_2777 | _EVAL_2150;
  assign _EVAL_4501 = _EVAL_1882 == 32'h63;
  assign _EVAL_1910 = _EVAL_5754 | _EVAL_4501;
  assign _EVAL_1255 = _EVAL_4743 & 32'h7f;
  assign _EVAL_2545 = _EVAL_1255 == 32'h6f;
  assign _EVAL_841 = _EVAL_1910 | _EVAL_2545;
  assign _EVAL_446 = _EVAL_4743 & 32'hffefffff;
  assign _EVAL_4572 = _EVAL_446 == 32'h73;
  assign _EVAL_5462 = _EVAL_841 | _EVAL_4572;
  assign _EVAL_3041 = _EVAL_4743 & 32'hfe00305f;
  assign _EVAL_662 = _EVAL_3041 == 32'h1013;
  assign _EVAL_1244 = _EVAL_5462 | _EVAL_662;
  assign _EVAL_2505 = _EVAL_4743 & 32'h705b;
  assign _EVAL_2782 = _EVAL_2505 == 32'h2003;
  assign _EVAL_5570 = _EVAL_1244 | _EVAL_2782;
  assign _EVAL_3538 = _EVAL_1184 == 32'h2013;
  assign _EVAL_463 = _EVAL_5570 | _EVAL_3538;
  assign _EVAL_322 = _EVAL_4743 & 32'h1800707f;
  assign _EVAL_4892 = _EVAL_322 == 32'h202f;
  assign _EVAL_2559 = _EVAL_463 | _EVAL_4892;
  assign _EVAL_5359 = _EVAL_1184 == 32'h2073;
  assign _EVAL_689 = _EVAL_2559 | _EVAL_5359;
  assign _EVAL_5420 = _EVAL_4743 & 32'hbe00705f;
  assign _EVAL_1560 = _EVAL_5420 == 32'h5013;
  assign _EVAL_377 = _EVAL_689 | _EVAL_1560;
  assign _EVAL_4808 = _EVAL_4743 & 32'he800707f;
  assign _EVAL_4208 = _EVAL_4808 == 32'h800202f;
  assign _EVAL_3157 = _EVAL_377 | _EVAL_4208;
  assign _EVAL_4482 = _EVAL_4743 & 32'hf9f0707f;
  assign _EVAL_3054 = _EVAL_4482 == 32'h1000202f;
  assign _EVAL_2785 = _EVAL_3157 | _EVAL_3054;
  assign _EVAL_480 = _EVAL_4743 & 32'hdfffffff;
  assign _EVAL_3970 = _EVAL_480 == 32'h10500073;
  assign _EVAL_1724 = _EVAL_2785 | _EVAL_3970;
  assign _EVAL_3608 = _EVAL_4743 & 32'hf600607f;
  assign _EVAL_5391 = _EVAL_3608 == 32'h20000053;
  assign _EVAL_4654 = _EVAL_1724 | _EVAL_5391;
  assign _EVAL_2947 = _EVAL_4743 & 32'h7e00607f;
  assign _EVAL_162 = _EVAL_2947 == 32'h20000053;
  assign _EVAL_4817 = _EVAL_4654 | _EVAL_162;
  assign _EVAL_2714 = _EVAL_4882 & 32'h90000034;
  assign _EVAL_4361 = _EVAL_3006 & 32'h18;
  assign _EVAL_2672 = _EVAL_4361 == 32'h0;
  assign _EVAL_197 = _EVAL_2837 == 2'h3;
  assign _EVAL_1525 = 1'h0 < _EVAL_197;
  assign _EVAL_5845 = _EVAL_5994 & _EVAL_1525;
  assign _EVAL_3010 = _EVAL_136[2:1];
  assign _EVAL_3528 = _EVAL_5648 ? _EVAL_3403 : _EVAL_3010;
  assign _EVAL_1371 = 2'h0 >= _EVAL_3528;
  assign _EVAL_5276 = _EVAL_5845 ? 1'h0 : _EVAL_1371;
  assign _EVAL_5833 = _EVAL_4728 == 2'h3;
  assign _EVAL_4360 = 1'h0 < _EVAL_5833;
  assign _EVAL_2513 = _EVAL_5276 & _EVAL_4360;
  assign _EVAL_1061 = 2'h1 >= _EVAL_3528;
  assign _EVAL_3052 = _EVAL_2513 ? 1'h0 : _EVAL_1061;
  assign _EVAL_3573 = _EVAL_3455[1:0];
  assign _EVAL_2970 = _EVAL_3573 == 2'h3;
  assign _EVAL_4887 = 1'h0 < _EVAL_2970;
  assign _EVAL_2051 = _EVAL_3052 & _EVAL_4887;
  assign _EVAL_3045 = 2'h2 >= _EVAL_3528;
  assign _EVAL_2142 = _EVAL_2051 ? 1'h0 : _EVAL_3045;
  assign _EVAL_2797 = _EVAL_2142 ? 2'h2 : 2'h3;
  assign _EVAL_4231 = _EVAL_3052 ? 2'h1 : _EVAL_2797;
  assign _EVAL_1213 = {_EVAL_1329,_EVAL_821,_EVAL_5340,2'h0};
  assign _EVAL_5685 = _EVAL_1213[6:5];
  assign _EVAL_2915 = _EVAL_1213[4:0];
  assign _EVAL_5067 = {_EVAL_5685,2'h1,_EVAL_5741,2'h1,_EVAL_1375,3'h2,_EVAL_2915,7'h27};
  assign _EVAL_2744 = {_EVAL_5685,2'h1,_EVAL_5741,2'h1,_EVAL_1375,3'h2,_EVAL_2915,7'h23};
  assign _EVAL_4236 = {_EVAL_3105,_EVAL_821,3'h0};
  assign _EVAL_1545 = _EVAL_4236[7:5];
  assign _EVAL_747 = _EVAL_4236[4:0];
  assign _EVAL_3951 = {_EVAL_1545,2'h1,_EVAL_5741,2'h1,_EVAL_1375,3'h3,_EVAL_747,7'h27};
  assign _EVAL_595 = {_EVAL_5685,2'h1,_EVAL_5741,2'h1,_EVAL_1375,3'h0,_EVAL_2915,7'h27};
  assign _EVAL_4337 = {_EVAL_1329,_EVAL_821,_EVAL_5340,2'h0,2'h1,_EVAL_1375,3'h2,2'h1,_EVAL_5741,7'h7};
  assign _EVAL_2622 = {_EVAL_1329,_EVAL_821,_EVAL_5340,2'h0,2'h1,_EVAL_1375,3'h2,2'h1,_EVAL_5741,7'h3};
  assign _EVAL_4314 = {_EVAL_3105,_EVAL_821,3'h0,2'h1,_EVAL_1375,3'h3,2'h1,_EVAL_5741,7'h7};
  assign _EVAL_667 = _EVAL_2666[10:7];
  assign _EVAL_3835 = _EVAL_2666[12:11];
  assign _EVAL_5603 = {_EVAL_667,_EVAL_3835,_EVAL_1329,_EVAL_5340,2'h0,5'h2,3'h0,2'h1,_EVAL_5741,7'h13};
  assign _EVAL_1544 = _EVAL_630 ? {{2'd0}, _EVAL_4314} : _EVAL_5603;
  assign _EVAL_3752 = _EVAL_1014 ? {{3'd0}, _EVAL_2622} : _EVAL_1544;
  assign _EVAL_6003 = _EVAL_4352 ? {{3'd0}, _EVAL_4337} : _EVAL_3752;
  assign _EVAL_3614 = _EVAL_4202 ? {{3'd0}, _EVAL_595} : _EVAL_6003;
  assign _EVAL_708 = _EVAL_2644 ? {{2'd0}, _EVAL_3951} : _EVAL_3614;
  assign _EVAL_5962 = _EVAL_5821 ? {{3'd0}, _EVAL_2744} : _EVAL_708;
  assign _EVAL_2878 = _EVAL_418 ? {{3'd0}, _EVAL_5067} : _EVAL_5962;
  assign _EVAL_3271 = {2'h0,_EVAL_2878};
  assign _EVAL_3897 = _EVAL_3271 & 32'h207f;
  assign _EVAL_2771 = _EVAL_3897 == 32'h3;
  assign _EVAL_2034 = _EVAL_3271 & 32'h607f;
  assign _EVAL_1077 = _EVAL_2034 == 32'hf;
  assign _EVAL_1079 = _EVAL_2771 | _EVAL_1077;
  assign _EVAL_6088 = _EVAL_3271 & 32'h5f;
  assign _EVAL_2192 = _EVAL_6088 == 32'h17;
  assign _EVAL_3280 = _EVAL_1079 | _EVAL_2192;
  assign _EVAL_205 = _EVAL_3271 & 32'hfc00007f;
  assign _EVAL_4368 = _EVAL_205 == 32'h33;
  assign _EVAL_3650 = _EVAL_3280 | _EVAL_4368;
  assign _EVAL_5535 = _EVAL_3271 & 32'hbe00707f;
  assign _EVAL_1855 = _EVAL_5535 == 32'h33;
  assign _EVAL_5970 = _EVAL_3650 | _EVAL_1855;
  assign _EVAL_1413 = _EVAL_3271 & 32'h6000073;
  assign _EVAL_4228 = _EVAL_1413 == 32'h43;
  assign _EVAL_5969 = _EVAL_5970 | _EVAL_4228;
  assign _EVAL_303 = _EVAL_3271 & 32'he600007f;
  assign _EVAL_4726 = _EVAL_303 == 32'h53;
  assign _EVAL_571 = _EVAL_5969 | _EVAL_4726;
  assign _EVAL_5115 = _EVAL_3271 & 32'h707b;
  assign _EVAL_1531 = _EVAL_5115 == 32'h63;
  assign _EVAL_5675 = _EVAL_571 | _EVAL_1531;
  assign _EVAL_3380 = _EVAL_3271 & 32'h7f;
  assign _EVAL_1328 = _EVAL_3380 == 32'h6f;
  assign _EVAL_3867 = _EVAL_5675 | _EVAL_1328;
  assign _EVAL_3678 = _EVAL_3271 & 32'hffefffff;
  assign _EVAL_1542 = _EVAL_3678 == 32'h73;
  assign _EVAL_683 = _EVAL_3867 | _EVAL_1542;
  assign _EVAL_3309 = _EVAL_3271 & 32'hfe00305f;
  assign _EVAL_2183 = _EVAL_3309 == 32'h1013;
  assign _EVAL_427 = _EVAL_683 | _EVAL_2183;
  assign _EVAL_5836 = _EVAL_3271 & 32'h705b;
  assign _EVAL_1971 = _EVAL_5836 == 32'h2003;
  assign _EVAL_2520 = _EVAL_427 | _EVAL_1971;
  assign _EVAL_3684 = _EVAL_3897 == 32'h2013;
  assign _EVAL_5190 = _EVAL_2520 | _EVAL_3684;
  assign _EVAL_3112 = _EVAL_3271 & 32'h1800707f;
  assign _EVAL_3118 = _EVAL_3112 == 32'h202f;
  assign _EVAL_2792 = _EVAL_5190 | _EVAL_3118;
  assign _EVAL_2156 = _EVAL_3897 == 32'h2073;
  assign _EVAL_4474 = _EVAL_2792 | _EVAL_2156;
  assign _EVAL_2391 = _EVAL_3271 & 32'hbe00705f;
  assign _EVAL_5695 = _EVAL_2391 == 32'h5013;
  assign _EVAL_3506 = _EVAL_4474 | _EVAL_5695;
  assign _EVAL_5860 = _EVAL_3271 & 32'he800707f;
  assign _EVAL_5543 = _EVAL_5860 == 32'h800202f;
  assign _EVAL_2892 = _EVAL_3506 | _EVAL_5543;
  assign _EVAL_401 = _EVAL_3271 & 32'hf9f0707f;
  assign _EVAL_1639 = _EVAL_401 == 32'h1000202f;
  assign _EVAL_1029 = _EVAL_2892 | _EVAL_1639;
  assign _EVAL_4878 = _EVAL_3271 & 32'hdfffffff;
  assign _EVAL_1075 = _EVAL_4878 == 32'h10500073;
  assign _EVAL_652 = _EVAL_1029 | _EVAL_1075;
  assign _EVAL_2078 = _EVAL_3271 & 32'hf600607f;
  assign _EVAL_3407 = _EVAL_2078 == 32'h20000053;
  assign _EVAL_775 = _EVAL_652 | _EVAL_3407;
  assign _EVAL_5930 = _EVAL_3271 & 32'h7e00607f;
  assign _EVAL_4946 = _EVAL_5930 == 32'h20000053;
  assign _EVAL_2930 = _EVAL_775 | _EVAL_4946;
  assign _EVAL_4219 = _EVAL_3271 & 32'h7e00507f;
  assign _EVAL_5687 = _EVAL_4219 == 32'h20000053;
  assign _EVAL_3584 = _EVAL_2930 | _EVAL_5687;
  assign _EVAL_1098 = _EVAL_3271 == 32'h30200073;
  assign _EVAL_3398 = _EVAL_3584 | _EVAL_1098;
  assign _EVAL_1731 = _EVAL_5133 & 32'h64;
  assign _EVAL_3850 = _EVAL_1731 == 32'h0;
  assign _EVAL_2680 = _EVAL_5133 & 32'h50;
  assign _EVAL_4875 = _EVAL_2680 == 32'h10;
  assign _EVAL_4025 = _EVAL_3850 | _EVAL_4875;
  assign _EVAL_1671 = _EVAL_5133 & 32'h2024;
  assign _EVAL_955 = _EVAL_1671 == 32'h24;
  assign _EVAL_909 = _EVAL_4025 | _EVAL_955;
  assign _EVAL_4554 = _EVAL_2837 == 2'h2;
  assign _EVAL_4968 = _EVAL_3078[19:15];
  assign _EVAL_1682 = _EVAL_5813[19:15];
  assign _EVAL_374 = _EVAL_1947[19:15];
  assign _EVAL_2057 = _EVAL_1958 ? _EVAL_1682 : _EVAL_374;
  assign _EVAL_4536 = _EVAL_4554 ? _EVAL_4968 : _EVAL_2057;
  assign _EVAL_4681 = _EVAL_3952 == 32'h40;
  assign _EVAL_2723 = _EVAL_5979 | _EVAL_4681;
  assign _EVAL_4164 = _EVAL_3006 & 32'h1040;
  assign _EVAL_3297 = _EVAL_4164 == 32'h1040;
  assign _EVAL_4256 = _EVAL_2723 | _EVAL_3297;
  assign _EVAL_4183 = _EVAL_4268 & 32'h2040;
  assign _EVAL_579 = _EVAL_4183 == 32'h2040;
  assign _EVAL_5311 = _EVAL_3455[31:0];
  assign _EVAL_5114 = _EVAL_5311 & 32'h2000040;
  assign _EVAL_607 = _EVAL_5114 == 32'h0;
  assign _EVAL_3979 = _EVAL_5311 & 32'h60;
  assign _EVAL_4530 = _EVAL_3979 == 32'h0;
  assign _EVAL_4748 = _EVAL_607 | _EVAL_4530;
  assign _EVAL_1733 = _EVAL_5311 & 32'h50;
  assign _EVAL_1483 = _EVAL_1733 == 32'h0;
  assign _EVAL_1650 = _EVAL_4748 | _EVAL_1483;
  assign _EVAL_3166 = _EVAL_5311 & 32'h44;
  assign _EVAL_2422 = _EVAL_3166 == 32'h4;
  assign _EVAL_4571 = _EVAL_1650 | _EVAL_2422;
  assign _EVAL_1805 = _EVAL_5311 & 32'h62003010;
  assign _EVAL_3361 = _EVAL_1805 == 32'h60000010;
  assign _EVAL_2304 = _EVAL_4571 | _EVAL_3361;
  assign _EVAL_3292 = _EVAL_2039 & 32'h2000040;
  assign _EVAL_373 = _EVAL_3292 == 32'h0;
  assign _EVAL_614 = _EVAL_2039 & 32'h60;
  assign _EVAL_3423 = _EVAL_614 == 32'h0;
  assign _EVAL_4345 = _EVAL_373 | _EVAL_3423;
  assign _EVAL_2681 = _EVAL_2445 == 32'h0;
  assign _EVAL_3641 = _EVAL_4345 | _EVAL_2681;
  assign _EVAL_3956 = _EVAL_2039 & 32'h44;
  assign _EVAL_570 = _EVAL_3956 == 32'h4;
  assign _EVAL_4059 = _EVAL_3641 | _EVAL_570;
  assign _EVAL_2030 = _EVAL_2039 & 32'h62003010;
  assign _EVAL_5532 = _EVAL_2030 == 32'h60000010;
  assign _EVAL_1817 = _EVAL_4059 | _EVAL_5532;
  assign _EVAL_5926 = _EVAL_3573 == 2'h2;
  assign _EVAL_1074 = _EVAL_3573 == 2'h1;
  assign _EVAL_4939 = _EVAL_1242 & 32'h2000040;
  assign _EVAL_4862 = _EVAL_4939 == 32'h0;
  assign _EVAL_777 = _EVAL_1242 & 32'h60;
  assign _EVAL_1961 = _EVAL_777 == 32'h0;
  assign _EVAL_4493 = _EVAL_4862 | _EVAL_1961;
  assign _EVAL_3076 = _EVAL_1242 & 32'h50;
  assign _EVAL_3260 = _EVAL_3076 == 32'h0;
  assign _EVAL_2902 = _EVAL_4493 | _EVAL_3260;
  assign _EVAL_2648 = _EVAL_1242 & 32'h44;
  assign _EVAL_2589 = _EVAL_2648 == 32'h4;
  assign _EVAL_2835 = _EVAL_2902 | _EVAL_2589;
  assign _EVAL_2190 = _EVAL_1242 & 32'h62003010;
  assign _EVAL_5292 = _EVAL_2190 == 32'h60000010;
  assign _EVAL_1367 = _EVAL_2835 | _EVAL_5292;
  assign _EVAL_4718 = _EVAL_2164 & 32'h2000040;
  assign _EVAL_4869 = _EVAL_4718 == 32'h0;
  assign _EVAL_852 = _EVAL_2164 & 32'h60;
  assign _EVAL_5171 = _EVAL_852 == 32'h0;
  assign _EVAL_5346 = _EVAL_4869 | _EVAL_5171;
  assign _EVAL_2438 = _EVAL_2164 & 32'h50;
  assign _EVAL_2471 = _EVAL_2438 == 32'h0;
  assign _EVAL_2698 = _EVAL_5346 | _EVAL_2471;
  assign _EVAL_2128 = _EVAL_2164 & 32'h44;
  assign _EVAL_577 = _EVAL_2128 == 32'h4;
  assign _EVAL_1157 = _EVAL_2698 | _EVAL_577;
  assign _EVAL_5674 = _EVAL_2164 & 32'h62003010;
  assign _EVAL_5127 = _EVAL_5674 == 32'h60000010;
  assign _EVAL_2025 = _EVAL_1157 | _EVAL_5127;
  assign _EVAL_2187 = _EVAL_1074 ? _EVAL_1367 : _EVAL_2025;
  assign _EVAL_3973 = _EVAL_5926 ? _EVAL_1817 : _EVAL_2187;
  assign _EVAL_5811 = _EVAL_2970 ? _EVAL_1817 : _EVAL_3973;
  assign _EVAL_4448 = _EVAL_2970 ? _EVAL_2304 : _EVAL_5811;
  assign _EVAL_3558 = _EVAL_5276 ? 2'h0 : _EVAL_4231;
  assign _EVAL_1720 = {_EVAL_3558, 1'h0};
  assign _EVAL_960 = {{29'd0}, _EVAL_1720};
  assign _EVAL_2463 = _EVAL_3078 & 32'heff0707f;
  assign _EVAL_3111 = _EVAL_386 & 32'h7e00507f;
  assign _EVAL_1679 = _EVAL_4897 == 32'h2013;
  assign _EVAL_4085 = _EVAL_3239 | _EVAL_1679;
  assign _EVAL_2965 = _EVAL_3078 & 32'h1800707f;
  assign _EVAL_2924 = _EVAL_2965 == 32'h202f;
  assign _EVAL_3087 = _EVAL_4085 | _EVAL_2924;
  assign _EVAL_2950 = _EVAL_4897 == 32'h2073;
  assign _EVAL_6059 = _EVAL_3087 | _EVAL_2950;
  assign _EVAL_5006 = _EVAL_3078 & 32'hbe00705f;
  assign _EVAL_259 = _EVAL_5006 == 32'h5013;
  assign _EVAL_1880 = _EVAL_6059 | _EVAL_259;
  assign _EVAL_5151 = _EVAL_3078 & 32'he800707f;
  assign _EVAL_1745 = _EVAL_5151 == 32'h800202f;
  assign _EVAL_1051 = _EVAL_1880 | _EVAL_1745;
  assign _EVAL_5320 = _EVAL_3078 & 32'hf9f0707f;
  assign _EVAL_5043 = _EVAL_5320 == 32'h1000202f;
  assign _EVAL_315 = _EVAL_1051 | _EVAL_5043;
  assign _EVAL_3607 = _EVAL_3078 & 32'hdfffffff;
  assign _EVAL_3925 = _EVAL_3607 == 32'h10500073;
  assign _EVAL_2577 = _EVAL_315 | _EVAL_3925;
  assign _EVAL_3644 = _EVAL_3078 & 32'hf600607f;
  assign _EVAL_2364 = _EVAL_3644 == 32'h20000053;
  assign _EVAL_1009 = _EVAL_2577 | _EVAL_2364;
  assign _EVAL_2451 = _EVAL_3078 & 32'h7e00607f;
  assign _EVAL_192 = _EVAL_2451 == 32'h20000053;
  assign _EVAL_536 = _EVAL_1009 | _EVAL_192;
  assign _EVAL_3391 = _EVAL_3078 & 32'h7e00507f;
  assign _EVAL_4651 = _EVAL_3391 == 32'h20000053;
  assign _EVAL_4297 = _EVAL_536 | _EVAL_4651;
  assign _EVAL_1830 = _EVAL_3078 == 32'h30200073;
  assign _EVAL_348 = _EVAL_4297 | _EVAL_1830;
  assign _EVAL_4430 = _EVAL_3078 & 32'hfff0007f;
  assign _EVAL_3744 = _EVAL_4430 == 32'h58000053;
  assign _EVAL_1034 = _EVAL_348 | _EVAL_3744;
  assign _EVAL_5088 = _EVAL_3078 == 32'h7b200073;
  assign _EVAL_1130 = _EVAL_1034 | _EVAL_5088;
  assign _EVAL_1201 = _EVAL_3078 & 32'hefe0007f;
  assign _EVAL_5066 = _EVAL_1201 == 32'hc0000053;
  assign _EVAL_3669 = _EVAL_1130 | _EVAL_5066;
  assign _EVAL_643 = _EVAL_3078 & 32'hfff0607f;
  assign _EVAL_4349 = _EVAL_643 == 32'he0000053;
  assign _EVAL_2001 = _EVAL_3669 | _EVAL_4349;
  assign _EVAL_2353 = _EVAL_2463 == 32'he0000053;
  assign _EVAL_1058 = _EVAL_2001 | _EVAL_2353;
  assign _EVAL_2248 = _EVAL_3078 & 32'hffd07fff;
  assign _EVAL_5789 = _EVAL_2248 == 32'hfc000073;
  assign _EVAL_3581 = _EVAL_1058 | _EVAL_5789;
  assign _EVAL_1591 = _EVAL_5133 & 32'h3c;
  assign _EVAL_1722 = _EVAL_1591 == 32'h4;
  assign _EVAL_3927 = _EVAL_5133 & 32'h80000060;
  assign _EVAL_4217 = _EVAL_3927 == 32'h40;
  assign _EVAL_2938 = _EVAL_1722 | _EVAL_4217;
  assign _EVAL_2827 = _EVAL_5133 & 32'h70;
  assign _EVAL_5949 = _EVAL_2827 == 32'h40;
  assign _EVAL_1078 = _EVAL_2938 | _EVAL_5949;
  assign _EVAL_4806 = _EVAL_5133 & 32'h306f;
  assign _EVAL_6045 = _EVAL_4806 == 32'h3;
  assign _EVAL_1647 = _EVAL_4268[1:0];
  assign _EVAL_5690 = _EVAL_1647 == 2'h3;
  assign _EVAL_1585 = _EVAL_3006 & 32'h80000060;
  assign _EVAL_2784 = _EVAL_1585 == 32'h40;
  assign _EVAL_878 = _EVAL_3006 & 32'h10000060;
  assign _EVAL_2221 = _EVAL_878 == 32'h40;
  assign _EVAL_3692 = _EVAL_2784 | _EVAL_2221;
  assign _EVAL_5004 = _EVAL_3006 & 32'h70;
  assign _EVAL_3390 = _EVAL_5004 == 32'h40;
  assign _EVAL_1908 = _EVAL_3692 | _EVAL_3390;
  assign _EVAL_2378 = _EVAL_1647 == 2'h2;
  assign _EVAL_2901 = _EVAL_1647 == 2'h1;
  assign _EVAL_2367 = _EVAL_4882 & 32'h80000060;
  assign _EVAL_5771 = _EVAL_2367 == 32'h40;
  assign _EVAL_5020 = _EVAL_4882 & 32'h10000060;
  assign _EVAL_4213 = _EVAL_5020 == 32'h40;
  assign _EVAL_3922 = _EVAL_5771 | _EVAL_4213;
  assign _EVAL_5539 = _EVAL_4882 & 32'h70;
  assign _EVAL_2101 = _EVAL_5539 == 32'h40;
  assign _EVAL_559 = _EVAL_3922 | _EVAL_2101;
  assign _EVAL_3986 = _EVAL_5133 & 32'h10000060;
  assign _EVAL_4419 = _EVAL_3986 == 32'h40;
  assign _EVAL_172 = _EVAL_4217 | _EVAL_4419;
  assign _EVAL_5327 = _EVAL_172 | _EVAL_5949;
  assign _EVAL_1270 = _EVAL_2901 ? _EVAL_559 : _EVAL_5327;
  assign _EVAL_3232 = _EVAL_2378 ? _EVAL_1908 : _EVAL_1270;
  assign _EVAL_4190 = _EVAL_5690 ? _EVAL_1908 : _EVAL_3232;
  assign _EVAL_3473 = _EVAL_60;
  assign _EVAL_4923 = _EVAL_39;
  assign _EVAL_5322 = {_EVAL_3473,1'h0,1'h0,_EVAL_4923};
  assign _EVAL_5959 = _EVAL_5322 >> _EVAL_4188;
  assign _EVAL_1644 = _EVAL_5959[0];
  assign _EVAL_2801 = _EVAL_5718 & _EVAL_1644;
  assign _EVAL_5244 = _EVAL_90;
  assign _EVAL_4115 = _EVAL_2801 & _EVAL_5244;
  assign _EVAL_519 = _EVAL_4177[1];
  assign _EVAL_5620 = _EVAL_1854 < _EVAL_5201;
  assign _EVAL_1295 = 3'h6 < _EVAL_1773;
  assign _EVAL_1972 = _EVAL_4226 & _EVAL_1295;
  assign _EVAL_2419 = _EVAL_5620 | _EVAL_1972;
  assign _EVAL_5527 = _EVAL_2419 == _EVAL_383;
  assign _EVAL_5012 = 4'h1 | _EVAL_3550;
  assign _EVAL_5541 = _EVAL_5012 == _EVAL_4784;
  assign _EVAL_2368 = _EVAL_4226 & _EVAL_5541;
  assign _EVAL_4079 = _EVAL_519 ? _EVAL_5527 : _EVAL_2368;
  assign _EVAL_3848 = _EVAL_4115 & _EVAL_4079;
  assign _EVAL_6064 = _EVAL_574 | _EVAL_1558;
  assign _EVAL_3955 = _EVAL_3848 & _EVAL_6064;
  assign _EVAL_2357 = _EVAL_48;
  assign _EVAL_527 = _EVAL_144;
  assign _EVAL_1086 = _EVAL_2110 & _EVAL_1928;
  assign _EVAL_2198 = 3'h6 < _EVAL_5107;
  assign _EVAL_3829 = _EVAL_5549 & _EVAL_2198;
  assign _EVAL_1595 = _EVAL_5844 | _EVAL_3829;
  assign _EVAL_1566 = _EVAL_1595 == _EVAL_3257;
  assign _EVAL_5606 = 4'h1 | _EVAL_3251;
  assign _EVAL_1022 = _EVAL_5606 == _EVAL_920;
  assign _EVAL_2021 = _EVAL_5549 & _EVAL_1022;
  assign _EVAL_2256 = _EVAL_5680 ? _EVAL_1566 : _EVAL_2021;
  assign _EVAL_3123 = _EVAL_977 & _EVAL_2256;
  assign _EVAL_5174 = _EVAL_5875 | _EVAL_3123;
  assign _EVAL_1660 = _EVAL_1086 & _EVAL_5174;
  assign _EVAL_3758 = _EVAL_49;
  assign _EVAL_5472 = _EVAL_5875 & _EVAL_3123;
  assign _EVAL_1048 = _EVAL_79;
  assign _EVAL_2053 = _EVAL_5472 ? _EVAL_1048 : 1'h0;
  assign _EVAL_2348 = _EVAL_1660 ? _EVAL_3758 : _EVAL_2053;
  assign _EVAL_5853 = _EVAL_1365 ? _EVAL_527 : _EVAL_2348;
  assign _EVAL_2383 = _EVAL_3955 ? _EVAL_2357 : _EVAL_5853;
  assign _EVAL_2374 = 3'h4 < _EVAL_1773;
  assign _EVAL_3377 = _EVAL_4226 & _EVAL_2374;
  assign _EVAL_991 = _EVAL_5620 | _EVAL_3377;
  assign _EVAL_5086 = _EVAL_991 == _EVAL_383;
  assign _EVAL_1278 = _EVAL_519 ? _EVAL_5086 : _EVAL_2968;
  assign _EVAL_3243 = _EVAL_4115 & _EVAL_1278;
  assign _EVAL_1555 = 3'h4 < _EVAL_3401;
  assign _EVAL_606 = _EVAL_584 & _EVAL_1555;
  assign _EVAL_2713 = _EVAL_1310 | _EVAL_606;
  assign _EVAL_2615 = _EVAL_2713 == _EVAL_1969;
  assign _EVAL_1602 = 4'h3 | _EVAL_4534;
  assign _EVAL_660 = _EVAL_1602 == _EVAL_3975;
  assign _EVAL_3832 = _EVAL_584 & _EVAL_660;
  assign _EVAL_5489 = _EVAL_4291 ? _EVAL_2615 : _EVAL_3832;
  assign _EVAL_5900 = _EVAL_5039 & _EVAL_5489;
  assign _EVAL_4138 = _EVAL_574 | _EVAL_5900;
  assign _EVAL_2917 = _EVAL_3243 & _EVAL_4138;
  assign _EVAL_704 = _EVAL_574 & _EVAL_5900;
  assign _EVAL_1777 = _EVAL_2110 | _EVAL_4867;
  assign _EVAL_409 = _EVAL_704 & _EVAL_1777;
  assign _EVAL_5454 = _EVAL_5875 & _EVAL_1006;
  assign _EVAL_4132 = _EVAL_5454 ? _EVAL_1048 : 1'h0;
  assign _EVAL_4295 = _EVAL_6001 ? _EVAL_3758 : _EVAL_4132;
  assign _EVAL_4428 = _EVAL_409 ? _EVAL_527 : _EVAL_4295;
  assign _EVAL_4168 = _EVAL_2917 ? _EVAL_2357 : _EVAL_4428;
  assign _EVAL_2223 = 3'h2 < _EVAL_1773;
  assign _EVAL_2945 = _EVAL_4226 & _EVAL_2223;
  assign _EVAL_1609 = _EVAL_5620 | _EVAL_2945;
  assign _EVAL_5937 = _EVAL_1609 == _EVAL_383;
  assign _EVAL_3364 = 4'h5 | _EVAL_3550;
  assign _EVAL_378 = _EVAL_3364 == _EVAL_4784;
  assign _EVAL_3437 = _EVAL_4226 & _EVAL_378;
  assign _EVAL_2707 = _EVAL_519 ? _EVAL_5937 : _EVAL_3437;
  assign _EVAL_3887 = _EVAL_4115 & _EVAL_2707;
  assign _EVAL_4484 = 3'h2 < _EVAL_3401;
  assign _EVAL_4389 = _EVAL_584 & _EVAL_4484;
  assign _EVAL_2062 = _EVAL_1310 | _EVAL_4389;
  assign _EVAL_5332 = _EVAL_2062 == _EVAL_1969;
  assign _EVAL_676 = 4'h5 | _EVAL_4534;
  assign _EVAL_5676 = _EVAL_676 == _EVAL_3975;
  assign _EVAL_3358 = _EVAL_584 & _EVAL_5676;
  assign _EVAL_1380 = _EVAL_4291 ? _EVAL_5332 : _EVAL_3358;
  assign _EVAL_202 = _EVAL_5039 & _EVAL_1380;
  assign _EVAL_6029 = _EVAL_574 | _EVAL_202;
  assign _EVAL_5373 = _EVAL_3887 & _EVAL_6029;
  assign _EVAL_2418 = _EVAL_574 & _EVAL_202;
  assign _EVAL_4959 = _EVAL_2127 & _EVAL_3370;
  assign _EVAL_1523 = _EVAL_4204 | _EVAL_4959;
  assign _EVAL_2498 = _EVAL_1523 == _EVAL_379;
  assign _EVAL_1629 = _EVAL_2127 & _EVAL_1323;
  assign _EVAL_3001 = _EVAL_4914 ? _EVAL_2498 : _EVAL_1629;
  assign _EVAL_1628 = _EVAL_5393 & _EVAL_3001;
  assign _EVAL_3658 = _EVAL_2110 | _EVAL_1628;
  assign _EVAL_3870 = _EVAL_2418 & _EVAL_3658;
  assign _EVAL_3444 = _EVAL_2110 & _EVAL_1628;
  assign _EVAL_680 = _EVAL_5549 & _EVAL_2371;
  assign _EVAL_2337 = _EVAL_5844 | _EVAL_680;
  assign _EVAL_859 = _EVAL_2337 == _EVAL_3257;
  assign _EVAL_5943 = _EVAL_5549 & _EVAL_2486;
  assign _EVAL_4043 = _EVAL_5680 ? _EVAL_859 : _EVAL_5943;
  assign _EVAL_5976 = _EVAL_977 & _EVAL_4043;
  assign _EVAL_6052 = _EVAL_5875 | _EVAL_5976;
  assign _EVAL_5135 = _EVAL_3444 & _EVAL_6052;
  assign _EVAL_5024 = _EVAL_5875 & _EVAL_5976;
  assign _EVAL_3967 = _EVAL_5024 ? _EVAL_1048 : 1'h0;
  assign _EVAL_803 = _EVAL_5135 ? _EVAL_3758 : _EVAL_3967;
  assign _EVAL_2105 = _EVAL_3870 ? _EVAL_527 : _EVAL_803;
  assign _EVAL_4401 = _EVAL_5373 ? _EVAL_2357 : _EVAL_2105;
  assign _EVAL_1385 = 3'h0 < _EVAL_1773;
  assign _EVAL_5430 = _EVAL_4226 & _EVAL_1385;
  assign _EVAL_5130 = _EVAL_5620 | _EVAL_5430;
  assign _EVAL_357 = _EVAL_5130 == _EVAL_383;
  assign _EVAL_4731 = 4'h7 | _EVAL_3550;
  assign _EVAL_2939 = _EVAL_4731 == _EVAL_4784;
  assign _EVAL_618 = _EVAL_4226 & _EVAL_2939;
  assign _EVAL_2732 = _EVAL_519 ? _EVAL_357 : _EVAL_618;
  assign _EVAL_2429 = _EVAL_4115 & _EVAL_2732;
  assign _EVAL_3876 = 3'h0 < _EVAL_3401;
  assign _EVAL_5725 = _EVAL_584 & _EVAL_3876;
  assign _EVAL_5423 = _EVAL_1310 | _EVAL_5725;
  assign _EVAL_4189 = _EVAL_5423 == _EVAL_1969;
  assign _EVAL_1462 = 4'h7 | _EVAL_4534;
  assign _EVAL_3445 = _EVAL_1462 == _EVAL_3975;
  assign _EVAL_2238 = _EVAL_584 & _EVAL_3445;
  assign _EVAL_4754 = _EVAL_4291 ? _EVAL_4189 : _EVAL_2238;
  assign _EVAL_3980 = _EVAL_5039 & _EVAL_4754;
  assign _EVAL_2949 = _EVAL_574 | _EVAL_3980;
  assign _EVAL_4716 = _EVAL_2429 & _EVAL_2949;
  assign _EVAL_4218 = _EVAL_574 & _EVAL_3980;
  assign _EVAL_1973 = _EVAL_2127 & _EVAL_2491;
  assign _EVAL_2216 = _EVAL_4204 | _EVAL_1973;
  assign _EVAL_3737 = _EVAL_2216 == _EVAL_379;
  assign _EVAL_3940 = _EVAL_2127 & _EVAL_3143;
  assign _EVAL_1478 = _EVAL_4914 ? _EVAL_3737 : _EVAL_3940;
  assign _EVAL_1422 = _EVAL_5393 & _EVAL_1478;
  assign _EVAL_4818 = _EVAL_2110 | _EVAL_1422;
  assign _EVAL_3070 = _EVAL_4218 & _EVAL_4818;
  assign _EVAL_2070 = _EVAL_2110 & _EVAL_1422;
  assign _EVAL_4848 = 3'h0 < _EVAL_5107;
  assign _EVAL_3141 = _EVAL_5549 & _EVAL_4848;
  assign _EVAL_3321 = _EVAL_5844 | _EVAL_3141;
  assign _EVAL_6090 = _EVAL_3321 == _EVAL_3257;
  assign _EVAL_5516 = 4'h7 | _EVAL_3251;
  assign _EVAL_2754 = _EVAL_5516 == _EVAL_920;
  assign _EVAL_1357 = _EVAL_5549 & _EVAL_2754;
  assign _EVAL_4826 = _EVAL_5680 ? _EVAL_6090 : _EVAL_1357;
  assign _EVAL_3337 = _EVAL_977 & _EVAL_4826;
  assign _EVAL_5388 = _EVAL_5875 | _EVAL_3337;
  assign _EVAL_1826 = _EVAL_2070 & _EVAL_5388;
  assign _EVAL_726 = _EVAL_5875 & _EVAL_3337;
  assign _EVAL_1597 = _EVAL_726 ? _EVAL_1048 : 1'h0;
  assign _EVAL_3272 = _EVAL_1826 ? _EVAL_3758 : _EVAL_1597;
  assign _EVAL_2706 = _EVAL_3070 ? _EVAL_527 : _EVAL_3272;
  assign _EVAL_2225 = _EVAL_4716 ? _EVAL_2357 : _EVAL_2706;
  assign _EVAL_1183 = {_EVAL_2383,_EVAL_4168,_EVAL_4401,_EVAL_2225};
  assign _EVAL_2389 = _EVAL_2666[1:0];
  assign _EVAL_1069 = _EVAL_2389 == 2'h3;
  assign _EVAL_4441 = 1'h0 < _EVAL_5690;
  assign _EVAL_1010 = _EVAL_2142 & _EVAL_4441;
  assign _EVAL_798 = _EVAL_1010 ? 1'h0 : 1'h1;
  assign _EVAL_3905 = _EVAL_1069 ? 1'h0 : _EVAL_798;
  assign _EVAL_5880 = _EVAL_5994 | _EVAL_5276;
  assign _EVAL_5422 = _EVAL_5880 | _EVAL_3052;
  assign _EVAL_4481 = _EVAL_5422 | _EVAL_2142;
  assign _EVAL_867 = _EVAL_4481 == 1'h0;
  assign _EVAL_1505 = _EVAL_3905 & _EVAL_867;
  assign _EVAL_5579 = _EVAL_1505 == 1'h0;
  assign _EVAL_5985 = _EVAL_3905 & _EVAL_5579;
  assign _EVAL_3676 = _EVAL_5422 == 1'h0;
  assign _EVAL_1613 = _EVAL_2142 & _EVAL_3676;
  assign _EVAL_258 = _EVAL_1613 == 1'h0;
  assign _EVAL_5337 = _EVAL_2142 & _EVAL_258;
  assign _EVAL_5777 = _EVAL_5880 == 1'h0;
  assign _EVAL_4994 = _EVAL_3052 & _EVAL_5777;
  assign _EVAL_3529 = _EVAL_4994 == 1'h0;
  assign _EVAL_1930 = _EVAL_3052 & _EVAL_3529;
  assign _EVAL_3904 = _EVAL_5994 == 1'h0;
  assign _EVAL_4772 = _EVAL_5276 & _EVAL_3904;
  assign _EVAL_6031 = _EVAL_4772 == 1'h0;
  assign _EVAL_1226 = _EVAL_5276 & _EVAL_6031;
  assign _EVAL_3219 = {_EVAL_5985,_EVAL_5337,_EVAL_1930,_EVAL_1226};
  assign _EVAL_1217 = _EVAL_3219[0];
  assign _EVAL_2765 = _EVAL_3219[1];
  assign _EVAL_1699 = _EVAL_3219[2];
  assign _EVAL_2002 = _EVAL_3219[3];
  assign _EVAL_5251 = _EVAL_2002 ? 4'h8 : 4'h0;
  assign _EVAL_907 = _EVAL_1699 ? 4'h4 : _EVAL_5251;
  assign _EVAL_2058 = _EVAL_2765 ? 4'h2 : _EVAL_907;
  assign _EVAL_4445 = _EVAL_1217 ? 4'h1 : _EVAL_2058;
  assign _EVAL_3266 = _EVAL_1183 & _EVAL_4445;
  assign _EVAL_232 = _EVAL_4882 & 32'h64;
  assign _EVAL_3554 = _EVAL_232 == 32'h0;
  assign _EVAL_1757 = _EVAL_4882 & 32'h50;
  assign _EVAL_360 = _EVAL_1757 == 32'h10;
  assign _EVAL_2867 = _EVAL_3554 | _EVAL_360;
  assign _EVAL_1291 = _EVAL_5311 & 32'h306f;
  assign _EVAL_4961 = ~ _EVAL_136;
  assign _EVAL_454 = _EVAL_4961 | 32'h7;
  assign _EVAL_532 = ~ _EVAL_454;
  assign _EVAL_4856 = _EVAL_3271 & 32'h2024;
  assign _EVAL_3893 = _EVAL_5311 & 32'h40000040;
  assign _EVAL_641 = _EVAL_3893 == 32'h40;
  assign _EVAL_2303 = _EVAL_5967 & _EVAL_2198;
  assign _EVAL_3103 = _EVAL_2293 | _EVAL_2303;
  assign _EVAL_3107 = _EVAL_3103 == _EVAL_3257;
  assign _EVAL_914 = _EVAL_5967 & _EVAL_1022;
  assign _EVAL_5770 = _EVAL_5680 ? _EVAL_3107 : _EVAL_914;
  assign _EVAL_432 = _EVAL_4063 & _EVAL_5770;
  assign _EVAL_5748 = _EVAL_5875 & _EVAL_432;
  assign _EVAL_3728 = _EVAL_6086 & _EVAL_5770;
  assign _EVAL_6011 = _EVAL_5875 & _EVAL_3728;
  assign _EVAL_391 = _EVAL_5748 ? 1'h1 : _EVAL_6011;
  assign _EVAL_740 = _EVAL_1362 & 32'hfff0007f;
  assign _EVAL_4622 = _EVAL_4882 & 32'h2000040;
  assign _EVAL_6009 = _EVAL_4622 == 32'h0;
  assign _EVAL_3996 = _EVAL_5813 & 32'h2000040;
  assign _EVAL_1191 = _EVAL_3996 == 32'h0;
  assign _EVAL_5801 = _EVAL_5813 & 32'h60;
  assign _EVAL_4737 = _EVAL_5801 == 32'h0;
  assign _EVAL_3387 = _EVAL_1191 | _EVAL_4737;
  assign _EVAL_3680 = _EVAL_5813 & 32'h50;
  assign _EVAL_4232 = _EVAL_3680 == 32'h0;
  assign _EVAL_1272 = _EVAL_3387 | _EVAL_4232;
  assign _EVAL_3618 = _EVAL_4702 & 32'h3c;
  assign _EVAL_1764 = _EVAL_3618 == 32'h4;
  assign _EVAL_4343 = _EVAL_4702 & 32'h80000060;
  assign _EVAL_1709 = _EVAL_4343 == 32'h40;
  assign _EVAL_3575 = _EVAL_1764 | _EVAL_1709;
  assign _EVAL_4930 = _EVAL_4702 & 32'h70;
  assign _EVAL_4636 = _EVAL_4930 == 32'h40;
  assign _EVAL_467 = _EVAL_3575 | _EVAL_4636;
  assign _EVAL_5820 = _EVAL_5133 & 32'h62003010;
  assign _EVAL_4227 = _EVAL_1242 & 32'heff0707f;
  assign _EVAL_362 = _EVAL_4268 & 32'h64;
  assign _EVAL_4434 = _EVAL_362 == 32'h0;
  assign _EVAL_2696 = _EVAL_4268 & 32'h50;
  assign _EVAL_426 = _EVAL_2696 == 32'h10;
  assign _EVAL_1845 = _EVAL_4434 | _EVAL_426;
  assign _EVAL_5778 = _EVAL_4268 & 32'h2024;
  assign _EVAL_3899 = _EVAL_5778 == 32'h24;
  assign _EVAL_968 = _EVAL_1845 | _EVAL_3899;
  assign _EVAL_4490 = _EVAL_2039[11:7];
  assign _EVAL_1621 = _EVAL_1242[11:7];
  assign _EVAL_3256 = _EVAL_2164[11:7];
  assign _EVAL_5155 = _EVAL_1074 ? _EVAL_1621 : _EVAL_3256;
  assign _EVAL_329 = _EVAL_5926 ? _EVAL_4490 : _EVAL_5155;
  assign _EVAL_880 = _EVAL_2970 ? _EVAL_4490 : _EVAL_329;
  assign _EVAL_2144 = _EVAL_4743 & 32'h70;
  assign _EVAL_1433 = _EVAL_2144 == 32'h40;
  assign _EVAL_4790 = _EVAL_386 & 32'h70;
  assign _EVAL_4271 = _EVAL_4790 == 32'h40;
  assign _EVAL_4136 = _EVAL_5952 ? _EVAL_1433 : _EVAL_4271;
  assign _EVAL_1361 = _EVAL_2648 == 32'h0;
  assign _EVAL_3654 = _EVAL_1242 & 32'h4024;
  assign _EVAL_2020 = _EVAL_3654 == 32'h20;
  assign _EVAL_3755 = _EVAL_1361 | _EVAL_2020;
  assign _EVAL_5191 = _EVAL_1242 & 32'h38;
  assign _EVAL_1781 = _EVAL_5191 == 32'h20;
  assign _EVAL_1975 = _EVAL_3755 | _EVAL_1781;
  assign _EVAL_2341 = _EVAL_5386[8:7];
  assign _EVAL_2439 = _EVAL_5386[12:9];
  assign _EVAL_1666 = {_EVAL_2341,_EVAL_2439,2'h0};
  assign _EVAL_462 = _EVAL_1666[7:5];
  assign _EVAL_772 = _EVAL_1666[4:0];
  assign _EVAL_4956 = {_EVAL_462,_EVAL_2272,5'h2,3'h2,_EVAL_772,7'h27};
  assign _EVAL_3193 = {_EVAL_462,_EVAL_2272,5'h2,3'h2,_EVAL_772,7'h23};
  assign _EVAL_1968 = {_EVAL_5546,_EVAL_688,3'h0};
  assign _EVAL_5604 = _EVAL_1968[8:5];
  assign _EVAL_3146 = _EVAL_1968[4:0];
  assign _EVAL_1926 = {_EVAL_5604,_EVAL_2272,5'h2,3'h3,_EVAL_3146,7'h27};
  assign _EVAL_3798 = _EVAL_2272 != 5'h0;
  assign _EVAL_2603 = {_EVAL_2272,_EVAL_4374,3'h0,_EVAL_4374,7'h33};
  assign _EVAL_5207 = _EVAL_4374 != 5'h0;
  assign _EVAL_4020 = {_EVAL_2272,_EVAL_4374,3'h0,12'he7};
  assign _EVAL_3416 = {_EVAL_2272,_EVAL_4374,3'h0,12'h67};
  assign _EVAL_1109 = _EVAL_3416[24:7];
  assign _EVAL_2325 = {_EVAL_1109,7'h73};
  assign _EVAL_4404 = _EVAL_2325 | 25'h100000;
  assign _EVAL_3939 = _EVAL_5207 ? _EVAL_4020 : _EVAL_4404;
  assign _EVAL_5815 = _EVAL_3798 ? _EVAL_2603 : _EVAL_3939;
  assign _EVAL_455 = {_EVAL_2272,5'h0,3'h4,_EVAL_4374,7'h33};
  assign _EVAL_3329 = _EVAL_3798 ? _EVAL_455 : _EVAL_3416;
  assign _EVAL_3768 = _EVAL_4111 ? _EVAL_5815 : _EVAL_3329;
  assign _EVAL_5183 = _EVAL_5386[3:2];
  assign _EVAL_1842 = _EVAL_5386[6:4];
  assign _EVAL_2215 = {_EVAL_5183,_EVAL_4111,_EVAL_1842,2'h0,5'h2,3'h2,_EVAL_4374,7'h7};
  assign _EVAL_3291 = {_EVAL_5183,_EVAL_4111,_EVAL_1842,2'h0,5'h2,3'h2,_EVAL_4374,7'h3};
  assign _EVAL_5363 = {_EVAL_1418,_EVAL_4111,_EVAL_5289,3'h0,5'h2,3'h3,_EVAL_4374,7'h7};
  assign _EVAL_4807 = {_EVAL_4111,_EVAL_2272,_EVAL_4374,3'h1,_EVAL_4374,7'h13};
  assign _EVAL_5785 = _EVAL_2175 ? _EVAL_5363 : {{3'd0}, _EVAL_4807};
  assign _EVAL_592 = _EVAL_179 ? {{1'd0}, _EVAL_3291} : _EVAL_5785;
  assign _EVAL_5203 = _EVAL_268 ? {{1'd0}, _EVAL_2215} : _EVAL_592;
  assign _EVAL_1663 = _EVAL_3261 ? {{4'd0}, _EVAL_3768} : _EVAL_5203;
  assign _EVAL_430 = _EVAL_3493 ? _EVAL_1926 : _EVAL_1663;
  assign _EVAL_2497 = _EVAL_4185 ? {{1'd0}, _EVAL_3193} : _EVAL_430;
  assign _EVAL_2440 = _EVAL_4999 ? {{1'd0}, _EVAL_4956} : _EVAL_2497;
  assign _EVAL_888 = {3'h0,_EVAL_2440};
  assign _EVAL_2898 = _EVAL_5311 & 32'h5f;
  assign _EVAL_6120 = _EVAL_2898 == 32'h17;
  assign _EVAL_5634 = {_EVAL_3620,_EVAL_3553};
  assign _EVAL_4843 = _EVAL_5634 != 12'h0;
  assign _EVAL_5966 = _EVAL_1743 ? _EVAL_4843 : 1'h1;
  assign _EVAL_526 = _EVAL_77;
  assign _EVAL_1986 = _EVAL_4492 & _EVAL_526;
  assign _EVAL_3164 = _EVAL_1242 & 32'h80000010;
  assign _EVAL_5713 = _EVAL_3164 == 32'h10;
  assign _EVAL_5504 = _EVAL_3076 == 32'h10;
  assign _EVAL_4711 = _EVAL_5713 | _EVAL_5504;
  assign _EVAL_3160 = _EVAL_1947 & 32'hffd07fff;
  assign _EVAL_1618 = _EVAL_4702 & 32'h2024;
  assign _EVAL_5724 = _EVAL_1618 == 32'h24;
  assign _EVAL_4982 = _EVAL_5813 & 32'h207f;
  assign _EVAL_1355 = _EVAL_4982 == 32'h3;
  assign _EVAL_1368 = _EVAL_5813 & 32'h607f;
  assign _EVAL_4987 = _EVAL_1368 == 32'hf;
  assign _EVAL_3046 = _EVAL_1355 | _EVAL_4987;
  assign _EVAL_1832 = _EVAL_5813 & 32'h5f;
  assign _EVAL_3545 = _EVAL_1832 == 32'h17;
  assign _EVAL_6105 = _EVAL_3046 | _EVAL_3545;
  assign _EVAL_5364 = _EVAL_5813 & 32'hfc00007f;
  assign _EVAL_5715 = _EVAL_5364 == 32'h33;
  assign _EVAL_2709 = _EVAL_6105 | _EVAL_5715;
  assign _EVAL_2690 = _EVAL_5813 & 32'hbe00707f;
  assign _EVAL_2063 = _EVAL_2690 == 32'h33;
  assign _EVAL_1638 = _EVAL_2709 | _EVAL_2063;
  assign _EVAL_4864 = _EVAL_5813 & 32'h6000073;
  assign _EVAL_1646 = _EVAL_4864 == 32'h43;
  assign _EVAL_1944 = _EVAL_1638 | _EVAL_1646;
  assign _EVAL_6022 = _EVAL_5813 & 32'he600007f;
  assign _EVAL_1864 = _EVAL_6022 == 32'h53;
  assign _EVAL_4810 = _EVAL_1944 | _EVAL_1864;
  assign _EVAL_3794 = _EVAL_5813 & 32'h707b;
  assign _EVAL_3645 = _EVAL_3794 == 32'h63;
  assign _EVAL_1651 = _EVAL_4810 | _EVAL_3645;
  assign _EVAL_3869 = _EVAL_5813 & 32'h7f;
  assign _EVAL_1853 = _EVAL_3869 == 32'h6f;
  assign _EVAL_1937 = _EVAL_1651 | _EVAL_1853;
  assign _EVAL_5219 = _EVAL_5813 & 32'hffefffff;
  assign _EVAL_1407 = _EVAL_5219 == 32'h73;
  assign _EVAL_5119 = _EVAL_1937 | _EVAL_1407;
  assign _EVAL_2029 = _EVAL_5813 & 32'hfe00305f;
  assign _EVAL_5661 = _EVAL_2029 == 32'h1013;
  assign _EVAL_5089 = _EVAL_5119 | _EVAL_5661;
  assign _EVAL_996 = _EVAL_5813 & 32'h705b;
  assign _EVAL_2936 = _EVAL_996 == 32'h2003;
  assign _EVAL_2048 = _EVAL_5089 | _EVAL_2936;
  assign _EVAL_5947 = _EVAL_4982 == 32'h2013;
  assign _EVAL_4237 = _EVAL_2048 | _EVAL_5947;
  assign _EVAL_5054 = _EVAL_5813 & 32'h1800707f;
  assign _EVAL_5253 = _EVAL_5054 == 32'h202f;
  assign _EVAL_2307 = _EVAL_4237 | _EVAL_5253;
  assign _EVAL_4658 = _EVAL_4982 == 32'h2073;
  assign _EVAL_1102 = _EVAL_2307 | _EVAL_4658;
  assign _EVAL_2456 = _EVAL_5813 & 32'hbe00705f;
  assign _EVAL_3439 = _EVAL_2456 == 32'h5013;
  assign _EVAL_2299 = _EVAL_1102 | _EVAL_3439;
  assign _EVAL_3954 = _EVAL_5813 & 32'he800707f;
  assign _EVAL_2780 = _EVAL_3954 == 32'h800202f;
  assign _EVAL_4823 = _EVAL_2299 | _EVAL_2780;
  assign _EVAL_5287 = _EVAL_5813 & 32'hf9f0707f;
  assign _EVAL_5596 = _EVAL_5287 == 32'h1000202f;
  assign _EVAL_887 = _EVAL_4823 | _EVAL_5596;
  assign _EVAL_1604 = _EVAL_5813 & 32'hdfffffff;
  assign _EVAL_5095 = _EVAL_1604 == 32'h10500073;
  assign _EVAL_5483 = _EVAL_887 | _EVAL_5095;
  assign _EVAL_3180 = _EVAL_5813 & 32'hf600607f;
  assign _EVAL_2016 = _EVAL_3180 == 32'h20000053;
  assign _EVAL_5231 = _EVAL_5483 | _EVAL_2016;
  assign _EVAL_2322 = _EVAL_5813 & 32'h7e00607f;
  assign _EVAL_5398 = _EVAL_2322 == 32'h20000053;
  assign _EVAL_4351 = _EVAL_5231 | _EVAL_5398;
  assign _EVAL_1956 = _EVAL_5813 & 32'h7e00507f;
  assign _EVAL_4665 = _EVAL_1956 == 32'h20000053;
  assign _EVAL_4663 = _EVAL_4351 | _EVAL_4665;
  assign _EVAL_601 = _EVAL_5813 == 32'h30200073;
  assign _EVAL_3119 = _EVAL_4663 | _EVAL_601;
  assign _EVAL_2627 = _EVAL_5813 & 32'hfff0007f;
  assign _EVAL_3020 = _EVAL_2627 == 32'h58000053;
  assign _EVAL_987 = _EVAL_3119 | _EVAL_3020;
  assign _EVAL_1045 = _EVAL_5813 == 32'h7b200073;
  assign _EVAL_5519 = _EVAL_987 | _EVAL_1045;
  assign _EVAL_3278 = _EVAL_5813 & 32'hefe0007f;
  assign _EVAL_1510 = _EVAL_3278 == 32'hc0000053;
  assign _EVAL_1239 = _EVAL_5519 | _EVAL_1510;
  assign _EVAL_4496 = _EVAL_4268 & 32'hbe00705f;
  assign _EVAL_2208 = _EVAL_4496 == 32'h5013;
  assign _EVAL_4931 = _EVAL_654[12:5];
  assign _EVAL_2558 = _EVAL_4931 != 8'h0;
  assign _EVAL_2979 = _EVAL_3016 ? 1'h1 : _EVAL_2558;
  assign _EVAL_4388 = _EVAL_5989 ? 1'h1 : _EVAL_2979;
  assign _EVAL_2179 = _EVAL_761 ? 1'h1 : _EVAL_4388;
  assign _EVAL_5305 = _EVAL_4440 ? 1'h1 : _EVAL_2179;
  assign _EVAL_2770 = _EVAL_1378 ? 1'h1 : _EVAL_5305;
  assign _EVAL_4950 = _EVAL_1978 & 32'h28;
  assign _EVAL_3379 = _EVAL_4950 == 32'h28;
  assign _EVAL_5665 = _EVAL_1947 & 32'h2010;
  assign _EVAL_2866 = _EVAL_5665 == 32'h2000;
  assign _EVAL_3255 = _EVAL_4268 & 32'hfe00305f;
  assign _EVAL_3985 = _EVAL_1947 & 32'hf9f0707f;
  assign _EVAL_389 = _EVAL_1362 & 32'h1800707f;
  assign _EVAL_3298 = _EVAL_4882 & 32'h207f;
  assign _EVAL_1702 = _EVAL_3298 == 32'h3;
  assign _EVAL_4821 = _EVAL_888 & 32'h64;
  assign _EVAL_1680 = _EVAL_4821 == 32'h20;
  assign _EVAL_6070 = _EVAL_888 & 32'h34;
  assign _EVAL_942 = _EVAL_6070 == 32'h20;
  assign _EVAL_1013 = _EVAL_1680 | _EVAL_942;
  assign _EVAL_1578 = _EVAL_5989 ? _EVAL_1360 : 1'h1;
  assign _EVAL_5323 = _EVAL_1978 & 32'h2040;
  assign _EVAL_3447 = _EVAL_5323 == 32'h2040;
  assign _EVAL_5575 = _EVAL_132;
  assign _EVAL_1458 = _EVAL_4702 & 32'h50;
  assign _EVAL_1974 = _EVAL_5311 & 32'h10000060;
  assign _EVAL_617 = _EVAL_1974 == 32'h10000040;
  assign _EVAL_621 = _EVAL_1947 & 32'h64;
  assign _EVAL_2449 = _EVAL_621 == 32'h0;
  assign _EVAL_1550 = _EVAL_1947 & 32'h50;
  assign _EVAL_4779 = _EVAL_1550 == 32'h10;
  assign _EVAL_3713 = _EVAL_2449 | _EVAL_4779;
  assign _EVAL_4301 = _EVAL_1947 & 32'h2040;
  assign _EVAL_1015 = _EVAL_3758 == 1'h0;
  assign _EVAL_5787 = _EVAL_1048 == 1'h0;
  assign _EVAL_3843 = _EVAL_5472 ? _EVAL_5787 : 1'h0;
  assign _EVAL_5164 = _EVAL_1660 ? _EVAL_1015 : _EVAL_3843;
  assign _EVAL_5854 = _EVAL_5386[31:0];
  assign _EVAL_6084 = _EVAL_5854 & 32'h64;
  assign _EVAL_2941 = _EVAL_6084 == 32'h20;
  assign _EVAL_1642 = _EVAL_5854 & 32'h34;
  assign _EVAL_4567 = _EVAL_1642 == 32'h20;
  assign _EVAL_2052 = _EVAL_2941 | _EVAL_4567;
  assign _EVAL_1804 = _EVAL_5854 & 32'h2048;
  assign _EVAL_6080 = _EVAL_1804 == 32'h2008;
  assign _EVAL_1829 = _EVAL_2052 | _EVAL_6080;
  assign _EVAL_1259 = _EVAL_2039 & 32'h64;
  assign _EVAL_787 = _EVAL_1259 == 32'h20;
  assign _EVAL_2678 = _EVAL_2039 & 32'h34;
  assign _EVAL_3715 = _EVAL_2678 == 32'h20;
  assign _EVAL_609 = _EVAL_787 | _EVAL_3715;
  assign _EVAL_2090 = _EVAL_2039 & 32'h2048;
  assign _EVAL_1197 = _EVAL_2090 == 32'h2008;
  assign _EVAL_1203 = _EVAL_609 | _EVAL_1197;
  assign _EVAL_540 = _EVAL_2039 & 32'h4003044;
  assign _EVAL_4403 = _EVAL_540 == 32'h4000040;
  assign _EVAL_3890 = _EVAL_1203 | _EVAL_4403;
  assign _EVAL_5072 = _EVAL_1362 & 32'h30;
  assign _EVAL_5400 = _EVAL_888 & 32'h207f;
  assign _EVAL_5224 = _EVAL_5400 == 32'h3;
  assign _EVAL_2130 = _EVAL_888 & 32'h607f;
  assign _EVAL_1448 = _EVAL_2130 == 32'hf;
  assign _EVAL_5899 = _EVAL_5224 | _EVAL_1448;
  assign _EVAL_3215 = _EVAL_1947[11:7];
  assign _EVAL_736 = _EVAL_5094[1:0];
  assign _EVAL_3722 = _EVAL_736 == 2'h3;
  assign _EVAL_3659 = _EVAL_3722 == 1'h0;
  assign _EVAL_4425 = _EVAL_3659 ? _EVAL_6019 : _EVAL_108;
  assign _EVAL_359 = _EVAL_3166 == 32'h0;
  assign _EVAL_4334 = _EVAL_5311 & 32'h4024;
  assign _EVAL_4045 = _EVAL_4334 == 32'h20;
  assign _EVAL_4858 = _EVAL_359 | _EVAL_4045;
  assign _EVAL_4602 = _EVAL_2164 & 32'h80000060;
  assign _EVAL_1634 = _EVAL_4602 == 32'h40;
  assign _EVAL_516 = _EVAL_2164 & 32'h10000060;
  assign _EVAL_3286 = _EVAL_516 == 32'h40;
  assign _EVAL_2154 = _EVAL_1634 | _EVAL_3286;
  assign _EVAL_3417 = _EVAL_4268 & 32'h40000040;
  assign _EVAL_4466 = _EVAL_3078 & 32'h2000040;
  assign _EVAL_4660 = _EVAL_3006 & 32'hfff0007f;
  assign _EVAL_1936 = _EVAL_4660 == 32'h58000053;
  assign _EVAL_4031 = _EVAL_2164 & 32'h80000010;
  assign _EVAL_975 = _EVAL_4031 == 32'h10;
  assign _EVAL_2233 = _EVAL_2438 == 32'h10;
  assign _EVAL_604 = _EVAL_975 | _EVAL_2233;
  assign _EVAL_5325 = _EVAL_2164 & 32'h40000040;
  assign _EVAL_2334 = _EVAL_5325 == 32'h40;
  assign _EVAL_3836 = _EVAL_604 | _EVAL_2334;
  assign _EVAL_5999 = _EVAL_3006 & 32'h207f;
  assign _EVAL_3098 = _EVAL_5999 == 32'h3;
  assign _EVAL_4355 = _EVAL_5386[12:2];
  assign _EVAL_2795 = _EVAL_4355 != 11'h0;
  assign _EVAL_1236 = _EVAL_179 ? _EVAL_5207 : 1'h1;
  assign _EVAL_1598 = _EVAL_268 ? 1'h1 : _EVAL_1236;
  assign _EVAL_4920 = _EVAL_3261 ? _EVAL_2795 : _EVAL_1598;
  assign _EVAL_5008 = _EVAL_3493 ? 1'h1 : _EVAL_4920;
  assign _EVAL_2116 = _EVAL_4185 ? 1'h1 : _EVAL_5008;
  assign _EVAL_846 = _EVAL_4999 ? 1'h1 : _EVAL_2116;
  assign _EVAL_4646 = _EVAL_5133 & 32'h80000010;
  assign _EVAL_2329 = _EVAL_4646 == 32'h10;
  assign _EVAL_1007 = _EVAL_2329 | _EVAL_4875;
  assign _EVAL_6137 = _EVAL_5133 & 32'h40000040;
  assign _EVAL_4639 = _EVAL_6137 == 32'h40;
  assign _EVAL_3310 = _EVAL_1007 | _EVAL_4639;
  assign _EVAL_5463 = _EVAL_5133 & 32'h20000040;
  assign _EVAL_5215 = _EVAL_5463 == 32'h40;
  assign _EVAL_3731 = _EVAL_3310 | _EVAL_5215;
  assign _EVAL_4244 = _EVAL_2680 == 32'h40;
  assign _EVAL_4239 = _EVAL_3731 | _EVAL_4244;
  assign _EVAL_4671 = _EVAL_5133 & 32'h1040;
  assign _EVAL_293 = _EVAL_4671 == 32'h1040;
  assign _EVAL_5268 = _EVAL_4239 | _EVAL_293;
  assign _EVAL_5622 = _EVAL_5133 & 32'h2040;
  assign _EVAL_2147 = _EVAL_5622 == 32'h2040;
  assign _EVAL_1652 = _EVAL_5268 | _EVAL_2147;
  assign _EVAL_4829 = _EVAL_597 ? _EVAL_863 : 1'h1;
  assign _EVAL_6006 = _EVAL_1674 ? 1'h1 : _EVAL_4829;
  assign _EVAL_4282 = _EVAL_936 ? _EVAL_3023 : _EVAL_6006;
  assign _EVAL_5384 = _EVAL_453 ? 1'h1 : _EVAL_4282;
  assign _EVAL_2669 = _EVAL_2288 ? 1'h1 : _EVAL_5384;
  assign _EVAL_1669 = _EVAL_4669 ? 1'h1 : _EVAL_2669;
  assign _EVAL_1537 = _EVAL_1669 == 1'h0;
  assign _EVAL_4583 = _EVAL_2039 & 32'heff0707f;
  assign _EVAL_5738 = _EVAL_4583 == 32'he0000053;
  assign _EVAL_1856 = _EVAL_1398 | _EVAL_5738;
  assign _EVAL_3133 = _EVAL_2039 & 32'hffd07fff;
  assign _EVAL_5912 = _EVAL_3133 == 32'hfc000073;
  assign _EVAL_3451 = _EVAL_1856 | _EVAL_5912;
  assign _EVAL_5582 = _EVAL_2039 & 32'h306f;
  assign _EVAL_2741 = _EVAL_5582 == 32'h1063;
  assign _EVAL_2296 = _EVAL_3451 | _EVAL_2741;
  assign _EVAL_939 = _EVAL_2039 & 32'h407f;
  assign _EVAL_4998 = _EVAL_939 == 32'h4063;
  assign _EVAL_1317 = _EVAL_2296 | _EVAL_4998;
  assign _EVAL_3609 = _EVAL_2039 & 32'h605f;
  assign _EVAL_2952 = _EVAL_3609 == 32'h3;
  assign _EVAL_2516 = _EVAL_1317 | _EVAL_2952;
  assign _EVAL_5756 = _EVAL_5582 == 32'h3;
  assign _EVAL_4004 = _EVAL_2516 | _EVAL_5756;
  assign _EVAL_5060 = _EVAL_1537 ? 1'h0 : _EVAL_4004;
  assign _EVAL_1912 = _EVAL_888 & 32'h5f;
  assign _EVAL_1027 = _EVAL_1912 == 32'h17;
  assign _EVAL_1541 = _EVAL_4882 & 32'h7e00507f;
  assign _EVAL_3323 = _EVAL_5875 | _EVAL_432;
  assign _EVAL_3018 = _EVAL_5854 & 32'hffd07fff;
  assign _EVAL_246 = _EVAL_4882 & 32'h4003044;
  assign _EVAL_715 = _EVAL_246 == 32'h4000040;
  assign _EVAL_5303 = _EVAL_3006[6:2];
  assign _EVAL_1163 = _EVAL_4882[6:2];
  assign _EVAL_1324 = _EVAL_5133[6:2];
  assign _EVAL_4638 = _EVAL_2901 ? _EVAL_1163 : _EVAL_1324;
  assign _EVAL_5452 = _EVAL_2378 ? _EVAL_5303 : _EVAL_4638;
  assign _EVAL_3003 = _EVAL_5690 ? _EVAL_5303 : _EVAL_5452;
  assign _EVAL_2570 = _EVAL_5690 ? _EVAL_3553 : _EVAL_3003;
  assign _EVAL_2405 = _EVAL_1242 & 32'hfff0007f;
  assign _EVAL_4978 = 29'h0 == _EVAL_5201;
  assign _EVAL_4462 = _EVAL_4978 & _EVAL_1385;
  assign _EVAL_2811 = _EVAL_4743 & 32'h7c;
  assign _EVAL_2858 = _EVAL_1242 & 32'h3c;
  assign _EVAL_624 = _EVAL_2858 == 32'h4;
  assign _EVAL_5670 = _EVAL_1242 & 32'h80000060;
  assign _EVAL_1868 = _EVAL_5670 == 32'h40;
  assign _EVAL_1356 = _EVAL_624 | _EVAL_1868;
  assign _EVAL_3194 = _EVAL_1242 & 32'h70;
  assign _EVAL_677 = _EVAL_3194 == 32'h40;
  assign _EVAL_213 = _EVAL_1356 | _EVAL_677;
  assign _EVAL_2500 = _EVAL_1242 & 32'h10000060;
  assign _EVAL_1846 = _EVAL_2500 == 32'h10000040;
  assign _EVAL_4206 = _EVAL_213 | _EVAL_1846;
  assign _EVAL_5908 = _EVAL_2164 & 32'h3c;
  assign _EVAL_950 = _EVAL_5908 == 32'h4;
  assign _EVAL_5438 = _EVAL_950 | _EVAL_1634;
  assign _EVAL_3088 = _EVAL_2164 & 32'h70;
  assign _EVAL_4890 = _EVAL_3088 == 32'h40;
  assign _EVAL_6037 = _EVAL_5438 | _EVAL_4890;
  assign _EVAL_2607 = _EVAL_516 == 32'h10000040;
  assign _EVAL_1464 = _EVAL_6037 | _EVAL_2607;
  assign _EVAL_2274 = _EVAL_1074 ? _EVAL_4206 : _EVAL_1464;
  assign _EVAL_1697 = _EVAL_1242 & 32'h2050;
  assign _EVAL_1327 = _EVAL_1697 == 32'h2000;
  assign _EVAL_397 = _EVAL_1975 | _EVAL_1327;
  assign _EVAL_5222 = _EVAL_1242 & 32'h90000034;
  assign _EVAL_4354 = _EVAL_5222 == 32'h90000010;
  assign _EVAL_270 = _EVAL_397 | _EVAL_4354;
  assign _EVAL_3413 = _EVAL_104;
  assign _EVAL_5525 = _EVAL_4492 & _EVAL_3413;
  assign _EVAL_5062 = 29'h0 < _EVAL_2382;
  assign _EVAL_1451 = 29'h0 == _EVAL_2382;
  assign _EVAL_4350 = _EVAL_1451 & _EVAL_4484;
  assign _EVAL_3426 = _EVAL_5062 | _EVAL_4350;
  assign _EVAL_2152 = _EVAL_3426 == _EVAL_1969;
  assign _EVAL_4510 = _EVAL_1451 & _EVAL_5676;
  assign _EVAL_351 = _EVAL_4291 ? _EVAL_2152 : _EVAL_4510;
  assign _EVAL_3787 = _EVAL_5525 & _EVAL_351;
  assign _EVAL_6131 = _EVAL_574 | _EVAL_3787;
  assign _EVAL_4373 = _EVAL_2039 & 32'h20000040;
  assign _EVAL_4084 = _EVAL_4373 == 32'h40;
  assign _EVAL_1985 = _EVAL_4286 | _EVAL_4084;
  assign _EVAL_5521 = _EVAL_2445 == 32'h40;
  assign _EVAL_3318 = _EVAL_1985 | _EVAL_5521;
  assign _EVAL_638 = _EVAL_2039 & 32'h1040;
  assign _EVAL_2879 = _EVAL_638 == 32'h1040;
  assign _EVAL_4528 = _EVAL_3318 | _EVAL_2879;
  assign _EVAL_6040 = _EVAL_2039 & 32'h2040;
  assign _EVAL_1264 = _EVAL_6040 == 32'h2040;
  assign _EVAL_5601 = _EVAL_4528 | _EVAL_1264;
  assign _EVAL_5495 = _EVAL_1242 & 32'h40000040;
  assign _EVAL_1205 = _EVAL_5495 == 32'h40;
  assign _EVAL_300 = _EVAL_4711 | _EVAL_1205;
  assign _EVAL_4504 = _EVAL_1242 & 32'h20000040;
  assign _EVAL_1399 = _EVAL_4504 == 32'h40;
  assign _EVAL_1219 = _EVAL_300 | _EVAL_1399;
  assign _EVAL_4055 = _EVAL_3076 == 32'h40;
  assign _EVAL_2692 = _EVAL_1219 | _EVAL_4055;
  assign _EVAL_6125 = _EVAL_1242 & 32'h1040;
  assign _EVAL_3435 = _EVAL_6125 == 32'h1040;
  assign _EVAL_3600 = _EVAL_2692 | _EVAL_3435;
  assign _EVAL_4596 = _EVAL_1242 & 32'h2040;
  assign _EVAL_2806 = _EVAL_4596 == 32'h2040;
  assign _EVAL_1005 = _EVAL_3600 | _EVAL_2806;
  assign _EVAL_5822 = _EVAL_2164 & 32'h20000040;
  assign _EVAL_445 = _EVAL_5822 == 32'h40;
  assign _EVAL_3931 = _EVAL_3836 | _EVAL_445;
  assign _EVAL_5432 = _EVAL_2438 == 32'h40;
  assign _EVAL_3732 = _EVAL_3931 | _EVAL_5432;
  assign _EVAL_1844 = _EVAL_2164 & 32'h1040;
  assign _EVAL_4209 = _EVAL_1844 == 32'h1040;
  assign _EVAL_2865 = _EVAL_3732 | _EVAL_4209;
  assign _EVAL_2843 = _EVAL_2164 & 32'h2040;
  assign _EVAL_6132 = _EVAL_2843 == 32'h2040;
  assign _EVAL_5326 = _EVAL_2865 | _EVAL_6132;
  assign _EVAL_5173 = _EVAL_1074 ? _EVAL_1005 : _EVAL_5326;
  assign _EVAL_2076 = _EVAL_5926 ? _EVAL_5601 : _EVAL_5173;
  assign _EVAL_2452 = _EVAL_4743 & 32'h605f;
  assign _EVAL_5193 = _EVAL_2452 == 32'h3;
  assign _EVAL_4704 = _EVAL_3271 & 32'h34;
  assign _EVAL_1955 = _EVAL_4704 == 32'h20;
  assign _EVAL_1879 = _EVAL_386 & 32'h207f;
  assign _EVAL_3770 = _EVAL_1879 == 32'h3;
  assign _EVAL_3911 = _EVAL_386 & 32'h607f;
  assign _EVAL_5611 = _EVAL_3911 == 32'hf;
  assign _EVAL_752 = _EVAL_3770 | _EVAL_5611;
  assign _EVAL_1515 = _EVAL_386 & 32'h5f;
  assign _EVAL_2895 = _EVAL_1515 == 32'h17;
  assign _EVAL_473 = _EVAL_752 | _EVAL_2895;
  assign _EVAL_1851 = _EVAL_386 & 32'hfc00007f;
  assign _EVAL_988 = _EVAL_1851 == 32'h33;
  assign _EVAL_1893 = _EVAL_473 | _EVAL_988;
  assign _EVAL_6075 = _EVAL_386 & 32'hbe00707f;
  assign _EVAL_247 = _EVAL_6075 == 32'h33;
  assign _EVAL_2875 = _EVAL_1893 | _EVAL_247;
  assign _EVAL_4548 = _EVAL_386 & 32'h6000073;
  assign _EVAL_1390 = _EVAL_4548 == 32'h43;
  assign _EVAL_3739 = _EVAL_2875 | _EVAL_1390;
  assign _EVAL_260 = _EVAL_386 & 32'he600007f;
  assign _EVAL_1819 = _EVAL_260 == 32'h53;
  assign _EVAL_340 = _EVAL_3739 | _EVAL_1819;
  assign _EVAL_4383 = _EVAL_386 & 32'h707b;
  assign _EVAL_3097 = _EVAL_4383 == 32'h63;
  assign _EVAL_1370 = _EVAL_340 | _EVAL_3097;
  assign _EVAL_1665 = _EVAL_386 & 32'h7f;
  assign _EVAL_4729 = _EVAL_1665 == 32'h6f;
  assign _EVAL_5876 = _EVAL_1370 | _EVAL_4729;
  assign _EVAL_2028 = _EVAL_386 & 32'hffefffff;
  assign _EVAL_3606 = _EVAL_2028 == 32'h73;
  assign _EVAL_1285 = _EVAL_5876 | _EVAL_3606;
  assign _EVAL_4174 = _EVAL_386 & 32'hfe00305f;
  assign _EVAL_4788 = _EVAL_4174 == 32'h1013;
  assign _EVAL_3711 = _EVAL_1285 | _EVAL_4788;
  assign _EVAL_518 = _EVAL_386 & 32'h705b;
  assign _EVAL_1511 = _EVAL_518 == 32'h2003;
  assign _EVAL_2229 = _EVAL_3711 | _EVAL_1511;
  assign _EVAL_2393 = _EVAL_1879 == 32'h2013;
  assign _EVAL_3214 = _EVAL_2229 | _EVAL_2393;
  assign _EVAL_5709 = _EVAL_386 & 32'h1800707f;
  assign _EVAL_5855 = _EVAL_5709 == 32'h202f;
  assign _EVAL_5745 = _EVAL_3214 | _EVAL_5855;
  assign _EVAL_4541 = _EVAL_1879 == 32'h2073;
  assign _EVAL_3211 = _EVAL_5745 | _EVAL_4541;
  assign _EVAL_1708 = _EVAL_386 & 32'hbe00705f;
  assign _EVAL_3784 = _EVAL_1708 == 32'h5013;
  assign _EVAL_5014 = _EVAL_3211 | _EVAL_3784;
  assign _EVAL_5058 = _EVAL_386 & 32'he800707f;
  assign _EVAL_3961 = _EVAL_5058 == 32'h800202f;
  assign _EVAL_1230 = _EVAL_5014 | _EVAL_3961;
  assign _EVAL_3605 = _EVAL_386 & 32'hf9f0707f;
  assign _EVAL_3419 = _EVAL_3605 == 32'h1000202f;
  assign _EVAL_3792 = _EVAL_1230 | _EVAL_3419;
  assign _EVAL_2338 = _EVAL_386 & 32'hdfffffff;
  assign _EVAL_1540 = _EVAL_2338 == 32'h10500073;
  assign _EVAL_546 = _EVAL_3792 | _EVAL_1540;
  assign _EVAL_4942 = _EVAL_386 & 32'hf600607f;
  assign _EVAL_2320 = _EVAL_4942 == 32'h20000053;
  assign _EVAL_710 = _EVAL_546 | _EVAL_2320;
  assign _EVAL_2587 = _EVAL_386 & 32'h7e00607f;
  assign _EVAL_5792 = _EVAL_2587 == 32'h20000053;
  assign _EVAL_731 = _EVAL_710 | _EVAL_5792;
  assign _EVAL_2980 = _EVAL_3111 == 32'h20000053;
  assign _EVAL_3700 = _EVAL_731 | _EVAL_2980;
  assign _EVAL_4980 = _EVAL_386 == 32'h30200073;
  assign _EVAL_5284 = _EVAL_3700 | _EVAL_4980;
  assign _EVAL_1374 = _EVAL_386 & 32'hfff0007f;
  assign _EVAL_1221 = _EVAL_1374 == 32'h58000053;
  assign _EVAL_3719 = _EVAL_5284 | _EVAL_1221;
  assign _EVAL_2578 = _EVAL_386 == 32'h7b200073;
  assign _EVAL_5482 = _EVAL_3719 | _EVAL_2578;
  assign _EVAL_5392 = _EVAL_386 & 32'hefe0007f;
  assign _EVAL_2571 = _EVAL_5392 == 32'hc0000053;
  assign _EVAL_3533 = _EVAL_5482 | _EVAL_2571;
  assign _EVAL_5464 = _EVAL_386 & 32'hfff0607f;
  assign _EVAL_4989 = _EVAL_5464 == 32'he0000053;
  assign _EVAL_5488 = _EVAL_3533 | _EVAL_4989;
  assign _EVAL_5584 = _EVAL_386 & 32'heff0707f;
  assign _EVAL_5784 = _EVAL_5584 == 32'he0000053;
  assign _EVAL_5234 = _EVAL_5488 | _EVAL_5784;
  assign _EVAL_503 = _EVAL_1978 & 32'h80000010;
  assign _EVAL_2783 = _EVAL_503 == 32'h10;
  assign _EVAL_596 = _EVAL_1978 & 32'h50;
  assign _EVAL_929 = _EVAL_596 == 32'h10;
  assign _EVAL_585 = _EVAL_2783 | _EVAL_929;
  assign _EVAL_6051 = _EVAL_1978 & 32'h40000040;
  assign _EVAL_848 = _EVAL_6051 == 32'h40;
  assign _EVAL_3063 = _EVAL_585 | _EVAL_848;
  assign _EVAL_4835 = _EVAL_1978 & 32'h20000040;
  assign _EVAL_2854 = _EVAL_4835 == 32'h40;
  assign _EVAL_891 = _EVAL_3063 | _EVAL_2854;
  assign _EVAL_5186 = _EVAL_596 == 32'h40;
  assign _EVAL_1151 = _EVAL_891 | _EVAL_5186;
  assign _EVAL_3071 = _EVAL_1978 & 32'h1040;
  assign _EVAL_5167 = _EVAL_3071 == 32'h1040;
  assign _EVAL_1822 = _EVAL_1151 | _EVAL_5167;
  assign _EVAL_4432 = _EVAL_4702 & 32'h44;
  assign _EVAL_4517 = _EVAL_4432 == 32'h0;
  assign _EVAL_5056 = _EVAL_5899 | _EVAL_1027;
  assign _EVAL_238 = _EVAL_888 & 32'hfc00007f;
  assign _EVAL_4657 = _EVAL_238 == 32'h33;
  assign _EVAL_4016 = _EVAL_5056 | _EVAL_4657;
  assign _EVAL_5664 = _EVAL_888 & 32'hbe00707f;
  assign _EVAL_1257 = _EVAL_5664 == 32'h33;
  assign _EVAL_2239 = _EVAL_4016 | _EVAL_1257;
  assign _EVAL_3074 = _EVAL_888 & 32'h6000073;
  assign _EVAL_5028 = _EVAL_3074 == 32'h43;
  assign _EVAL_3056 = _EVAL_2239 | _EVAL_5028;
  assign _EVAL_1590 = _EVAL_888 & 32'he600007f;
  assign _EVAL_2493 = _EVAL_1590 == 32'h53;
  assign _EVAL_4052 = _EVAL_3056 | _EVAL_2493;
  assign _EVAL_2244 = _EVAL_888 & 32'h707b;
  assign _EVAL_1420 = _EVAL_2244 == 32'h63;
  assign _EVAL_3515 = _EVAL_4052 | _EVAL_1420;
  assign _EVAL_3741 = _EVAL_888 & 32'h7f;
  assign _EVAL_1018 = _EVAL_3741 == 32'h6f;
  assign _EVAL_5898 = _EVAL_3515 | _EVAL_1018;
  assign _EVAL_2976 = _EVAL_888 & 32'hffefffff;
  assign _EVAL_2961 = _EVAL_2976 == 32'h73;
  assign _EVAL_484 = _EVAL_5898 | _EVAL_2961;
  assign _EVAL_1292 = _EVAL_888 & 32'hfe00305f;
  assign _EVAL_679 = _EVAL_1292 == 32'h1013;
  assign _EVAL_4151 = _EVAL_484 | _EVAL_679;
  assign _EVAL_6111 = _EVAL_888 & 32'h705b;
  assign _EVAL_297 = _EVAL_6111 == 32'h2003;
  assign _EVAL_2684 = _EVAL_4151 | _EVAL_297;
  assign _EVAL_564 = _EVAL_5400 == 32'h2013;
  assign _EVAL_3369 = _EVAL_2684 | _EVAL_564;
  assign _EVAL_279 = _EVAL_888 & 32'h1800707f;
  assign _EVAL_5446 = _EVAL_279 == 32'h202f;
  assign _EVAL_5232 = _EVAL_3369 | _EVAL_5446;
  assign _EVAL_4060 = _EVAL_5400 == 32'h2073;
  assign _EVAL_4171 = _EVAL_5232 | _EVAL_4060;
  assign _EVAL_4795 = _EVAL_888 & 32'hbe00705f;
  assign _EVAL_4409 = _EVAL_4795 == 32'h5013;
  assign _EVAL_5783 = _EVAL_4171 | _EVAL_4409;
  assign _EVAL_895 = _EVAL_888 & 32'he800707f;
  assign _EVAL_5491 = _EVAL_895 == 32'h800202f;
  assign _EVAL_2905 = _EVAL_5783 | _EVAL_5491;
  assign _EVAL_5776 = _EVAL_888 & 32'hfff0607f;
  assign _EVAL_4076 = _EVAL_2970 ? _EVAL_3655 : _EVAL_880;
  assign _EVAL_1224 = _EVAL_4743 & 32'h44;
  assign _EVAL_2759 = _EVAL_1224 == 32'h0;
  assign _EVAL_3693 = _EVAL_4743 & 32'h4024;
  assign _EVAL_1685 = _EVAL_3693 == 32'h20;
  assign _EVAL_5621 = _EVAL_2759 | _EVAL_1685;
  assign _EVAL_3729 = _EVAL_4743 & 32'h38;
  assign _EVAL_4415 = _EVAL_3729 == 32'h20;
  assign _EVAL_728 = _EVAL_5621 | _EVAL_4415;
  assign _EVAL_4263 = _EVAL_4743 & 32'h2050;
  assign _EVAL_3521 = _EVAL_4263 == 32'h2000;
  assign _EVAL_344 = _EVAL_728 | _EVAL_3521;
  assign _EVAL_273 = _EVAL_4743 & 32'h90000034;
  assign _EVAL_5494 = _EVAL_273 == 32'h90000010;
  assign _EVAL_5688 = _EVAL_344 | _EVAL_5494;
  assign _EVAL_3638 = _EVAL_1362 & 32'h5f;
  assign _EVAL_5978 = _EVAL_3638 == 32'h17;
  assign _EVAL_1501 = _EVAL_386 & 32'h2024;
  assign _EVAL_4468 = _EVAL_1501 == 32'h24;
  assign _EVAL_3806 = _EVAL_983 | _EVAL_4468;
  assign _EVAL_337 = _EVAL_386 & 32'h28;
  assign _EVAL_4269 = _EVAL_337 == 32'h28;
  assign _EVAL_1315 = _EVAL_3806 | _EVAL_4269;
  assign _EVAL_2148 = _EVAL_386 & 32'h30;
  assign _EVAL_1559 = _EVAL_2148 == 32'h30;
  assign _EVAL_1835 = _EVAL_1315 | _EVAL_1559;
  assign _EVAL_2685 = _EVAL_5311 & 32'h207f;
  assign _EVAL_5581 = _EVAL_2685 == 32'h3;
  assign _EVAL_499 = _EVAL_5311 & 32'h607f;
  assign _EVAL_497 = _EVAL_499 == 32'hf;
  assign _EVAL_2161 = _EVAL_5581 | _EVAL_497;
  assign _EVAL_4913 = _EVAL_2161 | _EVAL_6120;
  assign _EVAL_2530 = _EVAL_5311 & 32'hfc00007f;
  assign _EVAL_2697 = _EVAL_2530 == 32'h33;
  assign _EVAL_4142 = _EVAL_4913 | _EVAL_2697;
  assign _EVAL_2881 = _EVAL_5311 & 32'hbe00707f;
  assign _EVAL_4863 = _EVAL_2881 == 32'h33;
  assign _EVAL_4509 = _EVAL_4142 | _EVAL_4863;
  assign _EVAL_3208 = _EVAL_5311 & 32'h6000073;
  assign _EVAL_4512 = _EVAL_3208 == 32'h43;
  assign _EVAL_1126 = _EVAL_4509 | _EVAL_4512;
  assign _EVAL_2910 = _EVAL_5311 & 32'he600007f;
  assign _EVAL_4129 = _EVAL_2910 == 32'h53;
  assign _EVAL_3660 = _EVAL_1126 | _EVAL_4129;
  assign _EVAL_2574 = _EVAL_5311 & 32'h707b;
  assign _EVAL_3724 = _EVAL_2574 == 32'h63;
  assign _EVAL_3322 = _EVAL_3660 | _EVAL_3724;
  assign _EVAL_1068 = _EVAL_5311 & 32'h7f;
  assign _EVAL_5524 = _EVAL_1068 == 32'h6f;
  assign _EVAL_3264 = _EVAL_3322 | _EVAL_5524;
  assign _EVAL_739 = _EVAL_5311 & 32'hffefffff;
  assign _EVAL_3639 = _EVAL_739 == 32'h73;
  assign _EVAL_4644 = _EVAL_3264 | _EVAL_3639;
  assign _EVAL_2193 = _EVAL_5311 & 32'hfe00305f;
  assign _EVAL_5117 = _EVAL_2193 == 32'h1013;
  assign _EVAL_5749 = _EVAL_4644 | _EVAL_5117;
  assign _EVAL_5274 = _EVAL_5311 & 32'h705b;
  assign _EVAL_4725 = _EVAL_5274 == 32'h2003;
  assign _EVAL_5633 = _EVAL_5749 | _EVAL_4725;
  assign _EVAL_1057 = _EVAL_2685 == 32'h2013;
  assign _EVAL_5182 = _EVAL_5633 | _EVAL_1057;
  assign _EVAL_5919 = _EVAL_5311 & 32'h1800707f;
  assign _EVAL_5773 = _EVAL_5919 == 32'h202f;
  assign _EVAL_3040 = _EVAL_5182 | _EVAL_5773;
  assign _EVAL_3661 = _EVAL_2685 == 32'h2073;
  assign _EVAL_3184 = _EVAL_3040 | _EVAL_3661;
  assign _EVAL_3135 = _EVAL_5311 & 32'hbe00705f;
  assign _EVAL_1546 = _EVAL_3135 == 32'h5013;
  assign _EVAL_3734 = _EVAL_3184 | _EVAL_1546;
  assign _EVAL_3374 = _EVAL_5311 & 32'he800707f;
  assign _EVAL_1241 = _EVAL_3374 == 32'h800202f;
  assign _EVAL_2882 = _EVAL_3734 | _EVAL_1241;
  assign _EVAL_5646 = _EVAL_5311 & 32'hf9f0707f;
  assign _EVAL_495 = _EVAL_5646 == 32'h1000202f;
  assign _EVAL_1790 = _EVAL_2882 | _EVAL_495;
  assign _EVAL_2829 = _EVAL_5311 & 32'hdfffffff;
  assign _EVAL_5752 = _EVAL_2829 == 32'h10500073;
  assign _EVAL_4971 = _EVAL_1790 | _EVAL_5752;
  assign _EVAL_5240 = _EVAL_5311 & 32'hf600607f;
  assign _EVAL_1933 = _EVAL_5240 == 32'h20000053;
  assign _EVAL_2459 = _EVAL_4971 | _EVAL_1933;
  assign _EVAL_3522 = _EVAL_5311 & 32'h7e00607f;
  assign _EVAL_332 = _EVAL_3522 == 32'h20000053;
  assign _EVAL_354 = _EVAL_2459 | _EVAL_332;
  assign _EVAL_4973 = _EVAL_5311 & 32'h7e00507f;
  assign _EVAL_666 = _EVAL_4973 == 32'h20000053;
  assign _EVAL_4724 = _EVAL_354 | _EVAL_666;
  assign _EVAL_4668 = _EVAL_5311 == 32'h30200073;
  assign _EVAL_629 = _EVAL_4724 | _EVAL_4668;
  assign _EVAL_2074 = _EVAL_5311 & 32'hfff0007f;
  assign _EVAL_5479 = _EVAL_2074 == 32'h58000053;
  assign _EVAL_4859 = _EVAL_629 | _EVAL_5479;
  assign _EVAL_5105 = _EVAL_5311 == 32'h7b200073;
  assign _EVAL_5808 = _EVAL_4859 | _EVAL_5105;
  assign _EVAL_3686 = _EVAL_5311 & 32'hefe0007f;
  assign _EVAL_2196 = _EVAL_3686 == 32'hc0000053;
  assign _EVAL_5907 = _EVAL_5808 | _EVAL_2196;
  assign _EVAL_3696 = _EVAL_5311 & 32'hfff0607f;
  assign _EVAL_6077 = _EVAL_3696 == 32'he0000053;
  assign _EVAL_4977 = _EVAL_5907 | _EVAL_6077;
  assign _EVAL_1620 = _EVAL_5311 & 32'heff0707f;
  assign _EVAL_2386 = _EVAL_1620 == 32'he0000053;
  assign _EVAL_954 = _EVAL_4977 | _EVAL_2386;
  assign _EVAL_5029 = _EVAL_5311 & 32'hffd07fff;
  assign _EVAL_2185 = _EVAL_5029 == 32'hfc000073;
  assign _EVAL_3036 = _EVAL_954 | _EVAL_2185;
  assign _EVAL_962 = _EVAL_1291 == 32'h1063;
  assign _EVAL_504 = _EVAL_3036 | _EVAL_962;
  assign _EVAL_1300 = _EVAL_2164 & 32'h2010;
  assign _EVAL_3577 = _EVAL_3006 == 32'h30200073;
  assign _EVAL_4069 = _EVAL_4268 & 32'h3c;
  assign _EVAL_4074 = _EVAL_4069 == 32'h4;
  assign _EVAL_5170 = _EVAL_4268 & 32'h80000060;
  assign _EVAL_3788 = _EVAL_5170 == 32'h40;
  assign _EVAL_4451 = _EVAL_4074 | _EVAL_3788;
  assign _EVAL_2863 = _EVAL_4882 & 32'h607f;
  assign _EVAL_4965 = _EVAL_2863 == 32'hf;
  assign _EVAL_741 = _EVAL_1702 | _EVAL_4965;
  assign _EVAL_5883 = _EVAL_4882 & 32'h5f;
  assign _EVAL_4495 = _EVAL_5883 == 32'h17;
  assign _EVAL_450 = _EVAL_741 | _EVAL_4495;
  assign _EVAL_4604 = _EVAL_4882 & 32'hfc00007f;
  assign _EVAL_3222 = _EVAL_4604 == 32'h33;
  assign _EVAL_321 = _EVAL_450 | _EVAL_3222;
  assign _EVAL_1673 = _EVAL_4882 & 32'hbe00707f;
  assign _EVAL_3115 = _EVAL_1673 == 32'h33;
  assign _EVAL_4235 = _EVAL_321 | _EVAL_3115;
  assign _EVAL_4692 = _EVAL_4882 & 32'h6000073;
  assign _EVAL_4439 = _EVAL_4692 == 32'h43;
  assign _EVAL_460 = _EVAL_4235 | _EVAL_4439;
  assign _EVAL_3121 = _EVAL_4882 & 32'he600007f;
  assign _EVAL_4255 = _EVAL_3121 == 32'h53;
  assign _EVAL_911 = _EVAL_460 | _EVAL_4255;
  assign _EVAL_4708 = _EVAL_4882 & 32'h707b;
  assign _EVAL_5176 = _EVAL_4708 == 32'h63;
  assign _EVAL_4511 = _EVAL_911 | _EVAL_5176;
  assign _EVAL_2519 = _EVAL_4882 & 32'h7f;
  assign _EVAL_2612 = _EVAL_2519 == 32'h6f;
  assign _EVAL_1392 = _EVAL_4511 | _EVAL_2612;
  assign _EVAL_533 = _EVAL_4882 & 32'hffefffff;
  assign _EVAL_6117 = _EVAL_533 == 32'h73;
  assign _EVAL_5586 = _EVAL_1392 | _EVAL_6117;
  assign _EVAL_5990 = _EVAL_4882 & 32'hfe00305f;
  assign _EVAL_5637 = _EVAL_5990 == 32'h1013;
  assign _EVAL_5189 = _EVAL_5586 | _EVAL_5637;
  assign _EVAL_4739 = _EVAL_4882 & 32'h705b;
  assign _EVAL_3290 = _EVAL_4739 == 32'h2003;
  assign _EVAL_353 = _EVAL_5189 | _EVAL_3290;
  assign _EVAL_2868 = _EVAL_3298 == 32'h2013;
  assign _EVAL_4545 = _EVAL_353 | _EVAL_2868;
  assign _EVAL_4048 = _EVAL_4882 & 32'h1800707f;
  assign _EVAL_5585 = _EVAL_4048 == 32'h202f;
  assign _EVAL_1877 = _EVAL_4545 | _EVAL_5585;
  assign _EVAL_3851 = _EVAL_3298 == 32'h2073;
  assign _EVAL_1435 = _EVAL_1877 | _EVAL_3851;
  assign _EVAL_1732 = _EVAL_4882 & 32'hbe00705f;
  assign _EVAL_1417 = _EVAL_1732 == 32'h5013;
  assign _EVAL_404 = _EVAL_1435 | _EVAL_1417;
  assign _EVAL_4011 = _EVAL_4882 & 32'he800707f;
  assign _EVAL_985 = _EVAL_4011 == 32'h800202f;
  assign _EVAL_5590 = _EVAL_404 | _EVAL_985;
  assign _EVAL_6014 = _EVAL_4882 & 32'hf9f0707f;
  assign _EVAL_2431 = _EVAL_6014 == 32'h1000202f;
  assign _EVAL_5097 = _EVAL_5590 | _EVAL_2431;
  assign _EVAL_1989 = _EVAL_4882 & 32'hdfffffff;
  assign _EVAL_714 = _EVAL_1989 == 32'h10500073;
  assign _EVAL_2809 = _EVAL_5097 | _EVAL_714;
  assign _EVAL_368 = _EVAL_4882 & 32'hf600607f;
  assign _EVAL_3484 = _EVAL_368 == 32'h20000053;
  assign _EVAL_5316 = _EVAL_2809 | _EVAL_3484;
  assign _EVAL_1311 = _EVAL_4882 & 32'h7e00607f;
  assign _EVAL_857 = _EVAL_1311 == 32'h20000053;
  assign _EVAL_2623 = _EVAL_5316 | _EVAL_857;
  assign _EVAL_1099 = _EVAL_1541 == 32'h20000053;
  assign _EVAL_2473 = _EVAL_2623 | _EVAL_1099;
  assign _EVAL_3915 = _EVAL_4882 == 32'h30200073;
  assign _EVAL_2097 = _EVAL_2473 | _EVAL_3915;
  assign _EVAL_364 = _EVAL_4882 & 32'hfff0007f;
  assign _EVAL_615 = _EVAL_364 == 32'h58000053;
  assign _EVAL_5694 = _EVAL_2097 | _EVAL_615;
  assign _EVAL_5458 = _EVAL_4882 == 32'h7b200073;
  assign _EVAL_978 = _EVAL_5694 | _EVAL_5458;
  assign _EVAL_3549 = _EVAL_4882 & 32'hefe0007f;
  assign _EVAL_4857 = _EVAL_3549 == 32'hc0000053;
  assign _EVAL_1167 = _EVAL_978 | _EVAL_4857;
  assign _EVAL_1144 = _EVAL_2259 == 32'h20;
  assign _EVAL_637 = _EVAL_386 & 32'h34;
  assign _EVAL_993 = _EVAL_637 == 32'h20;
  assign _EVAL_236 = _EVAL_1144 | _EVAL_993;
  assign _EVAL_2694 = _EVAL_3271 & 32'h3c;
  assign _EVAL_4589 = _EVAL_5854 & 32'h2000040;
  assign _EVAL_4064 = _EVAL_3271 & 32'hffd07fff;
  assign _EVAL_4598 = _EVAL_4064 == 32'hfc000073;
  assign _EVAL_3487 = _EVAL_2901 ? _EVAL_2101 : _EVAL_5949;
  assign _EVAL_2851 = _EVAL_2378 ? _EVAL_3390 : _EVAL_3487;
  assign _EVAL_3415 = _EVAL_3078 & 32'h38;
  assign _EVAL_2344 = _EVAL_1978 & 32'h64;
  assign _EVAL_6074 = _EVAL_2344 == 32'h0;
  assign _EVAL_5772 = _EVAL_6074 | _EVAL_929;
  assign _EVAL_1960 = _EVAL_1978 & 32'h2024;
  assign _EVAL_1484 = _EVAL_1960 == 32'h24;
  assign _EVAL_2703 = _EVAL_5772 | _EVAL_1484;
  assign _EVAL_2460 = _EVAL_5133 & 32'hffd07fff;
  assign _EVAL_4159 = _EVAL_2164 & 32'h18;
  assign _EVAL_5558 = _EVAL_4159 == 32'h0;
  assign _EVAL_3785 = _EVAL_1300 == 32'h2000;
  assign _EVAL_394 = _EVAL_5558 | _EVAL_3785;
  assign _EVAL_5739 = _EVAL_2164 & 32'h8000040;
  assign _EVAL_4413 = _EVAL_5739 == 32'h8000040;
  assign _EVAL_2944 = _EVAL_394 | _EVAL_4413;
  assign _EVAL_3022 = _EVAL_4702 & 32'h607f;
  assign _EVAL_4606 = _EVAL_1242 & 32'hffd07fff;
  assign _EVAL_2069 = _EVAL_4606 == 32'hfc000073;
  assign _EVAL_730 = _EVAL_654[12:2];
  assign _EVAL_2844 = _EVAL_4702 & 32'he600007f;
  assign _EVAL_974 = _EVAL_411 == 32'h0;
  assign _EVAL_5691 = _EVAL_4882 & 32'h4024;
  assign _EVAL_2772 = _EVAL_5691 == 32'h20;
  assign _EVAL_767 = _EVAL_974 | _EVAL_2772;
  assign _EVAL_471 = _EVAL_4882 & 32'h38;
  assign _EVAL_567 = _EVAL_471 == 32'h20;
  assign _EVAL_5569 = _EVAL_767 | _EVAL_567;
  assign _EVAL_5350 = _EVAL_4882 & 32'h2050;
  assign _EVAL_628 = _EVAL_5350 == 32'h2000;
  assign _EVAL_3509 = _EVAL_5569 | _EVAL_628;
  assign _EVAL_4953 = _EVAL_2714 == 32'h90000010;
  assign _EVAL_889 = _EVAL_3509 | _EVAL_4953;
  assign _EVAL_6026 = _EVAL_1947 & 32'hf600607f;
  assign _EVAL_2064 = _EVAL_6026 == 32'h20000053;
  assign _EVAL_4941 = _EVAL_888 & 32'h70;
  assign _EVAL_697 = _EVAL_4941 == 32'h40;
  assign _EVAL_2853 = _EVAL_3570 ? _EVAL_697 : _EVAL_4136;
  assign _EVAL_4395 = _EVAL_5833 ? _EVAL_697 : _EVAL_2853;
  assign _EVAL_927 = _EVAL_5311 & 32'h34;
  assign _EVAL_1460 = _EVAL_927 == 32'h20;
  assign _EVAL_5297 = _EVAL_3078[11:7];
  assign _EVAL_4371 = _EVAL_5297 != 5'h0;
  assign _EVAL_5657 = _EVAL_3006 & 32'h38;
  assign _EVAL_5124 = _EVAL_3006 & 32'h607f;
  assign _EVAL_3635 = _EVAL_5124 == 32'hf;
  assign _EVAL_3029 = _EVAL_3098 | _EVAL_3635;
  assign _EVAL_1318 = _EVAL_3006 & 32'h5f;
  assign _EVAL_4749 = _EVAL_1318 == 32'h17;
  assign _EVAL_2509 = _EVAL_3029 | _EVAL_4749;
  assign _EVAL_4106 = _EVAL_3006 & 32'hfc00007f;
  assign _EVAL_1667 = _EVAL_4106 == 32'h33;
  assign _EVAL_653 = _EVAL_2509 | _EVAL_1667;
  assign _EVAL_267 = _EVAL_3006 & 32'hbe00707f;
  assign _EVAL_1693 = _EVAL_267 == 32'h33;
  assign _EVAL_3332 = _EVAL_653 | _EVAL_1693;
  assign _EVAL_4412 = _EVAL_3006 & 32'h6000073;
  assign _EVAL_3192 = _EVAL_4412 == 32'h43;
  assign _EVAL_4804 = _EVAL_3332 | _EVAL_3192;
  assign _EVAL_565 = _EVAL_3006 & 32'he600007f;
  assign _EVAL_5360 = _EVAL_565 == 32'h53;
  assign _EVAL_3790 = _EVAL_4804 | _EVAL_5360;
  assign _EVAL_5389 = _EVAL_3006 & 32'h707b;
  assign _EVAL_4187 = _EVAL_5389 == 32'h63;
  assign _EVAL_5194 = _EVAL_3790 | _EVAL_4187;
  assign _EVAL_3262 = _EVAL_3006 & 32'h7f;
  assign _EVAL_3963 = _EVAL_3262 == 32'h6f;
  assign _EVAL_2359 = _EVAL_5194 | _EVAL_3963;
  assign _EVAL_2825 = _EVAL_3006 & 32'hffefffff;
  assign _EVAL_5496 = _EVAL_2825 == 32'h73;
  assign _EVAL_2054 = _EVAL_2359 | _EVAL_5496;
  assign _EVAL_5531 = _EVAL_3006 & 32'hfe00305f;
  assign _EVAL_1866 = _EVAL_5531 == 32'h1013;
  assign _EVAL_634 = _EVAL_2054 | _EVAL_1866;
  assign _EVAL_2465 = _EVAL_3006 & 32'h705b;
  assign _EVAL_3428 = _EVAL_2465 == 32'h2003;
  assign _EVAL_5932 = _EVAL_634 | _EVAL_3428;
  assign _EVAL_4167 = _EVAL_5999 == 32'h2013;
  assign _EVAL_4450 = _EVAL_5932 | _EVAL_4167;
  assign _EVAL_2012 = _EVAL_3006 & 32'h1800707f;
  assign _EVAL_5896 = _EVAL_2012 == 32'h202f;
  assign _EVAL_5210 = _EVAL_4450 | _EVAL_5896;
  assign _EVAL_2476 = _EVAL_5999 == 32'h2073;
  assign _EVAL_3632 = _EVAL_5210 | _EVAL_2476;
  assign _EVAL_2191 = _EVAL_1947 & 32'h7e00507f;
  assign _EVAL_1635 = _EVAL_3006[24:20];
  assign _EVAL_1662 = _EVAL_4882[24:20];
  assign _EVAL_5293 = _EVAL_5133[24:20];
  assign _EVAL_2862 = _EVAL_2901 ? _EVAL_1662 : _EVAL_5293;
  assign _EVAL_1332 = _EVAL_2378 ? _EVAL_1635 : _EVAL_2862;
  assign _EVAL_3514 = _EVAL_2666[12:2];
  assign _EVAL_769 = _EVAL_3514 != 11'h0;
  assign _EVAL_1364 = _EVAL_1014 ? _EVAL_5924 : 1'h1;
  assign _EVAL_5923 = _EVAL_4352 ? 1'h1 : _EVAL_1364;
  assign _EVAL_5104 = _EVAL_4202 ? _EVAL_769 : _EVAL_5923;
  assign _EVAL_2464 = _EVAL_2644 ? 1'h1 : _EVAL_5104;
  assign _EVAL_1198 = _EVAL_5813 & 32'h407f;
  assign _EVAL_1935 = _EVAL_1242 & 32'h7c;
  assign _EVAL_1573 = {_EVAL_1746,_EVAL_2272};
  assign _EVAL_5245 = _EVAL_1573 != 12'h0;
  assign _EVAL_4002 = _EVAL_268 ? _EVAL_5245 : 1'h1;
  assign _EVAL_3675 = _EVAL_3261 ? 1'h1 : _EVAL_4002;
  assign _EVAL_922 = _EVAL_3493 ? 1'h1 : _EVAL_3675;
  assign _EVAL_1350 = _EVAL_4185 ? 1'h1 : _EVAL_922;
  assign _EVAL_5243 = _EVAL_4999 ? 1'h1 : _EVAL_1350;
  assign _EVAL_1405 = _EVAL_5243 == 1'h0;
  assign _EVAL_1263 = _EVAL_5311 & 32'h80000010;
  assign _EVAL_2411 = _EVAL_1263 == 32'h10;
  assign _EVAL_6083 = _EVAL_1733 == 32'h10;
  assign _EVAL_5925 = _EVAL_2411 | _EVAL_6083;
  assign _EVAL_2550 = _EVAL_5925 | _EVAL_641;
  assign _EVAL_2434 = _EVAL_5311 & 32'h20000040;
  assign _EVAL_524 = _EVAL_2434 == 32'h40;
  assign _EVAL_1800 = _EVAL_2550 | _EVAL_524;
  assign _EVAL_5300 = _EVAL_1733 == 32'h40;
  assign _EVAL_5589 = _EVAL_1800 | _EVAL_5300;
  assign _EVAL_2234 = _EVAL_5311 & 32'h1040;
  assign _EVAL_542 = _EVAL_2234 == 32'h1040;
  assign _EVAL_1820 = _EVAL_5589 | _EVAL_542;
  assign _EVAL_280 = _EVAL_5311 & 32'h2040;
  assign _EVAL_3976 = _EVAL_280 == 32'h2040;
  assign _EVAL_307 = _EVAL_1820 | _EVAL_3976;
  assign _EVAL_304 = {_EVAL_3905,_EVAL_2142,_EVAL_3052,_EVAL_5276};
  assign _EVAL_4463 = _EVAL_2164 & 32'h30;
  assign _EVAL_1495 = _EVAL_4463 == 32'h30;
  assign _EVAL_1995 = _EVAL_5133 & 32'h7c;
  assign _EVAL_5658 = _EVAL_1995 == 32'h24;
  assign _EVAL_3348 = _EVAL_2164 & 32'h7c;
  assign _EVAL_1728 = _EVAL_3348 == 32'h24;
  assign _EVAL_5528 = _EVAL_2164 & 32'h40000060;
  assign _EVAL_610 = _EVAL_5528 == 32'h40;
  assign _EVAL_2687 = _EVAL_1728 | _EVAL_610;
  assign _EVAL_4421 = _EVAL_2687 | _EVAL_4890;
  assign _EVAL_3499 = _EVAL_1947 & 32'h207f;
  assign _EVAL_850 = _EVAL_3499 == 32'h3;
  assign _EVAL_4118 = _EVAL_1947 & 32'h607f;
  assign _EVAL_1186 = _EVAL_4118 == 32'hf;
  assign _EVAL_345 = _EVAL_850 | _EVAL_1186;
  assign _EVAL_2287 = _EVAL_1947 & 32'h5f;
  assign _EVAL_528 = _EVAL_2287 == 32'h17;
  assign _EVAL_5202 = _EVAL_345 | _EVAL_528;
  assign _EVAL_2146 = _EVAL_1947 & 32'hfc00007f;
  assign _EVAL_5818 = _EVAL_2146 == 32'h33;
  assign _EVAL_1059 = _EVAL_5202 | _EVAL_5818;
  assign _EVAL_1083 = _EVAL_1947 & 32'hbe00707f;
  assign _EVAL_582 = _EVAL_1083 == 32'h33;
  assign _EVAL_758 = _EVAL_1059 | _EVAL_582;
  assign _EVAL_1942 = _EVAL_1947 & 32'h6000073;
  assign _EVAL_849 = _EVAL_1942 == 32'h43;
  assign _EVAL_4473 = _EVAL_758 | _EVAL_849;
  assign _EVAL_3424 = _EVAL_1947 & 32'he600007f;
  assign _EVAL_4197 = _EVAL_3424 == 32'h53;
  assign _EVAL_813 = _EVAL_4473 | _EVAL_4197;
  assign _EVAL_5348 = _EVAL_1947 & 32'h707b;
  assign _EVAL_4649 = _EVAL_5348 == 32'h63;
  assign _EVAL_4505 = _EVAL_813 | _EVAL_4649;
  assign _EVAL_2757 = _EVAL_1947 & 32'h7f;
  assign _EVAL_4860 = _EVAL_2757 == 32'h6f;
  assign _EVAL_1783 = _EVAL_4505 | _EVAL_4860;
  assign _EVAL_5501 = _EVAL_1947 & 32'hffefffff;
  assign _EVAL_2872 = _EVAL_5501 == 32'h73;
  assign _EVAL_5862 = _EVAL_1783 | _EVAL_2872;
  assign _EVAL_5877 = _EVAL_1947 & 32'hfe00305f;
  assign _EVAL_5280 = _EVAL_5877 == 32'h1013;
  assign _EVAL_2269 = _EVAL_5862 | _EVAL_5280;
  assign _EVAL_3796 = _EVAL_1947 & 32'h705b;
  assign _EVAL_2502 = _EVAL_3796 == 32'h2003;
  assign _EVAL_5233 = _EVAL_2269 | _EVAL_2502;
  assign _EVAL_177 = _EVAL_3499 == 32'h2013;
  assign _EVAL_3394 = _EVAL_5233 | _EVAL_177;
  assign _EVAL_2072 = _EVAL_1947 & 32'h1800707f;
  assign _EVAL_1261 = _EVAL_2072 == 32'h202f;
  assign _EVAL_2527 = _EVAL_3394 | _EVAL_1261;
  assign _EVAL_2748 = _EVAL_3499 == 32'h2073;
  assign _EVAL_2746 = _EVAL_2527 | _EVAL_2748;
  assign _EVAL_5144 = _EVAL_1947 & 32'hbe00705f;
  assign _EVAL_1104 = _EVAL_5144 == 32'h5013;
  assign _EVAL_5110 = _EVAL_2746 | _EVAL_1104;
  assign _EVAL_2083 = _EVAL_1947 & 32'he800707f;
  assign _EVAL_3599 = _EVAL_2083 == 32'h800202f;
  assign _EVAL_1442 = _EVAL_5110 | _EVAL_3599;
  assign _EVAL_623 = _EVAL_3985 == 32'h1000202f;
  assign _EVAL_2123 = _EVAL_1442 | _EVAL_623;
  assign _EVAL_3067 = _EVAL_4702 & 32'h2010;
  assign _EVAL_2859 = _EVAL_3067 == 32'h2000;
  assign _EVAL_4086 = _EVAL_2710 == 32'h3;
  assign _EVAL_2581 = _EVAL_1362 & 32'h607f;
  assign _EVAL_2201 = _EVAL_2581 == 32'hf;
  assign _EVAL_2507 = _EVAL_4086 | _EVAL_2201;
  assign _EVAL_1064 = _EVAL_3528 != 2'h3;
  assign _EVAL_915 = _EVAL_1069 == 1'h0;
  assign _EVAL_4192 = _EVAL_1064 | _EVAL_915;
  assign _EVAL_2485 = _EVAL_4192 == 1'h0;
  assign _EVAL_240 = _EVAL_888 & 32'h2048;
  assign _EVAL_6082 = _EVAL_240 == 32'h2008;
  assign _EVAL_5449 = _EVAL_4268 & 32'h7c;
  assign _EVAL_5033 = _EVAL_5449 == 32'h24;
  assign _EVAL_294 = _EVAL_4268 & 32'h40000060;
  assign _EVAL_5037 = _EVAL_294 == 32'h40;
  assign _EVAL_5905 = _EVAL_5033 | _EVAL_5037;
  assign _EVAL_5206 = _EVAL_386 & 32'h407f;
  assign _EVAL_333 = _EVAL_4268 & 32'h7e00607f;
  assign _EVAL_6032 = _EVAL_4882 & 32'h62003010;
  assign _EVAL_3769 = _EVAL_4743 & 32'h80000010;
  assign _EVAL_5641 = _EVAL_4268 & 32'h90000034;
  assign _EVAL_3130 = _EVAL_1242 == 32'h30200073;
  assign _EVAL_3892 = _EVAL_2344 == 32'h20;
  assign _EVAL_3057 = _EVAL_1978 & 32'h34;
  assign _EVAL_5733 = _EVAL_3057 == 32'h20;
  assign _EVAL_1668 = _EVAL_3892 | _EVAL_5733;
  assign _EVAL_3172 = _EVAL_5813 & 32'h80000010;
  assign _EVAL_5002 = _EVAL_4589 == 32'h0;
  assign _EVAL_1755 = _EVAL_5854 & 32'h60;
  assign _EVAL_4133 = _EVAL_1755 == 32'h0;
  assign _EVAL_1761 = _EVAL_5002 | _EVAL_4133;
  assign _EVAL_4562 = _EVAL_5854 & 32'h50;
  assign _EVAL_5786 = _EVAL_4562 == 32'h0;
  assign _EVAL_4141 = _EVAL_1761 | _EVAL_5786;
  assign _EVAL_4353 = _EVAL_5854 & 32'h44;
  assign _EVAL_4745 = _EVAL_4353 == 32'h4;
  assign _EVAL_4928 = _EVAL_4141 | _EVAL_4745;
  assign _EVAL_530 = _EVAL_5854 & 32'hfff0607f;
  assign _EVAL_3637 = _EVAL_386 & 32'h2000040;
  assign _EVAL_1506 = _EVAL_1978 & 32'h2048;
  assign _EVAL_5719 = _EVAL_1506 == 32'h2008;
  assign _EVAL_493 = _EVAL_1668 | _EVAL_5719;
  assign _EVAL_2640 = _EVAL_1978 & 32'h4003044;
  assign _EVAL_4398 = _EVAL_2640 == 32'h4000040;
  assign _EVAL_375 = _EVAL_493 | _EVAL_4398;
  assign _EVAL_3458 = _EVAL_4702 & 32'h8000040;
  assign _EVAL_4685 = _EVAL_3458 == 32'h8000040;
  assign _EVAL_3706 = _EVAL_3006 & 32'h2050;
  assign _EVAL_5720 = _EVAL_4702 & 32'h28;
  assign _EVAL_5790 = _EVAL_5720 == 32'h28;
  assign _EVAL_5283 = _EVAL_4743 & 32'h64;
  assign _EVAL_4382 = _EVAL_5283 == 32'h0;
  assign _EVAL_4601 = _EVAL_4743 & 32'h50;
  assign _EVAL_1250 = _EVAL_4601 == 32'h10;
  assign _EVAL_4696 = _EVAL_4382 | _EVAL_1250;
  assign _EVAL_2392 = _EVAL_4743 & 32'h2024;
  assign _EVAL_6054 = _EVAL_2392 == 32'h24;
  assign _EVAL_5000 = _EVAL_4696 | _EVAL_6054;
  assign _EVAL_3984 = _EVAL_4743 & 32'h28;
  assign _EVAL_1576 = _EVAL_3984 == 32'h28;
  assign _EVAL_1840 = _EVAL_5000 | _EVAL_1576;
  assign _EVAL_1200 = _EVAL_4743 & 32'h30;
  assign _EVAL_1607 = _EVAL_1200 == 32'h30;
  assign _EVAL_2639 = _EVAL_1840 | _EVAL_1607;
  assign _EVAL_6129 = _EVAL_4743 & 32'h90000010;
  assign _EVAL_5834 = _EVAL_6129 == 32'h80000010;
  assign _EVAL_2900 = _EVAL_2639 | _EVAL_5834;
  assign _EVAL_5863 = _EVAL_1173 & _EVAL_2646;
  assign _EVAL_4089 = _EVAL_5668 | _EVAL_5863;
  assign _EVAL_4558 = _EVAL_4089 == _EVAL_379;
  assign _EVAL_1437 = _EVAL_1173 & _EVAL_2874;
  assign _EVAL_1696 = _EVAL_4914 ? _EVAL_4558 : _EVAL_1437;
  assign _EVAL_5885 = _EVAL_4922 & _EVAL_1696;
  assign _EVAL_352 = _EVAL_2110 & _EVAL_5885;
  assign _EVAL_5302 = _EVAL_3078 & 32'h10000060;
  assign _EVAL_827 = _EVAL_5302 == 32'h10000040;
  assign _EVAL_1269 = _EVAL_3455[12:5];
  assign _EVAL_3854 = _EVAL_1269 != 8'h0;
  assign _EVAL_1920 = _EVAL_5755 ? 1'h1 : _EVAL_3854;
  assign _EVAL_2129 = _EVAL_597 ? 1'h1 : _EVAL_1920;
  assign _EVAL_5993 = _EVAL_1674 ? 1'h1 : _EVAL_2129;
  assign _EVAL_806 = _EVAL_3271 & 32'h28;
  assign _EVAL_1705 = _EVAL_806 == 32'h28;
  assign _EVAL_781 = _EVAL_3455[14];
  assign _EVAL_870 = _EVAL_1074 ? _EVAL_781 : _EVAL_781;
  assign _EVAL_2563 = _EVAL_5926 ? _EVAL_781 : _EVAL_870;
  assign _EVAL_3610 = _EVAL_2970 ? _EVAL_781 : _EVAL_2563;
  assign _EVAL_3253 = _EVAL_2970 ? 1'h0 : _EVAL_3610;
  assign _EVAL_1334 = _EVAL_4268[14];
  assign _EVAL_3328 = _EVAL_2901 ? _EVAL_1334 : _EVAL_1334;
  assign _EVAL_1471 = _EVAL_2378 ? _EVAL_1334 : _EVAL_3328;
  assign _EVAL_2841 = _EVAL_5690 ? _EVAL_1334 : _EVAL_1471;
  assign _EVAL_2521 = _EVAL_5690 ? 1'h0 : _EVAL_2841;
  assign _EVAL_4686 = _EVAL_2666[14];
  assign _EVAL_3050 = _EVAL_2389 == 2'h2;
  assign _EVAL_668 = _EVAL_2389 == 2'h1;
  assign _EVAL_3937 = _EVAL_668 ? _EVAL_4686 : _EVAL_4686;
  assign _EVAL_4570 = _EVAL_3050 ? _EVAL_4686 : _EVAL_3937;
  assign _EVAL_969 = _EVAL_1069 ? _EVAL_4686 : _EVAL_4570;
  assign _EVAL_4461 = _EVAL_5337 ? _EVAL_2521 : _EVAL_969;
  assign _EVAL_5328 = _EVAL_1930 ? _EVAL_3253 : _EVAL_4461;
  assign _EVAL_1262 = _EVAL_4882 & 32'h80000010;
  assign _EVAL_4909 = _EVAL_1262 == 32'h10;
  assign _EVAL_1388 = _EVAL_4909 | _EVAL_360;
  assign _EVAL_3845 = _EVAL_4882 & 32'h40000040;
  assign _EVAL_4047 = _EVAL_3845 == 32'h40;
  assign _EVAL_2611 = _EVAL_1388 | _EVAL_4047;
  assign _EVAL_3690 = _EVAL_4882 & 32'h20000040;
  assign _EVAL_2305 = _EVAL_3690 == 32'h40;
  assign _EVAL_1605 = _EVAL_2611 | _EVAL_2305;
  assign _EVAL_2919 = _EVAL_888 & 32'h2024;
  assign _EVAL_2258 = _EVAL_2919 == 32'h24;
  assign _EVAL_4017 = _EVAL_1978 & 32'h207f;
  assign _EVAL_2384 = _EVAL_4017 == 32'h3;
  assign _EVAL_3448 = _EVAL_1978 & 32'h607f;
  assign _EVAL_1414 = _EVAL_3448 == 32'hf;
  assign _EVAL_1499 = _EVAL_2384 | _EVAL_1414;
  assign _EVAL_295 = _EVAL_4366 == 32'h17;
  assign _EVAL_4816 = _EVAL_1499 | _EVAL_295;
  assign _EVAL_5469 = _EVAL_1978 & 32'hfc00007f;
  assign _EVAL_602 = _EVAL_5469 == 32'h33;
  assign _EVAL_905 = _EVAL_4816 | _EVAL_602;
  assign _EVAL_2102 = _EVAL_1978 & 32'hbe00707f;
  assign _EVAL_2346 = _EVAL_2102 == 32'h33;
  assign _EVAL_2625 = _EVAL_905 | _EVAL_2346;
  assign _EVAL_823 = _EVAL_1978 & 32'h6000073;
  assign _EVAL_1768 = _EVAL_823 == 32'h43;
  assign _EVAL_2552 = _EVAL_2625 | _EVAL_1768;
  assign _EVAL_1672 = _EVAL_1978 & 32'he600007f;
  assign _EVAL_4229 = _EVAL_1672 == 32'h53;
  assign _EVAL_1243 = _EVAL_2552 | _EVAL_4229;
  assign _EVAL_3099 = _EVAL_1978 & 32'h707b;
  assign _EVAL_1843 = _EVAL_3099 == 32'h63;
  assign _EVAL_4580 = _EVAL_1243 | _EVAL_1843;
  assign _EVAL_4627 = _EVAL_1978 & 32'h7f;
  assign _EVAL_5001 = _EVAL_4627 == 32'h6f;
  assign _EVAL_999 = _EVAL_4580 | _EVAL_5001;
  assign _EVAL_3472 = _EVAL_1978 & 32'hffefffff;
  assign _EVAL_274 = _EVAL_3472 == 32'h73;
  assign _EVAL_2923 = _EVAL_999 | _EVAL_274;
  assign _EVAL_5828 = _EVAL_1978 & 32'hfe00305f;
  assign _EVAL_4054 = _EVAL_5828 == 32'h1013;
  assign _EVAL_4752 = _EVAL_2923 | _EVAL_4054;
  assign _EVAL_924 = _EVAL_1978 & 32'h705b;
  assign _EVAL_253 = _EVAL_924 == 32'h2003;
  assign _EVAL_2885 = _EVAL_4752 | _EVAL_253;
  assign _EVAL_1209 = _EVAL_4017 == 32'h2013;
  assign _EVAL_5003 = _EVAL_2885 | _EVAL_1209;
  assign _EVAL_4487 = _EVAL_1978 & 32'h1800707f;
  assign _EVAL_466 = _EVAL_4487 == 32'h202f;
  assign _EVAL_5649 = _EVAL_5003 | _EVAL_466;
  assign _EVAL_725 = _EVAL_4017 == 32'h2073;
  assign _EVAL_2855 = _EVAL_5649 | _EVAL_725;
  assign _EVAL_4364 = _EVAL_1978 & 32'hbe00705f;
  assign _EVAL_879 = _EVAL_4364 == 32'h5013;
  assign _EVAL_3245 = _EVAL_2855 | _EVAL_879;
  assign _EVAL_2719 = _EVAL_1978 & 32'he800707f;
  assign _EVAL_4769 = _EVAL_2719 == 32'h800202f;
  assign _EVAL_4529 = _EVAL_3245 | _EVAL_4769;
  assign _EVAL_4744 = _EVAL_1978 & 32'hf9f0707f;
  assign _EVAL_2181 = _EVAL_4744 == 32'h1000202f;
  assign _EVAL_3885 = _EVAL_4529 | _EVAL_2181;
  assign _EVAL_2328 = _EVAL_1978 & 32'hdfffffff;
  assign _EVAL_2762 = _EVAL_2328 == 32'h10500073;
  assign _EVAL_4893 = _EVAL_3885 | _EVAL_2762;
  assign _EVAL_1653 = _EVAL_1978 & 32'hf600607f;
  assign _EVAL_1988 = _EVAL_1653 == 32'h20000053;
  assign _EVAL_5981 = _EVAL_4893 | _EVAL_1988;
  assign _EVAL_3386 = _EVAL_3271 & 32'h407f;
  assign _EVAL_3136 = _EVAL_3386 == 32'h4063;
  assign _EVAL_1984 = _EVAL_3455[14:12];
  assign _EVAL_4908 = _EVAL_2039[14:12];
  assign _EVAL_3849 = _EVAL_1242[14:12];
  assign _EVAL_2514 = _EVAL_2164[14:12];
  assign _EVAL_3125 = _EVAL_1074 ? _EVAL_3849 : _EVAL_2514;
  assign _EVAL_4634 = _EVAL_5926 ? _EVAL_4908 : _EVAL_3125;
  assign _EVAL_4698 = _EVAL_2970 ? _EVAL_4908 : _EVAL_4634;
  assign _EVAL_3351 = _EVAL_2970 ? _EVAL_1984 : _EVAL_4698;
  assign _EVAL_2112 = _EVAL_4268[14:12];
  assign _EVAL_5617 = _EVAL_3006[14:12];
  assign _EVAL_5842 = _EVAL_4882[14:12];
  assign _EVAL_1622 = _EVAL_5133[14:12];
  assign _EVAL_3513 = _EVAL_2901 ? _EVAL_5842 : _EVAL_1622;
  assign _EVAL_5806 = _EVAL_2378 ? _EVAL_5617 : _EVAL_3513;
  assign _EVAL_2151 = _EVAL_5690 ? _EVAL_5617 : _EVAL_5806;
  assign _EVAL_4798 = _EVAL_5690 ? _EVAL_2112 : _EVAL_2151;
  assign _EVAL_4608 = _EVAL_1978[14:12];
  assign _EVAL_5935 = _EVAL_1362[14:12];
  assign _EVAL_1977 = _EVAL_3271[14:12];
  assign _EVAL_5858 = _EVAL_668 ? _EVAL_5935 : _EVAL_1977;
  assign _EVAL_4722 = _EVAL_3050 ? _EVAL_4608 : _EVAL_5858;
  assign _EVAL_1486 = _EVAL_1069 ? _EVAL_4608 : _EVAL_4722;
  assign _EVAL_2656 = _EVAL_5337 ? _EVAL_4798 : _EVAL_1486;
  assign _EVAL_1363 = _EVAL_1930 ? _EVAL_3351 : _EVAL_2656;
  assign _EVAL_4262 = _EVAL_1978 & 32'h7c;
  assign _EVAL_4309 = _EVAL_4262 == 32'h24;
  assign _EVAL_1179 = _EVAL_1978 & 32'h40000060;
  assign _EVAL_1475 = _EVAL_1179 == 32'h40;
  assign _EVAL_1297 = _EVAL_4309 | _EVAL_1475;
  assign _EVAL_4126 = _EVAL_1978 & 32'h70;
  assign _EVAL_4329 = _EVAL_4126 == 32'h40;
  assign _EVAL_1040 = _EVAL_1297 | _EVAL_4329;
  assign _EVAL_4932 = _EVAL_1362 & 32'h7c;
  assign _EVAL_5331 = _EVAL_4932 == 32'h24;
  assign _EVAL_2427 = _EVAL_1362 & 32'h40000060;
  assign _EVAL_1450 = _EVAL_2427 == 32'h40;
  assign _EVAL_2566 = _EVAL_5331 | _EVAL_1450;
  assign _EVAL_3468 = _EVAL_1362 & 32'h70;
  assign _EVAL_4770 = _EVAL_3468 == 32'h40;
  assign _EVAL_2120 = _EVAL_2566 | _EVAL_4770;
  assign _EVAL_1921 = _EVAL_3271 & 32'h7c;
  assign _EVAL_4617 = _EVAL_1921 == 32'h24;
  assign _EVAL_1703 = _EVAL_3271 & 32'h40000060;
  assign _EVAL_2433 = _EVAL_1703 == 32'h40;
  assign _EVAL_782 = _EVAL_4617 | _EVAL_2433;
  assign _EVAL_456 = _EVAL_3271 & 32'h70;
  assign _EVAL_1739 = _EVAL_456 == 32'h40;
  assign _EVAL_3207 = _EVAL_782 | _EVAL_1739;
  assign _EVAL_4266 = _EVAL_668 ? _EVAL_2120 : _EVAL_3207;
  assign _EVAL_3224 = _EVAL_3050 ? _EVAL_1040 : _EVAL_4266;
  assign _EVAL_4733 = _EVAL_1069 ? _EVAL_1040 : _EVAL_3224;
  assign _EVAL_2027 = _EVAL_1242 & 32'hfc00007f;
  assign _EVAL_206 = _EVAL_1947 & 32'h306f;
  assign _EVAL_2475 = _EVAL_206 == 32'h1063;
  assign _EVAL_4027 = _EVAL_5133 & 32'h607f;
  assign _EVAL_2166 = _EVAL_3006 & 32'h7c;
  assign _EVAL_2833 = _EVAL_2166 == 32'h24;
  assign _EVAL_4945 = _EVAL_3006 & 32'h40000060;
  assign _EVAL_6063 = _EVAL_4945 == 32'h40;
  assign _EVAL_4524 = _EVAL_2833 | _EVAL_6063;
  assign _EVAL_407 = _EVAL_4524 | _EVAL_3390;
  assign _EVAL_3344 = _EVAL_4882 & 32'h7c;
  assign _EVAL_1698 = _EVAL_3344 == 32'h24;
  assign _EVAL_3432 = _EVAL_4882 & 32'h40000060;
  assign _EVAL_3308 = _EVAL_3432 == 32'h40;
  assign _EVAL_3932 = _EVAL_1698 | _EVAL_3308;
  assign _EVAL_5168 = _EVAL_3932 | _EVAL_2101;
  assign _EVAL_3203 = _EVAL_5133 & 32'h40000060;
  assign _EVAL_2247 = _EVAL_3203 == 32'h40;
  assign _EVAL_5597 = _EVAL_5658 | _EVAL_2247;
  assign _EVAL_1337 = _EVAL_5597 | _EVAL_5949;
  assign _EVAL_1333 = _EVAL_2901 ? _EVAL_5168 : _EVAL_1337;
  assign _EVAL_3198 = _EVAL_2378 ? _EVAL_407 : _EVAL_1333;
  assign _EVAL_3170 = _EVAL_5690 ? _EVAL_407 : _EVAL_3198;
  assign _EVAL_4370 = _EVAL_4743 & 32'h18;
  assign _EVAL_1412 = _EVAL_4370 == 32'h0;
  assign _EVAL_3179 = _EVAL_4743 & 32'h2010;
  assign _EVAL_4546 = _EVAL_3179 == 32'h2000;
  assign _EVAL_2282 = _EVAL_1412 | _EVAL_4546;
  assign _EVAL_1874 = _EVAL_4743 & 32'h8000040;
  assign _EVAL_5204 = _EVAL_1874 == 32'h8000040;
  assign _EVAL_2261 = _EVAL_2282 | _EVAL_5204;
  assign _EVAL_1496 = _EVAL_386 & 32'h18;
  assign _EVAL_4507 = _EVAL_1496 == 32'h0;
  assign _EVAL_3204 = _EVAL_386 & 32'h2010;
  assign _EVAL_3640 = _EVAL_3204 == 32'h2000;
  assign _EVAL_1857 = _EVAL_4507 | _EVAL_3640;
  assign _EVAL_3301 = _EVAL_386 & 32'h8000040;
  assign _EVAL_2428 = _EVAL_3301 == 32'h8000040;
  assign _EVAL_3541 = _EVAL_1857 | _EVAL_2428;
  assign _EVAL_6133 = _EVAL_5952 ? _EVAL_2261 : _EVAL_3541;
  assign _EVAL_2626 = _EVAL_3078 & 32'h44;
  assign _EVAL_4061 = _EVAL_2626 == 32'h0;
  assign _EVAL_4023 = _EVAL_3078 & 32'h4024;
  assign _EVAL_3212 = _EVAL_4023 == 32'h20;
  assign _EVAL_1146 = _EVAL_4061 | _EVAL_3212;
  assign _EVAL_2649 = _EVAL_3415 == 32'h20;
  assign _EVAL_3727 = _EVAL_1146 | _EVAL_2649;
  assign _EVAL_5902 = _EVAL_3078 & 32'h2050;
  assign _EVAL_3517 = _EVAL_5902 == 32'h2000;
  assign _EVAL_1172 = _EVAL_3727 | _EVAL_3517;
  assign _EVAL_1000 = _EVAL_3078 & 32'h90000034;
  assign _EVAL_3896 = _EVAL_1000 == 32'h90000010;
  assign _EVAL_5779 = _EVAL_1172 | _EVAL_3896;
  assign _EVAL_3824 = _EVAL_4702 & 32'h4024;
  assign _EVAL_3305 = _EVAL_3824 == 32'h20;
  assign _EVAL_3879 = _EVAL_4517 | _EVAL_3305;
  assign _EVAL_4181 = _EVAL_4702 & 32'h38;
  assign _EVAL_311 = _EVAL_4181 == 32'h20;
  assign _EVAL_1603 = _EVAL_3879 | _EVAL_311;
  assign _EVAL_4363 = _EVAL_4702 & 32'h2050;
  assign _EVAL_3902 = _EVAL_4363 == 32'h2000;
  assign _EVAL_2302 = _EVAL_1603 | _EVAL_3902;
  assign _EVAL_5881 = _EVAL_4702 & 32'h90000034;
  assign _EVAL_5677 = _EVAL_5881 == 32'h90000010;
  assign _EVAL_561 = _EVAL_2302 | _EVAL_5677;
  assign _EVAL_1149 = _EVAL_5813 & 32'h44;
  assign _EVAL_4838 = _EVAL_1149 == 32'h0;
  assign _EVAL_5796 = _EVAL_5813 & 32'h4024;
  assign _EVAL_1287 = _EVAL_5796 == 32'h20;
  assign _EVAL_5758 = _EVAL_4838 | _EVAL_1287;
  assign _EVAL_4344 = _EVAL_5813 & 32'h38;
  assign _EVAL_2301 = _EVAL_4344 == 32'h20;
  assign _EVAL_4760 = _EVAL_5758 | _EVAL_2301;
  assign _EVAL_3446 = _EVAL_5813 & 32'h2050;
  assign _EVAL_831 = _EVAL_3446 == 32'h2000;
  assign _EVAL_3730 = _EVAL_4760 | _EVAL_831;
  assign _EVAL_2876 = _EVAL_5813 & 32'h90000034;
  assign _EVAL_3617 = _EVAL_2876 == 32'h90000010;
  assign _EVAL_2284 = _EVAL_3730 | _EVAL_3617;
  assign _EVAL_2583 = _EVAL_1947 & 32'h44;
  assign _EVAL_3557 = _EVAL_2583 == 32'h0;
  assign _EVAL_1719 = _EVAL_1947 & 32'h4024;
  assign _EVAL_4839 = _EVAL_1719 == 32'h20;
  assign _EVAL_2091 = _EVAL_3557 | _EVAL_4839;
  assign _EVAL_2794 = _EVAL_1947 & 32'h38;
  assign _EVAL_4166 = _EVAL_2794 == 32'h20;
  assign _EVAL_509 = _EVAL_2091 | _EVAL_4166;
  assign _EVAL_2297 = _EVAL_1947 & 32'h2050;
  assign _EVAL_2932 = _EVAL_2297 == 32'h2000;
  assign _EVAL_2312 = _EVAL_509 | _EVAL_2932;
  assign _EVAL_1153 = _EVAL_1947 & 32'h90000034;
  assign _EVAL_3895 = _EVAL_1153 == 32'h90000010;
  assign _EVAL_5082 = _EVAL_2312 | _EVAL_3895;
  assign _EVAL_5252 = _EVAL_1958 ? _EVAL_2284 : _EVAL_5082;
  assign _EVAL_1922 = _EVAL_4554 ? _EVAL_5779 : _EVAL_5252;
  assign _EVAL_4632 = _EVAL_197 ? _EVAL_5779 : _EVAL_1922;
  assign _EVAL_4356 = _EVAL_197 ? _EVAL_561 : _EVAL_4632;
  assign _EVAL_188 = _EVAL_3271 & 32'h64;
  assign _EVAL_4822 = _EVAL_188 == 32'h0;
  assign _EVAL_4387 = _EVAL_3271 & 32'h50;
  assign _EVAL_3764 = _EVAL_4387 == 32'h10;
  assign _EVAL_3465 = _EVAL_4822 | _EVAL_3764;
  assign _EVAL_2104 = _EVAL_4856 == 32'h24;
  assign _EVAL_3847 = _EVAL_3465 | _EVAL_2104;
  assign _EVAL_3726 = _EVAL_3847 | _EVAL_1705;
  assign _EVAL_1212 = _EVAL_3271 & 32'h30;
  assign _EVAL_3027 = _EVAL_1212 == 32'h30;
  assign _EVAL_2326 = _EVAL_3726 | _EVAL_3027;
  assign _EVAL_5057 = _EVAL_888[11:7];
  assign _EVAL_4574 = _EVAL_3712 ? 1'h1 : _EVAL_5966;
  assign _EVAL_842 = _EVAL_2321 ? 1'h1 : _EVAL_4574;
  assign _EVAL_1120 = _EVAL_5053 ? 1'h1 : _EVAL_842;
  assign _EVAL_2370 = _EVAL_5623 ? 1'h1 : _EVAL_1120;
  assign _EVAL_2115 = _EVAL_2370 == 1'h0;
  assign _EVAL_1567 = _EVAL_4882 & 32'hfff0607f;
  assign _EVAL_1504 = _EVAL_1567 == 32'he0000053;
  assign _EVAL_5500 = _EVAL_1167 | _EVAL_1504;
  assign _EVAL_1282 = _EVAL_4882 & 32'heff0707f;
  assign _EVAL_4550 = _EVAL_1282 == 32'he0000053;
  assign _EVAL_4026 = _EVAL_5500 | _EVAL_4550;
  assign _EVAL_5732 = _EVAL_4882 & 32'hffd07fff;
  assign _EVAL_2441 = _EVAL_5732 == 32'hfc000073;
  assign _EVAL_807 = _EVAL_4026 | _EVAL_2441;
  assign _EVAL_3520 = _EVAL_4882 & 32'h306f;
  assign _EVAL_754 = _EVAL_3520 == 32'h1063;
  assign _EVAL_1915 = _EVAL_807 | _EVAL_754;
  assign _EVAL_1925 = _EVAL_4882 & 32'h407f;
  assign _EVAL_1729 = _EVAL_1925 == 32'h4063;
  assign _EVAL_2056 = _EVAL_1915 | _EVAL_1729;
  assign _EVAL_5354 = _EVAL_4882 & 32'h605f;
  assign _EVAL_3559 = _EVAL_5354 == 32'h3;
  assign _EVAL_6005 = _EVAL_2056 | _EVAL_3559;
  assign _EVAL_3978 = _EVAL_3520 == 32'h3;
  assign _EVAL_4041 = _EVAL_6005 | _EVAL_3978;
  assign _EVAL_1899 = _EVAL_2115 ? 1'h0 : _EVAL_4041;
  assign _EVAL_632 = _EVAL_4268[12:5];
  assign _EVAL_5213 = _EVAL_632 != 8'h0;
  assign _EVAL_1684 = _EVAL_5573 ? 1'h1 : _EVAL_5213;
  assign _EVAL_250 = _EVAL_4038 ? 1'h1 : _EVAL_1684;
  assign _EVAL_4242 = _EVAL_1743 ? 1'h1 : _EVAL_250;
  assign _EVAL_5693 = _EVAL_3712 ? 1'h1 : _EVAL_4242;
  assign _EVAL_5178 = _EVAL_2321 ? 1'h1 : _EVAL_5693;
  assign _EVAL_1564 = _EVAL_5053 ? 1'h1 : _EVAL_5178;
  assign _EVAL_1825 = _EVAL_5623 ? 1'h1 : _EVAL_1564;
  assign _EVAL_1601 = _EVAL_1825 == 1'h0;
  assign _EVAL_1571 = _EVAL_5133 & 32'h207f;
  assign _EVAL_4458 = _EVAL_1571 == 32'h3;
  assign _EVAL_5402 = _EVAL_4027 == 32'hf;
  assign _EVAL_3142 = _EVAL_4458 | _EVAL_5402;
  assign _EVAL_457 = _EVAL_5133 & 32'h5f;
  assign _EVAL_2487 = _EVAL_457 == 32'h17;
  assign _EVAL_972 = _EVAL_3142 | _EVAL_2487;
  assign _EVAL_4553 = _EVAL_5133 & 32'hfc00007f;
  assign _EVAL_1997 = _EVAL_4553 == 32'h33;
  assign _EVAL_898 = _EVAL_972 | _EVAL_1997;
  assign _EVAL_5196 = _EVAL_5133 & 32'hbe00707f;
  assign _EVAL_5448 = _EVAL_5196 == 32'h33;
  assign _EVAL_5075 = _EVAL_898 | _EVAL_5448;
  assign _EVAL_2084 = _EVAL_5133 & 32'h6000073;
  assign _EVAL_1979 = _EVAL_2084 == 32'h43;
  assign _EVAL_2467 = _EVAL_5075 | _EVAL_1979;
  assign _EVAL_2904 = _EVAL_5133 & 32'he600007f;
  assign _EVAL_6021 = _EVAL_2904 == 32'h53;
  assign _EVAL_4436 = _EVAL_2467 | _EVAL_6021;
  assign _EVAL_2347 = _EVAL_5133 & 32'h707b;
  assign _EVAL_1894 = _EVAL_2347 == 32'h63;
  assign _EVAL_1411 = _EVAL_4436 | _EVAL_1894;
  assign _EVAL_2232 = _EVAL_5133 & 32'h7f;
  assign _EVAL_1439 = _EVAL_2232 == 32'h6f;
  assign _EVAL_1423 = _EVAL_1411 | _EVAL_1439;
  assign _EVAL_5071 = _EVAL_5133 & 32'hffefffff;
  assign _EVAL_875 = _EVAL_5071 == 32'h73;
  assign _EVAL_1849 = _EVAL_1423 | _EVAL_875;
  assign _EVAL_3580 = _EVAL_5133 & 32'hfe00305f;
  assign _EVAL_6038 = _EVAL_3580 == 32'h1013;
  assign _EVAL_5625 = _EVAL_1849 | _EVAL_6038;
  assign _EVAL_3101 = _EVAL_5133 & 32'h705b;
  assign _EVAL_3578 = _EVAL_3101 == 32'h2003;
  assign _EVAL_3702 = _EVAL_5625 | _EVAL_3578;
  assign _EVAL_1549 = _EVAL_1571 == 32'h2013;
  assign _EVAL_2554 = _EVAL_3702 | _EVAL_1549;
  assign _EVAL_3360 = _EVAL_5133 & 32'h1800707f;
  assign _EVAL_3750 = _EVAL_3360 == 32'h202f;
  assign _EVAL_2846 = _EVAL_2554 | _EVAL_3750;
  assign _EVAL_1016 = _EVAL_1571 == 32'h2073;
  assign _EVAL_4537 = _EVAL_2846 | _EVAL_1016;
  assign _EVAL_5632 = _EVAL_5133 & 32'hbe00705f;
  assign _EVAL_6139 = _EVAL_5632 == 32'h5013;
  assign _EVAL_4081 = _EVAL_4537 | _EVAL_6139;
  assign _EVAL_2332 = _EVAL_5133 & 32'he800707f;
  assign _EVAL_3903 = _EVAL_2332 == 32'h800202f;
  assign _EVAL_5017 = _EVAL_4081 | _EVAL_3903;
  assign _EVAL_1788 = _EVAL_5133 & 32'hf9f0707f;
  assign _EVAL_4014 = _EVAL_1788 == 32'h1000202f;
  assign _EVAL_1581 = _EVAL_5017 | _EVAL_4014;
  assign _EVAL_3999 = _EVAL_5133 & 32'hdfffffff;
  assign _EVAL_4717 = _EVAL_3999 == 32'h10500073;
  assign _EVAL_820 = _EVAL_1581 | _EVAL_4717;
  assign _EVAL_874 = _EVAL_5133 & 32'hf600607f;
  assign _EVAL_4763 = _EVAL_874 == 32'h20000053;
  assign _EVAL_1798 = _EVAL_820 | _EVAL_4763;
  assign _EVAL_494 = _EVAL_5133 & 32'h7e00607f;
  assign _EVAL_1929 = _EVAL_494 == 32'h20000053;
  assign _EVAL_4153 = _EVAL_1798 | _EVAL_1929;
  assign _EVAL_1331 = _EVAL_5133 & 32'h7e00507f;
  assign _EVAL_1249 = _EVAL_1331 == 32'h20000053;
  assign _EVAL_4037 = _EVAL_4153 | _EVAL_1249;
  assign _EVAL_4418 = _EVAL_5133 == 32'h30200073;
  assign _EVAL_5064 = _EVAL_4037 | _EVAL_4418;
  assign _EVAL_4119 = _EVAL_5133 & 32'hfff0007f;
  assign _EVAL_1721 = _EVAL_4119 == 32'h58000053;
  assign _EVAL_903 = _EVAL_5064 | _EVAL_1721;
  assign _EVAL_1394 = _EVAL_5133 == 32'h7b200073;
  assign _EVAL_3233 = _EVAL_903 | _EVAL_1394;
  assign _EVAL_3749 = _EVAL_5133 & 32'hefe0007f;
  assign _EVAL_3965 = _EVAL_3749 == 32'hc0000053;
  assign _EVAL_3622 = _EVAL_3233 | _EVAL_3965;
  assign _EVAL_1557 = _EVAL_5133 & 32'hfff0607f;
  assign _EVAL_3662 = _EVAL_1557 == 32'he0000053;
  assign _EVAL_3275 = _EVAL_3622 | _EVAL_3662;
  assign _EVAL_5555 = _EVAL_5133 & 32'heff0707f;
  assign _EVAL_5692 = _EVAL_5555 == 32'he0000053;
  assign _EVAL_5163 = _EVAL_3275 | _EVAL_5692;
  assign _EVAL_1953 = _EVAL_2460 == 32'hfc000073;
  assign _EVAL_2009 = _EVAL_5163 | _EVAL_1953;
  assign _EVAL_560 = _EVAL_4806 == 32'h1063;
  assign _EVAL_5816 = _EVAL_2009 | _EVAL_560;
  assign _EVAL_2579 = _EVAL_5133 & 32'h407f;
  assign _EVAL_2222 = _EVAL_2579 == 32'h4063;
  assign _EVAL_3543 = _EVAL_5816 | _EVAL_2222;
  assign _EVAL_5401 = _EVAL_5133 & 32'h605f;
  assign _EVAL_5958 = _EVAL_5401 == 32'h3;
  assign _EVAL_4911 = _EVAL_3543 | _EVAL_5958;
  assign _EVAL_3090 = _EVAL_4911 | _EVAL_6045;
  assign _EVAL_1751 = _EVAL_1601 ? 1'h0 : _EVAL_3090;
  assign _EVAL_5894 = _EVAL_2901 ? _EVAL_1899 : _EVAL_1751;
  assign _EVAL_520 = _EVAL_4702 & 32'h306f;
  assign _EVAL_1990 = _EVAL_520 == 32'h3;
  assign _EVAL_320 = _EVAL_5386[14];
  assign _EVAL_4289 = _EVAL_5952 ? _EVAL_320 : _EVAL_320;
  assign _EVAL_1881 = _EVAL_3570 ? _EVAL_320 : _EVAL_4289;
  assign _EVAL_1175 = _EVAL_5833 ? _EVAL_320 : _EVAL_1881;
  assign _EVAL_6050 = _EVAL_5833 ? 1'h0 : _EVAL_1175;
  assign _EVAL_5729 = _EVAL_5854 & 32'h4003044;
  assign _EVAL_656 = _EVAL_5729 == 32'h4000040;
  assign _EVAL_805 = {_EVAL_2007,_EVAL_2075};
  assign _EVAL_6046 = _EVAL_805 != 12'h0;
  assign _EVAL_2609 = _EVAL_1674 ? _EVAL_6046 : 1'h1;
  assign _EVAL_1142 = _EVAL_936 ? 1'h1 : _EVAL_2609;
  assign _EVAL_640 = _EVAL_453 ? 1'h1 : _EVAL_1142;
  assign _EVAL_3355 = _EVAL_2288 ? 1'h1 : _EVAL_640;
  assign _EVAL_800 = _EVAL_4669 ? 1'h1 : _EVAL_3355;
  assign _EVAL_5563 = _EVAL_800 == 1'h0;
  assign _EVAL_4687 = _EVAL_4268 & 32'h2000040;
  assign _EVAL_576 = _EVAL_4687 == 32'h0;
  assign _EVAL_4937 = _EVAL_4268 & 32'h60;
  assign _EVAL_5812 = _EVAL_4937 == 32'h0;
  assign _EVAL_1532 = _EVAL_576 | _EVAL_5812;
  assign _EVAL_4592 = _EVAL_2696 == 32'h0;
  assign _EVAL_4641 = _EVAL_1532 | _EVAL_4592;
  assign _EVAL_1718 = _EVAL_4268 & 32'h44;
  assign _EVAL_4001 = _EVAL_1718 == 32'h4;
  assign _EVAL_5697 = _EVAL_4641 | _EVAL_4001;
  assign _EVAL_2654 = _EVAL_888 & 32'h40000060;
  assign _EVAL_776 = _EVAL_2654 == 32'h40;
  assign _EVAL_562 = _EVAL_5020 == 32'h10000040;
  assign _EVAL_2017 = _EVAL_2164 == 32'h30200073;
  assign _EVAL_1366 = _EVAL_2362 | _EVAL_2017;
  assign _EVAL_3418 = _EVAL_2164 & 32'hfff0007f;
  assign _EVAL_5568 = _EVAL_3418 == 32'h58000053;
  assign _EVAL_5453 = _EVAL_1366 | _EVAL_5568;
  assign _EVAL_4306 = _EVAL_936 ? 1'h1 : _EVAL_5993;
  assign _EVAL_865 = _EVAL_5854 & 32'h80000010;
  assign _EVAL_3781 = _EVAL_865 == 32'h10;
  assign _EVAL_164 = _EVAL_4562 == 32'h10;
  assign _EVAL_5548 = _EVAL_3781 | _EVAL_164;
  assign _EVAL_4427 = _EVAL_5854 & 32'h40000040;
  assign _EVAL_5478 = _EVAL_4427 == 32'h40;
  assign _EVAL_963 = _EVAL_5548 | _EVAL_5478;
  assign _EVAL_1035 = _EVAL_5854 & 32'h20000040;
  assign _EVAL_4661 = _EVAL_1035 == 32'h40;
  assign _EVAL_2880 = _EVAL_963 | _EVAL_4661;
  assign _EVAL_5857 = _EVAL_5813 & 32'h8000040;
  assign _EVAL_2106 = _EVAL_5857 == 32'h8000040;
  assign _EVAL_3338 = _EVAL_4702 & 32'h80000010;
  assign _EVAL_5829 = _EVAL_3338 == 32'h10;
  assign _EVAL_2170 = _EVAL_1458 == 32'h10;
  assign _EVAL_1789 = _EVAL_5829 | _EVAL_2170;
  assign _EVAL_1614 = _EVAL_4702 & 32'h40000040;
  assign _EVAL_4070 = _EVAL_1614 == 32'h40;
  assign _EVAL_1994 = _EVAL_1789 | _EVAL_4070;
  assign _EVAL_1113 = _EVAL_4702 & 32'h20000040;
  assign _EVAL_1967 = _EVAL_1113 == 32'h40;
  assign _EVAL_810 = _EVAL_1994 | _EVAL_1967;
  assign _EVAL_5208 = _EVAL_1458 == 32'h40;
  assign _EVAL_5909 = _EVAL_810 | _EVAL_5208;
  assign _EVAL_1982 = _EVAL_1451 & _EVAL_979;
  assign _EVAL_1325 = _EVAL_5062 | _EVAL_1982;
  assign _EVAL_3623 = _EVAL_1325 == _EVAL_1969;
  assign _EVAL_4542 = _EVAL_5854 & 32'h207f;
  assign _EVAL_1876 = _EVAL_4542 == 32'h3;
  assign _EVAL_5109 = _EVAL_5854 & 32'h607f;
  assign _EVAL_1816 = _EVAL_5109 == 32'hf;
  assign _EVAL_3285 = _EVAL_1876 | _EVAL_1816;
  assign _EVAL_544 = _EVAL_5854 & 32'h5f;
  assign _EVAL_1811 = _EVAL_544 == 32'h17;
  assign _EVAL_4480 = _EVAL_3285 | _EVAL_1811;
  assign _EVAL_6096 = _EVAL_5854 & 32'hfc00007f;
  assign _EVAL_1382 = _EVAL_6096 == 32'h33;
  assign _EVAL_1381 = _EVAL_4480 | _EVAL_1382;
  assign _EVAL_5314 = _EVAL_5854 & 32'hbe00707f;
  assign _EVAL_3149 = _EVAL_5314 == 32'h33;
  assign _EVAL_2289 = _EVAL_1381 | _EVAL_3149;
  assign _EVAL_5195 = _EVAL_5854 & 32'h6000073;
  assign _EVAL_5794 = _EVAL_5195 == 32'h43;
  assign _EVAL_3315 = _EVAL_2289 | _EVAL_5794;
  assign _EVAL_4740 = _EVAL_5854 & 32'he600007f;
  assign _EVAL_3579 = _EVAL_4740 == 32'h53;
  assign _EVAL_1780 = _EVAL_3315 | _EVAL_3579;
  assign _EVAL_1600 = _EVAL_5854 & 32'h707b;
  assign _EVAL_214 = _EVAL_1600 == 32'h63;
  assign _EVAL_1026 = _EVAL_1780 | _EVAL_214;
  assign _EVAL_501 = _EVAL_5854 & 32'h7f;
  assign _EVAL_5817 = _EVAL_501 == 32'h6f;
  assign _EVAL_3908 = _EVAL_1026 | _EVAL_5817;
  assign _EVAL_1951 = _EVAL_5854 & 32'hffefffff;
  assign _EVAL_1795 = _EVAL_1951 == 32'h73;
  assign _EVAL_3228 = _EVAL_3908 | _EVAL_1795;
  assign _EVAL_5065 = _EVAL_5854 & 32'hfe00305f;
  assign _EVAL_703 = _EVAL_5065 == 32'h1013;
  assign _EVAL_1535 = _EVAL_3228 | _EVAL_703;
  assign _EVAL_3306 = _EVAL_5854 & 32'h705b;
  assign _EVAL_5007 = _EVAL_3306 == 32'h2003;
  assign _EVAL_3187 = _EVAL_1535 | _EVAL_5007;
  assign _EVAL_1123 = _EVAL_4542 == 32'h2013;
  assign _EVAL_2262 = _EVAL_3187 | _EVAL_1123;
  assign _EVAL_4078 = _EVAL_5854 & 32'h1800707f;
  assign _EVAL_1812 = _EVAL_4078 == 32'h202f;
  assign _EVAL_4926 = _EVAL_2262 | _EVAL_1812;
  assign _EVAL_5511 = _EVAL_4542 == 32'h2073;
  assign _EVAL_3837 = _EVAL_4926 | _EVAL_5511;
  assign _EVAL_4042 = _EVAL_5854 & 32'hbe00705f;
  assign _EVAL_2665 = _EVAL_4042 == 32'h5013;
  assign _EVAL_2182 = _EVAL_3837 | _EVAL_2665;
  assign _EVAL_4385 = _EVAL_5854 & 32'he800707f;
  assign _EVAL_2292 = _EVAL_4385 == 32'h800202f;
  assign _EVAL_3738 = _EVAL_2182 | _EVAL_2292;
  assign _EVAL_4080 = _EVAL_5854 & 32'hf9f0707f;
  assign _EVAL_1246 = _EVAL_4080 == 32'h1000202f;
  assign _EVAL_1892 = _EVAL_3738 | _EVAL_1246;
  assign _EVAL_2987 = _EVAL_1242 & 32'hfff0607f;
  assign _EVAL_2006 = _EVAL_2987 == 32'he0000053;
  assign _EVAL_1980 = _EVAL_100 == 3'h0;
  assign _EVAL_2250 = {_EVAL_1980,_EVAL_100};
  assign _EVAL_3461 = _EVAL_2250[3:1];
  assign _EVAL_919 = _EVAL_5337 ? 2'h2 : 2'h3;
  assign _EVAL_4832 = _EVAL_1930 ? 2'h1 : _EVAL_919;
  assign _EVAL_2822 = _EVAL_1226 ? 2'h0 : _EVAL_4832;
  assign _EVAL_858 = {_EVAL_2822, 1'h0};
  assign _EVAL_3083 = _EVAL_5311 & 32'h3c;
  assign _EVAL_4088 = _EVAL_3083 == 32'h4;
  assign _EVAL_2260 = {_EVAL_815,_EVAL_372,_EVAL_3526,_EVAL_5165};
  assign _EVAL_4577 = _EVAL_2260 != 4'h0;
  assign _EVAL_5600 = _EVAL_4577 | _EVAL_3659;
  assign _EVAL_2086 = _EVAL_2357 == 1'h0;
  assign _EVAL_5417 = _EVAL_527 == 1'h0;
  assign _EVAL_1904 = _EVAL_1365 ? _EVAL_5417 : _EVAL_5164;
  assign _EVAL_1114 = _EVAL_3955 ? _EVAL_2086 : _EVAL_1904;
  assign _EVAL_5217 = _EVAL_5454 ? _EVAL_5787 : 1'h0;
  assign _EVAL_4758 = _EVAL_6001 ? _EVAL_1015 : _EVAL_5217;
  assign _EVAL_964 = _EVAL_409 ? _EVAL_5417 : _EVAL_4758;
  assign _EVAL_5918 = _EVAL_2917 ? _EVAL_2086 : _EVAL_964;
  assign _EVAL_2526 = _EVAL_5024 ? _EVAL_5787 : 1'h0;
  assign _EVAL_3544 = _EVAL_5135 ? _EVAL_1015 : _EVAL_2526;
  assign _EVAL_5298 = _EVAL_3870 ? _EVAL_5417 : _EVAL_3544;
  assign _EVAL_2245 = _EVAL_5373 ? _EVAL_2086 : _EVAL_5298;
  assign _EVAL_965 = _EVAL_726 ? _EVAL_5787 : 1'h0;
  assign _EVAL_3376 = _EVAL_1826 ? _EVAL_1015 : _EVAL_965;
  assign _EVAL_2645 = _EVAL_3070 ? _EVAL_5417 : _EVAL_3376;
  assign _EVAL_4879 = _EVAL_4716 ? _EVAL_2086 : _EVAL_2645;
  assign _EVAL_1330 = {_EVAL_1114,_EVAL_5918,_EVAL_2245,_EVAL_4879};
  assign _EVAL_5788 = _EVAL_304[0];
  assign _EVAL_1299 = _EVAL_304[1];
  assign _EVAL_2956 = _EVAL_304[2];
  assign _EVAL_3196 = _EVAL_304[3];
  assign _EVAL_1809 = _EVAL_3196 ? 4'h8 : 4'h0;
  assign _EVAL_2031 = _EVAL_2956 ? 4'h4 : _EVAL_1809;
  assign _EVAL_4375 = _EVAL_1299 ? 4'h2 : _EVAL_2031;
  assign _EVAL_4170 = _EVAL_5788 ? 4'h1 : _EVAL_4375;
  assign _EVAL_4984 = _EVAL_5994 ? 4'h0 : _EVAL_4170;
  assign _EVAL_5671 = _EVAL_1330 & _EVAL_4984;
  assign _EVAL_5588 = _EVAL_5671 != 4'h0;
  assign _EVAL_4426 = _EVAL_5600 ? _EVAL_3526 : _EVAL_5588;
  assign _EVAL_4087 = _EVAL_4702 & 32'h18;
  assign _EVAL_5282 = _EVAL_3455[31:25];
  assign _EVAL_515 = _EVAL_2164 & 32'h306f;
  assign _EVAL_5631 = _EVAL_515 == 32'h1063;
  assign _EVAL_4741 = _EVAL_4268 & 32'h80000010;
  assign _EVAL_6023 = _EVAL_4741 == 32'h10;
  assign _EVAL_2602 = _EVAL_6023 | _EVAL_426;
  assign _EVAL_6016 = _EVAL_3417 == 32'h40;
  assign _EVAL_590 = _EVAL_2602 | _EVAL_6016;
  assign _EVAL_292 = _EVAL_5854 & 32'h28;
  assign _EVAL_2387 = _EVAL_1947 & 32'h30;
  assign _EVAL_5882 = _EVAL_2387 == 32'h30;
  assign _EVAL_3186 = _EVAL_4268 & 32'h207f;
  assign _EVAL_161 = _EVAL_3186 == 32'h3;
  assign _EVAL_4066 = _EVAL_4268 & 32'h607f;
  assign _EVAL_989 = _EVAL_4066 == 32'hf;
  assign _EVAL_4175 = _EVAL_161 | _EVAL_989;
  assign _EVAL_3247 = _EVAL_4268 & 32'h5f;
  assign _EVAL_2693 = _EVAL_3247 == 32'h17;
  assign _EVAL_1129 = _EVAL_4175 | _EVAL_2693;
  assign _EVAL_5166 = _EVAL_4268 & 32'hfc00007f;
  assign _EVAL_310 = _EVAL_5166 == 32'h33;
  assign _EVAL_961 = _EVAL_1129 | _EVAL_310;
  assign _EVAL_2206 = _EVAL_4268 & 32'hbe00707f;
  assign _EVAL_2264 = _EVAL_2206 == 32'h33;
  assign _EVAL_223 = _EVAL_961 | _EVAL_2264;
  assign _EVAL_3612 = _EVAL_4268 & 32'h6000073;
  assign _EVAL_2584 = _EVAL_3612 == 32'h43;
  assign _EVAL_3327 = _EVAL_223 | _EVAL_2584;
  assign _EVAL_5376 = _EVAL_4268 & 32'he600007f;
  assign _EVAL_1409 = _EVAL_5376 == 32'h53;
  assign _EVAL_5512 = _EVAL_3327 | _EVAL_1409;
  assign _EVAL_2773 = _EVAL_4268 & 32'h707b;
  assign _EVAL_1888 = _EVAL_2773 == 32'h63;
  assign _EVAL_1617 = _EVAL_5512 | _EVAL_1888;
  assign _EVAL_678 = _EVAL_4268 & 32'h7f;
  assign _EVAL_3281 = _EVAL_678 == 32'h6f;
  assign _EVAL_3284 = _EVAL_1617 | _EVAL_3281;
  assign _EVAL_6010 = _EVAL_4268 & 32'hffefffff;
  assign _EVAL_1837 = _EVAL_6010 == 32'h73;
  assign _EVAL_5835 = _EVAL_3284 | _EVAL_1837;
  assign _EVAL_2249 = _EVAL_3255 == 32'h1013;
  assign _EVAL_3333 = _EVAL_5835 | _EVAL_2249;
  assign _EVAL_5197 = _EVAL_4268 & 32'h705b;
  assign _EVAL_3147 = _EVAL_5197 == 32'h2003;
  assign _EVAL_1734 = _EVAL_3333 | _EVAL_3147;
  assign _EVAL_1611 = _EVAL_3186 == 32'h2013;
  assign _EVAL_3393 = _EVAL_1734 | _EVAL_1611;
  assign _EVAL_408 = _EVAL_4268 & 32'h1800707f;
  assign _EVAL_3695 = _EVAL_408 == 32'h202f;
  assign _EVAL_783 = _EVAL_3393 | _EVAL_3695;
  assign _EVAL_1474 = _EVAL_3186 == 32'h2073;
  assign _EVAL_1949 = _EVAL_783 | _EVAL_1474;
  assign _EVAL_5717 = _EVAL_1949 | _EVAL_2208;
  assign _EVAL_6121 = _EVAL_4268 & 32'he800707f;
  assign _EVAL_2542 = _EVAL_6121 == 32'h800202f;
  assign _EVAL_2948 = _EVAL_5717 | _EVAL_2542;
  assign _EVAL_3930 = _EVAL_4268 & 32'hf9f0707f;
  assign _EVAL_3995 = _EVAL_3930 == 32'h1000202f;
  assign _EVAL_750 = _EVAL_2948 | _EVAL_3995;
  assign _EVAL_5209 = _EVAL_4268 & 32'hdfffffff;
  assign _EVAL_420 = _EVAL_5209 == 32'h10500073;
  assign _EVAL_1082 = _EVAL_750 | _EVAL_420;
  assign _EVAL_1993 = _EVAL_4268 & 32'hf600607f;
  assign _EVAL_3454 = _EVAL_1993 == 32'h20000053;
  assign _EVAL_1216 = _EVAL_1082 | _EVAL_3454;
  assign _EVAL_2401 = _EVAL_333 == 32'h20000053;
  assign _EVAL_1245 = _EVAL_1216 | _EVAL_2401;
  assign _EVAL_1502 = _EVAL_4268 & 32'h7e00507f;
  assign _EVAL_2077 = _EVAL_1502 == 32'h20000053;
  assign _EVAL_2750 = _EVAL_1245 | _EVAL_2077;
  assign _EVAL_5351 = _EVAL_4268 == 32'h30200073;
  assign _EVAL_2972 = _EVAL_2750 | _EVAL_5351;
  assign _EVAL_981 = _EVAL_4268 & 32'hfff0007f;
  assign _EVAL_3667 = _EVAL_981 == 32'h58000053;
  assign _EVAL_6008 = _EVAL_2972 | _EVAL_3667;
  assign _EVAL_1030 = _EVAL_4268 == 32'h7b200073;
  assign _EVAL_4201 = _EVAL_6008 | _EVAL_1030;
  assign _EVAL_2891 = _EVAL_3078 & 32'h64;
  assign _EVAL_3673 = _EVAL_2891 == 32'h20;
  assign _EVAL_4581 = _EVAL_3078 & 32'h34;
  assign _EVAL_2999 = _EVAL_4581 == 32'h20;
  assign _EVAL_5063 = _EVAL_3673 | _EVAL_2999;
  assign _EVAL_1656 = _EVAL_3078 & 32'h2048;
  assign _EVAL_3707 = _EVAL_1656 == 32'h2008;
  assign _EVAL_3363 = _EVAL_5063 | _EVAL_3707;
  assign _EVAL_3202 = _EVAL_3078 & 32'h4003044;
  assign _EVAL_670 = _EVAL_3202 == 32'h4000040;
  assign _EVAL_3459 = _EVAL_3363 | _EVAL_670;
  assign _EVAL_3168 = _EVAL_888 & 32'h4003044;
  assign _EVAL_219 = _EVAL_888 & 32'h2040;
  assign _EVAL_1023 = _EVAL_3078 & 32'h605f;
  assign _EVAL_2008 = _EVAL_3659 ? _EVAL_717 : _EVAL_127;
  assign _EVAL_3682 = _EVAL_3271 & 32'h44;
  assign _EVAL_5567 = _EVAL_3682 == 32'h0;
  assign _EVAL_1645 = _EVAL_3271 & 32'h4024;
  assign _EVAL_1688 = _EVAL_1645 == 32'h20;
  assign _EVAL_4483 = _EVAL_5567 | _EVAL_1688;
  assign _EVAL_3163 = _EVAL_1362 & 32'h34;
  assign _EVAL_4642 = _EVAL_3006 & 32'h306f;
  assign _EVAL_1284 = _EVAL_4642 == 32'h3;
  assign _EVAL_5667 = _EVAL_2110 | _EVAL_2093;
  assign _EVAL_5847 = _EVAL_4702 & 32'h605f;
  assign _EVAL_6123 = _EVAL_1362 & 32'h18;
  assign _EVAL_1917 = _EVAL_6123 == 32'h0;
  assign _EVAL_587 = _EVAL_1362 & 32'h2010;
  assign _EVAL_4640 = _EVAL_587 == 32'h2000;
  assign _EVAL_3691 = _EVAL_1917 | _EVAL_4640;
  assign _EVAL_2909 = _EVAL_1362 & 32'h8000040;
  assign _EVAL_4525 = _EVAL_2909 == 32'h8000040;
  assign _EVAL_4670 = _EVAL_3691 | _EVAL_4525;
  assign _EVAL_3759 = _EVAL_3271 & 32'h18;
  assign _EVAL_1032 = _EVAL_3759 == 32'h0;
  assign _EVAL_3068 = _EVAL_3271 & 32'h2010;
  assign _EVAL_5339 = _EVAL_3068 == 32'h2000;
  assign _EVAL_3037 = _EVAL_1032 | _EVAL_5339;
  assign _EVAL_1440 = _EVAL_3271 & 32'h8000040;
  assign _EVAL_4457 = _EVAL_1440 == 32'h8000040;
  assign _EVAL_4072 = _EVAL_3037 | _EVAL_4457;
  assign _EVAL_3611 = _EVAL_668 ? _EVAL_4670 : _EVAL_4072;
  assign _EVAL_4161 = _EVAL_4562 == 32'h40;
  assign _EVAL_2856 = _EVAL_2880 | _EVAL_4161;
  assign _EVAL_5795 = _EVAL_1242 & 32'hbe00705f;
  assign _EVAL_2253 = _EVAL_2039 & 32'h3c;
  assign _EVAL_1716 = _EVAL_2253 == 32'h4;
  assign _EVAL_4825 = _EVAL_888 & 32'h10000060;
  assign _EVAL_2973 = _EVAL_4825 == 32'h40;
  assign _EVAL_2647 = _EVAL_3271 & 32'h38;
  assign _EVAL_4316 = _EVAL_2647 == 32'h20;
  assign _EVAL_5285 = _EVAL_4483 | _EVAL_4316;
  assign _EVAL_2955 = _EVAL_3271 & 32'h2050;
  assign _EVAL_5011 = _EVAL_2955 == 32'h2000;
  assign _EVAL_4974 = _EVAL_5285 | _EVAL_5011;
  assign _EVAL_3480 = _EVAL_5854 & 32'h7c;
  assign _EVAL_4853 = _EVAL_3480 == 32'h24;
  assign _EVAL_4963 = _EVAL_5854 & 32'h40000060;
  assign _EVAL_3131 = _EVAL_4963 == 32'h40;
  assign _EVAL_2816 = _EVAL_4853 | _EVAL_3131;
  assign _EVAL_2610 = _EVAL_5813 & 32'h7c;
  assign _EVAL_3875 = _EVAL_5133 & 32'h44;
  assign _EVAL_5102 = _EVAL_3875 == 32'h0;
  assign _EVAL_5318 = _EVAL_5102 | _EVAL_5723;
  assign _EVAL_2079 = _EVAL_5133 & 32'h38;
  assign _EVAL_4500 = _EVAL_2079 == 32'h20;
  assign _EVAL_4499 = _EVAL_5318 | _EVAL_4500;
  assign _EVAL_845 = _EVAL_5133 & 32'h2050;
  assign _EVAL_580 = _EVAL_845 == 32'h2000;
  assign _EVAL_2404 = _EVAL_4499 | _EVAL_580;
  assign _EVAL_5565 = _EVAL_1242 & 32'h5f;
  assign _EVAL_2335 = _EVAL_5565 == 32'h17;
  assign _EVAL_608 = _EVAL_888 & 32'h306f;
  assign _EVAL_682 = _EVAL_608 == 32'h3;
  assign _EVAL_2786 = _EVAL_5386[19:15];
  assign _EVAL_2745 = _EVAL_888[19:15];
  assign _EVAL_3449 = _EVAL_4743[19:15];
  assign _EVAL_897 = _EVAL_386[19:15];
  assign _EVAL_2511 = _EVAL_5952 ? _EVAL_3449 : _EVAL_897;
  assign _EVAL_5080 = _EVAL_3570 ? _EVAL_2745 : _EVAL_2511;
  assign _EVAL_3929 = _EVAL_5833 ? _EVAL_2745 : _EVAL_5080;
  assign _EVAL_5607 = _EVAL_5833 ? _EVAL_2786 : _EVAL_3929;
  assign _EVAL_3882 = _EVAL_3455[19:15];
  assign _EVAL_5734 = _EVAL_2039[19:15];
  assign _EVAL_4781 = _EVAL_1242[19:15];
  assign _EVAL_2958 = _EVAL_2164[19:15];
  assign _EVAL_5295 = _EVAL_1074 ? _EVAL_4781 : _EVAL_2958;
  assign _EVAL_1093 = _EVAL_5926 ? _EVAL_5734 : _EVAL_5295;
  assign _EVAL_4800 = _EVAL_2970 ? _EVAL_5734 : _EVAL_1093;
  assign _EVAL_4753 = _EVAL_2970 ? _EVAL_3882 : _EVAL_4800;
  assign _EVAL_3340 = _EVAL_4268[19:15];
  assign _EVAL_1907 = _EVAL_3006[19:15];
  assign _EVAL_1296 = _EVAL_4882[19:15];
  assign _EVAL_5577 = _EVAL_5133[19:15];
  assign _EVAL_1431 = _EVAL_2901 ? _EVAL_1296 : _EVAL_5577;
  assign _EVAL_627 = _EVAL_2378 ? _EVAL_1907 : _EVAL_1431;
  assign _EVAL_308 = _EVAL_5690 ? _EVAL_1907 : _EVAL_627;
  assign _EVAL_531 = _EVAL_5690 ? _EVAL_3340 : _EVAL_308;
  assign _EVAL_945 = _EVAL_1978[19:15];
  assign _EVAL_3026 = _EVAL_1362[19:15];
  assign _EVAL_3857 = _EVAL_3271[19:15];
  assign _EVAL_285 = _EVAL_668 ? _EVAL_3026 : _EVAL_3857;
  assign _EVAL_458 = _EVAL_3050 ? _EVAL_945 : _EVAL_285;
  assign _EVAL_5797 = _EVAL_1069 ? _EVAL_945 : _EVAL_458;
  assign _EVAL_5226 = _EVAL_2142 ? _EVAL_531 : _EVAL_5797;
  assign _EVAL_4180 = _EVAL_3052 ? _EVAL_4753 : _EVAL_5226;
  assign _EVAL_3983 = _EVAL_5276 ? _EVAL_5607 : _EVAL_4180;
  assign _EVAL_1465 = _EVAL_1978 & 32'h62003010;
  assign _EVAL_5442 = _EVAL_1465 == 32'h60000010;
  assign _EVAL_1723 = _EVAL_4702 & 32'h5f;
  assign _EVAL_3656 = _EVAL_1723 == 32'h17;
  assign _EVAL_5255 = _EVAL_5472 ? 1'h1 : _EVAL_391;
  assign _EVAL_1004 = _EVAL_5875 & _EVAL_165;
  assign _EVAL_6055 = _EVAL_5875 & _EVAL_4214;
  assign _EVAL_1081 = _EVAL_1004 ? 1'h1 : _EVAL_6055;
  assign _EVAL_1630 = _EVAL_5454 ? 1'h1 : _EVAL_1081;
  assign _EVAL_2510 = _EVAL_5875 & _EVAL_2194;
  assign _EVAL_3508 = _EVAL_6086 & _EVAL_952;
  assign _EVAL_3950 = _EVAL_5875 & _EVAL_3508;
  assign _EVAL_183 = _EVAL_2510 ? 1'h1 : _EVAL_3950;
  assign _EVAL_5841 = _EVAL_5024 ? 1'h1 : _EVAL_183;
  assign _EVAL_5136 = _EVAL_5967 & _EVAL_4848;
  assign _EVAL_4573 = _EVAL_2293 | _EVAL_5136;
  assign _EVAL_4294 = _EVAL_4573 == _EVAL_3257;
  assign _EVAL_1903 = _EVAL_5967 & _EVAL_2754;
  assign _EVAL_2594 = _EVAL_5680 ? _EVAL_4294 : _EVAL_1903;
  assign _EVAL_5140 = _EVAL_4063 & _EVAL_2594;
  assign _EVAL_283 = _EVAL_5875 & _EVAL_5140;
  assign _EVAL_239 = _EVAL_6086 & _EVAL_2594;
  assign _EVAL_4880 = _EVAL_5875 & _EVAL_239;
  assign _EVAL_5583 = _EVAL_283 ? 1'h1 : _EVAL_4880;
  assign _EVAL_5473 = _EVAL_726 ? 1'h1 : _EVAL_5583;
  assign _EVAL_2385 = {_EVAL_5255,_EVAL_1630,_EVAL_5841,_EVAL_5473};
  assign _EVAL_3012 = _EVAL_2385 & _EVAL_4984;
  assign _EVAL_2394 = _EVAL_5854 & 32'hfff0007f;
  assign _EVAL_4044 = _EVAL_5813 & 32'h3c;
  assign _EVAL_5480 = _EVAL_4044 == 32'h4;
  assign _EVAL_1897 = _EVAL_5813 & 32'h80000060;
  assign _EVAL_5933 = _EVAL_1897 == 32'h40;
  assign _EVAL_4734 = _EVAL_5480 | _EVAL_5933;
  assign _EVAL_224 = _EVAL_5813 & 32'h70;
  assign _EVAL_2596 = _EVAL_224 == 32'h40;
  assign _EVAL_4836 = _EVAL_4734 | _EVAL_2596;
  assign _EVAL_2839 = _EVAL_5133[11:7];
  assign _EVAL_3396 = _EVAL_5854 & 32'h80000060;
  assign _EVAL_1267 = _EVAL_3396 == 32'h40;
  assign _EVAL_2470 = _EVAL_4743 & 32'h306f;
  assign _EVAL_1606 = _EVAL_2470 == 32'h1063;
  assign _EVAL_4677 = _EVAL_4882 & 32'h60;
  assign _EVAL_675 = _EVAL_4677 == 32'h0;
  assign _EVAL_2911 = _EVAL_6009 | _EVAL_675;
  assign _EVAL_1582 = _EVAL_888 & 32'hdfffffff;
  assign _EVAL_290 = _EVAL_1757 == 32'h40;
  assign _EVAL_4625 = _EVAL_1605 | _EVAL_290;
  assign _EVAL_5158 = _EVAL_4882 & 32'h1040;
  assign _EVAL_1553 = _EVAL_5158 == 32'h1040;
  assign _EVAL_3137 = _EVAL_4625 | _EVAL_1553;
  assign _EVAL_1415 = _EVAL_2694 == 32'h4;
  assign _EVAL_388 = _EVAL_3006 & 32'he800707f;
  assign _EVAL_5540 = _EVAL_388 == 32'h800202f;
  assign _EVAL_3295 = _EVAL_5854 & 32'hefe0007f;
  assign _EVAL_5188 = _EVAL_3295 == 32'hc0000053;
  assign _EVAL_4402 = _EVAL_4702 & 32'hfff0607f;
  assign _EVAL_2653 = _EVAL_4702 & 32'h64;
  assign _EVAL_4225 = _EVAL_2653 == 32'h20;
  assign _EVAL_4662 = _EVAL_4702 & 32'h34;
  assign _EVAL_4868 = _EVAL_4662 == 32'h20;
  assign _EVAL_598 = _EVAL_4225 | _EVAL_4868;
  assign _EVAL_498 = _EVAL_4702 & 32'h2048;
  assign _EVAL_4134 = _EVAL_498 == 32'h2008;
  assign _EVAL_3583 = _EVAL_598 | _EVAL_4134;
  assign _EVAL_959 = _EVAL_5854 == 32'h30200073;
  assign _EVAL_2228 = _EVAL_5854 & 32'h1040;
  assign _EVAL_2540 = _EVAL_2228 == 32'h1040;
  assign _EVAL_5156 = _EVAL_2856 | _EVAL_2540;
  assign _EVAL_5408 = _EVAL_5854 & 32'h2040;
  assign _EVAL_2323 = _EVAL_5408 == 32'h2040;
  assign _EVAL_3081 = _EVAL_5156 | _EVAL_2323;
  assign _EVAL_1592 = _EVAL_5813[11:7];
  assign _EVAL_181 = _EVAL_1958 ? _EVAL_1592 : _EVAL_3215;
  assign _EVAL_2311 = _EVAL_888 & 32'h7c;
  assign _EVAL_2479 = _EVAL_1242 & 32'h407f;
  assign _EVAL_286 = _EVAL_1362 & 32'h7f;
  assign _EVAL_3942 = _EVAL_1362 & 32'h80000060;
  assign _EVAL_3482 = _EVAL_3942 == 32'h40;
  assign _EVAL_3898 = _EVAL_1362 & 32'h10000060;
  assign _EVAL_2455 = _EVAL_3898 == 32'h40;
  assign _EVAL_884 = _EVAL_3482 | _EVAL_2455;
  assign _EVAL_4248 = _EVAL_884 | _EVAL_4770;
  assign _EVAL_2702 = _EVAL_3271 & 32'h80000060;
  assign _EVAL_3564 = _EVAL_2702 == 32'h40;
  assign _EVAL_3842 = _EVAL_3271 & 32'h10000060;
  assign _EVAL_2236 = _EVAL_3842 == 32'h40;
  assign _EVAL_1661 = _EVAL_3564 | _EVAL_2236;
  assign _EVAL_2798 = _EVAL_1661 | _EVAL_1739;
  assign _EVAL_4969 = _EVAL_668 ? _EVAL_4248 : _EVAL_2798;
  assign _EVAL_4290 = _EVAL_3271 & 32'hefe0007f;
  assign _EVAL_778 = _EVAL_4290 == 32'hc0000053;
  assign _EVAL_4332 = _EVAL_1978 == 32'h7b200073;
  assign _EVAL_1446 = _EVAL_5133 & 32'h90000010;
  assign _EVAL_5229 = _EVAL_1446 == 32'h80000010;
  assign _EVAL_4960 = _EVAL_5133 & 32'h34;
  assign _EVAL_1524 = _EVAL_4960 == 32'h20;
  assign _EVAL_4674 = _EVAL_4743 & 32'h20000040;
  assign _EVAL_1891 = _EVAL_4674 == 32'h40;
  assign _EVAL_4278 = _EVAL_2507 | _EVAL_5978;
  assign _EVAL_451 = _EVAL_1362 & 32'hfc00007f;
  assign _EVAL_5988 = _EVAL_451 == 32'h33;
  assign _EVAL_3009 = _EVAL_4278 | _EVAL_5988;
  assign _EVAL_2088 = _EVAL_1362 & 32'hbe00707f;
  assign _EVAL_4683 = _EVAL_2088 == 32'h33;
  assign _EVAL_1071 = _EVAL_3009 | _EVAL_4683;
  assign _EVAL_2708 = _EVAL_1362 & 32'h6000073;
  assign _EVAL_2033 = _EVAL_2708 == 32'h43;
  assign _EVAL_3809 = _EVAL_1071 | _EVAL_2033;
  assign _EVAL_4910 = _EVAL_1362 & 32'he600007f;
  assign _EVAL_3486 = _EVAL_4910 == 32'h53;
  assign _EVAL_2907 = _EVAL_3809 | _EVAL_3486;
  assign _EVAL_1312 = _EVAL_1362 & 32'h707b;
  assign _EVAL_5946 = _EVAL_1312 == 32'h63;
  assign _EVAL_789 = _EVAL_2907 | _EVAL_5946;
  assign _EVAL_3886 = _EVAL_286 == 32'h6f;
  assign _EVAL_5382 = _EVAL_789 | _EVAL_3886;
  assign _EVAL_429 = _EVAL_1362 & 32'hffefffff;
  assign _EVAL_2888 = _EVAL_429 == 32'h73;
  assign _EVAL_5260 = _EVAL_5382 | _EVAL_2888;
  assign _EVAL_6101 = _EVAL_1362 & 32'hfe00305f;
  assign _EVAL_3060 = _EVAL_6101 == 32'h1013;
  assign _EVAL_3586 = _EVAL_5260 | _EVAL_3060;
  assign _EVAL_2316 = _EVAL_1362 & 32'h705b;
  assign _EVAL_5116 = _EVAL_2316 == 32'h2003;
  assign _EVAL_2533 = _EVAL_3586 | _EVAL_5116;
  assign _EVAL_4628 = _EVAL_2710 == 32'h2013;
  assign _EVAL_2489 = _EVAL_2533 | _EVAL_4628;
  assign _EVAL_5544 = _EVAL_389 == 32'h202f;
  assign _EVAL_6110 = _EVAL_2489 | _EVAL_5544;
  assign _EVAL_1053 = _EVAL_6110 | _EVAL_4647;
  assign _EVAL_3034 = _EVAL_1362 & 32'hbe00705f;
  assign _EVAL_1814 = _EVAL_3034 == 32'h5013;
  assign _EVAL_4018 = _EVAL_1053 | _EVAL_1814;
  assign _EVAL_6130 = _EVAL_1362 & 32'he800707f;
  assign _EVAL_2421 = _EVAL_6130 == 32'h800202f;
  assign _EVAL_4559 = _EVAL_4018 | _EVAL_2421;
  assign _EVAL_2138 = _EVAL_1362 & 32'hf9f0707f;
  assign _EVAL_5470 = _EVAL_2138 == 32'h1000202f;
  assign _EVAL_5895 = _EVAL_4559 | _EVAL_5470;
  assign _EVAL_1938 = _EVAL_1362 & 32'hdfffffff;
  assign _EVAL_2118 = _EVAL_1938 == 32'h10500073;
  assign _EVAL_1214 = _EVAL_5895 | _EVAL_2118;
  assign _EVAL_437 = _EVAL_1362 & 32'hf600607f;
  assign _EVAL_3346 = _EVAL_437 == 32'h20000053;
  assign _EVAL_1202 = _EVAL_1214 | _EVAL_3346;
  assign _EVAL_5879 = _EVAL_1362 & 32'h7e00607f;
  assign _EVAL_1400 = _EVAL_5879 == 32'h20000053;
  assign _EVAL_5929 = _EVAL_1202 | _EVAL_1400;
  assign _EVAL_1218 = _EVAL_1362 & 32'h7e00507f;
  assign _EVAL_3777 = _EVAL_1218 == 32'h20000053;
  assign _EVAL_5643 = _EVAL_5929 | _EVAL_3777;
  assign _EVAL_3152 = _EVAL_1362 == 32'h30200073;
  assign _EVAL_1463 = _EVAL_5643 | _EVAL_3152;
  assign _EVAL_5049 = _EVAL_740 == 32'h58000053;
  assign _EVAL_3924 = _EVAL_1463 | _EVAL_5049;
  assign _EVAL_2580 = _EVAL_1362 == 32'h7b200073;
  assign _EVAL_657 = _EVAL_3924 | _EVAL_2580;
  assign _EVAL_4108 = _EVAL_3271 == 32'h7b200073;
  assign _EVAL_1543 = _EVAL_2039 & 32'h18;
  assign _EVAL_1107 = _EVAL_1543 == 32'h0;
  assign _EVAL_5380 = _EVAL_888 & 32'h80000010;
  assign _EVAL_4288 = _EVAL_5380 == 32'h10;
  assign _EVAL_4471 = _EVAL_888 & 32'h50;
  assign _EVAL_5272 = _EVAL_4471 == 32'h10;
  assign _EVAL_3008 = _EVAL_4288 | _EVAL_5272;
  assign _EVAL_3086 = _EVAL_888 & 32'h40000040;
  assign _EVAL_5419 = _EVAL_3086 == 32'h40;
  assign _EVAL_1577 = _EVAL_3008 | _EVAL_5419;
  assign _EVAL_1793 = _EVAL_888 & 32'h20000040;
  assign _EVAL_4367 = _EVAL_1793 == 32'h40;
  assign _EVAL_2538 = _EVAL_1577 | _EVAL_4367;
  assign _EVAL_3231 = _EVAL_4743 & 32'h80000060;
  assign _EVAL_4714 = _EVAL_3231 == 32'h40;
  assign _EVAL_4925 = _EVAL_4743 & 32'h10000060;
  assign _EVAL_1072 = _EVAL_4925 == 32'h40;
  assign _EVAL_838 = _EVAL_4714 | _EVAL_1072;
  assign _EVAL_3238 = _EVAL_838 | _EVAL_1433;
  assign _EVAL_591 = _EVAL_4702 & 32'h7c;
  assign _EVAL_5466 = _EVAL_5854 & 32'hdfffffff;
  assign _EVAL_2309 = _EVAL_5466 == 32'h10500073;
  assign _EVAL_3783 = _EVAL_1892 | _EVAL_2309;
  assign _EVAL_549 = _EVAL_5854 & 32'hf600607f;
  assign _EVAL_5262 = _EVAL_549 == 32'h20000053;
  assign _EVAL_4712 = _EVAL_3783 | _EVAL_5262;
  assign _EVAL_1631 = _EVAL_5854 & 32'h7e00607f;
  assign _EVAL_2061 = _EVAL_1631 == 32'h20000053;
  assign _EVAL_4783 = _EVAL_4712 | _EVAL_2061;
  assign _EVAL_5814 = _EVAL_5854 & 32'h7e00507f;
  assign _EVAL_5451 = _EVAL_5814 == 32'h20000053;
  assign _EVAL_182 = _EVAL_4783 | _EVAL_5451;
  assign _EVAL_946 = _EVAL_182 | _EVAL_959;
  assign _EVAL_393 = _EVAL_2394 == 32'h58000053;
  assign _EVAL_4109 = _EVAL_946 | _EVAL_393;
  assign _EVAL_1063 = _EVAL_5854 == 32'h7b200073;
  assign _EVAL_1810 = _EVAL_4109 | _EVAL_1063;
  assign _EVAL_3069 = _EVAL_1810 | _EVAL_5188;
  assign _EVAL_4410 = _EVAL_530 == 32'he0000053;
  assign _EVAL_3077 = _EVAL_3069 | _EVAL_4410;
  assign _EVAL_4701 = _EVAL_5854 & 32'heff0707f;
  assign _EVAL_4756 = _EVAL_4701 == 32'he0000053;
  assign _EVAL_2667 = _EVAL_3077 | _EVAL_4756;
  assign _EVAL_3268 = _EVAL_3018 == 32'hfc000073;
  assign _EVAL_1019 = _EVAL_2667 | _EVAL_3268;
  assign _EVAL_2582 = _EVAL_5854 & 32'h306f;
  assign _EVAL_1717 = _EVAL_2582 == 32'h1063;
  assign _EVAL_2735 = _EVAL_1019 | _EVAL_1717;
  assign _EVAL_2826 = _EVAL_5854 & 32'h407f;
  assign _EVAL_4948 = _EVAL_2826 == 32'h4063;
  assign _EVAL_558 = _EVAL_2735 | _EVAL_4948;
  assign _EVAL_5538 = _EVAL_5854 & 32'h605f;
  assign _EVAL_299 = _EVAL_5538 == 32'h3;
  assign _EVAL_2400 = _EVAL_558 | _EVAL_299;
  assign _EVAL_4506 = _EVAL_2582 == 32'h3;
  assign _EVAL_4918 = _EVAL_2400 | _EVAL_4506;
  assign _EVAL_2349 = _EVAL_846 == 1'h0;
  assign _EVAL_1875 = _EVAL_888 & 32'hf9f0707f;
  assign _EVAL_1273 = _EVAL_1875 == 32'h1000202f;
  assign _EVAL_2857 = _EVAL_2905 | _EVAL_1273;
  assign _EVAL_2899 = _EVAL_1582 == 32'h10500073;
  assign _EVAL_3457 = _EVAL_2857 | _EVAL_2899;
  assign _EVAL_2055 = _EVAL_888 & 32'hf600607f;
  assign _EVAL_3516 = _EVAL_2055 == 32'h20000053;
  assign _EVAL_5727 = _EVAL_3457 | _EVAL_3516;
  assign _EVAL_3024 = _EVAL_888 & 32'h7e00607f;
  assign _EVAL_3775 = _EVAL_3024 == 32'h20000053;
  assign _EVAL_2840 = _EVAL_5727 | _EVAL_3775;
  assign _EVAL_5405 = _EVAL_888 & 32'h7e00507f;
  assign _EVAL_2512 = _EVAL_5405 == 32'h20000053;
  assign _EVAL_2099 = _EVAL_2840 | _EVAL_2512;
  assign _EVAL_3948 = _EVAL_888 == 32'h30200073;
  assign _EVAL_3279 = _EVAL_2099 | _EVAL_3948;
  assign _EVAL_1736 = _EVAL_888 & 32'hfff0007f;
  assign _EVAL_1534 = _EVAL_1736 == 32'h58000053;
  assign _EVAL_3943 = _EVAL_3279 | _EVAL_1534;
  assign _EVAL_3017 = _EVAL_888 == 32'h7b200073;
  assign _EVAL_438 = _EVAL_3943 | _EVAL_3017;
  assign _EVAL_1469 = _EVAL_888 & 32'hefe0007f;
  assign _EVAL_4526 = _EVAL_1469 == 32'hc0000053;
  assign _EVAL_163 = _EVAL_438 | _EVAL_4526;
  assign _EVAL_3760 = _EVAL_5776 == 32'he0000053;
  assign _EVAL_4854 = _EVAL_163 | _EVAL_3760;
  assign _EVAL_5608 = _EVAL_888 & 32'heff0707f;
  assign _EVAL_331 = _EVAL_5608 == 32'he0000053;
  assign _EVAL_6092 = _EVAL_4854 | _EVAL_331;
  assign _EVAL_5277 = _EVAL_888 & 32'hffd07fff;
  assign _EVAL_3576 = _EVAL_5277 == 32'hfc000073;
  assign _EVAL_2023 = _EVAL_6092 | _EVAL_3576;
  assign _EVAL_5347 = _EVAL_608 == 32'h1063;
  assign _EVAL_1775 = _EVAL_2023 | _EVAL_5347;
  assign _EVAL_474 = _EVAL_888 & 32'h407f;
  assign _EVAL_2066 = _EVAL_474 == 32'h4063;
  assign _EVAL_3028 = _EVAL_1775 | _EVAL_2066;
  assign _EVAL_4392 = _EVAL_888 & 32'h605f;
  assign _EVAL_4891 = _EVAL_4392 == 32'h3;
  assign _EVAL_2501 = _EVAL_3028 | _EVAL_4891;
  assign _EVAL_3831 = _EVAL_2501 | _EVAL_682;
  assign _EVAL_4303 = _EVAL_2349 ? 1'h0 : _EVAL_3831;
  assign _EVAL_3596 = _EVAL_4743 & 32'h7e00507f;
  assign _EVAL_5556 = _EVAL_3596 == 32'h20000053;
  assign _EVAL_3803 = _EVAL_4817 | _EVAL_5556;
  assign _EVAL_4117 = _EVAL_4743 == 32'h30200073;
  assign _EVAL_366 = _EVAL_3803 | _EVAL_4117;
  assign _EVAL_2522 = _EVAL_4743 & 32'hfff0007f;
  assign _EVAL_795 = _EVAL_2522 == 32'h58000053;
  assign _EVAL_2960 = _EVAL_366 | _EVAL_795;
  assign _EVAL_2189 = _EVAL_4743 == 32'h7b200073;
  assign _EVAL_4678 = _EVAL_2960 | _EVAL_2189;
  assign _EVAL_1467 = _EVAL_4743 & 32'hefe0007f;
  assign _EVAL_2599 = _EVAL_1467 == 32'hc0000053;
  assign _EVAL_6044 = _EVAL_4678 | _EVAL_2599;
  assign _EVAL_1792 = _EVAL_4743 & 32'hfff0607f;
  assign _EVAL_3425 = _EVAL_1792 == 32'he0000053;
  assign _EVAL_251 = _EVAL_6044 | _EVAL_3425;
  assign _EVAL_6043 = _EVAL_4743 & 32'heff0707f;
  assign _EVAL_3165 = _EVAL_6043 == 32'he0000053;
  assign _EVAL_4995 = _EVAL_251 | _EVAL_3165;
  assign _EVAL_1452 = _EVAL_4743 & 32'hffd07fff;
  assign _EVAL_5036 = _EVAL_1452 == 32'hfc000073;
  assign _EVAL_6073 = _EVAL_4995 | _EVAL_5036;
  assign _EVAL_944 = _EVAL_6073 | _EVAL_1606;
  assign _EVAL_2544 = _EVAL_4743 & 32'h407f;
  assign _EVAL_5934 = _EVAL_2544 == 32'h4063;
  assign _EVAL_2481 = _EVAL_944 | _EVAL_5934;
  assign _EVAL_665 = _EVAL_2481 | _EVAL_5193;
  assign _EVAL_3627 = _EVAL_2470 == 32'h3;
  assign _EVAL_2454 = _EVAL_665 | _EVAL_3627;
  assign _EVAL_5296 = _EVAL_1405 ? 1'h0 : _EVAL_2454;
  assign _EVAL_3830 = _EVAL_5386[12:5];
  assign _EVAL_2092 = _EVAL_3830 != 8'h0;
  assign _EVAL_2635 = _EVAL_2175 ? 1'h1 : _EVAL_2092;
  assign _EVAL_2408 = _EVAL_179 ? 1'h1 : _EVAL_2635;
  assign _EVAL_3371 = _EVAL_268 ? 1'h1 : _EVAL_2408;
  assign _EVAL_5100 = _EVAL_3261 ? 1'h1 : _EVAL_3371;
  assign _EVAL_1193 = _EVAL_3493 ? 1'h1 : _EVAL_5100;
  assign _EVAL_3671 = _EVAL_4185 ? 1'h1 : _EVAL_1193;
  assign _EVAL_2453 = _EVAL_4999 ? 1'h1 : _EVAL_3671;
  assign _EVAL_2425 = _EVAL_2453 == 1'h0;
  assign _EVAL_6056 = _EVAL_386 & 32'hffd07fff;
  assign _EVAL_4003 = _EVAL_6056 == 32'hfc000073;
  assign _EVAL_4082 = _EVAL_5234 | _EVAL_4003;
  assign _EVAL_2149 = _EVAL_386 & 32'h306f;
  assign _EVAL_696 = _EVAL_2149 == 32'h1063;
  assign _EVAL_1039 = _EVAL_4082 | _EVAL_696;
  assign _EVAL_658 = _EVAL_5206 == 32'h4063;
  assign _EVAL_2171 = _EVAL_1039 | _EVAL_658;
  assign _EVAL_5762 = _EVAL_386 & 32'h605f;
  assign _EVAL_6124 = _EVAL_5762 == 32'h3;
  assign _EVAL_3058 = _EVAL_2171 | _EVAL_6124;
  assign _EVAL_825 = _EVAL_2149 == 32'h3;
  assign _EVAL_5508 = _EVAL_3058 | _EVAL_825;
  assign _EVAL_4780 = _EVAL_2425 ? 1'h0 : _EVAL_5508;
  assign _EVAL_4446 = _EVAL_5952 ? _EVAL_5296 : _EVAL_4780;
  assign _EVAL_4284 = _EVAL_3570 ? _EVAL_4303 : _EVAL_4446;
  assign _EVAL_4147 = _EVAL_5833 ? _EVAL_4303 : _EVAL_4284;
  assign _EVAL_4296 = _EVAL_5833 ? _EVAL_4918 : _EVAL_4147;
  assign _EVAL_2971 = _EVAL_5311 & 32'h407f;
  assign _EVAL_5083 = _EVAL_2971 == 32'h4063;
  assign _EVAL_1494 = _EVAL_504 | _EVAL_5083;
  assign _EVAL_2137 = _EVAL_5311 & 32'h605f;
  assign _EVAL_3582 = _EVAL_2137 == 32'h3;
  assign _EVAL_3365 = _EVAL_1494 | _EVAL_3582;
  assign _EVAL_1125 = _EVAL_1291 == 32'h3;
  assign _EVAL_2432 = _EVAL_3365 | _EVAL_1125;
  assign _EVAL_5799 = _EVAL_1242 & 32'h207f;
  assign _EVAL_4814 = _EVAL_5799 == 32'h3;
  assign _EVAL_4747 = _EVAL_1242 & 32'h607f;
  assign _EVAL_6013 = _EVAL_4747 == 32'hf;
  assign _EVAL_753 = _EVAL_4814 | _EVAL_6013;
  assign _EVAL_1821 = _EVAL_753 | _EVAL_2335;
  assign _EVAL_2180 = _EVAL_2027 == 32'h33;
  assign _EVAL_276 = _EVAL_1821 | _EVAL_2180;
  assign _EVAL_4212 = _EVAL_1242 & 32'hbe00707f;
  assign _EVAL_1834 = _EVAL_4212 == 32'h33;
  assign _EVAL_2492 = _EVAL_276 | _EVAL_1834;
  assign _EVAL_1569 = _EVAL_1242 & 32'h6000073;
  assign _EVAL_733 = _EVAL_1569 == 32'h43;
  assign _EVAL_1676 = _EVAL_2492 | _EVAL_733;
  assign _EVAL_4405 = _EVAL_1242 & 32'he600007f;
  assign _EVAL_720 = _EVAL_4405 == 32'h53;
  assign _EVAL_4502 = _EVAL_1676 | _EVAL_720;
  assign _EVAL_433 = _EVAL_1242 & 32'h707b;
  assign _EVAL_3162 = _EVAL_433 == 32'h63;
  assign _EVAL_4962 = _EVAL_4502 | _EVAL_3162;
  assign _EVAL_1787 = _EVAL_1242 & 32'h7f;
  assign _EVAL_3765 = _EVAL_1787 == 32'h6f;
  assign _EVAL_1389 = _EVAL_4962 | _EVAL_3765;
  assign _EVAL_5866 = _EVAL_1242 & 32'hffefffff;
  assign _EVAL_3120 = _EVAL_5866 == 32'h73;
  assign _EVAL_3109 = _EVAL_1389 | _EVAL_3120;
  assign _EVAL_2306 = _EVAL_1242 & 32'hfe00305f;
  assign _EVAL_1987 = _EVAL_2306 == 32'h1013;
  assign _EVAL_1379 = _EVAL_3109 | _EVAL_1987;
  assign _EVAL_5246 = _EVAL_1379 | _EVAL_1280;
  assign _EVAL_1155 = _EVAL_5799 == 32'h2013;
  assign _EVAL_5139 = _EVAL_5246 | _EVAL_1155;
  assign _EVAL_2098 = _EVAL_1242 & 32'h1800707f;
  assign _EVAL_5185 = _EVAL_2098 == 32'h202f;
  assign _EVAL_5662 = _EVAL_5139 | _EVAL_5185;
  assign _EVAL_5499 = _EVAL_5799 == 32'h2073;
  assign _EVAL_4207 = _EVAL_5662 | _EVAL_5499;
  assign _EVAL_4746 = _EVAL_5795 == 32'h5013;
  assign _EVAL_2643 = _EVAL_4207 | _EVAL_4746;
  assign _EVAL_2082 = _EVAL_1242 & 32'he800707f;
  assign _EVAL_1227 = _EVAL_2082 == 32'h800202f;
  assign _EVAL_3005 = _EVAL_2643 | _EVAL_1227;
  assign _EVAL_2992 = _EVAL_1242 & 32'hf9f0707f;
  assign _EVAL_3779 = _EVAL_2992 == 32'h1000202f;
  assign _EVAL_734 = _EVAL_3005 | _EVAL_3779;
  assign _EVAL_3776 = _EVAL_1242 & 32'hdfffffff;
  assign _EVAL_1251 = _EVAL_3776 == 32'h10500073;
  assign _EVAL_1207 = _EVAL_734 | _EVAL_1251;
  assign _EVAL_1108 = _EVAL_1242 & 32'hf600607f;
  assign _EVAL_1965 = _EVAL_1108 == 32'h20000053;
  assign _EVAL_1293 = _EVAL_1207 | _EVAL_1965;
  assign _EVAL_934 = _EVAL_1242 & 32'h7e00607f;
  assign _EVAL_3497 = _EVAL_934 == 32'h20000053;
  assign _EVAL_1432 = _EVAL_1293 | _EVAL_3497;
  assign _EVAL_4285 = _EVAL_1242 & 32'h7e00507f;
  assign _EVAL_3634 = _EVAL_4285 == 32'h20000053;
  assign _EVAL_1744 = _EVAL_1432 | _EVAL_3634;
  assign _EVAL_6066 = _EVAL_1744 | _EVAL_3130;
  assign _EVAL_900 = _EVAL_2405 == 32'h58000053;
  assign _EVAL_5160 = _EVAL_6066 | _EVAL_900;
  assign _EVAL_4954 = _EVAL_1242 == 32'h7b200073;
  assign _EVAL_1305 = _EVAL_5160 | _EVAL_4954;
  assign _EVAL_2659 = _EVAL_1242 & 32'hefe0007f;
  assign _EVAL_4336 = _EVAL_2659 == 32'hc0000053;
  assign _EVAL_4160 = _EVAL_1305 | _EVAL_4336;
  assign _EVAL_5181 = _EVAL_4160 | _EVAL_2006;
  assign _EVAL_3354 = _EVAL_4227 == 32'he0000053;
  assign _EVAL_3504 = _EVAL_5181 | _EVAL_3354;
  assign _EVAL_4637 = _EVAL_3504 | _EVAL_2069;
  assign _EVAL_1060 = _EVAL_1242 & 32'h306f;
  assign _EVAL_5522 = _EVAL_1060 == 32'h1063;
  assign _EVAL_3888 = _EVAL_4637 | _EVAL_5522;
  assign _EVAL_3933 = _EVAL_2479 == 32'h4063;
  assign _EVAL_1067 = _EVAL_3888 | _EVAL_3933;
  assign _EVAL_2733 = _EVAL_1242 & 32'h605f;
  assign _EVAL_5502 = _EVAL_2733 == 32'h3;
  assign _EVAL_3225 = _EVAL_1067 | _EVAL_5502;
  assign _EVAL_2842 = _EVAL_1060 == 32'h3;
  assign _EVAL_3381 = _EVAL_3225 | _EVAL_2842;
  assign _EVAL_5050 = _EVAL_5563 ? 1'h0 : _EVAL_3381;
  assign _EVAL_2100 = _EVAL_453 ? 1'h1 : _EVAL_4306;
  assign _EVAL_3699 = _EVAL_2288 ? 1'h1 : _EVAL_2100;
  assign _EVAL_3747 = _EVAL_4669 ? 1'h1 : _EVAL_3699;
  assign _EVAL_5264 = _EVAL_3747 == 1'h0;
  assign _EVAL_5523 = _EVAL_2164 == 32'h7b200073;
  assign _EVAL_3397 = _EVAL_5453 | _EVAL_5523;
  assign _EVAL_5172 = _EVAL_2164 & 32'hefe0007f;
  assign _EVAL_215 = _EVAL_5172 == 32'hc0000053;
  assign _EVAL_2046 = _EVAL_3397 | _EVAL_215;
  assign _EVAL_3709 = _EVAL_2164 & 32'hfff0607f;
  assign _EVAL_5887 = _EVAL_3709 == 32'he0000053;
  assign _EVAL_1192 = _EVAL_2046 | _EVAL_5887;
  assign _EVAL_4699 = _EVAL_2164 & 32'heff0707f;
  assign _EVAL_5610 = _EVAL_4699 == 32'he0000053;
  assign _EVAL_4767 = _EVAL_1192 | _EVAL_5610;
  assign _EVAL_1485 = _EVAL_2164 & 32'hffd07fff;
  assign _EVAL_2734 = _EVAL_1485 == 32'hfc000073;
  assign _EVAL_4030 = _EVAL_4767 | _EVAL_2734;
  assign _EVAL_5653 = _EVAL_4030 | _EVAL_5631;
  assign _EVAL_3797 = _EVAL_2164 & 32'h407f;
  assign _EVAL_5301 = _EVAL_3797 == 32'h4063;
  assign _EVAL_5868 = _EVAL_5653 | _EVAL_5301;
  assign _EVAL_4631 = _EVAL_2164 & 32'h605f;
  assign _EVAL_2675 = _EVAL_4631 == 32'h3;
  assign _EVAL_5137 = _EVAL_5868 | _EVAL_2675;
  assign _EVAL_338 = _EVAL_515 == 32'h3;
  assign _EVAL_766 = _EVAL_5137 | _EVAL_338;
  assign _EVAL_756 = _EVAL_5264 ? 1'h0 : _EVAL_766;
  assign _EVAL_5294 = _EVAL_1074 ? _EVAL_5050 : _EVAL_756;
  assign _EVAL_5319 = _EVAL_5926 ? _EVAL_5060 : _EVAL_5294;
  assign _EVAL_2403 = _EVAL_2970 ? _EVAL_5060 : _EVAL_5319;
  assign _EVAL_6030 = _EVAL_2970 ? _EVAL_2432 : _EVAL_2403;
  assign _EVAL_228 = _EVAL_4268 & 32'hefe0007f;
  assign _EVAL_2616 = _EVAL_228 == 32'hc0000053;
  assign _EVAL_2807 = _EVAL_4201 | _EVAL_2616;
  assign _EVAL_1640 = _EVAL_4268 & 32'hfff0607f;
  assign _EVAL_4317 = _EVAL_1640 == 32'he0000053;
  assign _EVAL_3267 = _EVAL_2807 | _EVAL_4317;
  assign _EVAL_2068 = _EVAL_4268 & 32'heff0707f;
  assign _EVAL_2701 = _EVAL_2068 == 32'he0000053;
  assign _EVAL_2285 = _EVAL_3267 | _EVAL_2701;
  assign _EVAL_2270 = _EVAL_4268 & 32'hffd07fff;
  assign _EVAL_1141 = _EVAL_2270 == 32'hfc000073;
  assign _EVAL_4803 = _EVAL_2285 | _EVAL_1141;
  assign _EVAL_1349 = _EVAL_4268 & 32'h306f;
  assign _EVAL_557 = _EVAL_1349 == 32'h1063;
  assign _EVAL_4417 = _EVAL_4803 | _EVAL_557;
  assign _EVAL_4833 = _EVAL_4268 & 32'h407f;
  assign _EVAL_4040 = _EVAL_4833 == 32'h4063;
  assign _EVAL_1911 = _EVAL_4417 | _EVAL_4040;
  assign _EVAL_2237 = _EVAL_4268 & 32'h605f;
  assign _EVAL_296 = _EVAL_2237 == 32'h3;
  assign _EVAL_2804 = _EVAL_1911 | _EVAL_296;
  assign _EVAL_2676 = _EVAL_1349 == 32'h3;
  assign _EVAL_3921 = _EVAL_2804 | _EVAL_2676;
  assign _EVAL_4924 = _EVAL_4268[12:2];
  assign _EVAL_4075 = _EVAL_4924 != 11'h0;
  assign _EVAL_3766 = _EVAL_4038 ? _EVAL_3685 : 1'h1;
  assign _EVAL_288 = _EVAL_1743 ? 1'h1 : _EVAL_3766;
  assign _EVAL_1369 = _EVAL_3712 ? _EVAL_4075 : _EVAL_288;
  assign _EVAL_563 = _EVAL_2321 ? 1'h1 : _EVAL_1369;
  assign _EVAL_3774 = _EVAL_5053 ? 1'h1 : _EVAL_563;
  assign _EVAL_1122 = _EVAL_5623 ? 1'h1 : _EVAL_3774;
  assign _EVAL_843 = _EVAL_1122 == 1'h0;
  assign _EVAL_2870 = _EVAL_3006 & 32'hbe00705f;
  assign _EVAL_1677 = _EVAL_2870 == 32'h5013;
  assign _EVAL_5595 = _EVAL_3632 | _EVAL_1677;
  assign _EVAL_4988 = _EVAL_5595 | _EVAL_5540;
  assign _EVAL_613 = _EVAL_3006 & 32'hf9f0707f;
  assign _EVAL_4590 = _EVAL_613 == 32'h1000202f;
  assign _EVAL_3089 = _EVAL_4988 | _EVAL_4590;
  assign _EVAL_1225 = _EVAL_3006 & 32'hdfffffff;
  assign _EVAL_1352 = _EVAL_1225 == 32'h10500073;
  assign _EVAL_413 = _EVAL_3089 | _EVAL_1352;
  assign _EVAL_3462 = _EVAL_3006 & 32'hf600607f;
  assign _EVAL_839 = _EVAL_3462 == 32'h20000053;
  assign _EVAL_3772 = _EVAL_413 | _EVAL_839;
  assign _EVAL_3075 = _EVAL_3006 & 32'h7e00607f;
  assign _EVAL_3501 = _EVAL_3075 == 32'h20000053;
  assign _EVAL_1090 = _EVAL_3772 | _EVAL_3501;
  assign _EVAL_403 = _EVAL_3006 & 32'h7e00507f;
  assign _EVAL_906 = _EVAL_403 == 32'h20000053;
  assign _EVAL_5026 = _EVAL_1090 | _EVAL_906;
  assign _EVAL_5254 = _EVAL_5026 | _EVAL_3577;
  assign _EVAL_3721 = _EVAL_5254 | _EVAL_1936;
  assign _EVAL_1089 = _EVAL_3006 == 32'h7b200073;
  assign _EVAL_2674 = _EVAL_3721 | _EVAL_1089;
  assign _EVAL_4993 = _EVAL_3006 & 32'hefe0007f;
  assign _EVAL_211 = _EVAL_4993 == 32'hc0000053;
  assign _EVAL_1461 = _EVAL_2674 | _EVAL_211;
  assign _EVAL_770 = _EVAL_3006 & 32'hfff0607f;
  assign _EVAL_4871 = _EVAL_770 == 32'he0000053;
  assign _EVAL_1948 = _EVAL_1461 | _EVAL_4871;
  assign _EVAL_3441 = _EVAL_3006 & 32'heff0707f;
  assign _EVAL_2379 = _EVAL_3441 == 32'he0000053;
  assign _EVAL_2921 = _EVAL_1948 | _EVAL_2379;
  assign _EVAL_5514 = _EVAL_3006 & 32'hffd07fff;
  assign _EVAL_406 = _EVAL_5514 == 32'hfc000073;
  assign _EVAL_6072 = _EVAL_2921 | _EVAL_406;
  assign _EVAL_2109 = _EVAL_4642 == 32'h1063;
  assign _EVAL_5048 = _EVAL_6072 | _EVAL_2109;
  assign _EVAL_4929 = _EVAL_3006 & 32'h407f;
  assign _EVAL_4101 = _EVAL_4929 == 32'h4063;
  assign _EVAL_2045 = _EVAL_5048 | _EVAL_4101;
  assign _EVAL_885 = _EVAL_3006 & 32'h605f;
  assign _EVAL_3254 = _EVAL_885 == 32'h3;
  assign _EVAL_231 = _EVAL_2045 | _EVAL_3254;
  assign _EVAL_4552 = _EVAL_231 | _EVAL_1284;
  assign _EVAL_4393 = _EVAL_843 ? 1'h0 : _EVAL_4552;
  assign _EVAL_3916 = _EVAL_2378 ? _EVAL_4393 : _EVAL_5894;
  assign _EVAL_1916 = _EVAL_5690 ? _EVAL_4393 : _EVAL_3916;
  assign _EVAL_3108 = _EVAL_5690 ? _EVAL_3921 : _EVAL_1916;
  assign _EVAL_545 = _EVAL_5821 ? 1'h1 : _EVAL_2464;
  assign _EVAL_6004 = _EVAL_418 ? 1'h1 : _EVAL_545;
  assign _EVAL_1459 = _EVAL_6004 == 1'h0;
  assign _EVAL_699 = _EVAL_1978 & 32'h7e00607f;
  assign _EVAL_817 = _EVAL_699 == 32'h20000053;
  assign _EVAL_3567 = _EVAL_5981 | _EVAL_817;
  assign _EVAL_1031 = _EVAL_1978 & 32'h7e00507f;
  assign _EVAL_3236 = _EVAL_1031 == 32'h20000053;
  assign _EVAL_5509 = _EVAL_3567 | _EVAL_3236;
  assign _EVAL_3490 = _EVAL_1978 == 32'h30200073;
  assign _EVAL_2217 = _EVAL_5509 | _EVAL_3490;
  assign _EVAL_2019 = _EVAL_1978 & 32'hfff0007f;
  assign _EVAL_5142 = _EVAL_2019 == 32'h58000053;
  assign _EVAL_4904 = _EVAL_2217 | _EVAL_5142;
  assign _EVAL_4607 = _EVAL_4904 | _EVAL_4332;
  assign _EVAL_2420 = _EVAL_1978 & 32'hefe0007f;
  assign _EVAL_539 = _EVAL_2420 == 32'hc0000053;
  assign _EVAL_3154 = _EVAL_4607 | _EVAL_539;
  assign _EVAL_1335 = _EVAL_1978 & 32'hfff0607f;
  assign _EVAL_2738 = _EVAL_1335 == 32'he0000053;
  assign _EVAL_3532 = _EVAL_3154 | _EVAL_2738;
  assign _EVAL_2435 = _EVAL_1978 & 32'heff0707f;
  assign _EVAL_5551 = _EVAL_2435 == 32'he0000053;
  assign _EVAL_700 = _EVAL_3532 | _EVAL_5551;
  assign _EVAL_3657 = _EVAL_1978 & 32'hffd07fff;
  assign _EVAL_2342 = _EVAL_3657 == 32'hfc000073;
  assign _EVAL_4313 = _EVAL_700 | _EVAL_2342;
  assign _EVAL_1281 = _EVAL_1978 & 32'h306f;
  assign _EVAL_4073 = _EVAL_1281 == 32'h1063;
  assign _EVAL_4776 = _EVAL_4313 | _EVAL_4073;
  assign _EVAL_1196 = _EVAL_1978 & 32'h407f;
  assign _EVAL_1204 = _EVAL_1196 == 32'h4063;
  assign _EVAL_2499 = _EVAL_4776 | _EVAL_1204;
  assign _EVAL_1776 = _EVAL_1978 & 32'h605f;
  assign _EVAL_2633 = _EVAL_1776 == 32'h3;
  assign _EVAL_3649 = _EVAL_2499 | _EVAL_2633;
  assign _EVAL_4497 = _EVAL_1281 == 32'h3;
  assign _EVAL_424 = _EVAL_3649 | _EVAL_4497;
  assign _EVAL_4886 = _EVAL_1459 ? 1'h0 : _EVAL_424;
  assign _EVAL_4407 = {_EVAL_2409,_EVAL_4489};
  assign _EVAL_4539 = _EVAL_4407 != 12'h0;
  assign _EVAL_6091 = _EVAL_4352 ? _EVAL_4539 : 1'h1;
  assign _EVAL_774 = _EVAL_4202 ? 1'h1 : _EVAL_6091;
  assign _EVAL_2774 = _EVAL_2644 ? 1'h1 : _EVAL_774;
  assign _EVAL_5444 = _EVAL_5821 ? 1'h1 : _EVAL_2774;
  assign _EVAL_3571 = _EVAL_418 ? 1'h1 : _EVAL_5444;
  assign _EVAL_6039 = _EVAL_3571 == 1'h0;
  assign _EVAL_5343 = _EVAL_1362 & 32'hefe0007f;
  assign _EVAL_1132 = _EVAL_5343 == 32'hc0000053;
  assign _EVAL_5890 = _EVAL_657 | _EVAL_1132;
  assign _EVAL_940 = _EVAL_1362 & 32'hfff0607f;
  assign _EVAL_4408 = _EVAL_940 == 32'he0000053;
  assign _EVAL_3325 = _EVAL_5890 | _EVAL_4408;
  assign _EVAL_1712 = _EVAL_1362 & 32'heff0707f;
  assign _EVAL_3409 = _EVAL_1712 == 32'he0000053;
  assign _EVAL_5371 = _EVAL_3325 | _EVAL_3409;
  assign _EVAL_5288 = _EVAL_1362 & 32'hffd07fff;
  assign _EVAL_4149 = _EVAL_5288 == 32'hfc000073;
  assign _EVAL_1256 = _EVAL_5371 | _EVAL_4149;
  assign _EVAL_4881 = _EVAL_1362 & 32'h306f;
  assign _EVAL_5635 = _EVAL_4881 == 32'h1063;
  assign _EVAL_809 = _EVAL_1256 | _EVAL_5635;
  assign _EVAL_1785 = _EVAL_1362 & 32'h407f;
  assign _EVAL_5940 = _EVAL_1785 == 32'h4063;
  assign _EVAL_5200 = _EVAL_809 | _EVAL_5940;
  assign _EVAL_4609 = _EVAL_1362 & 32'h605f;
  assign _EVAL_4707 = _EVAL_4609 == 32'h3;
  assign _EVAL_3025 = _EVAL_5200 | _EVAL_4707;
  assign _EVAL_4785 = _EVAL_4881 == 32'h3;
  assign _EVAL_4238 = _EVAL_3025 | _EVAL_4785;
  assign _EVAL_4990 = _EVAL_6039 ? 1'h0 : _EVAL_4238;
  assign _EVAL_500 = _EVAL_2666[12:5];
  assign _EVAL_5914 = _EVAL_500 != 8'h0;
  assign _EVAL_1909 = _EVAL_630 ? 1'h1 : _EVAL_5914;
  assign _EVAL_2632 = _EVAL_1014 ? 1'h1 : _EVAL_1909;
  assign _EVAL_2474 = _EVAL_4352 ? 1'h1 : _EVAL_2632;
  assign _EVAL_5256 = _EVAL_4202 ? 1'h1 : _EVAL_2474;
  assign _EVAL_326 = _EVAL_2644 ? 1'h1 : _EVAL_5256;
  assign _EVAL_902 = _EVAL_5821 ? 1'h1 : _EVAL_326;
  assign _EVAL_3055 = _EVAL_418 ? 1'h1 : _EVAL_902;
  assign _EVAL_1833 = _EVAL_3055 == 1'h0;
  assign _EVAL_5134 = _EVAL_3271 & 32'hfff0007f;
  assign _EVAL_5682 = _EVAL_5134 == 32'h58000053;
  assign _EVAL_4477 = _EVAL_3398 | _EVAL_5682;
  assign _EVAL_4705 = _EVAL_4477 | _EVAL_4108;
  assign _EVAL_847 = _EVAL_4705 | _EVAL_778;
  assign _EVAL_4527 = _EVAL_3271 & 32'hfff0607f;
  assign _EVAL_5921 = _EVAL_4527 == 32'he0000053;
  assign _EVAL_1354 = _EVAL_847 | _EVAL_5921;
  assign _EVAL_547 = _EVAL_3271 & 32'heff0707f;
  assign _EVAL_4102 = _EVAL_547 == 32'he0000053;
  assign _EVAL_3663 = _EVAL_1354 | _EVAL_4102;
  assign _EVAL_1741 = _EVAL_3663 | _EVAL_4598;
  assign _EVAL_5757 = _EVAL_3271 & 32'h306f;
  assign _EVAL_3725 = _EVAL_5757 == 32'h1063;
  assign _EVAL_2136 = _EVAL_1741 | _EVAL_3725;
  assign _EVAL_5782 = _EVAL_2136 | _EVAL_3136;
  assign _EVAL_2426 = _EVAL_3271 & 32'h605f;
  assign _EVAL_5791 = _EVAL_2426 == 32'h3;
  assign _EVAL_4253 = _EVAL_5782 | _EVAL_5791;
  assign _EVAL_1873 = _EVAL_5757 == 32'h3;
  assign _EVAL_2085 = _EVAL_4253 | _EVAL_1873;
  assign _EVAL_2871 = _EVAL_1833 ? 1'h0 : _EVAL_2085;
  assign _EVAL_6127 = _EVAL_668 ? _EVAL_4990 : _EVAL_2871;
  assign _EVAL_1952 = _EVAL_3050 ? _EVAL_4886 : _EVAL_6127;
  assign _EVAL_5619 = _EVAL_1069 ? _EVAL_4886 : _EVAL_1952;
  assign _EVAL_178 = _EVAL_2142 ? _EVAL_3108 : _EVAL_5619;
  assign _EVAL_2300 = _EVAL_3052 ? _EVAL_6030 : _EVAL_178;
  assign _EVAL_1750 = _EVAL_5276 ? _EVAL_4296 : _EVAL_2300;
  assign _EVAL_2508 = _EVAL_1362 & 32'h40000040;
  assign _EVAL_4865 = _EVAL_2039 & 32'h28;
  assign _EVAL_2126 = _EVAL_4865 == 32'h28;
  assign _EVAL_5131 = _EVAL_5133 & 32'h2000040;
  assign _EVAL_1037 = _EVAL_5131 == 32'h0;
  assign _EVAL_3527 = _EVAL_5133 & 32'h60;
  assign _EVAL_1608 = _EVAL_3527 == 32'h0;
  assign _EVAL_4438 = _EVAL_1037 | _EVAL_1608;
  assign _EVAL_1704 = _EVAL_2680 == 32'h0;
  assign _EVAL_1304 = _EVAL_4438 | _EVAL_1704;
  assign _EVAL_3936 = _EVAL_3875 == 32'h4;
  assign _EVAL_4222 = _EVAL_1304 | _EVAL_3936;
  assign _EVAL_5052 = _EVAL_52 & _EVAL_26;
  assign _EVAL_1850 = _EVAL_1362 & 32'h20000040;
  assign _EVAL_792 = {_EVAL_1802,_EVAL_1321};
  assign _EVAL_4765 = _EVAL_2039[6:2];
  assign _EVAL_3551 = _EVAL_1242[6:2];
  assign _EVAL_1847 = _EVAL_2164[6:2];
  assign _EVAL_421 = _EVAL_1074 ? _EVAL_3551 : _EVAL_1847;
  assign _EVAL_3913 = _EVAL_5926 ? _EVAL_4765 : _EVAL_421;
  assign _EVAL_1710 = _EVAL_2970 ? _EVAL_4765 : _EVAL_3913;
  assign _EVAL_698 = _EVAL_2970 ? _EVAL_2075 : _EVAL_1710;
  assign _EVAL_1434 = _EVAL_3524 & _EVAL_5187;
  assign _EVAL_5378 = _EVAL_2110 & _EVAL_1434;
  assign _EVAL_4579 = _EVAL_6084 == 32'h0;
  assign _EVAL_612 = _EVAL_4821 == 32'h0;
  assign _EVAL_198 = _EVAL_612 | _EVAL_5272;
  assign _EVAL_6078 = _EVAL_198 | _EVAL_2258;
  assign _EVAL_1945 = _EVAL_888 & 32'h28;
  assign _EVAL_2119 = _EVAL_1945 == 32'h28;
  assign _EVAL_1782 = _EVAL_6078 | _EVAL_2119;
  assign _EVAL_6109 = _EVAL_888 & 32'h30;
  assign _EVAL_4610 = _EVAL_6109 == 32'h30;
  assign _EVAL_729 = _EVAL_1782 | _EVAL_4610;
  assign _EVAL_4870 = _EVAL_888 & 32'h90000010;
  assign _EVAL_4735 = _EVAL_4870 == 32'h80000010;
  assign _EVAL_4019 = _EVAL_729 | _EVAL_4735;
  assign _EVAL_1174 = _EVAL_5057 != 5'h0;
  assign _EVAL_1492 = _EVAL_4019 & _EVAL_1174;
  assign _EVAL_5878 = _EVAL_4743[11:7];
  assign _EVAL_1797 = _EVAL_5878 != 5'h0;
  assign _EVAL_1340 = _EVAL_2900 & _EVAL_1797;
  assign _EVAL_1248 = _EVAL_386 & 32'h90000010;
  assign _EVAL_425 = _EVAL_1248 == 32'h80000010;
  assign _EVAL_1828 = _EVAL_1835 | _EVAL_425;
  assign _EVAL_6087 = _EVAL_386[11:7];
  assign _EVAL_4955 = _EVAL_6087 != 5'h0;
  assign _EVAL_541 = _EVAL_1828 & _EVAL_4955;
  assign _EVAL_3563 = _EVAL_5952 ? _EVAL_1340 : _EVAL_541;
  assign _EVAL_1827 = _EVAL_3570 ? _EVAL_1492 : _EVAL_3563;
  assign _EVAL_4454 = _EVAL_5833 ? _EVAL_1492 : _EVAL_1827;
  assign _EVAL_4416 = _EVAL_3461 >= 3'h4;
  assign _EVAL_1105 = _EVAL_1226 | _EVAL_1930;
  assign _EVAL_465 = _EVAL_1105 | _EVAL_5337;
  assign _EVAL_1185 = _EVAL_465 | _EVAL_5985;
  assign _EVAL_4381 = 1'h1 + _EVAL_5833;
  assign _EVAL_5481 = {{1'd0}, _EVAL_2970};
  assign _EVAL_3299 = 2'h2 + _EVAL_5481;
  assign _EVAL_2638 = {{1'd0}, _EVAL_5690};
  assign _EVAL_298 = 2'h3 + _EVAL_2638;
  assign _EVAL_184 = _EVAL_5337 ? {{1'd0}, _EVAL_298} : 4'h4;
  assign _EVAL_3061 = _EVAL_1930 ? {{1'd0}, _EVAL_3299} : _EVAL_184;
  assign _EVAL_1472 = _EVAL_1226 ? {{2'd0}, _EVAL_4381} : _EVAL_3061;
  assign _EVAL_722 = {{1'd0}, _EVAL_197};
  assign _EVAL_2791 = _EVAL_2142 ? {{1'd0}, _EVAL_298} : 4'h4;
  assign _EVAL_712 = _EVAL_3052 ? {{1'd0}, _EVAL_3299} : _EVAL_2791;
  assign _EVAL_6085 = _EVAL_5276 ? {{2'd0}, _EVAL_4381} : _EVAL_712;
  assign _EVAL_2943 = _EVAL_5994 ? {{2'd0}, _EVAL_722} : _EVAL_6085;
  assign _EVAL_693 = _EVAL_1185 ? _EVAL_1472 : _EVAL_2943;
  assign _EVAL_358 = _EVAL_693 == 4'h3;
  assign _EVAL_5859 = _EVAL_4416 & _EVAL_358;
  assign _EVAL_3810 = _EVAL_2485 | _EVAL_5859;
  assign _EVAL_5126 = _EVAL_5854 & 32'h10000060;
  assign _EVAL_1616 = _EVAL_5126 == 32'h40;
  assign _EVAL_2543 = _EVAL_1267 | _EVAL_1616;
  assign _EVAL_511 = _EVAL_1978 & 32'h3c;
  assign _EVAL_1449 = _EVAL_511 == 32'h4;
  assign _EVAL_2588 = _EVAL_1978 & 32'h80000060;
  assign _EVAL_4051 = _EVAL_2588 == 32'h40;
  assign _EVAL_2230 = _EVAL_1449 | _EVAL_4051;
  assign _EVAL_2767 = _EVAL_2230 | _EVAL_4329;
  assign _EVAL_2931 = _EVAL_1978 & 32'h10000060;
  assign _EVAL_2704 = _EVAL_2931 == 32'h10000040;
  assign _EVAL_3258 = _EVAL_2767 | _EVAL_2704;
  assign _EVAL_5486 = _EVAL_1362 & 32'h3c;
  assign _EVAL_4251 = _EVAL_5486 == 32'h4;
  assign _EVAL_417 = _EVAL_4251 | _EVAL_3482;
  assign _EVAL_4058 = _EVAL_417 | _EVAL_4770;
  assign _EVAL_2376 = _EVAL_3898 == 32'h10000040;
  assign _EVAL_3626 = _EVAL_4058 | _EVAL_2376;
  assign _EVAL_1487 = _EVAL_1415 | _EVAL_3564;
  assign _EVAL_5650 = _EVAL_1487 | _EVAL_1739;
  assign _EVAL_4508 = _EVAL_3842 == 32'h10000040;
  assign _EVAL_3716 = _EVAL_5650 | _EVAL_4508;
  assign _EVAL_3878 = _EVAL_668 ? _EVAL_3626 : _EVAL_3716;
  assign _EVAL_2345 = _EVAL_3050 ? _EVAL_3258 : _EVAL_3878;
  assign _EVAL_5027 = _EVAL_3065 == 32'h20;
  assign _EVAL_3934 = _EVAL_3006 & 32'h34;
  assign _EVAL_4249 = _EVAL_3934 == 32'h20;
  assign _EVAL_325 = _EVAL_5027 | _EVAL_4249;
  assign _EVAL_2689 = _EVAL_4702 & 32'hf600607f;
  assign _EVAL_5290 = _EVAL_2689 == 32'h20000053;
  assign _EVAL_3540 = _EVAL_1362 & 32'h2040;
  assign _EVAL_3384 = _EVAL_3540 == 32'h2040;
  assign _EVAL_1180 = _EVAL_4402 == 32'he0000053;
  assign _EVAL_1659 = _EVAL_3078 & 32'h50;
  assign _EVAL_2747 = _EVAL_1659 == 32'h40;
  assign _EVAL_4736 = _EVAL_352 & _EVAL_3323;
  assign _EVAL_2569 = _EVAL_3524 & _EVAL_1696;
  assign _EVAL_3566 = _EVAL_2110 & _EVAL_2569;
  assign _EVAL_5333 = _EVAL_5875 | _EVAL_3728;
  assign _EVAL_5518 = _EVAL_3566 & _EVAL_5333;
  assign _EVAL_811 = _EVAL_4736 ? 1'h1 : _EVAL_5518;
  assign _EVAL_4682 = _EVAL_1660 ? 1'h1 : _EVAL_811;
  assign _EVAL_3740 = _EVAL_5813 & 32'h64;
  assign _EVAL_3167 = _EVAL_3740 == 32'h20;
  assign _EVAL_318 = _EVAL_5813 & 32'h34;
  assign _EVAL_2049 = _EVAL_318 == 32'h20;
  assign _EVAL_1529 = _EVAL_3167 | _EVAL_2049;
  assign _EVAL_339 = _EVAL_5813 & 32'h2048;
  assign _EVAL_1156 = _EVAL_339 == 32'h2008;
  assign _EVAL_2823 = _EVAL_1529 | _EVAL_1156;
  assign _EVAL_5735 = _EVAL_5813 & 32'h4003044;
  assign _EVAL_4792 = _EVAL_5735 == 32'h4000040;
  assign _EVAL_1148 = _EVAL_2823 | _EVAL_4792;
  assign _EVAL_4898 = _EVAL_621 == 32'h20;
  assign _EVAL_4384 = _EVAL_1947 & 32'h34;
  assign _EVAL_5838 = _EVAL_4384 == 32'h20;
  assign _EVAL_669 = _EVAL_4898 | _EVAL_5838;
  assign _EVAL_1426 = _EVAL_1947 & 32'h2048;
  assign _EVAL_1964 = _EVAL_1426 == 32'h2008;
  assign _EVAL_4376 = _EVAL_669 | _EVAL_1964;
  assign _EVAL_1143 = _EVAL_1947 & 32'h4003044;
  assign _EVAL_2661 = _EVAL_1143 == 32'h4000040;
  assign _EVAL_4778 = _EVAL_4376 | _EVAL_2661;
  assign _EVAL_2812 = _EVAL_1958 ? _EVAL_1148 : _EVAL_4778;
  assign _EVAL_835 = _EVAL_4268 & 32'h62003010;
  assign _EVAL_5954 = _EVAL_835 == 32'h60000010;
  assign _EVAL_5161 = _EVAL_5697 | _EVAL_5954;
  assign _EVAL_2226 = _EVAL_3006 & 32'h2000040;
  assign _EVAL_4690 = _EVAL_2226 == 32'h0;
  assign _EVAL_323 = _EVAL_3006 & 32'h60;
  assign _EVAL_1998 = _EVAL_323 == 32'h0;
  assign _EVAL_4797 = _EVAL_4690 | _EVAL_1998;
  assign _EVAL_4196 = _EVAL_3952 == 32'h0;
  assign _EVAL_1271 = _EVAL_4797 | _EVAL_4196;
  assign _EVAL_6093 = _EVAL_3006 & 32'h44;
  assign _EVAL_1806 = _EVAL_6093 == 32'h4;
  assign _EVAL_1232 = _EVAL_1271 | _EVAL_1806;
  assign _EVAL_4957 = _EVAL_3006 & 32'h62003010;
  assign _EVAL_4091 = _EVAL_4957 == 32'h60000010;
  assign _EVAL_3763 = _EVAL_1232 | _EVAL_4091;
  assign _EVAL_4245 = _EVAL_1757 == 32'h0;
  assign _EVAL_3274 = _EVAL_2911 | _EVAL_4245;
  assign _EVAL_4029 = _EVAL_3274 | _EVAL_3011;
  assign _EVAL_3912 = _EVAL_6032 == 32'h60000010;
  assign _EVAL_5599 = _EVAL_4029 | _EVAL_3912;
  assign _EVAL_3542 = _EVAL_5820 == 32'h60000010;
  assign _EVAL_1396 = _EVAL_4222 | _EVAL_3542;
  assign _EVAL_992 = _EVAL_2901 ? _EVAL_5599 : _EVAL_1396;
  assign _EVAL_1238 = _EVAL_2378 ? _EVAL_3763 : _EVAL_992;
  assign _EVAL_1234 = _EVAL_5690 ? _EVAL_3763 : _EVAL_1238;
  assign _EVAL_953 = _EVAL_5690 ? _EVAL_5161 : _EVAL_1234;
  assign _EVAL_1976 = _EVAL_1978 & 32'h2000040;
  assign _EVAL_4028 = _EVAL_1976 == 32'h0;
  assign _EVAL_2537 = _EVAL_1978 & 32'h60;
  assign _EVAL_395 = _EVAL_2537 == 32'h0;
  assign _EVAL_6067 = _EVAL_4028 | _EVAL_395;
  assign _EVAL_5798 = _EVAL_596 == 32'h0;
  assign _EVAL_671 = _EVAL_6067 | _EVAL_5798;
  assign _EVAL_6079 = _EVAL_1978 & 32'h44;
  assign _EVAL_5025 = _EVAL_6079 == 32'h4;
  assign _EVAL_5425 = _EVAL_671 | _EVAL_5025;
  assign _EVAL_195 = _EVAL_5425 | _EVAL_5442;
  assign _EVAL_982 = _EVAL_1362 & 32'h2000040;
  assign _EVAL_3201 = _EVAL_982 == 32'h0;
  assign _EVAL_916 = _EVAL_1362 & 32'h60;
  assign _EVAL_5407 = _EVAL_916 == 32'h0;
  assign _EVAL_2549 = _EVAL_3201 | _EVAL_5407;
  assign _EVAL_3813 = _EVAL_1362 & 32'h50;
  assign _EVAL_5263 = _EVAL_3813 == 32'h0;
  assign _EVAL_3536 = _EVAL_2549 | _EVAL_5263;
  assign _EVAL_3084 = _EVAL_1096 == 32'h4;
  assign _EVAL_5683 = _EVAL_3536 | _EVAL_3084;
  assign _EVAL_4819 = _EVAL_1362 & 32'h62003010;
  assign _EVAL_3317 = _EVAL_4819 == 32'h60000010;
  assign _EVAL_4272 = _EVAL_5683 | _EVAL_3317;
  assign _EVAL_5513 = _EVAL_3271 & 32'h2000040;
  assign _EVAL_5856 = _EVAL_5513 == 32'h0;
  assign _EVAL_552 = _EVAL_3271 & 32'h60;
  assign _EVAL_2753 = _EVAL_552 == 32'h0;
  assign _EVAL_5108 = _EVAL_5856 | _EVAL_2753;
  assign _EVAL_2165 = _EVAL_4387 == 32'h0;
  assign _EVAL_5587 = _EVAL_5108 | _EVAL_2165;
  assign _EVAL_3687 = _EVAL_3682 == 32'h4;
  assign _EVAL_6061 = _EVAL_5587 | _EVAL_3687;
  assign _EVAL_5963 = _EVAL_3271 & 32'h62003010;
  assign _EVAL_2729 = _EVAL_5963 == 32'h60000010;
  assign _EVAL_1738 = _EVAL_6061 | _EVAL_2729;
  assign _EVAL_4949 = _EVAL_668 ? _EVAL_4272 : _EVAL_1738;
  assign _EVAL_5764 = _EVAL_3050 ? _EVAL_195 : _EVAL_4949;
  assign _EVAL_5129 = _EVAL_1069 ? _EVAL_195 : _EVAL_5764;
  assign _EVAL_5299 = _EVAL_5337 ? _EVAL_953 : _EVAL_5129;
  assign _EVAL_4861 = _EVAL_3006 & 32'h3c;
  assign _EVAL_3085 = _EVAL_4861 == 32'h4;
  assign _EVAL_5819 = _EVAL_5854 & 32'h70;
  assign _EVAL_2953 = _EVAL_5819 == 32'h40;
  assign _EVAL_2682 = _EVAL_2543 | _EVAL_2953;
  assign _EVAL_2828 = _EVAL_888 & 32'h80000060;
  assign _EVAL_3007 = _EVAL_2828 == 32'h40;
  assign _EVAL_655 = _EVAL_3007 | _EVAL_2973;
  assign _EVAL_6099 = _EVAL_655 | _EVAL_697;
  assign _EVAL_4519 = _EVAL_386 & 32'h80000060;
  assign _EVAL_2158 = _EVAL_4519 == 32'h40;
  assign _EVAL_4274 = _EVAL_386 & 32'h10000060;
  assign _EVAL_3191 = _EVAL_4274 == 32'h40;
  assign _EVAL_4156 = _EVAL_2158 | _EVAL_3191;
  assign _EVAL_226 = _EVAL_4156 | _EVAL_4271;
  assign _EVAL_5850 = _EVAL_5952 ? _EVAL_3238 : _EVAL_226;
  assign _EVAL_5460 = _EVAL_3570 ? _EVAL_6099 : _EVAL_5850;
  assign _EVAL_3368 = _EVAL_5833 ? _EVAL_6099 : _EVAL_5460;
  assign _EVAL_5955 = _EVAL_5833 ? _EVAL_2682 : _EVAL_3368;
  assign _EVAL_853 = _EVAL_5311 & 32'h80000060;
  assign _EVAL_2679 = _EVAL_853 == 32'h40;
  assign _EVAL_4566 = _EVAL_1974 == 32'h40;
  assign _EVAL_6100 = _EVAL_2679 | _EVAL_4566;
  assign _EVAL_3714 = _EVAL_5311 & 32'h70;
  assign _EVAL_5728 = _EVAL_3714 == 32'h40;
  assign _EVAL_1596 = _EVAL_6100 | _EVAL_5728;
  assign _EVAL_3977 = _EVAL_2039 & 32'h80000060;
  assign _EVAL_3476 = _EVAL_3977 == 32'h40;
  assign _EVAL_5526 = _EVAL_2039 & 32'h10000060;
  assign _EVAL_5598 = _EVAL_5526 == 32'h40;
  assign _EVAL_434 = _EVAL_3476 | _EVAL_5598;
  assign _EVAL_3825 = _EVAL_2039 & 32'h70;
  assign _EVAL_3653 = _EVAL_3825 == 32'h40;
  assign _EVAL_3555 = _EVAL_434 | _EVAL_3653;
  assign _EVAL_3316 = _EVAL_2500 == 32'h40;
  assign _EVAL_4520 = _EVAL_1868 | _EVAL_3316;
  assign _EVAL_220 = _EVAL_4520 | _EVAL_677;
  assign _EVAL_2094 = _EVAL_2154 | _EVAL_4890;
  assign _EVAL_4672 = _EVAL_1074 ? _EVAL_220 : _EVAL_2094;
  assign _EVAL_1943 = _EVAL_5926 ? _EVAL_3555 : _EVAL_4672;
  assign _EVAL_3181 = _EVAL_2970 ? _EVAL_3555 : _EVAL_1943;
  assign _EVAL_2565 = _EVAL_2970 ? _EVAL_1596 : _EVAL_3181;
  assign _EVAL_4757 = _EVAL_4268 & 32'h10000060;
  assign _EVAL_2065 = _EVAL_4757 == 32'h40;
  assign _EVAL_385 = _EVAL_3788 | _EVAL_2065;
  assign _EVAL_1872 = _EVAL_4268 & 32'h70;
  assign _EVAL_4912 = _EVAL_1872 == 32'h40;
  assign _EVAL_3185 = _EVAL_385 | _EVAL_4912;
  assign _EVAL_1561 = _EVAL_5690 ? _EVAL_3185 : _EVAL_4190;
  assign _EVAL_4549 = _EVAL_2931 == 32'h40;
  assign _EVAL_3773 = _EVAL_4051 | _EVAL_4549;
  assign _EVAL_1932 = _EVAL_3773 | _EVAL_4329;
  assign _EVAL_5177 = _EVAL_3050 ? _EVAL_1932 : _EVAL_4969;
  assign _EVAL_2395 = _EVAL_1069 ? _EVAL_1932 : _EVAL_5177;
  assign _EVAL_235 = _EVAL_2142 ? _EVAL_1561 : _EVAL_2395;
  assign _EVAL_3601 = _EVAL_3052 ? _EVAL_2565 : _EVAL_235;
  assign _EVAL_4378 = _EVAL_5276 ? _EVAL_5955 : _EVAL_3601;
  assign _EVAL_3161 = _EVAL_5641 == 32'h90000010;
  assign _EVAL_5436 = _EVAL_386 & 32'h40000060;
  assign _EVAL_5751 = _EVAL_5875 | _EVAL_3508;
  assign _EVAL_2227 = _EVAL_5378 & _EVAL_5751;
  assign _EVAL_4981 = _EVAL_3460 ? 1'h1 : _EVAL_2227;
  assign _EVAL_3664 = _EVAL_5135 ? 1'h1 : _EVAL_4981;
  assign _EVAL_984 = _EVAL_4922 & _EVAL_2213;
  assign _EVAL_5018 = _EVAL_2110 & _EVAL_984;
  assign _EVAL_5169 = _EVAL_5875 | _EVAL_5140;
  assign _EVAL_5148 = _EVAL_5018 & _EVAL_5169;
  assign _EVAL_2562 = _EVAL_5875 | _EVAL_239;
  assign _EVAL_3176 = _EVAL_1342 & _EVAL_2562;
  assign _EVAL_1626 = _EVAL_5148 ? 1'h1 : _EVAL_3176;
  assign _EVAL_727 = _EVAL_1826 ? 1'h1 : _EVAL_1626;
  assign _EVAL_3900 = {_EVAL_4682,_EVAL_881,_EVAL_3664,_EVAL_727};
  assign _EVAL_5125 = _EVAL_3900 & _EVAL_4984;
  assign _EVAL_1020 = _EVAL_730 != 11'h0;
  assign _EVAL_3804 = _EVAL_761 ? 1'h1 : _EVAL_1578;
  assign _EVAL_773 = _EVAL_4440 ? _EVAL_1020 : _EVAL_3804;
  assign _EVAL_917 = _EVAL_1378 ? 1'h1 : _EVAL_773;
  assign _EVAL_275 = _EVAL_537 ? 1'h1 : _EVAL_917;
  assign _EVAL_1427 = _EVAL_1088 ? 1'h1 : _EVAL_275;
  assign _EVAL_4095 = _EVAL_1427 == 1'h0;
  assign _EVAL_4794 = _EVAL_1259 == 32'h0;
  assign _EVAL_631 = _EVAL_4794 | _EVAL_1275;
  assign _EVAL_5911 = _EVAL_2039 & 32'h2024;
  assign _EVAL_1562 = _EVAL_5911 == 32'h24;
  assign _EVAL_1774 = _EVAL_631 | _EVAL_1562;
  assign _EVAL_556 = _EVAL_1774 | _EVAL_2126;
  assign _EVAL_910 = _EVAL_1659 == 32'h10;
  assign _EVAL_5865 = _EVAL_888 & 32'h8000040;
  assign _EVAL_444 = _EVAL_5865 == 32'h8000040;
  assign _EVAL_3647 = _EVAL_386 & 32'h20000040;
  assign _EVAL_507 = _EVAL_3647 == 32'h40;
  assign _EVAL_217 = _EVAL_232 == 32'h20;
  assign _EVAL_2472 = _EVAL_4882 & 32'h34;
  assign _EVAL_1509 = _EVAL_2472 == 32'h20;
  assign _EVAL_5307 = _EVAL_217 | _EVAL_1509;
  assign _EVAL_5073 = 3'h0 < _EVAL_3461;
  assign _EVAL_3805 = _EVAL_1226 & _EVAL_5073;
  assign _EVAL_3269 = 3'h1 < _EVAL_3461;
  assign _EVAL_5704 = _EVAL_1930 & _EVAL_3269;
  assign _EVAL_799 = _EVAL_3805 | _EVAL_5704;
  assign _EVAL_225 = _EVAL_1978 & 32'h8000040;
  assign _EVAL_4479 = _EVAL_2970 ? _EVAL_5601 : _EVAL_2076;
  assign _EVAL_4975 = _EVAL_1947 & 32'h2024;
  assign _EVAL_1344 = _EVAL_4975 == 32'h24;
  assign _EVAL_793 = _EVAL_3713 | _EVAL_1344;
  assign _EVAL_3227 = _EVAL_1947 & 32'h2000040;
  assign _EVAL_2504 = _EVAL_3227 == 32'h0;
  assign _EVAL_1404 = _EVAL_1947 & 32'h60;
  assign _EVAL_4907 = _EVAL_1404 == 32'h0;
  assign _EVAL_3220 = _EVAL_2504 | _EVAL_4907;
  assign _EVAL_5091 = _EVAL_1550 == 32'h0;
  assign _EVAL_2787 = _EVAL_3220 | _EVAL_5091;
  assign _EVAL_1410 = _EVAL_2583 == 32'h4;
  assign _EVAL_1139 = _EVAL_2787 | _EVAL_1410;
  assign _EVAL_5974 = _EVAL_5311 & 32'h64;
  assign _EVAL_956 = _EVAL_5974 == 32'h20;
  assign _EVAL_5098 = _EVAL_956 | _EVAL_1460;
  assign _EVAL_1796 = _EVAL_5311 & 32'h2048;
  assign _EVAL_5571 = _EVAL_1796 == 32'h2008;
  assign _EVAL_3603 = _EVAL_5098 | _EVAL_5571;
  assign _EVAL_967 = _EVAL_4882 & 32'h2040;
  assign _EVAL_6115 = _EVAL_136 | 32'h6;
  assign _EVAL_3289 = _EVAL_2801 & _EVAL_5575;
  assign _EVAL_5399 = 29'h0 < _EVAL_5201;
  assign _EVAL_1373 = _EVAL_4978 & _EVAL_2374;
  assign _EVAL_2705 = _EVAL_5399 | _EVAL_1373;
  assign _EVAL_3353 = _EVAL_2705 == _EVAL_383;
  assign _EVAL_3938 = _EVAL_4978 & _EVAL_5997;
  assign _EVAL_2124 = _EVAL_519 ? _EVAL_3353 : _EVAL_3938;
  assign _EVAL_3283 = _EVAL_3289 & _EVAL_2124;
  assign _EVAL_5090 = _EVAL_2164 & 32'h64;
  assign _EVAL_1258 = _EVAL_5090 == 32'h0;
  assign _EVAL_4270 = _EVAL_1258 | _EVAL_2233;
  assign _EVAL_851 = _EVAL_2164 & 32'h2024;
  assign _EVAL_4331 = _EVAL_851 == 32'h24;
  assign _EVAL_4850 = _EVAL_4270 | _EVAL_4331;
  assign _EVAL_2861 = _EVAL_2164 & 32'h28;
  assign _EVAL_3110 = _EVAL_2861 == 32'h28;
  assign _EVAL_4165 = _EVAL_4850 | _EVAL_3110;
  assign _EVAL_2041 = _EVAL_4165 | _EVAL_1495;
  assign _EVAL_5471 = _EVAL_2164 & 32'h90000010;
  assign _EVAL_4124 = _EVAL_5471 == 32'h80000010;
  assign _EVAL_3683 = _EVAL_2041 | _EVAL_4124;
  assign _EVAL_5267 = _EVAL_3256 != 5'h0;
  assign _EVAL_3633 = _EVAL_3683 & _EVAL_5267;
  assign _EVAL_4684 = _EVAL_4743 & 32'h62003010;
  assign _EVAL_2133 = _EVAL_4684 == 32'h60000010;
  assign _EVAL_1253 = _EVAL_888 & 32'h2000040;
  assign _EVAL_1359 = _EVAL_1253 == 32'h0;
  assign _EVAL_4341 = _EVAL_888 & 32'h60;
  assign _EVAL_4121 = _EVAL_4341 == 32'h0;
  assign _EVAL_4287 = _EVAL_1359 | _EVAL_4121;
  assign _EVAL_3512 = _EVAL_4471 == 32'h0;
  assign _EVAL_4921 = _EVAL_4287 | _EVAL_3512;
  assign _EVAL_3145 = _EVAL_3078 & 32'h7c;
  assign _EVAL_6057 = _EVAL_3145 == 32'h24;
  assign _EVAL_2024 = _EVAL_3078 & 32'h40000060;
  assign _EVAL_1220 = _EVAL_2024 == 32'h40;
  assign _EVAL_6062 = _EVAL_6057 | _EVAL_1220;
  assign _EVAL_1223 = _EVAL_3078 & 32'h70;
  assign _EVAL_2310 = _EVAL_1223 == 32'h40;
  assign _EVAL_616 = _EVAL_6062 | _EVAL_2310;
  assign _EVAL_2103 = _EVAL_2610 == 32'h24;
  assign _EVAL_1457 = _EVAL_5813 & 32'h40000060;
  assign _EVAL_242 = _EVAL_1457 == 32'h40;
  assign _EVAL_361 = _EVAL_2103 | _EVAL_242;
  assign _EVAL_469 = _EVAL_361 | _EVAL_2596;
  assign _EVAL_370 = _EVAL_1947 & 32'h7c;
  assign _EVAL_2756 = _EVAL_370 == 32'h24;
  assign _EVAL_1042 = _EVAL_1947 & 32'h40000060;
  assign _EVAL_2636 = _EVAL_1042 == 32'h40;
  assign _EVAL_369 = _EVAL_2756 | _EVAL_2636;
  assign _EVAL_2212 = _EVAL_1947 & 32'h70;
  assign _EVAL_160 = _EVAL_2212 == 32'h40;
  assign _EVAL_2836 = _EVAL_369 | _EVAL_160;
  assign _EVAL_4614 = _EVAL_1958 ? _EVAL_469 : _EVAL_2836;
  assign _EVAL_3651 = _EVAL_4554 ? _EVAL_616 : _EVAL_4614;
  assign _EVAL_4258 = _EVAL_197 ? _EVAL_616 : _EVAL_3651;
  assign _EVAL_1919 = _EVAL_4743 & 32'h2040;
  assign _EVAL_648 = _EVAL_2703 | _EVAL_3379;
  assign _EVAL_4369 = _EVAL_1978 & 32'h30;
  assign _EVAL_1735 = _EVAL_4369 == 32'h30;
  assign _EVAL_1878 = _EVAL_648 | _EVAL_1735;
  assign _EVAL_1228 = _EVAL_1978 & 32'h90000010;
  assign _EVAL_4811 = _EVAL_1228 == 32'h80000010;
  assign _EVAL_302 = _EVAL_1878 | _EVAL_4811;
  assign _EVAL_3589 = _EVAL_4087 == 32'h0;
  assign _EVAL_5341 = _EVAL_1978 & 32'h38;
  assign _EVAL_2276 = _EVAL_386 & 32'h38;
  assign _EVAL_768 = _EVAL_2276 == 32'h20;
  assign _EVAL_1222 = _EVAL_1451 & _EVAL_3876;
  assign _EVAL_2590 = _EVAL_5062 | _EVAL_1222;
  assign _EVAL_5361 = _EVAL_2590 == _EVAL_1969;
  assign _EVAL_2951 = _EVAL_1451 & _EVAL_3445;
  assign _EVAL_2963 = _EVAL_4291 ? _EVAL_5361 : _EVAL_2951;
  assign _EVAL_254 = _EVAL_1986 & _EVAL_2963;
  assign _EVAL_2211 = _EVAL_574 | _EVAL_254;
  assign _EVAL_5410 = _EVAL_3271 & 32'h90000010;
  assign _EVAL_1730 = _EVAL_5410 == 32'h80000010;
  assign _EVAL_4906 = _EVAL_2326 | _EVAL_1730;
  assign _EVAL_872 = _EVAL_4268 & 32'h4003044;
  assign _EVAL_3958 = _EVAL_5283 == 32'h20;
  assign _EVAL_2224 = _EVAL_4743 & 32'h34;
  assign _EVAL_2339 = _EVAL_2224 == 32'h20;
  assign _EVAL_6135 = _EVAL_3958 | _EVAL_2339;
  assign _EVAL_1981 = _EVAL_4743 & 32'h2048;
  assign _EVAL_4406 = _EVAL_1981 == 32'h2008;
  assign _EVAL_1772 = _EVAL_6135 | _EVAL_4406;
  assign _EVAL_4469 = _EVAL_888[31:25];
  assign _EVAL_3817 = _EVAL_4743[31:25];
  assign _EVAL_2894 = _EVAL_386[31:25];
  assign _EVAL_5628 = _EVAL_5952 ? _EVAL_3817 : _EVAL_2894;
  assign _EVAL_3488 = _EVAL_3570 ? _EVAL_4469 : _EVAL_5628;
  assign _EVAL_2929 = _EVAL_5854 & 32'h3c;
  assign _EVAL_3994 = _EVAL_2039 & 32'h30;
  assign _EVAL_3866 = _EVAL_3994 == 32'h30;
  assign _EVAL_5630 = _EVAL_556 | _EVAL_3866;
  assign _EVAL_1654 = _EVAL_2039 & 32'h90000010;
  assign _EVAL_1931 = _EVAL_1654 == 32'h80000010;
  assign _EVAL_864 = _EVAL_5630 | _EVAL_1931;
  assign _EVAL_490 = _EVAL_2164[31:25];
  assign _EVAL_3042 = _EVAL_5813 & 32'h20000040;
  assign _EVAL_4787 = _EVAL_3042 == 32'h40;
  assign _EVAL_4057 = _EVAL_362 == 32'h20;
  assign _EVAL_1313 = _EVAL_4268 & 32'h34;
  assign _EVAL_330 = _EVAL_1313 == 32'h20;
  assign _EVAL_2000 = _EVAL_4057 | _EVAL_330;
  assign _EVAL_1133 = _EVAL_4268 & 32'h2048;
  assign _EVAL_5927 = _EVAL_1133 == 32'h2008;
  assign _EVAL_5269 = _EVAL_2000 | _EVAL_5927;
  assign _EVAL_2662 = _EVAL_872 == 32'h4000040;
  assign _EVAL_3666 = _EVAL_5269 | _EVAL_2662;
  assign _EVAL_4056 = _EVAL_3065 == 32'h0;
  assign _EVAL_3745 = _EVAL_4056 | _EVAL_4113;
  assign _EVAL_3800 = _EVAL_3006 & 32'h2024;
  assign _EVAL_6076 = _EVAL_3800 == 32'h24;
  assign _EVAL_5431 = _EVAL_3745 | _EVAL_6076;
  assign _EVAL_2365 = _EVAL_3006 & 32'h28;
  assign _EVAL_4157 = _EVAL_2365 == 32'h28;
  assign _EVAL_4688 = _EVAL_5431 | _EVAL_4157;
  assign _EVAL_1260 = _EVAL_3006 & 32'h30;
  assign _EVAL_3964 = _EVAL_1260 == 32'h30;
  assign _EVAL_1648 = _EVAL_4688 | _EVAL_3964;
  assign _EVAL_760 = _EVAL_3006 & 32'h90000010;
  assign _EVAL_4629 = _EVAL_760 == 32'h80000010;
  assign _EVAL_3537 = _EVAL_1648 | _EVAL_4629;
  assign _EVAL_2406 = _EVAL_3271 & 32'h4003044;
  assign _EVAL_1655 = _EVAL_2406 == 32'h4000040;
  assign _EVAL_4934 = _EVAL_5399 | _EVAL_4462;
  assign _EVAL_826 = _EVAL_4934 == _EVAL_383;
  assign _EVAL_2071 = _EVAL_4978 & _EVAL_2939;
  assign _EVAL_3047 = _EVAL_519 ? _EVAL_826 : _EVAL_2071;
  assign _EVAL_2641 = _EVAL_3289 & _EVAL_3047;
  assign _EVAL_201 = _EVAL_2641 & _EVAL_2211;
  assign _EVAL_1070 = _EVAL_1947 & 32'h18;
  assign _EVAL_4653 = _EVAL_1070 == 32'h0;
  assign _EVAL_4322 = _EVAL_4653 | _EVAL_2866;
  assign _EVAL_5406 = _EVAL_1947 & 32'h8000040;
  assign _EVAL_3031 = _EVAL_5406 == 32'h8000040;
  assign _EVAL_6136 = _EVAL_4322 | _EVAL_3031;
  assign _EVAL_4340 = _EVAL_1958 ? _EVAL_2596 : _EVAL_160;
  assign _EVAL_1538 = _EVAL_4554 ? _EVAL_2310 : _EVAL_4340;
  assign _EVAL_3173 = _EVAL_5525 & _EVAL_2963;
  assign _EVAL_4773 = _EVAL_574 | _EVAL_3173;
  assign _EVAL_1168 = _EVAL_1947 & 32'h28;
  assign _EVAL_2884 = _EVAL_1168 == 32'h28;
  assign _EVAL_2766 = _EVAL_793 | _EVAL_2884;
  assign _EVAL_3992 = _EVAL_693[1:0];
  assign _EVAL_5574 = _EVAL_3461[1:0];
  assign _EVAL_3080 = _EVAL_3992 >= _EVAL_5574;
  assign _EVAL_2458 = _EVAL_2508 == 32'h40;
  assign _EVAL_5418 = _EVAL_888 & 32'h3c;
  assign _EVAL_4470 = _EVAL_5386[24:20];
  assign _EVAL_5153 = _EVAL_888[24:20];
  assign _EVAL_5261 = _EVAL_3570 ? _EVAL_5153 : _EVAL_5074;
  assign _EVAL_4919 = _EVAL_5833 ? _EVAL_5153 : _EVAL_5261;
  assign _EVAL_2141 = _EVAL_5833 ? _EVAL_4470 : _EVAL_4919;
  assign _EVAL_3703 = _EVAL_3455[24:20];
  assign _EVAL_2336 = _EVAL_2039[24:20];
  assign _EVAL_4223 = _EVAL_1242[24:20];
  assign _EVAL_2388 = _EVAL_2164[24:20];
  assign _EVAL_1276 = _EVAL_1074 ? _EVAL_4223 : _EVAL_2388;
  assign _EVAL_1593 = _EVAL_5926 ? _EVAL_2336 : _EVAL_1276;
  assign _EVAL_5377 = _EVAL_2970 ? _EVAL_2336 : _EVAL_1593;
  assign _EVAL_3104 = _EVAL_2970 ? _EVAL_3703 : _EVAL_5377;
  assign _EVAL_4491 = _EVAL_4268[24:20];
  assign _EVAL_794 = _EVAL_5690 ? _EVAL_1635 : _EVAL_1332;
  assign _EVAL_4846 = _EVAL_5690 ? _EVAL_4491 : _EVAL_794;
  assign _EVAL_3594 = _EVAL_1978[24:20];
  assign _EVAL_261 = _EVAL_1362[24:20];
  assign _EVAL_166 = _EVAL_3271[24:20];
  assign _EVAL_5965 = _EVAL_668 ? _EVAL_261 : _EVAL_166;
  assign _EVAL_5128 = _EVAL_3050 ? _EVAL_3594 : _EVAL_5965;
  assign _EVAL_3548 = _EVAL_1069 ? _EVAL_3594 : _EVAL_5128;
  assign _EVAL_5492 = _EVAL_2142 ? _EVAL_4846 : _EVAL_3548;
  assign _EVAL_1028 = _EVAL_3052 ? _EVAL_3104 : _EVAL_5492;
  assign _EVAL_2343 = _EVAL_5276 ? _EVAL_2141 : _EVAL_1028;
  assign _EVAL_639 = _EVAL_3271[6:2];
  assign _EVAL_4486 = _EVAL_1947 & 32'h1040;
  assign _EVAL_317 = _EVAL_4486 == 32'h1040;
  assign _EVAL_3969 = _EVAL_2929 == 32'h4;
  assign _EVAL_4339 = _EVAL_3969 | _EVAL_1267;
  assign _EVAL_5572 = _EVAL_4339 | _EVAL_2953;
  assign _EVAL_4585 = _EVAL_1242 & 32'h8000040;
  assign _EVAL_5247 = _EVAL_4978 & _EVAL_1295;
  assign _EVAL_3259 = _EVAL_3006[11:7];
  assign _EVAL_2496 = _EVAL_4882[11:7];
  assign _EVAL_5520 = _EVAL_2901 ? _EVAL_2496 : _EVAL_2839;
  assign _EVAL_3059 = _EVAL_2378 ? _EVAL_3259 : _EVAL_5520;
  assign _EVAL_3828 = _EVAL_4702 & 32'hfff0007f;
  assign _EVAL_1887 = _EVAL_4268 & 32'h18;
  assign _EVAL_400 = _EVAL_1887 == 32'h0;
  assign _EVAL_3140 = _EVAL_4268 & 32'h2010;
  assign _EVAL_2139 = _EVAL_3140 == 32'h2000;
  assign _EVAL_229 = _EVAL_400 | _EVAL_2139;
  assign _EVAL_1338 = _EVAL_4268 & 32'h8000040;
  assign _EVAL_381 = _EVAL_1338 == 32'h8000040;
  assign _EVAL_4320 = _EVAL_229 | _EVAL_381;
  assign _EVAL_928 = _EVAL_2891 == 32'h0;
  assign _EVAL_2717 = _EVAL_928 | _EVAL_910;
  assign _EVAL_3404 = _EVAL_3078 & 32'h2024;
  assign _EVAL_2986 = _EVAL_3404 == 32'h24;
  assign _EVAL_534 = _EVAL_2717 | _EVAL_2986;
  assign _EVAL_5397 = _EVAL_3078 & 32'h28;
  assign _EVAL_1424 = _EVAL_5397 == 32'h28;
  assign _EVAL_4476 = _EVAL_534 | _EVAL_1424;
  assign _EVAL_5016 = _EVAL_3078 & 32'h30;
  assign _EVAL_2906 = _EVAL_5016 == 32'h30;
  assign _EVAL_2631 = _EVAL_4476 | _EVAL_2906;
  assign _EVAL_3629 = _EVAL_3078 & 32'h90000010;
  assign _EVAL_832 = _EVAL_3629 == 32'h80000010;
  assign _EVAL_489 = _EVAL_2631 | _EVAL_832;
  assign _EVAL_4254 = _EVAL_489 & _EVAL_4371;
  assign _EVAL_5986 = _EVAL_3740 == 32'h0;
  assign _EVAL_3248 = _EVAL_3680 == 32'h10;
  assign _EVAL_5445 = _EVAL_5986 | _EVAL_3248;
  assign _EVAL_514 = _EVAL_5813 & 32'h2024;
  assign _EVAL_5157 = _EVAL_514 == 32'h24;
  assign _EVAL_2355 = _EVAL_5445 | _EVAL_5157;
  assign _EVAL_5906 = _EVAL_5813 & 32'h28;
  assign _EVAL_2763 = _EVAL_5906 == 32'h28;
  assign _EVAL_1518 = _EVAL_2355 | _EVAL_2763;
  assign _EVAL_4144 = _EVAL_5813 & 32'h30;
  assign _EVAL_749 = _EVAL_4144 == 32'h30;
  assign _EVAL_4346 = _EVAL_1518 | _EVAL_749;
  assign _EVAL_1017 = _EVAL_5813 & 32'h90000010;
  assign _EVAL_5306 = _EVAL_1017 == 32'h80000010;
  assign _EVAL_4840 = _EVAL_4346 | _EVAL_5306;
  assign _EVAL_893 = _EVAL_1592 != 5'h0;
  assign _EVAL_5150 = _EVAL_4840 & _EVAL_893;
  assign _EVAL_3450 = _EVAL_2766 | _EVAL_5882;
  assign _EVAL_194 = _EVAL_1947 & 32'h90000010;
  assign _EVAL_2220 = _EVAL_194 == 32'h80000010;
  assign _EVAL_5374 = _EVAL_3450 | _EVAL_2220;
  assign _EVAL_3155 = _EVAL_3215 != 5'h0;
  assign _EVAL_5022 = _EVAL_5374 & _EVAL_3155;
  assign _EVAL_1043 = _EVAL_1958 ? _EVAL_5150 : _EVAL_5022;
  assign _EVAL_4877 = _EVAL_4554 ? _EVAL_4254 : _EVAL_1043;
  assign _EVAL_174 = _EVAL_5133 & 32'h90000034;
  assign _EVAL_412 = _EVAL_174 == 32'h90000010;
  assign _EVAL_4766 = _EVAL_2404 | _EVAL_412;
  assign _EVAL_5032 = _EVAL_386 & 32'h2050;
  assign _EVAL_2591 = _EVAL_5032 == 32'h2000;
  assign _EVAL_441 = _EVAL_1242 & 32'h2024;
  assign _EVAL_4328 = _EVAL_1362 & 32'h28;
  assign _EVAL_2317 = _EVAL_4328 == 32'h28;
  assign _EVAL_4252 = _EVAL_1242 & 32'h18;
  assign _EVAL_3799 = _EVAL_4252 == 32'h0;
  assign _EVAL_196 = _EVAL_1242 & 32'h2010;
  assign _EVAL_2038 = _EVAL_196 == 32'h2000;
  assign _EVAL_3282 = _EVAL_3799 | _EVAL_2038;
  assign _EVAL_4365 = _EVAL_4585 == 32'h8000040;
  assign _EVAL_1691 = _EVAL_3282 | _EVAL_4365;
  assign _EVAL_384 = _EVAL_1074 ? _EVAL_1691 : _EVAL_2944;
  assign _EVAL_5678 = _EVAL_5311 & 32'h4003044;
  assign _EVAL_5230 = _EVAL_5678 == 32'h4000040;
  assign _EVAL_566 = _EVAL_3603 | _EVAL_5230;
  assign _EVAL_4623 = _EVAL_386 & 32'h44;
  assign _EVAL_4243 = _EVAL_4623 == 32'h0;
  assign _EVAL_4442 = _EVAL_386 & 32'h4024;
  assign _EVAL_6106 = _EVAL_4442 == 32'h20;
  assign _EVAL_204 = _EVAL_4243 | _EVAL_6106;
  assign _EVAL_5980 = _EVAL_204 | _EVAL_768;
  assign _EVAL_1658 = _EVAL_5813 & 32'h18;
  assign _EVAL_1923 = _EVAL_1658 == 32'h0;
  assign _EVAL_2488 = _EVAL_5813 & 32'h2010;
  assign _EVAL_281 = _EVAL_2488 == 32'h2000;
  assign _EVAL_2415 = _EVAL_1923 | _EVAL_281;
  assign _EVAL_3273 = _EVAL_2415 | _EVAL_2106;
  assign _EVAL_3244 = _EVAL_3271 & 32'h80000010;
  assign _EVAL_2620 = _EVAL_3244 == 32'h10;
  assign _EVAL_2815 = _EVAL_2620 | _EVAL_3764;
  assign _EVAL_3856 = _EVAL_3271 & 32'h40000040;
  assign _EVAL_1445 = _EVAL_3856 == 32'h40;
  assign _EVAL_5059 = _EVAL_2815 | _EVAL_1445;
  assign _EVAL_3865 = _EVAL_3271 & 32'h20000040;
  assign _EVAL_2803 = _EVAL_3865 == 32'h40;
  assign _EVAL_5968 = _EVAL_5059 | _EVAL_2803;
  assign _EVAL_5972 = _EVAL_4387 == 32'h40;
  assign _EVAL_521 = _EVAL_5968 | _EVAL_5972;
  assign _EVAL_1343 = _EVAL_4490 != 5'h0;
  assign _EVAL_4315 = _EVAL_864 & _EVAL_1343;
  assign _EVAL_3313 = _EVAL_1242 & 32'h64;
  assign _EVAL_5310 = _EVAL_3313 == 32'h0;
  assign _EVAL_6122 = _EVAL_5310 | _EVAL_5504;
  assign _EVAL_4032 = _EVAL_441 == 32'h24;
  assign _EVAL_4090 = _EVAL_6122 | _EVAL_4032;
  assign _EVAL_1901 = _EVAL_1242 & 32'h28;
  assign _EVAL_4035 = _EVAL_1901 == 32'h28;
  assign _EVAL_5871 = _EVAL_4090 | _EVAL_4035;
  assign _EVAL_5146 = _EVAL_1242 & 32'h30;
  assign _EVAL_737 = _EVAL_5146 == 32'h30;
  assign _EVAL_5235 = _EVAL_5871 | _EVAL_737;
  assign _EVAL_1625 = _EVAL_1242 & 32'h90000010;
  assign _EVAL_1714 = _EVAL_1625 == 32'h80000010;
  assign _EVAL_248 = _EVAL_5235 | _EVAL_1714;
  assign _EVAL_2366 = _EVAL_1621 != 5'h0;
  assign _EVAL_1548 = _EVAL_248 & _EVAL_2366;
  assign _EVAL_1966 = _EVAL_1074 ? _EVAL_1548 : _EVAL_3633;
  assign _EVAL_1401 = _EVAL_5926 ? _EVAL_4315 : _EVAL_1966;
  assign _EVAL_6024 = _EVAL_1947 & 32'hdfffffff;
  assign _EVAL_2450 = _EVAL_6024 == 32'h10500073;
  assign _EVAL_4498 = _EVAL_2123 | _EVAL_2450;
  assign _EVAL_5827 = _EVAL_3078 & 32'h306f;
  assign _EVAL_535 = _EVAL_5827 == 32'h1063;
  assign _EVAL_5805 = _EVAL_3581 | _EVAL_535;
  assign _EVAL_3092 = _EVAL_3078 & 32'h407f;
  assign _EVAL_1288 = _EVAL_3092 == 32'h4063;
  assign _EVAL_599 = _EVAL_5805 | _EVAL_1288;
  assign _EVAL_4298 = _EVAL_1023 == 32'h3;
  assign _EVAL_4158 = _EVAL_599 | _EVAL_4298;
  assign _EVAL_5447 = _EVAL_197 ? _EVAL_4968 : _EVAL_4536;
  assign _EVAL_5767 = _EVAL_5436 == 32'h40;
  assign _EVAL_2995 = _EVAL_1362 & 32'h64;
  assign _EVAL_573 = _EVAL_2995 == 32'h0;
  assign _EVAL_2650 = _EVAL_3813 == 32'h10;
  assign _EVAL_5726 = _EVAL_573 | _EVAL_2650;
  assign _EVAL_995 = _EVAL_1362 & 32'h2024;
  assign _EVAL_3511 = _EVAL_995 == 32'h24;
  assign _EVAL_1397 = _EVAL_5726 | _EVAL_3511;
  assign _EVAL_305 = _EVAL_1397 | _EVAL_2317;
  assign _EVAL_2331 = _EVAL_5072 == 32'h30;
  assign _EVAL_1999 = _EVAL_305 | _EVAL_2331;
  assign _EVAL_5803 = _EVAL_1362 & 32'h90000010;
  assign _EVAL_4900 = _EVAL_5803 == 32'h80000010;
  assign _EVAL_5742 = _EVAL_1999 | _EVAL_4900;
  assign _EVAL_190 = _EVAL_1362[11:7];
  assign _EVAL_266 = _EVAL_190 != 5'h0;
  assign _EVAL_4377 = _EVAL_5742 & _EVAL_266;
  assign _EVAL_4706 = _EVAL_2653 == 32'h0;
  assign _EVAL_3197 = _EVAL_4706 | _EVAL_2170;
  assign _EVAL_572 = _EVAL_3197 | _EVAL_5724;
  assign _EVAL_6114 = _EVAL_572 | _EVAL_5790;
  assign _EVAL_2402 = _EVAL_4702 & 32'h30;
  assign _EVAL_4307 = _EVAL_2402 == 32'h30;
  assign _EVAL_5873 = _EVAL_6114 | _EVAL_4307;
  assign _EVAL_2155 = _EVAL_4702 & 32'h90000010;
  assign _EVAL_5084 = _EVAL_2155 == 32'h80000010;
  assign _EVAL_5468 = _EVAL_5873 | _EVAL_5084;
  assign _EVAL_1237 = _EVAL_5468 & _EVAL_1360;
  assign _EVAL_4555 = _EVAL_197 ? _EVAL_4254 : _EVAL_4877;
  assign _EVAL_3205 = _EVAL_197 ? _EVAL_1237 : _EVAL_4555;
  assign _EVAL_5507 = _EVAL_4882 & 32'h8000040;
  assign _EVAL_4130 = _EVAL_5507 == 32'h8000040;
  assign _EVAL_2832 = _EVAL_4268 & 32'h28;
  assign _EVAL_1786 = _EVAL_2832 == 32'h28;
  assign _EVAL_4195 = _EVAL_968 | _EVAL_1786;
  assign _EVAL_5035 = _EVAL_4268 & 32'h30;
  assign _EVAL_4616 = _EVAL_5035 == 32'h30;
  assign _EVAL_3427 = _EVAL_4195 | _EVAL_4616;
  assign _EVAL_3688 = _EVAL_4268 & 32'h90000010;
  assign _EVAL_5910 = _EVAL_3688 == 32'h80000010;
  assign _EVAL_1584 = _EVAL_3427 | _EVAL_5910;
  assign _EVAL_216 = _EVAL_1584 & _EVAL_3685;
  assign _EVAL_1055 = _EVAL_3259 != 5'h0;
  assign _EVAL_2716 = _EVAL_3537 & _EVAL_1055;
  assign _EVAL_4205 = _EVAL_4882 & 32'h2024;
  assign _EVAL_3442 = _EVAL_4205 == 32'h24;
  assign _EVAL_428 = _EVAL_2867 | _EVAL_3442;
  assign _EVAL_4005 = _EVAL_4882 & 32'h28;
  assign _EVAL_5545 = _EVAL_4005 == 32'h28;
  assign _EVAL_3171 = _EVAL_428 | _EVAL_5545;
  assign _EVAL_5950 = _EVAL_4882 & 32'h30;
  assign _EVAL_1480 = _EVAL_5950 == 32'h30;
  assign _EVAL_2978 = _EVAL_3171 | _EVAL_1480;
  assign _EVAL_3652 = _EVAL_4882 & 32'h90000010;
  assign _EVAL_3565 = _EVAL_3652 == 32'h80000010;
  assign _EVAL_784 = _EVAL_2978 | _EVAL_3565;
  assign _EVAL_589 = _EVAL_2496 != 5'h0;
  assign _EVAL_1308 = _EVAL_784 & _EVAL_589;
  assign _EVAL_625 = _EVAL_5133 & 32'h28;
  assign _EVAL_4721 = _EVAL_625 == 32'h28;
  assign _EVAL_4010 = _EVAL_909 | _EVAL_4721;
  assign _EVAL_3252 = _EVAL_5133 & 32'h30;
  assign _EVAL_819 = _EVAL_3252 == 32'h30;
  assign _EVAL_4851 = _EVAL_4010 | _EVAL_819;
  assign _EVAL_4007 = _EVAL_4851 | _EVAL_5229;
  assign _EVAL_3159 = _EVAL_2839 != 5'h0;
  assign _EVAL_3858 = _EVAL_4007 & _EVAL_3159;
  assign _EVAL_1517 = _EVAL_2901 ? _EVAL_1308 : _EVAL_3858;
  assign _EVAL_3568 = _EVAL_2378 ? _EVAL_2716 : _EVAL_1517;
  assign _EVAL_485 = _EVAL_5690 ? _EVAL_2716 : _EVAL_3568;
  assign _EVAL_5180 = _EVAL_5690 ? _EVAL_216 : _EVAL_485;
  assign _EVAL_4150 = _EVAL_1978[11:7];
  assign _EVAL_844 = _EVAL_4150 != 5'h0;
  assign _EVAL_862 = _EVAL_302 & _EVAL_844;
  assign _EVAL_488 = _EVAL_3271[11:7];
  assign _EVAL_3791 = _EVAL_488 != 5'h0;
  assign _EVAL_4611 = _EVAL_4906 & _EVAL_3791;
  assign _EVAL_5103 = _EVAL_668 ? _EVAL_4377 : _EVAL_4611;
  assign _EVAL_4424 = _EVAL_3050 ? _EVAL_862 : _EVAL_5103;
  assign _EVAL_4015 = _EVAL_1069 ? _EVAL_862 : _EVAL_4424;
  assign _EVAL_4259 = _EVAL_2142 ? _EVAL_5180 : _EVAL_4015;
  assign _EVAL_958 = _EVAL_2164 & 32'h38;
  assign _EVAL_5370 = _EVAL_3078 & 32'h80000010;
  assign _EVAL_2446 = _EVAL_5370 == 32'h10;
  assign _EVAL_5279 = _EVAL_2446 | _EVAL_910;
  assign _EVAL_4599 = _EVAL_3078 & 32'h40000040;
  assign _EVAL_5085 = _EVAL_4599 == 32'h40;
  assign _EVAL_1913 = _EVAL_5279 | _EVAL_5085;
  assign _EVAL_5747 = _EVAL_3078 & 32'h20000040;
  assign _EVAL_189 = _EVAL_5747 == 32'h40;
  assign _EVAL_523 = _EVAL_1913 | _EVAL_189;
  assign _EVAL_2695 = _EVAL_523 | _EVAL_2747;
  assign _EVAL_5241 = _EVAL_3078 & 32'h1040;
  assign _EVAL_931 = _EVAL_5241 == 32'h1040;
  assign _EVAL_4943 = _EVAL_2695 | _EVAL_931;
  assign _EVAL_2700 = _EVAL_1395 == 32'h10000040;
  assign _EVAL_3304 = _EVAL_4836 | _EVAL_2700;
  assign _EVAL_319 = _EVAL_1947 & 32'h3c;
  assign _EVAL_1298 = _EVAL_319 == 32'h4;
  assign _EVAL_4423 = _EVAL_1947 & 32'h80000060;
  assign _EVAL_1946 = _EVAL_4423 == 32'h40;
  assign _EVAL_419 = _EVAL_1298 | _EVAL_1946;
  assign _EVAL_4516 = _EVAL_419 | _EVAL_160;
  assign _EVAL_4899 = _EVAL_1947 & 32'h10000060;
  assign _EVAL_840 = _EVAL_4899 == 32'h10000040;
  assign _EVAL_3122 = _EVAL_4516 | _EVAL_840;
  assign _EVAL_3422 = _EVAL_1958 ? _EVAL_3304 : _EVAL_3122;
  assign _EVAL_5626 = _EVAL_1362 & 32'h4024;
  assign _EVAL_3230 = _EVAL_5626 == 32'h20;
  assign _EVAL_3375 = _EVAL_1451 & _EVAL_3373;
  assign _EVAL_3981 = _EVAL_4291 ? _EVAL_3623 : _EVAL_3375;
  assign _EVAL_3044 = _EVAL_5525 & _EVAL_3981;
  assign _EVAL_221 = _EVAL_574 & _EVAL_3044;
  assign _EVAL_1615 = _EVAL_2110 | _EVAL_5885;
  assign _EVAL_314 = _EVAL_221 & _EVAL_1615;
  assign _EVAL_2760 = _EVAL_1986 & _EVAL_3981;
  assign _EVAL_475 = _EVAL_574 & _EVAL_2760;
  assign _EVAL_2593 = _EVAL_2110 | _EVAL_2569;
  assign _EVAL_5852 = _EVAL_475 & _EVAL_2593;
  assign _EVAL_4240 = _EVAL_314 ? 1'h1 : _EVAL_5852;
  assign _EVAL_5450 = _EVAL_1947 & 32'h80000010;
  assign _EVAL_4844 = _EVAL_5450 == 32'h10;
  assign _EVAL_3697 = _EVAL_4844 | _EVAL_4779;
  assign _EVAL_4414 = _EVAL_1947 & 32'h40000040;
  assign _EVAL_4569 = _EVAL_4414 == 32'h40;
  assign _EVAL_6036 = _EVAL_3697 | _EVAL_4569;
  assign _EVAL_786 = _EVAL_1947 & 32'h20000040;
  assign _EVAL_2793 = _EVAL_786 == 32'h40;
  assign _EVAL_1632 = _EVAL_6036 | _EVAL_2793;
  assign _EVAL_899 = _EVAL_3006 & 32'h2040;
  assign _EVAL_686 = _EVAL_899 == 32'h2040;
  assign _EVAL_5218 = _EVAL_4256 | _EVAL_686;
  assign _EVAL_1522 = _EVAL_967 == 32'h2040;
  assign _EVAL_5353 = _EVAL_3137 | _EVAL_1522;
  assign _EVAL_4983 = _EVAL_2901 ? _EVAL_5353 : _EVAL_1652;
  assign _EVAL_743 = _EVAL_2378 ? _EVAL_5218 : _EVAL_4983;
  assign _EVAL_2824 = _EVAL_1365 ? 1'h1 : _EVAL_4240;
  assign _EVAL_2927 = _EVAL_1451 & _EVAL_1555;
  assign _EVAL_4837 = _EVAL_5062 | _EVAL_2927;
  assign _EVAL_4323 = _EVAL_4837 == _EVAL_1969;
  assign _EVAL_4300 = _EVAL_1451 & _EVAL_660;
  assign _EVAL_2730 = _EVAL_4291 ? _EVAL_4323 : _EVAL_4300;
  assign _EVAL_3668 = _EVAL_5525 & _EVAL_2730;
  assign _EVAL_2495 = _EVAL_574 & _EVAL_3668;
  assign _EVAL_5257 = _EVAL_2495 & _EVAL_5667;
  assign _EVAL_6025 = _EVAL_1986 & _EVAL_2730;
  assign _EVAL_2162 = _EVAL_574 & _EVAL_6025;
  assign _EVAL_5996 = _EVAL_2110 | _EVAL_209;
  assign _EVAL_2637 = _EVAL_2162 & _EVAL_5996;
  assign _EVAL_3151 = _EVAL_5257 ? 1'h1 : _EVAL_2637;
  assign _EVAL_663 = _EVAL_409 ? 1'h1 : _EVAL_3151;
  assign _EVAL_186 = _EVAL_574 & _EVAL_3787;
  assign _EVAL_3742 = _EVAL_2110 | _EVAL_935;
  assign _EVAL_2160 = _EVAL_186 & _EVAL_3742;
  assign _EVAL_1094 = _EVAL_1986 & _EVAL_351;
  assign _EVAL_1619 = _EVAL_574 & _EVAL_1094;
  assign _EVAL_5824 = _EVAL_2110 | _EVAL_1434;
  assign _EVAL_4676 = _EVAL_1619 & _EVAL_5824;
  assign _EVAL_1038 = _EVAL_2160 ? 1'h1 : _EVAL_4676;
  assign _EVAL_4068 = _EVAL_3870 ? 1'h1 : _EVAL_1038;
  assign _EVAL_399 = _EVAL_574 & _EVAL_3173;
  assign _EVAL_4472 = _EVAL_2110 | _EVAL_984;
  assign _EVAL_2728 = _EVAL_399 & _EVAL_4472;
  assign _EVAL_2966 = _EVAL_574 & _EVAL_254;
  assign _EVAL_716 = _EVAL_2110 | _EVAL_3402;
  assign _EVAL_2169 = _EVAL_2966 & _EVAL_716;
  assign _EVAL_2413 = _EVAL_2728 ? 1'h1 : _EVAL_2169;
  assign _EVAL_2925 = _EVAL_3070 ? 1'h1 : _EVAL_2413;
  assign _EVAL_1889 = {_EVAL_2824,_EVAL_663,_EVAL_4068,_EVAL_2925};
  assign _EVAL_4595 = _EVAL_1889 & _EVAL_4984;
  assign _EVAL_4006 = _EVAL_4595 != 4'h0;
  assign _EVAL_2447 = _EVAL_1171 ? 1'h1 : _EVAL_4006;
  assign _EVAL_2218 = _EVAL_4702 & 32'h4003044;
  assign _EVAL_2942 = _EVAL_2218 == 32'h4000040;
  assign _EVAL_2990 = _EVAL_3583 | _EVAL_2942;
  assign _EVAL_692 = _EVAL_4554 ? _EVAL_3459 : _EVAL_2812;
  assign _EVAL_816 = _EVAL_197 ? _EVAL_3459 : _EVAL_692;
  assign _EVAL_4849 = _EVAL_197 ? _EVAL_2990 : _EVAL_816;
  assign _EVAL_1178 = _EVAL_3313 == 32'h20;
  assign _EVAL_1240 = _EVAL_1242 & 32'h34;
  assign _EVAL_2095 = _EVAL_1240 == 32'h20;
  assign _EVAL_5536 = _EVAL_1178 | _EVAL_2095;
  assign _EVAL_5358 = _EVAL_1242 & 32'h2048;
  assign _EVAL_4169 = _EVAL_5358 == 32'h2008;
  assign _EVAL_1818 = _EVAL_5536 | _EVAL_4169;
  assign _EVAL_5730 = _EVAL_1242 & 32'h4003044;
  assign _EVAL_866 = _EVAL_5730 == 32'h4000040;
  assign _EVAL_4162 = _EVAL_1818 | _EVAL_866;
  assign _EVAL_349 = _EVAL_5090 == 32'h20;
  assign _EVAL_2254 = _EVAL_2164 & 32'h34;
  assign _EVAL_1683 = _EVAL_2254 == 32'h20;
  assign _EVAL_3464 = _EVAL_349 | _EVAL_1683;
  assign _EVAL_1046 = _EVAL_2164 & 32'h2048;
  assign _EVAL_3226 = _EVAL_1046 == 32'h2008;
  assign _EVAL_4464 = _EVAL_3464 | _EVAL_3226;
  assign _EVAL_5485 = _EVAL_2164 & 32'h4003044;
  assign _EVAL_2688 = _EVAL_5485 == 32'h4000040;
  assign _EVAL_2893 = _EVAL_4464 | _EVAL_2688;
  assign _EVAL_5412 = _EVAL_1074 ? _EVAL_4162 : _EVAL_2893;
  assign _EVAL_5647 = _EVAL_5926 ? _EVAL_3890 : _EVAL_5412;
  assign _EVAL_4279 = _EVAL_2970 ? _EVAL_3890 : _EVAL_5647;
  assign _EVAL_5554 = _EVAL_2970 ? _EVAL_566 : _EVAL_4279;
  assign _EVAL_5917 = _EVAL_3006 & 32'h2048;
  assign _EVAL_2356 = _EVAL_5917 == 32'h2008;
  assign _EVAL_4523 = _EVAL_325 | _EVAL_2356;
  assign _EVAL_3556 = _EVAL_3006 & 32'h4003044;
  assign _EVAL_5936 = _EVAL_3556 == 32'h4000040;
  assign _EVAL_3127 = _EVAL_4523 | _EVAL_5936;
  assign _EVAL_2536 = _EVAL_365 == 32'h2008;
  assign _EVAL_1252 = _EVAL_5307 | _EVAL_2536;
  assign _EVAL_5592 = _EVAL_1252 | _EVAL_715;
  assign _EVAL_176 = _EVAL_1731 == 32'h20;
  assign _EVAL_2601 = _EVAL_176 | _EVAL_1524;
  assign _EVAL_4312 = _EVAL_5133 & 32'h2048;
  assign _EVAL_1533 = _EVAL_4312 == 32'h2008;
  assign _EVAL_869 = _EVAL_2601 | _EVAL_1533;
  assign _EVAL_5467 = _EVAL_5133 & 32'h4003044;
  assign _EVAL_5922 = _EVAL_5467 == 32'h4000040;
  assign _EVAL_1229 = _EVAL_869 | _EVAL_5922;
  assign _EVAL_2518 = _EVAL_2901 ? _EVAL_5592 : _EVAL_1229;
  assign _EVAL_6142 = _EVAL_2378 ? _EVAL_3127 : _EVAL_2518;
  assign _EVAL_5266 = _EVAL_5690 ? _EVAL_3127 : _EVAL_6142;
  assign _EVAL_3132 = _EVAL_5690 ? _EVAL_3666 : _EVAL_5266;
  assign _EVAL_5763 = _EVAL_2995 == 32'h20;
  assign _EVAL_5040 = _EVAL_3163 == 32'h20;
  assign _EVAL_5395 = _EVAL_5763 | _EVAL_5040;
  assign _EVAL_529 = _EVAL_1362 & 32'h2048;
  assign _EVAL_5106 = _EVAL_529 == 32'h2008;
  assign _EVAL_2686 = _EVAL_5395 | _EVAL_5106;
  assign _EVAL_5627 = _EVAL_1362 & 32'h4003044;
  assign _EVAL_3429 = _EVAL_5627 == 32'h4000040;
  assign _EVAL_4761 = _EVAL_2686 | _EVAL_3429;
  assign _EVAL_1767 = _EVAL_188 == 32'h20;
  assign _EVAL_5457 = _EVAL_1767 | _EVAL_1955;
  assign _EVAL_3095 = _EVAL_3271 & 32'h2048;
  assign _EVAL_5184 = _EVAL_3095 == 32'h2008;
  assign _EVAL_873 = _EVAL_5457 | _EVAL_5184;
  assign _EVAL_5349 = _EVAL_873 | _EVAL_1655;
  assign _EVAL_3237 = _EVAL_668 ? _EVAL_4761 : _EVAL_5349;
  assign _EVAL_1147 = _EVAL_3050 ? _EVAL_375 : _EVAL_3237;
  assign _EVAL_3569 = _EVAL_1069 ? _EVAL_375 : _EVAL_1147;
  assign _EVAL_4600 = _EVAL_2142 ? _EVAL_3132 : _EVAL_3569;
  assign _EVAL_2634 = _EVAL_3052 ? _EVAL_5554 : _EVAL_4600;
  assign _EVAL_2630 = _EVAL_1550 == 32'h40;
  assign _EVAL_5984 = _EVAL_1632 | _EVAL_2630;
  assign _EVAL_5706 = _EVAL_3078 & 32'h3c;
  assign _EVAL_3743 = _EVAL_5706 == 32'h4;
  assign _EVAL_5681 = _EVAL_3078 & 32'h80000060;
  assign _EVAL_199 = _EVAL_5681 == 32'h40;
  assign _EVAL_2852 = _EVAL_3743 | _EVAL_199;
  assign _EVAL_2764 = _EVAL_2852 | _EVAL_2310;
  assign _EVAL_4053 = _EVAL_2764 | _EVAL_827;
  assign _EVAL_5684 = _EVAL_4554 ? _EVAL_4053 : _EVAL_3422;
  assign _EVAL_1497 = _EVAL_197 ? _EVAL_4053 : _EVAL_5684;
  assign _EVAL_1012 = _EVAL_3078 & 32'h8000040;
  assign _EVAL_711 = _EVAL_1012 == 32'h8000040;
  assign _EVAL_990 = _EVAL_4978 & _EVAL_2223;
  assign _EVAL_1011 = _EVAL_5399 | _EVAL_990;
  assign _EVAL_170 = _EVAL_1011 == _EVAL_383;
  assign _EVAL_3019 = _EVAL_1718 == 32'h0;
  assign _EVAL_2286 = _EVAL_4268 & 32'h4024;
  assign _EVAL_5031 = _EVAL_2286 == 32'h20;
  assign _EVAL_933 = _EVAL_3019 | _EVAL_5031;
  assign _EVAL_765 = _EVAL_4268 & 32'h38;
  assign _EVAL_713 = _EVAL_765 == 32'h20;
  assign _EVAL_4650 = _EVAL_933 | _EVAL_713;
  assign _EVAL_1301 = _EVAL_4268 & 32'h2050;
  assign _EVAL_4459 = _EVAL_1301 == 32'h2000;
  assign _EVAL_5998 = _EVAL_4650 | _EVAL_4459;
  assign _EVAL_4380 = _EVAL_591 == 32'h24;
  assign _EVAL_3505 = _EVAL_4702 & 32'h40000060;
  assign _EVAL_3195 = _EVAL_3505 == 32'h40;
  assign _EVAL_3547 = _EVAL_4380 | _EVAL_3195;
  assign _EVAL_622 = _EVAL_3547 | _EVAL_4636;
  assign _EVAL_2553 = _EVAL_197 ? _EVAL_622 : _EVAL_4258;
  assign _EVAL_2974 = _EVAL_5337 ? _EVAL_1561 : _EVAL_2395;
  assign _EVAL_5710 = _EVAL_3271 & 32'h90000034;
  assign _EVAL_912 = _EVAL_5710 == 32'h90000010;
  assign _EVAL_4958 = _EVAL_4974 | _EVAL_912;
  assign _EVAL_3771 = _EVAL_1330 & _EVAL_4445;
  assign _EVAL_4675 = _EVAL_5994 | _EVAL_4192;
  assign _EVAL_4411 = _EVAL_4702 & 32'h207f;
  assign _EVAL_5111 = _EVAL_4411 == 32'h3;
  assign _EVAL_1637 = _EVAL_3022 == 32'hf;
  assign _EVAL_5030 = _EVAL_5111 | _EVAL_1637;
  assign _EVAL_1841 = _EVAL_5030 | _EVAL_3656;
  assign _EVAL_2298 = _EVAL_4702 & 32'hfc00007f;
  assign _EVAL_723 = _EVAL_2298 == 32'h33;
  assign _EVAL_4093 = _EVAL_1841 | _EVAL_723;
  assign _EVAL_2922 = _EVAL_4702 & 32'hbe00707f;
  assign _EVAL_1024 = _EVAL_2922 == 32'h33;
  assign _EVAL_208 = _EVAL_4093 | _EVAL_1024;
  assign _EVAL_3615 = _EVAL_4702 & 32'h6000073;
  assign _EVAL_4938 = _EVAL_3615 == 32'h43;
  assign _EVAL_3889 = _EVAL_208 | _EVAL_4938;
  assign _EVAL_3572 = _EVAL_2844 == 32'h53;
  assign _EVAL_2478 = _EVAL_3889 | _EVAL_3572;
  assign _EVAL_802 = _EVAL_4702 & 32'h707b;
  assign _EVAL_4046 = _EVAL_802 == 32'h63;
  assign _EVAL_5982 = _EVAL_2478 | _EVAL_4046;
  assign _EVAL_5639 = _EVAL_4702 & 32'h7f;
  assign _EVAL_2560 = _EVAL_5639 == 32'h6f;
  assign _EVAL_1838 = _EVAL_5982 | _EVAL_2560;
  assign _EVAL_5983 = _EVAL_4702 & 32'hffefffff;
  assign _EVAL_1503 = _EVAL_5983 == 32'h73;
  assign _EVAL_2369 = _EVAL_1838 | _EVAL_1503;
  assign _EVAL_3523 = _EVAL_4702 & 32'hfe00305f;
  assign _EVAL_2354 = _EVAL_3523 == 32'h1013;
  assign _EVAL_2810 = _EVAL_2369 | _EVAL_2354;
  assign _EVAL_508 = _EVAL_4702 & 32'h705b;
  assign _EVAL_1815 = _EVAL_508 == 32'h2003;
  assign _EVAL_1195 = _EVAL_2810 | _EVAL_1815;
  assign _EVAL_1347 = _EVAL_4411 == 32'h2013;
  assign _EVAL_1885 = _EVAL_1195 | _EVAL_1347;
  assign _EVAL_2775 = _EVAL_4702 & 32'h1800707f;
  assign _EVAL_949 = _EVAL_2775 == 32'h202f;
  assign _EVAL_482 = _EVAL_1885 | _EVAL_949;
  assign _EVAL_3539 = _EVAL_4411 == 32'h2073;
  assign _EVAL_1001 = _EVAL_482 | _EVAL_3539;
  assign _EVAL_2660 = _EVAL_4702 & 32'hbe00705f;
  assign _EVAL_6095 = _EVAL_2660 == 32'h5013;
  assign _EVAL_1664 = _EVAL_1001 | _EVAL_6095;
  assign _EVAL_4433 = _EVAL_4702 & 32'he800707f;
  assign _EVAL_4107 = _EVAL_4433 == 32'h800202f;
  assign _EVAL_3362 = _EVAL_1664 | _EVAL_4107;
  assign _EVAL_664 = _EVAL_4702 & 32'hf9f0707f;
  assign _EVAL_3124 = _EVAL_664 == 32'h1000202f;
  assign _EVAL_244 = _EVAL_3362 | _EVAL_3124;
  assign _EVAL_6060 = _EVAL_4702 & 32'hdfffffff;
  assign _EVAL_4215 = _EVAL_6060 == 32'h10500073;
  assign _EVAL_5152 = _EVAL_244 | _EVAL_4215;
  assign _EVAL_2361 = _EVAL_5152 | _EVAL_5290;
  assign _EVAL_2283 = _EVAL_4125 == 32'h20000053;
  assign _EVAL_5839 = _EVAL_2361 | _EVAL_2283;
  assign _EVAL_6058 = _EVAL_4702 & 32'h7e00507f;
  assign _EVAL_930 = _EVAL_6058 == 32'h20000053;
  assign _EVAL_5046 = _EVAL_5839 | _EVAL_930;
  assign _EVAL_313 = _EVAL_4702 == 32'h30200073;
  assign _EVAL_3158 = _EVAL_5046 | _EVAL_313;
  assign _EVAL_230 = _EVAL_3828 == 32'h58000053;
  assign _EVAL_442 = _EVAL_3158 | _EVAL_230;
  assign _EVAL_4310 = _EVAL_4702 == 32'h7b200073;
  assign _EVAL_2015 = _EVAL_442 | _EVAL_4310;
  assign _EVAL_387 = _EVAL_4702 & 32'hefe0007f;
  assign _EVAL_1049 = _EVAL_387 == 32'hc0000053;
  assign _EVAL_4357 = _EVAL_2015 | _EVAL_1049;
  assign _EVAL_1725 = _EVAL_4357 | _EVAL_1180;
  assign _EVAL_3592 = _EVAL_4702 & 32'heff0707f;
  assign _EVAL_2363 = _EVAL_3592 == 32'he0000053;
  assign _EVAL_1514 = _EVAL_1725 | _EVAL_2363;
  assign _EVAL_3357 = _EVAL_4702 & 32'hffd07fff;
  assign _EVAL_4299 = _EVAL_3357 == 32'hfc000073;
  assign _EVAL_925 = _EVAL_1514 | _EVAL_4299;
  assign _EVAL_1895 = _EVAL_520 == 32'h1063;
  assign _EVAL_1770 = _EVAL_925 | _EVAL_1895;
  assign _EVAL_4582 = _EVAL_4702 & 32'h407f;
  assign _EVAL_5205 = _EVAL_4582 == 32'h4063;
  assign _EVAL_1154 = _EVAL_1770 | _EVAL_5205;
  assign _EVAL_3342 = _EVAL_1947 & 32'h605f;
  assign _EVAL_2813 = _EVAL_3342 == 32'h3;
  assign _EVAL_4824 = _EVAL_1362[31:25];
  assign _EVAL_5192 = _EVAL_1978[6:2];
  assign _EVAL_4605 = _EVAL_1362[6:2];
  assign _EVAL_2873 = _EVAL_668 ? _EVAL_4605 : _EVAL_639;
  assign _EVAL_5849 = _EVAL_3050 ? _EVAL_5192 : _EVAL_2873;
  assign _EVAL_3754 = _EVAL_1069 ? _EVAL_5192 : _EVAL_5849;
  assign _EVAL_1188 = _EVAL_4978 & _EVAL_5541;
  assign _EVAL_791 = _EVAL_5311 & 32'h7c;
  assign _EVAL_5317 = _EVAL_791 == 32'h24;
  assign _EVAL_2864 = _EVAL_5311 & 32'h40000060;
  assign _EVAL_271 = _EVAL_2864 == 32'h40;
  assign _EVAL_6134 = _EVAL_5317 | _EVAL_271;
  assign _EVAL_1294 = _EVAL_3078[6:2];
  assign _EVAL_4624 = _EVAL_1183 & _EVAL_4984;
  assign _EVAL_586 = _EVAL_2385 & _EVAL_4445;
  assign _EVAL_5793 = _EVAL_5952 ? _EVAL_5878 : _EVAL_6087;
  assign _EVAL_3033 = _EVAL_3570 ? _EVAL_5057 : _EVAL_5793;
  assign _EVAL_3689 = _EVAL_5833 ? _EVAL_5057 : _EVAL_3033;
  assign _EVAL_3456 = _EVAL_5833 ? _EVAL_4374 : _EVAL_3689;
  assign _EVAL_2294 = _EVAL_5690 ? _EVAL_3259 : _EVAL_3059;
  assign _EVAL_1692 = _EVAL_5690 ? _EVAL_932 : _EVAL_2294;
  assign _EVAL_4612 = _EVAL_668 ? _EVAL_190 : _EVAL_488;
  assign _EVAL_1091 = _EVAL_3050 ? _EVAL_4150 : _EVAL_4612;
  assign _EVAL_390 = _EVAL_1069 ? _EVAL_4150 : _EVAL_1091;
  assign _EVAL_5248 = _EVAL_2142 ? _EVAL_1692 : _EVAL_390;
  assign _EVAL_5312 = _EVAL_3052 ? _EVAL_4076 : _EVAL_5248;
  assign _EVAL_2291 = _EVAL_5276 ? _EVAL_3456 : _EVAL_5312;
  assign _EVAL_2273 = _EVAL_5974 == 32'h0;
  assign _EVAL_1002 = _EVAL_2273 | _EVAL_6083;
  assign _EVAL_3389 = _EVAL_5311 & 32'h2024;
  assign _EVAL_191 = _EVAL_3389 == 32'h24;
  assign _EVAL_1438 = _EVAL_1002 | _EVAL_191;
  assign _EVAL_3335 = _EVAL_5311 & 32'h28;
  assign _EVAL_1345 = _EVAL_3335 == 32'h28;
  assign _EVAL_3388 = _EVAL_1438 | _EVAL_1345;
  assign _EVAL_5154 = _EVAL_5311 & 32'h30;
  assign _EVAL_1247 = _EVAL_5154 == 32'h30;
  assign _EVAL_2333 = _EVAL_3388 | _EVAL_1247;
  assign _EVAL_3093 = _EVAL_5311 & 32'h90000010;
  assign _EVAL_4564 = _EVAL_3093 == 32'h80000010;
  assign _EVAL_1902 = _EVAL_2333 | _EVAL_4564;
  assign _EVAL_4888 = _EVAL_1902 & _EVAL_863;
  assign _EVAL_3868 = _EVAL_2970 ? _EVAL_4315 : _EVAL_1401;
  assign _EVAL_5830 = _EVAL_2970 ? _EVAL_4888 : _EVAL_3868;
  assign _EVAL_1403 = _EVAL_5337 ? _EVAL_5180 : _EVAL_4015;
  assign _EVAL_3998 = _EVAL_1930 ? _EVAL_5830 : _EVAL_1403;
  assign _EVAL_3665 = _EVAL_386 & 32'h90000034;
  assign _EVAL_398 = _EVAL_3665 == 32'h90000010;
  assign _EVAL_487 = _EVAL_3160 == 32'hfc000073;
  assign _EVAL_4379 = _EVAL_2128 == 32'h0;
  assign _EVAL_1306 = _EVAL_2164 & 32'h4024;
  assign _EVAL_363 = _EVAL_1306 == 32'h20;
  assign _EVAL_3993 = _EVAL_4379 | _EVAL_363;
  assign _EVAL_1801 = _EVAL_958 == 32'h20;
  assign _EVAL_555 = _EVAL_3993 | _EVAL_1801;
  assign _EVAL_3156 = _EVAL_2164 & 32'h2050;
  assign _EVAL_941 = _EVAL_3156 == 32'h2000;
  assign _EVAL_3175 = _EVAL_555 | _EVAL_941;
  assign _EVAL_5055 = _EVAL_2164 & 32'h90000034;
  assign _EVAL_5366 = _EVAL_5055 == 32'h90000010;
  assign _EVAL_2768 = _EVAL_3175 | _EVAL_5366;
  assign _EVAL_2195 = _EVAL_1074 ? _EVAL_270 : _EVAL_2768;
  assign _EVAL_2985 = _EVAL_4268 & 32'h20000040;
  assign _EVAL_3552 = _EVAL_2985 == 32'h40;
  assign _EVAL_1512 = _EVAL_590 | _EVAL_3552;
  assign _EVAL_2448 = _EVAL_2696 == 32'h40;
  assign _EVAL_5092 = _EVAL_1512 | _EVAL_2448;
  assign _EVAL_3350 = _EVAL_4268 & 32'h1040;
  assign _EVAL_3919 = _EVAL_3350 == 32'h1040;
  assign _EVAL_443 = _EVAL_5092 | _EVAL_3919;
  assign _EVAL_1117 = _EVAL_443 | _EVAL_579;
  assign _EVAL_1521 = _EVAL_5690 ? _EVAL_5218 : _EVAL_743;
  assign _EVAL_459 = _EVAL_5690 ? _EVAL_1117 : _EVAL_1521;
  assign _EVAL_2946 = _EVAL_1822 | _EVAL_3447;
  assign _EVAL_5199 = _EVAL_1362 & 32'h80000010;
  assign _EVAL_3753 = _EVAL_5199 == 32'h10;
  assign _EVAL_4666 = _EVAL_3753 | _EVAL_2650;
  assign _EVAL_980 = _EVAL_4666 | _EVAL_2458;
  assign _EVAL_2726 = _EVAL_1850 == 32'h40;
  assign _EVAL_828 = _EVAL_980 | _EVAL_2726;
  assign _EVAL_472 = _EVAL_3813 == 32'h40;
  assign _EVAL_3894 = _EVAL_828 | _EVAL_472;
  assign _EVAL_3780 = _EVAL_1362 & 32'h1040;
  assign _EVAL_5068 = _EVAL_3780 == 32'h1040;
  assign _EVAL_5901 = _EVAL_3894 | _EVAL_5068;
  assign _EVAL_3174 = _EVAL_5901 | _EVAL_3384;
  assign _EVAL_4246 = _EVAL_3271 & 32'h1040;
  assign _EVAL_1963 = _EVAL_4246 == 32'h1040;
  assign _EVAL_4456 = _EVAL_521 | _EVAL_1963;
  assign _EVAL_2243 = _EVAL_3271 & 32'h2040;
  assign _EVAL_2424 = _EVAL_2243 == 32'h2040;
  assign _EVAL_4565 = _EVAL_4456 | _EVAL_2424;
  assign _EVAL_5861 = _EVAL_668 ? _EVAL_3174 : _EVAL_4565;
  assign _EVAL_342 = _EVAL_3050 ? _EVAL_2946 : _EVAL_5861;
  assign _EVAL_901 = _EVAL_1069 ? _EVAL_2946 : _EVAL_342;
  assign _EVAL_1861 = _EVAL_5337 ? _EVAL_459 : _EVAL_901;
  assign _EVAL_3188 = _EVAL_3659 ? _EVAL_1726 : _EVAL_73;
  assign _EVAL_681 = _EVAL_3078 & 32'h2010;
  assign _EVAL_833 = _EVAL_154;
  assign _EVAL_5121 = _EVAL_2801 & _EVAL_833;
  assign _EVAL_4619 = _EVAL_5399 | _EVAL_5247;
  assign _EVAL_3366 = _EVAL_4619 == _EVAL_383;
  assign _EVAL_3217 = _EVAL_519 ? _EVAL_3366 : _EVAL_1188;
  assign _EVAL_2988 = _EVAL_5121 & _EVAL_3217;
  assign _EVAL_3270 = _EVAL_574 | _EVAL_3044;
  assign _EVAL_661 = _EVAL_2988 & _EVAL_3270;
  assign _EVAL_233 = _EVAL_3289 & _EVAL_3217;
  assign _EVAL_2436 = _EVAL_574 | _EVAL_2760;
  assign _EVAL_4700 = _EVAL_233 & _EVAL_2436;
  assign _EVAL_1870 = _EVAL_661 ? 1'h1 : _EVAL_4700;
  assign _EVAL_5846 = _EVAL_3955 ? 1'h1 : _EVAL_1870;
  assign _EVAL_890 = _EVAL_5121 & _EVAL_2124;
  assign _EVAL_4889 = _EVAL_574 | _EVAL_3668;
  assign _EVAL_3367 = _EVAL_890 & _EVAL_4889;
  assign _EVAL_3604 = _EVAL_574 | _EVAL_6025;
  assign _EVAL_5221 = _EVAL_3283 & _EVAL_3604;
  assign _EVAL_3597 = _EVAL_3367 ? 1'h1 : _EVAL_5221;
  assign _EVAL_478 = _EVAL_2917 ? 1'h1 : _EVAL_3597;
  assign _EVAL_4723 = _EVAL_4978 & _EVAL_378;
  assign _EVAL_2168 = _EVAL_519 ? _EVAL_170 : _EVAL_4723;
  assign _EVAL_742 = _EVAL_5121 & _EVAL_2168;
  assign _EVAL_1886 = _EVAL_742 & _EVAL_6131;
  assign _EVAL_6069 = _EVAL_3289 & _EVAL_2168;
  assign _EVAL_5566 = _EVAL_574 | _EVAL_1094;
  assign _EVAL_2340 = _EVAL_6069 & _EVAL_5566;
  assign _EVAL_603 = _EVAL_1886 ? 1'h1 : _EVAL_2340;
  assign _EVAL_4241 = _EVAL_5373 ? 1'h1 : _EVAL_603;
  assign _EVAL_2918 = _EVAL_5121 & _EVAL_3047;
  assign _EVAL_1436 = _EVAL_2918 & _EVAL_4773;
  assign _EVAL_1087 = _EVAL_1436 ? 1'h1 : _EVAL_201;
  assign _EVAL_814 = _EVAL_4716 ? 1'h1 : _EVAL_1087;
  assign _EVAL_2089 = {_EVAL_5846,_EVAL_478,_EVAL_4241,_EVAL_814};
  assign _EVAL_1554 = _EVAL_1149 == 32'h4;
  assign _EVAL_1165 = _EVAL_1272 | _EVAL_1554;
  assign _EVAL_973 = _EVAL_5600 ? _EVAL_815 : _EVAL_29;
  assign _EVAL_525 = _EVAL_386 & 32'h7c;
  assign _EVAL_918 = _EVAL_525 == 32'h24;
  assign _EVAL_2652 = _EVAL_5337 ? _EVAL_1692 : _EVAL_390;
  assign _EVAL_5414 = _EVAL_46 & _EVAL_52;
  assign _EVAL_4615 = _EVAL_386 & 32'h3c;
  assign _EVAL_994 = _EVAL_4615 == 32'h4;
  assign _EVAL_4587 = _EVAL_994 | _EVAL_2158;
  assign _EVAL_883 = _EVAL_4587 | _EVAL_4271;
  assign _EVAL_3199 = _EVAL_1829 | _EVAL_656;
  assign _EVAL_3625 = _EVAL_5980 | _EVAL_2591;
  assign _EVAL_4710 = _EVAL_1458 == 32'h0;
  assign _EVAL_2381 = _EVAL_4624 != 4'h0;
  assign _EVAL_1145 = _EVAL_4466 == 32'h0;
  assign _EVAL_3153 = _EVAL_3078 & 32'h60;
  assign _EVAL_4105 = _EVAL_3153 == 32'h0;
  assign _EVAL_4679 = _EVAL_1145 | _EVAL_4105;
  assign _EVAL_2586 = _EVAL_1659 == 32'h0;
  assign _EVAL_5506 = _EVAL_4679 | _EVAL_2586;
  assign _EVAL_5655 = _EVAL_2626 == 32'h4;
  assign _EVAL_3525 = _EVAL_5506 | _EVAL_5655;
  assign _EVAL_1386 = _EVAL_3078 & 32'h62003010;
  assign _EVAL_1756 = _EVAL_1386 == 32'h60000010;
  assign _EVAL_4873 = _EVAL_3525 | _EVAL_1756;
  assign _EVAL_1468 = _EVAL_888 & 32'h2050;
  assign _EVAL_2998 = _EVAL_5125 != 4'h0;
  assign _EVAL_3144 = _EVAL_2241 ? 1'h1 : _EVAL_2998;
  assign _EVAL_1574 = _EVAL_5133 & 32'h8000040;
  assign _EVAL_2267 = _EVAL_2970 ? _EVAL_307 : _EVAL_4479;
  assign _EVAL_5237 = _EVAL_1930 ? _EVAL_4076 : _EVAL_2652;
  assign _EVAL_5250 = _EVAL_6093 == 32'h0;
  assign _EVAL_249 = _EVAL_3006 & 32'h4024;
  assign _EVAL_4621 = _EVAL_249 == 32'h20;
  assign _EVAL_336 = _EVAL_5250 | _EVAL_4621;
  assign _EVAL_619 = _EVAL_5657 == 32'h20;
  assign _EVAL_2619 = _EVAL_336 | _EVAL_619;
  assign _EVAL_2319 = _EVAL_3706 == 32'h2000;
  assign _EVAL_2677 = _EVAL_2619 | _EVAL_2319;
  assign _EVAL_4915 = _EVAL_5854 & 32'h18;
  assign _EVAL_517 = _EVAL_4915 == 32'h0;
  assign _EVAL_4597 = _EVAL_5854 & 32'h2010;
  assign _EVAL_4275 = _EVAL_4597 == 32'h2000;
  assign _EVAL_4000 = _EVAL_517 | _EVAL_4275;
  assign _EVAL_1794 = _EVAL_5854 & 32'h8000040;
  assign _EVAL_5120 = _EVAL_1794 == 32'h8000040;
  assign _EVAL_1865 = _EVAL_4000 | _EVAL_5120;
  assign _EVAL_2172 = _EVAL_5311 & 32'h38;
  assign _EVAL_2928 = _EVAL_2172 == 32'h20;
  assign _EVAL_4514 = _EVAL_4858 | _EVAL_2928;
  assign _EVAL_1159 = _EVAL_5311 & 32'h2050;
  assign _EVAL_4986 = _EVAL_1159 == 32'h2000;
  assign _EVAL_1883 = _EVAL_4514 | _EVAL_4986;
  assign _EVAL_2265 = _EVAL_5311 & 32'h90000034;
  assign _EVAL_2416 = _EVAL_2265 == 32'h90000010;
  assign _EVAL_2814 = _EVAL_1883 | _EVAL_2416;
  assign _EVAL_6141 = _EVAL_3956 == 32'h0;
  assign _EVAL_1303 = _EVAL_2039 & 32'h4024;
  assign _EVAL_649 = _EVAL_1303 == 32'h20;
  assign _EVAL_1599 = _EVAL_6141 | _EVAL_649;
  assign _EVAL_2969 = _EVAL_2039 & 32'h38;
  assign _EVAL_414 = _EVAL_2969 == 32'h20;
  assign _EVAL_3717 = _EVAL_1599 | _EVAL_414;
  assign _EVAL_3704 = _EVAL_2039 & 32'h2050;
  assign _EVAL_2983 = _EVAL_3704 == 32'h2000;
  assign _EVAL_1372 = _EVAL_3717 | _EVAL_2983;
  assign _EVAL_3038 = _EVAL_2039 & 32'h90000034;
  assign _EVAL_492 = _EVAL_3038 == 32'h90000010;
  assign _EVAL_2755 = _EVAL_1372 | _EVAL_492;
  assign _EVAL_3982 = _EVAL_5926 ? _EVAL_2755 : _EVAL_2195;
  assign _EVAL_4568 = _EVAL_2970 ? _EVAL_2755 : _EVAL_3982;
  assign _EVAL_5198 = _EVAL_2970 ? _EVAL_2814 : _EVAL_4568;
  assign _EVAL_207 = _EVAL_4702 & 32'h1040;
  assign _EVAL_1941 = _EVAL_207 == 32'h1040;
  assign _EVAL_4952 = _EVAL_5909 | _EVAL_1941;
  assign _EVAL_3303 = _EVAL_5421 | _EVAL_3230;
  assign _EVAL_790 = _EVAL_1362 & 32'h38;
  assign _EVAL_5550 = _EVAL_790 == 32'h20;
  assign _EVAL_4137 = _EVAL_3303 | _EVAL_5550;
  assign _EVAL_4789 = _EVAL_1362 & 32'h2050;
  assign _EVAL_5021 = _EVAL_4789 == 32'h2000;
  assign _EVAL_4805 = _EVAL_4137 | _EVAL_5021;
  assign _EVAL_2731 = _EVAL_1362 & 32'h90000034;
  assign _EVAL_5216 = _EVAL_2731 == 32'h90000010;
  assign _EVAL_886 = _EVAL_4805 | _EVAL_5216;
  assign _EVAL_5321 = _EVAL_668 ? _EVAL_886 : _EVAL_4958;
  assign _EVAL_3968 = _EVAL_888 & 32'h44;
  assign _EVAL_2159 = _EVAL_3968 == 32'h0;
  assign _EVAL_3114 = _EVAL_888 & 32'h4024;
  assign _EVAL_2954 = _EVAL_3114 == 32'h20;
  assign _EVAL_2573 = _EVAL_2159 | _EVAL_2954;
  assign _EVAL_3221 = _EVAL_888 & 32'h38;
  assign _EVAL_3530 = _EVAL_3221 == 32'h20;
  assign _EVAL_1508 = _EVAL_2573 | _EVAL_3530;
  assign _EVAL_5433 = _EVAL_1947 == 32'h7b200073;
  assign _EVAL_3276 = _EVAL_5827 == 32'h3;
  assign _EVAL_1274 = _EVAL_4158 | _EVAL_3276;
  assign _EVAL_1547 = _EVAL_4095 ? 1'h0 : _EVAL_1274;
  assign _EVAL_2081 = _EVAL_792 != 12'h0;
  assign _EVAL_5703 = _EVAL_761 ? _EVAL_2081 : 1'h1;
  assign _EVAL_3718 = _EVAL_4440 ? 1'h1 : _EVAL_5703;
  assign _EVAL_1898 = _EVAL_1378 ? 1'h1 : _EVAL_3718;
  assign _EVAL_636 = _EVAL_537 ? 1'h1 : _EVAL_1898;
  assign _EVAL_5987 = _EVAL_1088 ? 1'h1 : _EVAL_636;
  assign _EVAL_2605 = _EVAL_5987 == 1'h0;
  assign _EVAL_5118 = _EVAL_5813 & 32'hfff0607f;
  assign _EVAL_5673 = _EVAL_5118 == 32'he0000053;
  assign _EVAL_3510 = _EVAL_1239 | _EVAL_5673;
  assign _EVAL_1231 = _EVAL_5813 & 32'heff0707f;
  assign _EVAL_2556 = _EVAL_1231 == 32'he0000053;
  assign _EVAL_2275 = _EVAL_3510 | _EVAL_2556;
  assign _EVAL_5939 = _EVAL_5813 & 32'hffd07fff;
  assign _EVAL_1580 = _EVAL_5939 == 32'hfc000073;
  assign _EVAL_491 = _EVAL_2275 | _EVAL_1580;
  assign _EVAL_1309 = _EVAL_5813 & 32'h306f;
  assign _EVAL_4768 = _EVAL_1309 == 32'h1063;
  assign _EVAL_5576 = _EVAL_491 | _EVAL_4768;
  assign _EVAL_5973 = _EVAL_1198 == 32'h4063;
  assign _EVAL_4556 = _EVAL_5576 | _EVAL_5973;
  assign _EVAL_2121 = _EVAL_5813 & 32'h605f;
  assign _EVAL_423 = _EVAL_2121 == 32'h3;
  assign _EVAL_5345 = _EVAL_4556 | _EVAL_423;
  assign _EVAL_237 = _EVAL_1309 == 32'h3;
  assign _EVAL_3479 = _EVAL_5345 | _EVAL_237;
  assign _EVAL_5557 = _EVAL_2605 ? 1'h0 : _EVAL_3479;
  assign _EVAL_3066 = _EVAL_537 ? 1'h1 : _EVAL_2770;
  assign _EVAL_3989 = _EVAL_1088 ? 1'h1 : _EVAL_3066;
  assign _EVAL_6035 = _EVAL_3989 == 1'h0;
  assign _EVAL_5746 = _EVAL_4498 | _EVAL_2064;
  assign _EVAL_2059 = _EVAL_1947 & 32'h7e00607f;
  assign _EVAL_5614 = _EVAL_2059 == 32'h20000053;
  assign _EVAL_5645 = _EVAL_5746 | _EVAL_5614;
  assign _EVAL_5889 = _EVAL_2191 == 32'h20000053;
  assign _EVAL_1454 = _EVAL_5645 | _EVAL_5889;
  assign _EVAL_4452 = _EVAL_1947 == 32'h30200073;
  assign _EVAL_5840 = _EVAL_1454 | _EVAL_4452;
  assign _EVAL_3331 = _EVAL_1947 & 32'hfff0007f;
  assign _EVAL_6107 = _EVAL_3331 == 32'h58000053;
  assign _EVAL_6103 = _EVAL_5840 | _EVAL_6107;
  assign _EVAL_1760 = _EVAL_6103 | _EVAL_5433;
  assign _EVAL_2018 = _EVAL_1947 & 32'hefe0007f;
  assign _EVAL_1441 = _EVAL_2018 == 32'hc0000053;
  assign _EVAL_5424 = _EVAL_1760 | _EVAL_1441;
  assign _EVAL_2604 = _EVAL_1947 & 32'hfff0607f;
  assign _EVAL_751 = _EVAL_2604 == 32'he0000053;
  assign _EVAL_3485 = _EVAL_5424 | _EVAL_751;
  assign _EVAL_2184 = _EVAL_1947 & 32'heff0707f;
  assign _EVAL_5659 = _EVAL_2184 == 32'he0000053;
  assign _EVAL_2523 = _EVAL_3485 | _EVAL_5659;
  assign _EVAL_3723 = _EVAL_2523 | _EVAL_487;
  assign _EVAL_2278 = _EVAL_3723 | _EVAL_2475;
  assign _EVAL_4422 = _EVAL_1947 & 32'h407f;
  assign _EVAL_4143 = _EVAL_4422 == 32'h4063;
  assign _EVAL_2352 = _EVAL_2278 | _EVAL_4143;
  assign _EVAL_1482 = _EVAL_2352 | _EVAL_2813;
  assign _EVAL_5942 = _EVAL_206 == 32'h3;
  assign _EVAL_5737 = _EVAL_1482 | _EVAL_5942;
  assign _EVAL_684 = _EVAL_6035 ? 1'h0 : _EVAL_5737;
  assign _EVAL_452 = _EVAL_1958 ? _EVAL_5557 : _EVAL_684;
  assign _EVAL_4883 = _EVAL_4554 ? _EVAL_1547 : _EVAL_452;
  assign _EVAL_3433 = _EVAL_3659 ? _EVAL_718 : _EVAL_12;
  assign _EVAL_5916 = _EVAL_5133 & 32'h18;
  assign _EVAL_1589 = _EVAL_5916 == 32'h0;
  assign _EVAL_1623 = _EVAL_5133 & 32'h2010;
  assign _EVAL_496 = _EVAL_1623 == 32'h2000;
  assign _EVAL_2850 = _EVAL_1589 | _EVAL_496;
  assign _EVAL_2761 = _EVAL_386 & 32'h2048;
  assign _EVAL_5038 = _EVAL_386 & 32'h80000010;
  assign _EVAL_3782 = _EVAL_5038 == 32'h10;
  assign _EVAL_3974 = _EVAL_3782 | _EVAL_706;
  assign _EVAL_904 = _EVAL_386 & 32'h40000040;
  assign _EVAL_2670 = _EVAL_904 == 32'h40;
  assign _EVAL_3039 = _EVAL_3974 | _EVAL_2670;
  assign _EVAL_1624 = _EVAL_3039 | _EVAL_507;
  assign _EVAL_1737 = _EVAL_1473 == 32'h40;
  assign _EVAL_5475 = _EVAL_1624 | _EVAL_1737;
  assign _EVAL_1791 = _EVAL_3078 & 32'h18;
  assign _EVAL_4304 = _EVAL_888[6:2];
  assign _EVAL_3720 = _EVAL_4743[6:2];
  assign _EVAL_6138 = _EVAL_386[6:2];
  assign _EVAL_5843 = _EVAL_5952 ? _EVAL_3720 : _EVAL_6138;
  assign _EVAL_2561 = _EVAL_3570 ? _EVAL_4304 : _EVAL_5843;
  assign _EVAL_2313 = _EVAL_5854 & 32'h2050;
  assign _EVAL_4852 = _EVAL_2313 == 32'h2000;
  assign _EVAL_1489 = _EVAL_3006 & 32'h2010;
  assign _EVAL_2737 = _EVAL_1489 == 32'h2000;
  assign _EVAL_3735 = _EVAL_2672 | _EVAL_2737;
  assign _EVAL_1588 = _EVAL_3006 & 32'h8000040;
  assign _EVAL_324 = _EVAL_1588 == 32'h8000040;
  assign _EVAL_4435 = _EVAL_3735 | _EVAL_324;
  assign _EVAL_3481 = _EVAL_4882 & 32'h18;
  assign _EVAL_3535 = _EVAL_3481 == 32'h0;
  assign _EVAL_6049 = _EVAL_4882 & 32'h2010;
  assign _EVAL_3349 = _EVAL_6049 == 32'h2000;
  assign _EVAL_5019 = _EVAL_3535 | _EVAL_3349;
  assign _EVAL_5042 = _EVAL_5019 | _EVAL_4130;
  assign _EVAL_4976 = _EVAL_1574 == 32'h8000040;
  assign _EVAL_986 = _EVAL_2850 | _EVAL_4976;
  assign _EVAL_402 = _EVAL_2901 ? _EVAL_5042 : _EVAL_986;
  assign _EVAL_2683 = _EVAL_2378 ? _EVAL_4435 : _EVAL_402;
  assign _EVAL_4135 = _EVAL_5690 ? _EVAL_4435 : _EVAL_2683;
  assign _EVAL_5147 = _EVAL_2039 & 32'h7c;
  assign _EVAL_4198 = _EVAL_5147 == 32'h24;
  assign _EVAL_1594 = _EVAL_4825 == 32'h10000040;
  assign _EVAL_3178 = _EVAL_1978 & 32'h90000034;
  assign _EVAL_5081 = _EVAL_2311 == 32'h24;
  assign _EVAL_4557 = _EVAL_5081 | _EVAL_776;
  assign _EVAL_5888 = _EVAL_4557 | _EVAL_697;
  assign _EVAL_5652 = _EVAL_2811 == 32'h24;
  assign _EVAL_1208 = _EVAL_4743 & 32'h40000060;
  assign _EVAL_5768 = _EVAL_1208 == 32'h40;
  assign _EVAL_5975 = _EVAL_5652 | _EVAL_5768;
  assign _EVAL_4184 = _EVAL_5975 | _EVAL_1433;
  assign _EVAL_3420 = _EVAL_918 | _EVAL_5767;
  assign _EVAL_5394 = _EVAL_3420 | _EVAL_4271;
  assign _EVAL_3624 = _EVAL_5952 ? _EVAL_4184 : _EVAL_5394;
  assign _EVAL_4902 = _EVAL_3570 ? _EVAL_5888 : _EVAL_3624;
  assign _EVAL_3002 = _EVAL_4743 & 32'h2000040;
  assign _EVAL_5336 = _EVAL_1978 & 32'h2050;
  assign _EVAL_5497 = _EVAL_5813 & 32'h62003010;
  assign _EVAL_2916 = _EVAL_5497 == 32'h60000010;
  assign _EVAL_4970 = _EVAL_1165 | _EVAL_2916;
  assign _EVAL_1047 = _EVAL_1947 & 32'h62003010;
  assign _EVAL_4828 = _EVAL_1047 == 32'h60000010;
  assign _EVAL_1319 = _EVAL_1139 | _EVAL_4828;
  assign _EVAL_4485 = _EVAL_1958 ? _EVAL_4970 : _EVAL_1319;
  assign _EVAL_3079 = _EVAL_4554 ? _EVAL_4873 : _EVAL_4485;
  assign _EVAL_4667 = _EVAL_197 ? _EVAL_4873 : _EVAL_3079;
  assign _EVAL_721 = _EVAL_5311 & 32'h18;
  assign _EVAL_1762 = _EVAL_721 == 32'h0;
  assign _EVAL_4802 = _EVAL_5311 & 32'h2010;
  assign _EVAL_1513 = _EVAL_4802 == 32'h2000;
  assign _EVAL_5807 = _EVAL_1762 | _EVAL_1513;
  assign _EVAL_3694 = _EVAL_5311 & 32'h8000040;
  assign _EVAL_1490 = _EVAL_3694 == 32'h8000040;
  assign _EVAL_4173 = _EVAL_5807 | _EVAL_1490;
  assign _EVAL_1097 = _EVAL_2039 & 32'h2010;
  assign _EVAL_824 = _EVAL_1097 == 32'h2000;
  assign _EVAL_3495 = _EVAL_1107 | _EVAL_824;
  assign _EVAL_4691 = _EVAL_2039 & 32'h8000040;
  assign _EVAL_3751 = _EVAL_4691 == 32'h8000040;
  assign _EVAL_5413 = _EVAL_3495 | _EVAL_3751;
  assign _EVAL_277 = _EVAL_5926 ? _EVAL_5413 : _EVAL_384;
  assign _EVAL_2722 = _EVAL_2970 ? _EVAL_5413 : _EVAL_277;
  assign _EVAL_4145 = _EVAL_2970 ? _EVAL_4173 : _EVAL_2722;
  assign _EVAL_860 = _EVAL_888 & 32'h18;
  assign _EVAL_4049 = _EVAL_860 == 32'h0;
  assign _EVAL_5884 = _EVAL_888 & 32'h2010;
  assign _EVAL_5239 = _EVAL_5884 == 32'h2000;
  assign _EVAL_3917 = _EVAL_4049 | _EVAL_5239;
  assign _EVAL_2131 = _EVAL_3917 | _EVAL_444;
  assign _EVAL_289 = _EVAL_3659 == 1'h0;
  assign _EVAL_854 = _EVAL_5994 & _EVAL_289;
  assign _EVAL_5660 = _EVAL_4664 + 32'h2;
  assign _EVAL_659 = _EVAL_5660 != _EVAL_136;
  assign _EVAL_5957 = _EVAL_854 & _EVAL_659;
  assign _EVAL_5537 = _EVAL_1468 == 32'h2000;
  assign _EVAL_5605 = _EVAL_1508 | _EVAL_5537;
  assign _EVAL_2271 = _EVAL_888 & 32'h90000034;
  assign _EVAL_1991 = _EVAL_2271 == 32'h90000010;
  assign _EVAL_5162 = _EVAL_5605 | _EVAL_1991;
  assign _EVAL_4024 = _EVAL_3625 | _EVAL_398;
  assign _EVAL_2257 = _EVAL_5952 ? _EVAL_5688 : _EVAL_4024;
  assign _EVAL_3438 = _EVAL_3570 ? _EVAL_5162 : _EVAL_2257;
  assign _EVAL_4656 = _EVAL_3637 == 32'h0;
  assign _EVAL_2280 = _EVAL_386 & 32'h60;
  assign _EVAL_513 = _EVAL_2280 == 32'h0;
  assign _EVAL_5362 = _EVAL_4656 | _EVAL_513;
  assign _EVAL_1519 = _EVAL_1473 == 32'h0;
  assign _EVAL_2789 = _EVAL_5362 | _EVAL_1519;
  assign _EVAL_2042 = _EVAL_1013 | _EVAL_6082;
  assign _EVAL_2834 = _EVAL_3168 == 32'h4000040;
  assign _EVAL_5461 = _EVAL_2042 | _EVAL_2834;
  assign _EVAL_1527 = _EVAL_5813[31:25];
  assign _EVAL_2295 = _EVAL_2039[31:25];
  assign _EVAL_4576 = _EVAL_1242[31:25];
  assign _EVAL_1419 = _EVAL_1074 ? _EVAL_4576 : _EVAL_490;
  assign _EVAL_5848 = _EVAL_5926 ? _EVAL_2295 : _EVAL_1419;
  assign _EVAL_5915 = _EVAL_2970 ? _EVAL_2295 : _EVAL_5848;
  assign _EVAL_4759 = _EVAL_2970 ? _EVAL_5282 : _EVAL_5915;
  assign _EVAL_2967 = _EVAL_4268[31:25];
  assign _EVAL_594 = _EVAL_3006[31:25];
  assign _EVAL_4694 = _EVAL_4882[31:25];
  assign _EVAL_3762 = _EVAL_5133[31:25];
  assign _EVAL_1836 = _EVAL_2901 ? _EVAL_4694 : _EVAL_3762;
  assign _EVAL_5800 = _EVAL_2378 ? _EVAL_594 : _EVAL_1836;
  assign _EVAL_3430 = _EVAL_5690 ? _EVAL_594 : _EVAL_5800;
  assign _EVAL_2324 = _EVAL_5690 ? _EVAL_2967 : _EVAL_3430;
  assign _EVAL_1918 = _EVAL_1978[31:25];
  assign _EVAL_4009 = _EVAL_3271[31:25];
  assign _EVAL_4152 = _EVAL_668 ? _EVAL_4824 : _EVAL_4009;
  assign _EVAL_1552 = _EVAL_3050 ? _EVAL_1918 : _EVAL_4152;
  assign _EVAL_1066 = _EVAL_1069 ? _EVAL_1918 : _EVAL_1552;
  assign _EVAL_1353 = _EVAL_2142 ? _EVAL_2324 : _EVAL_1066;
  assign _EVAL_468 = _EVAL_3052 ? _EVAL_4759 : _EVAL_1353;
  assign _EVAL_797 = _EVAL_1958 ? _EVAL_3273 : _EVAL_6136;
  assign _EVAL_575 = _EVAL_3006 & 32'h90000034;
  assign _EVAL_4643 = _EVAL_575 == 32'h90000010;
  assign _EVAL_1753 = _EVAL_2677 | _EVAL_4643;
  assign _EVAL_2715 = _EVAL_2901 ? _EVAL_889 : _EVAL_4766;
  assign _EVAL_3812 = _EVAL_2378 ? _EVAL_1753 : _EVAL_2715;
  assign _EVAL_5941 = _EVAL_5690 ? _EVAL_1753 : _EVAL_3812;
  assign _EVAL_926 = _EVAL_3172 == 32'h10;
  assign _EVAL_6000 = _EVAL_926 | _EVAL_3248;
  assign _EVAL_3953 = _EVAL_5813 & 32'h40000040;
  assign _EVAL_461 = _EVAL_3953 == 32'h40;
  assign _EVAL_4855 = _EVAL_6000 | _EVAL_461;
  assign _EVAL_2818 = _EVAL_4855 | _EVAL_4787;
  assign _EVAL_3681 = _EVAL_3680 == 32'h40;
  assign _EVAL_4083 = _EVAL_2818 | _EVAL_3681;
  assign _EVAL_779 = _EVAL_5813 & 32'h1040;
  assign _EVAL_3746 = _EVAL_779 == 32'h1040;
  assign _EVAL_4885 = _EVAL_4083 | _EVAL_3746;
  assign _EVAL_3860 = _EVAL_5813 & 32'h2040;
  assign _EVAL_4540 = _EVAL_3860 == 32'h2040;
  assign _EVAL_3347 = _EVAL_4885 | _EVAL_4540;
  assign _EVAL_5547 = _EVAL_5847 == 32'h3;
  assign _EVAL_3814 = _EVAL_1154 | _EVAL_5547;
  assign _EVAL_5995 = _EVAL_3814 | _EVAL_1990;
  assign _EVAL_6007 = _EVAL_197 ? _EVAL_1547 : _EVAL_4883;
  assign _EVAL_2567 = _EVAL_197 ? _EVAL_5995 : _EVAL_6007;
  assign _EVAL_4182 = _EVAL_1074 ? _EVAL_677 : _EVAL_4890;
  assign _EVAL_316 = _EVAL_5926 ? _EVAL_3653 : _EVAL_4182;
  assign _EVAL_5122 = _EVAL_2970 ? _EVAL_3653 : _EVAL_316;
  assign _EVAL_5273 = _EVAL_3085 | _EVAL_2784;
  assign _EVAL_2035 = _EVAL_5273 | _EVAL_3390;
  assign _EVAL_5951 = _EVAL_5600 ? _EVAL_372 : _EVAL_143;
  assign _EVAL_1402 = _EVAL_5854 & 32'h62003010;
  assign _EVAL_2529 = _EVAL_1402 == 32'h60000010;
  assign _EVAL_5517 = _EVAL_5854 & 32'h38;
  assign _EVAL_5352 = _EVAL_2142 ? _EVAL_2570 : _EVAL_3754;
  assign _EVAL_2330 = _EVAL_3002 == 32'h0;
  assign _EVAL_1556 = _EVAL_4301 == 32'h2040;
  assign _EVAL_3990 = _EVAL_5337 ? _EVAL_2570 : _EVAL_3754;
  assign _EVAL_748 = _EVAL_1930 ? _EVAL_698 : _EVAL_3990;
  assign _EVAL_6017 = _EVAL_4471 == 32'h40;
  assign _EVAL_3352 = _EVAL_2538 | _EVAL_6017;
  assign _EVAL_2443 = _EVAL_888 & 32'h1040;
  assign _EVAL_2468 = _EVAL_2443 == 32'h1040;
  assign _EVAL_3491 = _EVAL_3352 | _EVAL_2468;
  assign _EVAL_855 = _EVAL_219 == 32'h2040;
  assign _EVAL_1326 = _EVAL_3491 | _EVAL_855;
  assign _EVAL_5711 = _EVAL_3769 == 32'h10;
  assign _EVAL_1268 = _EVAL_5711 | _EVAL_1250;
  assign _EVAL_2490 = _EVAL_4743 & 32'h40000040;
  assign _EVAL_3502 = _EVAL_2490 == 32'h40;
  assign _EVAL_1769 = _EVAL_1268 | _EVAL_3502;
  assign _EVAL_1586 = _EVAL_1769 | _EVAL_1891;
  assign _EVAL_3030 = _EVAL_4601 == 32'h40;
  assign _EVAL_3189 = _EVAL_1586 | _EVAL_3030;
  assign _EVAL_3855 = _EVAL_4743 & 32'h1040;
  assign _EVAL_5249 = _EVAL_3855 == 32'h1040;
  assign _EVAL_3670 = _EVAL_3189 | _EVAL_5249;
  assign _EVAL_2800 = _EVAL_1919 == 32'h2040;
  assign _EVAL_2060 = _EVAL_3670 | _EVAL_2800;
  assign _EVAL_3631 = _EVAL_386 & 32'h1040;
  assign _EVAL_5096 = _EVAL_3631 == 32'h1040;
  assign _EVAL_5640 = _EVAL_5475 | _EVAL_5096;
  assign _EVAL_2658 = _EVAL_386 & 32'h2040;
  assign _EVAL_2043 = _EVAL_2658 == 32'h2040;
  assign _EVAL_291 = _EVAL_5640 | _EVAL_2043;
  assign _EVAL_2318 = _EVAL_5952 ? _EVAL_2060 : _EVAL_291;
  assign _EVAL_3288 = _EVAL_3570 ? _EVAL_1326 : _EVAL_2318;
  assign _EVAL_4443 = _EVAL_4579 | _EVAL_164;
  assign _EVAL_6002 = _EVAL_5854 & 32'h2024;
  assign _EVAL_2177 = _EVAL_6002 == 32'h24;
  assign _EVAL_856 = _EVAL_4443 | _EVAL_2177;
  assign _EVAL_3265 = _EVAL_3570 ? _EVAL_2131 : _EVAL_6133;
  assign _EVAL_971 = _EVAL_5833 ? _EVAL_2131 : _EVAL_3265;
  assign _EVAL_2718 = _EVAL_5418 == 32'h4;
  assign _EVAL_5275 = _EVAL_2718 | _EVAL_3007;
  assign _EVAL_2621 = _EVAL_5275 | _EVAL_697;
  assign _EVAL_2358 = _EVAL_878 == 32'h10000040;
  assign _EVAL_6028 = _EVAL_2035 | _EVAL_2358;
  assign _EVAL_1377 = _EVAL_4882 & 32'h3c;
  assign _EVAL_3816 = _EVAL_1377 == 32'h4;
  assign _EVAL_1421 = _EVAL_3816 | _EVAL_5771;
  assign _EVAL_5179 = _EVAL_1421 | _EVAL_2101;
  assign _EVAL_265 = _EVAL_5179 | _EVAL_562;
  assign _EVAL_2140 = _EVAL_3986 == 32'h10000040;
  assign _EVAL_3872 = _EVAL_1078 | _EVAL_2140;
  assign _EVAL_3884 = _EVAL_2901 ? _EVAL_265 : _EVAL_3872;
  assign _EVAL_2886 = _EVAL_2378 ? _EVAL_6028 : _EVAL_3884;
  assign _EVAL_3619 = _EVAL_5690 ? _EVAL_6028 : _EVAL_2886;
  assign _EVAL_633 = _EVAL_5337 ? _EVAL_4846 : _EVAL_3548;
  assign _EVAL_5368 = _EVAL_1930 ? _EVAL_3104 : _EVAL_633;
  assign _EVAL_976 = _EVAL_4088 | _EVAL_2679;
  assign _EVAL_3503 = _EVAL_976 | _EVAL_5728;
  assign _EVAL_1062 = _EVAL_3503 | _EVAL_617;
  assign _EVAL_5434 = _EVAL_1716 | _EVAL_3476;
  assign _EVAL_5498 = _EVAL_5434 | _EVAL_3653;
  assign _EVAL_3819 = _EVAL_5526 == 32'h10000040;
  assign _EVAL_5594 = _EVAL_5498 | _EVAL_3819;
  assign _EVAL_2820 = _EVAL_5926 ? _EVAL_5594 : _EVAL_2274;
  assign _EVAL_5651 = _EVAL_2970 ? _EVAL_5594 : _EVAL_2820;
  assign _EVAL_2117 = _EVAL_2970 ? _EVAL_1062 : _EVAL_5651;
  assign _EVAL_1470 = _EVAL_4451 | _EVAL_4912;
  assign _EVAL_4635 = _EVAL_4757 == 32'h10000040;
  assign _EVAL_5047 = _EVAL_1470 | _EVAL_4635;
  assign _EVAL_672 = _EVAL_5690 ? _EVAL_5047 : _EVAL_3619;
  assign _EVAL_4997 = _EVAL_1069 ? _EVAL_3258 : _EVAL_2345;
  assign _EVAL_2203 = _EVAL_2142 ? _EVAL_672 : _EVAL_4997;
  assign _EVAL_4326 = _EVAL_3052 ? _EVAL_2117 : _EVAL_2203;
  assign _EVAL_5291 = _EVAL_3078[24:20];
  assign _EVAL_1054 = _EVAL_5813[24:20];
  assign _EVAL_4067 = _EVAL_1947[24:20];
  assign _EVAL_1852 = _EVAL_1958 ? _EVAL_1054 : _EVAL_4067;
  assign _EVAL_5484 = _EVAL_4554 ? _EVAL_5291 : _EVAL_1852;
  assign _EVAL_3945 = _EVAL_197 ? _EVAL_5291 : _EVAL_5484;
  assign _EVAL_3314 = _EVAL_3659 ? _EVAL_5225 : _EVAL_152;
  assign _EVAL_4116 = _EVAL_1978 & 32'h18;
  assign _EVAL_3294 = _EVAL_4116 == 32'h0;
  assign _EVAL_4896 = _EVAL_1978 & 32'h2010;
  assign _EVAL_4727 = _EVAL_4896 == 32'h2000;
  assign _EVAL_3672 = _EVAL_3294 | _EVAL_4727;
  assign _EVAL_1871 = _EVAL_225 == 32'h8000040;
  assign _EVAL_1957 = _EVAL_3672 | _EVAL_1871;
  assign _EVAL_1341 = _EVAL_3050 ? _EVAL_1957 : _EVAL_3611;
  assign _EVAL_2145 = _EVAL_668 ? _EVAL_4770 : _EVAL_1739;
  assign _EVAL_1085 = _EVAL_3050 ? _EVAL_4329 : _EVAL_2145;
  assign _EVAL_2186 = _EVAL_1069 ? _EVAL_4329 : _EVAL_1085;
  assign _EVAL_1033 = _EVAL_693 >= 4'h3;
  assign _EVAL_2531 = _EVAL_2485 | _EVAL_1033;
  assign _EVAL_3944 = _EVAL_3461 < 3'h4;
  assign _EVAL_3648 = _EVAL_3944 & _EVAL_3080;
  assign _EVAL_1959 = _EVAL_2531 | _EVAL_3648;
  assign _EVAL_1106 = _EVAL_2761 == 32'h2008;
  assign _EVAL_2799 = _EVAL_236 | _EVAL_1106;
  assign _EVAL_691 = _EVAL_4274 == 32'h10000040;
  assign _EVAL_6015 = _EVAL_883 | _EVAL_691;
  assign _EVAL_2205 = _EVAL_3968 == 32'h4;
  assign _EVAL_1080 = _EVAL_4921 | _EVAL_2205;
  assign _EVAL_1579 = _EVAL_888 & 32'h62003010;
  assign _EVAL_3585 = _EVAL_1579 == 32'h60000010;
  assign _EVAL_6018 = _EVAL_1080 | _EVAL_3585;
  assign _EVAL_3463 = _EVAL_4743 & 32'h60;
  assign _EVAL_1695 = _EVAL_3463 == 32'h0;
  assign _EVAL_5708 = _EVAL_2330 | _EVAL_1695;
  assign _EVAL_4992 = _EVAL_4601 == 32'h0;
  assign _EVAL_4652 = _EVAL_5708 | _EVAL_4992;
  assign _EVAL_5559 = _EVAL_1224 == 32'h4;
  assign _EVAL_1176 = _EVAL_4652 | _EVAL_5559;
  assign _EVAL_1150 = _EVAL_1176 | _EVAL_2133;
  assign _EVAL_4895 = _EVAL_4623 == 32'h4;
  assign _EVAL_5886 = _EVAL_2789 | _EVAL_4895;
  assign _EVAL_1488 = _EVAL_386 & 32'h62003010;
  assign _EVAL_1376 = _EVAL_1488 == 32'h60000010;
  assign _EVAL_187 = _EVAL_5886 | _EVAL_1376;
  assign _EVAL_5013 = _EVAL_5952 ? _EVAL_1150 : _EVAL_187;
  assign _EVAL_1044 = _EVAL_3570 ? _EVAL_6018 : _EVAL_5013;
  assign _EVAL_6048 = _EVAL_6079 == 32'h0;
  assign _EVAL_1539 = _EVAL_292 == 32'h28;
  assign _EVAL_2044 = _EVAL_654[14:12];
  assign _EVAL_3021 = _EVAL_3078[14:12];
  assign _EVAL_3546 = _EVAL_5813[14:12];
  assign _EVAL_4234 = _EVAL_1947[14:12];
  assign _EVAL_1266 = _EVAL_1958 ? _EVAL_3546 : _EVAL_4234;
  assign _EVAL_5656 = _EVAL_4554 ? _EVAL_3021 : _EVAL_1266;
  assign _EVAL_1391 = _EVAL_197 ? _EVAL_3021 : _EVAL_5656;
  assign _EVAL_3249 = _EVAL_197 ? _EVAL_2044 : _EVAL_1391;
  assign _EVAL_347 = _EVAL_4353 == 32'h0;
  assign _EVAL_2484 = _EVAL_5854 & 32'h4024;
  assign _EVAL_2207 = _EVAL_2484 == 32'h20;
  assign _EVAL_3411 = _EVAL_347 | _EVAL_2207;
  assign _EVAL_483 = _EVAL_5517 == 32'h20;
  assign _EVAL_4775 = _EVAL_3411 | _EVAL_483;
  assign _EVAL_5330 = _EVAL_4775 | _EVAL_4852;
  assign _EVAL_3901 = _EVAL_5854 & 32'h90000034;
  assign _EVAL_3116 = _EVAL_3901 == 32'h90000010;
  assign _EVAL_4146 = _EVAL_5330 | _EVAL_3116;
  assign _EVAL_1476 = _EVAL_5337 ? _EVAL_672 : _EVAL_4997;
  assign _EVAL_4283 = _EVAL_2970 ? 1'h0 : 1'h1;
  assign _EVAL_2617 = _EVAL_5690 ? 1'h0 : 1'h1;
  assign _EVAL_5553 = _EVAL_5337 ? _EVAL_2617 : 1'h1;
  assign _EVAL_2377 = _EVAL_1930 ? _EVAL_4283 : _EVAL_5553;
  assign _EVAL_168 = _EVAL_4743 & 32'h4003044;
  assign _EVAL_3475 = _EVAL_3052 ? _EVAL_5830 : _EVAL_4259;
  assign _EVAL_3852 = _EVAL_386[14:12];
  assign _EVAL_1983 = _EVAL_3052 ? _EVAL_698 : _EVAL_5352;
  assign _EVAL_551 = _EVAL_654[14];
  assign _EVAL_3646 = _EVAL_5905 | _EVAL_4912;
  assign _EVAL_2751 = _EVAL_5386[14:12];
  assign _EVAL_382 = _EVAL_888[14:12];
  assign _EVAL_3246 = _EVAL_4743[14:12];
  assign _EVAL_5960 = _EVAL_5952 ? _EVAL_3246 : _EVAL_3852;
  assign _EVAL_3064 = _EVAL_3570 ? _EVAL_382 : _EVAL_5960;
  assign _EVAL_538 = _EVAL_5833 ? _EVAL_382 : _EVAL_3064;
  assign _EVAL_4455 = _EVAL_5833 ? _EVAL_2751 : _EVAL_538;
  assign _EVAL_245 = _EVAL_5957 ? 1'h1 : _EVAL_95;
  assign _EVAL_908 = _EVAL_3012 != 4'h0;
  assign _EVAL_2896 = _EVAL_2142 ? _EVAL_2617 : 1'h1;
  assign _EVAL_4131 = _EVAL_3052 ? _EVAL_4283 : _EVAL_2896;
  assign _EVAL_4543 = _EVAL_1930 ? _EVAL_2117 : _EVAL_1476;
  assign _EVAL_301 = _EVAL_2816 | _EVAL_2953;
  assign _EVAL_3452 = _EVAL_5833 ? 1'h0 : 1'h1;
  assign _EVAL_3421 = _EVAL_5690 ? _EVAL_3390 : _EVAL_2851;
  assign _EVAL_3789 = _EVAL_5690 ? _EVAL_4912 : _EVAL_3421;
  assign _EVAL_3928 = _EVAL_2142 ? _EVAL_3789 : _EVAL_2186;
  assign _EVAL_5010 = _EVAL_5337 ? _EVAL_3108 : _EVAL_5619;
  assign _EVAL_5051 = _EVAL_1930 ? _EVAL_6030 : _EVAL_5010;
  assign _EVAL_3949 = _EVAL_4928 | _EVAL_2529;
  assign _EVAL_256 = _EVAL_5833 ? _EVAL_6018 : _EVAL_1044;
  assign _EVAL_1279 = _EVAL_5833 ? _EVAL_3949 : _EVAL_256;
  assign _EVAL_4820 = _EVAL_2142 ? _EVAL_953 : _EVAL_5129;
  assign _EVAL_2399 = _EVAL_3052 ? _EVAL_4448 : _EVAL_4820;
  assign _EVAL_5642 = _EVAL_5276 ? _EVAL_1279 : _EVAL_2399;
  assign _EVAL_4972 = _EVAL_2039 & 32'h40000060;
  assign _EVAL_3190 = _EVAL_4972 == 32'h40;
  assign _EVAL_405 = _EVAL_4198 | _EVAL_3190;
  assign _EVAL_1307 = _EVAL_405 | _EVAL_3653;
  assign _EVAL_674 = _EVAL_1935 == 32'h24;
  assign _EVAL_5700 = _EVAL_1242 & 32'h40000060;
  assign _EVAL_2994 = _EVAL_5700 == 32'h40;
  assign _EVAL_1823 = _EVAL_674 | _EVAL_2994;
  assign _EVAL_2551 = _EVAL_1823 | _EVAL_677;
  assign _EVAL_3431 = _EVAL_1074 ? _EVAL_2551 : _EVAL_4421;
  assign _EVAL_3971 = _EVAL_5926 ? _EVAL_1307 : _EVAL_3431;
  assign _EVAL_1115 = _EVAL_2970 ? _EVAL_1307 : _EVAL_3971;
  assign _EVAL_4358 = _EVAL_2142 ? _EVAL_2521 : _EVAL_969;
  assign _EVAL_4342 = _EVAL_3052 ? _EVAL_3253 : _EVAL_4358;
  assign _EVAL_1752 = _EVAL_5833 ? _EVAL_1326 : _EVAL_3288;
  assign _EVAL_4588 = _EVAL_5833 ? _EVAL_3081 : _EVAL_1752;
  assign _EVAL_3531 = _EVAL_2142 ? _EVAL_459 : _EVAL_901;
  assign _EVAL_4139 = _EVAL_3052 ? _EVAL_2267 : _EVAL_3531;
  assign _EVAL_1351 = _EVAL_5276 ? _EVAL_4588 : _EVAL_4139;
  assign _EVAL_2727 = _EVAL_5690 ? _EVAL_3646 : _EVAL_3170;
  assign _EVAL_1166 = _EVAL_5337 ? _EVAL_2727 : _EVAL_4733;
  assign _EVAL_3914 = _EVAL_386 & 32'h4003044;
  assign _EVAL_4311 = _EVAL_3078 & 32'h2040;
  assign _EVAL_1867 = _EVAL_5833 ? _EVAL_2953 : _EVAL_4395;
  assign _EVAL_5427 = _EVAL_2970 ? _EVAL_5728 : _EVAL_5122;
  assign _EVAL_1254 = _EVAL_3052 ? _EVAL_5427 : _EVAL_3928;
  assign _EVAL_2080 = _EVAL_5276 ? _EVAL_1867 : _EVAL_1254;
  assign _EVAL_5780 = _EVAL_6134 | _EVAL_5728;
  assign _EVAL_1500 = _EVAL_2970 ? _EVAL_5780 : _EVAL_1115;
  assign _EVAL_605 = _EVAL_1930 ? _EVAL_1500 : _EVAL_1166;
  assign _EVAL_416 = _EVAL_2277 == 32'h0;
  assign _EVAL_2981 = _EVAL_4702 & 32'h60;
  assign _EVAL_6041 = _EVAL_2981 == 32'h0;
  assign _EVAL_5774 = _EVAL_416 | _EVAL_6041;
  assign _EVAL_732 = _EVAL_5774 | _EVAL_4710;
  assign _EVAL_3587 = _EVAL_4432 == 32'h4;
  assign _EVAL_5367 = _EVAL_732 | _EVAL_3587;
  assign _EVAL_4979 = _EVAL_4702 & 32'h62003010;
  assign _EVAL_435 = _EVAL_4979 == 32'h60000010;
  assign _EVAL_312 = _EVAL_5367 | _EVAL_435;
  assign _EVAL_804 = _EVAL_197 ? _EVAL_312 : _EVAL_4667;
  assign _EVAL_3838 = _EVAL_5854 & 32'h30;
  assign _EVAL_396 = _EVAL_3838 == 32'h30;
  assign _EVAL_4586 = _EVAL_856 | _EVAL_1539;
  assign _EVAL_355 = _EVAL_4586 | _EVAL_396;
  assign _EVAL_4782 = _EVAL_5854 & 32'h90000010;
  assign _EVAL_3302 = _EVAL_4782 == 32'h80000010;
  assign _EVAL_921 = _EVAL_355 | _EVAL_3302;
  assign _EVAL_3489 = _EVAL_921 & _EVAL_5207;
  assign _EVAL_4203 = _EVAL_5833 ? _EVAL_3489 : _EVAL_4454;
  assign _EVAL_1466 = _EVAL_5998 | _EVAL_3161;
  assign _EVAL_4488 = _EVAL_5690 ? _EVAL_1466 : _EVAL_5941;
  assign _EVAL_1862 = _EVAL_1978 & 32'h4024;
  assign _EVAL_3786 = _EVAL_1862 == 32'h20;
  assign _EVAL_2125 = _EVAL_6048 | _EVAL_3786;
  assign _EVAL_4786 = _EVAL_5341 == 32'h20;
  assign _EVAL_2548 = _EVAL_2125 | _EVAL_4786;
  assign _EVAL_3356 = _EVAL_5336 == 32'h2000;
  assign _EVAL_4713 = _EVAL_2548 | _EVAL_3356;
  assign _EVAL_1687 = _EVAL_3178 == 32'h90000010;
  assign _EVAL_2515 = _EVAL_4713 | _EVAL_1687;
  assign _EVAL_3177 = _EVAL_3050 ? _EVAL_2515 : _EVAL_5321;
  assign _EVAL_834 = _EVAL_1069 ? _EVAL_2515 : _EVAL_3177;
  assign _EVAL_4127 = _EVAL_5337 ? _EVAL_4488 : _EVAL_834;
  assign _EVAL_2535 = _EVAL_5302 == 32'h40;
  assign _EVAL_5761 = _EVAL_1958 ? _EVAL_551 : _EVAL_551;
  assign _EVAL_3873 = _EVAL_4554 ? _EVAL_551 : _EVAL_5761;
  assign _EVAL_4276 = _EVAL_197 ? _EVAL_551 : _EVAL_3873;
  assign _EVAL_5644 = _EVAL_197 ? 1'h0 : _EVAL_4276;
  assign _EVAL_2073 = _EVAL_197 ? _EVAL_2310 : _EVAL_1538;
  assign _EVAL_3833 = _EVAL_5690 ? _EVAL_4320 : _EVAL_4135;
  assign _EVAL_4874 = _EVAL_4899 == 32'h40;
  assign _EVAL_1233 = _EVAL_4311 == 32'h2040;
  assign _EVAL_3494 = _EVAL_4943 | _EVAL_1233;
  assign _EVAL_3941 = _EVAL_5984 | _EVAL_317;
  assign _EVAL_3561 = _EVAL_3941 | _EVAL_1556;
  assign _EVAL_3492 = _EVAL_1958 ? _EVAL_3347 : _EVAL_3561;
  assign _EVAL_3400 = _EVAL_4554 ? _EVAL_3494 : _EVAL_3492;
  assign _EVAL_3818 = _EVAL_5833 ? _EVAL_5162 : _EVAL_3438;
  assign _EVAL_1118 = _EVAL_3659 ? _EVAL_4273 : _EVAL_92;
  assign _EVAL_2889 = _EVAL_2142 ? _EVAL_2727 : _EVAL_4733;
  assign _EVAL_5242 = _EVAL_3052 ? _EVAL_1500 : _EVAL_2889;
  assign _EVAL_3853 = _EVAL_4743 & 32'h3c;
  assign _EVAL_3312 = _EVAL_3853 == 32'h4;
  assign _EVAL_702 = _EVAL_3312 | _EVAL_4714;
  assign _EVAL_4940 = _EVAL_702 | _EVAL_1433;
  assign _EVAL_4742 = _EVAL_5337 ? _EVAL_531 : _EVAL_5797;
  assign _EVAL_2037 = _EVAL_1930 ? _EVAL_4753 : _EVAL_4742;
  assign _EVAL_2830 = 3'h2 < _EVAL_3461;
  assign _EVAL_6104 = _EVAL_4793 ? 1'h1 : _EVAL_908;
  assign _EVAL_2957 = _EVAL_4702 & 32'h10000060;
  assign _EVAL_2847 = _EVAL_2957 == 32'h10000040;
  assign _EVAL_2903 = _EVAL_467 | _EVAL_2847;
  assign _EVAL_5837 = _EVAL_197 ? _EVAL_2903 : _EVAL_1497;
  assign _EVAL_2691 = _EVAL_3589 | _EVAL_2859;
  assign _EVAL_2423 = _EVAL_2691 | _EVAL_4685;
  assign _EVAL_309 = _EVAL_1791 == 32'h0;
  assign _EVAL_1138 = _EVAL_681 == 32'h2000;
  assign _EVAL_1425 = _EVAL_309 | _EVAL_1138;
  assign _EVAL_1444 = _EVAL_1425 | _EVAL_711;
  assign _EVAL_1706 = _EVAL_4554 ? _EVAL_1444 : _EVAL_797;
  assign _EVAL_3935 = _EVAL_197 ? _EVAL_1444 : _EVAL_1706;
  assign _EVAL_1387 = _EVAL_197 ? _EVAL_2423 : _EVAL_3935;
  assign _EVAL_4494 = _EVAL_197 ? _EVAL_3494 : _EVAL_3400;
  assign _EVAL_943 = _EVAL_4702 & 32'h2040;
  assign _EVAL_4866 = _EVAL_943 == 32'h2040;
  assign _EVAL_3756 = _EVAL_4952 | _EVAL_4866;
  assign _EVAL_506 = _EVAL_5337 ? _EVAL_3789 : _EVAL_2186;
  assign _EVAL_5552 = _EVAL_3659 ? _EVAL_701 : _EVAL_43;
  assign _EVAL_4720 = _EVAL_168 == 32'h4000040;
  assign _EVAL_5669 = _EVAL_1772 | _EVAL_4720;
  assign _EVAL_3733 = _EVAL_3914 == 32'h4000040;
  assign _EVAL_5769 = _EVAL_2799 | _EVAL_3733;
  assign _EVAL_5534 = _EVAL_5952 ? _EVAL_5669 : _EVAL_5769;
  assign _EVAL_5409 = _EVAL_3570 ? _EVAL_5461 : _EVAL_5534;
  assign _EVAL_966 = _EVAL_1946 | _EVAL_4874;
  assign _EVAL_6033 = _EVAL_4554 ? _EVAL_5297 : _EVAL_181;
  assign _EVAL_4847 = _EVAL_197 ? _EVAL_5297 : _EVAL_6033;
  assign _EVAL_3223 = _EVAL_197 ? _EVAL_4094 : _EVAL_4847;
  assign _EVAL_2167 = _EVAL_1889 & _EVAL_4445;
  assign _EVAL_5722 = {{29'd0}, _EVAL_858};
  assign _EVAL_3793 = _EVAL_3078[31:25];
  assign _EVAL_5869 = _EVAL_1947[31:25];
  assign _EVAL_829 = _EVAL_1958 ? _EVAL_1527 : _EVAL_5869;
  assign _EVAL_1906 = _EVAL_4554 ? _EVAL_3793 : _EVAL_829;
  assign _EVAL_796 = _EVAL_3659 ? _EVAL_3907 : _EVAL_47;
  assign _EVAL_2199 = _EVAL_1930 ? _EVAL_2267 : _EVAL_1861;
  assign _EVAL_2564 = _EVAL_5276 ? _EVAL_4203 : _EVAL_3475;
  assign _EVAL_1572 = _EVAL_1069 ? _EVAL_1957 : _EVAL_1341;
  assign _EVAL_5372 = _EVAL_5337 ? _EVAL_3833 : _EVAL_1572;
  assign _EVAL_3960 = _EVAL_2142 ? _EVAL_4798 : _EVAL_1486;
  assign _EVAL_4321 = _EVAL_3052 ? _EVAL_3351 : _EVAL_3960;
  assign _EVAL_4703 = _EVAL_4554 ? _EVAL_1294 : _EVAL_3562;
  assign _EVAL_5953 = _EVAL_197 ? _EVAL_1294 : _EVAL_4703;
  assign _EVAL_4738 = _EVAL_5833 ? _EVAL_4146 : _EVAL_3818;
  assign _EVAL_3035 = _EVAL_2957 == 32'h40;
  assign _EVAL_4917 = _EVAL_654[19:15];
  assign _EVAL_4884 = _EVAL_4925 == 32'h10000040;
  assign _EVAL_4584 = _EVAL_4940 | _EVAL_4884;
  assign _EVAL_4178 = _EVAL_199 | _EVAL_2535;
  assign _EVAL_2040 = _EVAL_2142 ? _EVAL_4488 : _EVAL_834;
  assign _EVAL_3469 = _EVAL_3052 ? _EVAL_5198 : _EVAL_2040;
  assign _EVAL_1711 = _EVAL_5276 ? _EVAL_4738 : _EVAL_3469;
  assign _EVAL_4475 = _EVAL_5833 ? _EVAL_5461 : _EVAL_5409;
  assign _EVAL_3698 = _EVAL_5833 ? _EVAL_3199 : _EVAL_4475;
  assign _EVAL_2959 = _EVAL_654[24:20];
  assign _EVAL_685 = _EVAL_197 ? _EVAL_2959 : _EVAL_3945;
  assign _EVAL_1884 = _EVAL_5337 & _EVAL_2830;
  assign _EVAL_4099 = _EVAL_799 | _EVAL_1884;
  assign _EVAL_3072 = _EVAL_5386[31:25];
  assign _EVAL_588 = _EVAL_654[31:25];
  assign _EVAL_3500 = _EVAL_197 ? _EVAL_3793 : _EVAL_1906;
  assign _EVAL_3240 = _EVAL_197 ? _EVAL_588 : _EVAL_3500;
  assign _EVAL_2796 = _EVAL_2089 & _EVAL_4984;
  assign _EVAL_1406 = _EVAL_5600 ? 1'h0 : _EVAL_245;
  assign _EVAL_4097 = _EVAL_4774 ? 1'h1 : _EVAL_1406;
  assign _EVAL_2010 = _EVAL_1930 ? _EVAL_5198 : _EVAL_4127;
  assign _EVAL_3339 = _EVAL_2796 != 4'h0;
  assign _EVAL_1052 = _EVAL_5335 ? 1'h1 : _EVAL_3339;
  assign _EVAL_200 = _EVAL_5276 ? _EVAL_4455 : _EVAL_4321;
  assign _EVAL_4179 = _EVAL_5126 == 32'h10000040;
  assign _EVAL_257 = _EVAL_5572 | _EVAL_4179;
  assign _EVAL_709 = _EVAL_5833 ? _EVAL_4469 : _EVAL_3488;
  assign _EVAL_1456 = _EVAL_5833 ? _EVAL_3072 : _EVAL_709;
  assign _EVAL_5765 = _EVAL_5276 ? _EVAL_1456 : _EVAL_468;
  assign _EVAL_6116 = _EVAL_966 | _EVAL_160;
  assign _EVAL_2887 = _EVAL_5337 ? _EVAL_2324 : _EVAL_1066;
  assign _EVAL_2575 = _EVAL_1930 ? _EVAL_4759 : _EVAL_2887;
  assign _EVAL_5079 = _EVAL_5276 ? _EVAL_3452 : _EVAL_4131;
  assign _EVAL_3128 = _EVAL_5833 ? _EVAL_5888 : _EVAL_4902;
  assign _EVAL_611 = _EVAL_5833 ? _EVAL_301 : _EVAL_3128;
  assign _EVAL_4996 = _EVAL_2621 | _EVAL_1594;
  assign _EVAL_4522 = _EVAL_5952 ? _EVAL_4584 : _EVAL_6015;
  assign _EVAL_4280 = _EVAL_3570 ? _EVAL_4996 : _EVAL_4522;
  assign _EVAL_422 = _EVAL_5833 ? _EVAL_4996 : _EVAL_4280;
  assign _EVAL_5707 = _EVAL_5833 ? _EVAL_257 : _EVAL_422;
  assign _EVAL_1530 = _EVAL_3659 ? _EVAL_2740 : _EVAL_117;
  assign _EVAL_3383 = _EVAL_5833 ? _EVAL_4304 : _EVAL_2561;
  assign _EVAL_2004 = _EVAL_3659 ? _EVAL_4123 : _EVAL_122;
  assign _EVAL_818 = _EVAL_1930 ? _EVAL_4448 : _EVAL_5299;
  assign _EVAL_4967 = _EVAL_4178 | _EVAL_2310;
  assign _EVAL_1740 = _EVAL_5833 ? _EVAL_1865 : _EVAL_971;
  assign _EVAL_4265 = _EVAL_3900 & _EVAL_4445;
  assign _EVAL_2997 = _EVAL_1395 == 32'h40;
  assign _EVAL_4335 = _EVAL_5933 | _EVAL_2997;
  assign _EVAL_4033 = _EVAL_3659 ? _EVAL_5701 : _EVAL_1;
  assign _EVAL_4431 = _EVAL_1709 | _EVAL_3035;
  assign _EVAL_5379 = _EVAL_4335 | _EVAL_2596;
  assign _EVAL_4077 = _EVAL_1958 ? _EVAL_5379 : _EVAL_6116;
  assign _EVAL_2380 = _EVAL_4554 ? _EVAL_4967 : _EVAL_4077;
  assign _EVAL_3862 = _EVAL_197 ? _EVAL_4967 : _EVAL_2380;
  assign _EVAL_1127 = 3'h3 < _EVAL_3461;
  assign _EVAL_5308 = _EVAL_5833 ? _EVAL_2272 : _EVAL_3383;
  assign _EVAL_1190 = _EVAL_5276 ? _EVAL_5308 : _EVAL_1983;
  assign _EVAL_3073 = _EVAL_1930 ? _EVAL_4145 : _EVAL_5372;
  assign _EVAL_1813 = _EVAL_3659 ? _EVAL_1563 : _EVAL_13;
  assign _EVAL_1447 = _EVAL_197 ? _EVAL_4636 : _EVAL_2073;
  assign _EVAL_1748 = _EVAL_2142 ? _EVAL_3833 : _EVAL_1572;
  assign _EVAL_3324 = _EVAL_3052 ? _EVAL_4145 : _EVAL_1748;
  assign _EVAL_4122 = _EVAL_5337 ? _EVAL_3132 : _EVAL_3569;
  assign _EVAL_5666 = _EVAL_1930 ? _EVAL_5554 : _EVAL_4122;
  assign _EVAL_970 = _EVAL_197 ? _EVAL_1321 : _EVAL_5953;
  assign _EVAL_6102 = _EVAL_3659 ? _EVAL_2281 : _EVAL_8;
  assign _EVAL_3959 = _EVAL_197 ? _EVAL_4917 : _EVAL_5447;
  assign _EVAL_4966 = _EVAL_3659 ? _EVAL_4261 : _EVAL_61;
  assign _EVAL_1765 = _EVAL_5276 ? _EVAL_1740 : _EVAL_3324;
  assign _EVAL_2721 = _EVAL_5276 ? _EVAL_3698 : _EVAL_2634;
  assign _EVAL_1758 = _EVAL_5276 ? _EVAL_5707 : _EVAL_4326;
  assign _EVAL_5591 = _EVAL_4431 | _EVAL_4636;
  assign _EVAL_5045 = _EVAL_3659 ? _EVAL_2135 : _EVAL_75;
  assign _EVAL_724 = _EVAL_1930 ? _EVAL_2565 : _EVAL_2974;
  assign _EVAL_1158 = _EVAL_5276 ? _EVAL_6050 : _EVAL_4342;
  assign _EVAL_3801 = _EVAL_197 ? _EVAL_3756 : _EVAL_4494;
  assign _EVAL_440 = _EVAL_197 ? 1'h0 : 1'h1;
  assign _EVAL_4533 = _EVAL_532 + _EVAL_960;
  assign _EVAL_6098 = _EVAL_3659 ? _EVAL_2202 : _EVAL_110;
  assign _EVAL_2743 = _EVAL_5276 ? _EVAL_611 : _EVAL_5242;
  assign _EVAL_3918 = _EVAL_5985 & _EVAL_1127;
  assign _EVAL_1694 = _EVAL_197 ? _EVAL_5591 : _EVAL_3862;
  assign _EVAL_1896 = _EVAL_1930 ? _EVAL_5427 : _EVAL_506;
  assign _EVAL_3359 = _EVAL_5600 ? 1'h0 : 1'h1;
  assign _EVAL_5212 = _EVAL_113 ? _EVAL_693 : {{2'd0}, _EVAL_3403};
  assign _EVAL_2869 = _EVAL_2089 & _EVAL_4445;
  assign _EVAL_2724 = _EVAL_3659 ? _EVAL_788 : _EVAL_42;
  assign _EVAL_2962 = _EVAL_5600 ? _EVAL_5165 : _EVAL_2381;
  assign _EVAL_21 = _EVAL_5994 ? _EVAL_1052 : _EVAL_3339;
  assign _EVAL_87 = _EVAL_5994 ? _EVAL_2553 : _EVAL_2743;
  assign _EVAL_96 = _EVAL_5994 ? _EVAL_3223 : _EVAL_2291;
  assign _EVAL_7 = _EVAL_2869 != 4'h0;
  assign _EVAL_20 = _EVAL_5994 ? _EVAL_6098 : _EVAL_110;
  assign _EVAL_105 = _EVAL_1226 ? _EVAL_5707 : _EVAL_4543;
  assign _EVAL_157 = _EVAL_5994 ? _EVAL_6104 : _EVAL_908;
  assign _EVAL_138 = _EVAL_5994 ? _EVAL_2962 : _EVAL_2381;
  assign _EVAL_129 = _EVAL_5994 ? _EVAL_3205 : _EVAL_2564;
  assign _EVAL_111 = _EVAL_5994 ? _EVAL_3959 : _EVAL_3983;
  assign _EVAL_23 = _EVAL_586 != 4'h0;
  assign _EVAL_78 = _EVAL_5994 ? _EVAL_4966 : _EVAL_61;
  assign _EVAL_118 = _EVAL_5994 ? _EVAL_5837 : _EVAL_1758;
  assign _EVAL_58 = _EVAL_75;
  assign _EVAL_85 = _EVAL_5994 ? _EVAL_4426 : _EVAL_5588;
  assign _EVAL_97 = _EVAL_1226 ? _EVAL_1279 : _EVAL_818;
  assign _EVAL_80 = _EVAL_5994 ? _EVAL_4425 : _EVAL_108;
  assign _EVAL_124 = _EVAL_5994 ? _EVAL_5644 : _EVAL_1158;
  assign _EVAL_114 = _EVAL_5994 ? _EVAL_1387 : _EVAL_1765;
  assign _EVAL_68 = _EVAL_1226 ? _EVAL_4296 : _EVAL_5051;
  assign _EVAL_116 = _EVAL_5994 ? _EVAL_3188 : _EVAL_73;
  assign _EVAL_140 = _EVAL_5994 ? _EVAL_440 : _EVAL_5079;
  assign _EVAL_159 = _EVAL_1226 ? _EVAL_4738 : _EVAL_2010;
  assign _EVAL_18 = _EVAL_13;
  assign _EVAL_151 = _EVAL_143;
  assign _EVAL_94 = _EVAL_8;
  assign _EVAL_103 = _EVAL_4265 != 4'h0;
  assign _EVAL_109 = _EVAL_73;
  assign _EVAL_101 = _EVAL_5994 ? _EVAL_973 : _EVAL_29;
  assign _EVAL_30 = _EVAL_5994 ? _EVAL_1118 : _EVAL_92;
  assign _EVAL_36 = _EVAL_5994 ? _EVAL_2724 : _EVAL_42;
  assign _EVAL = _EVAL_5994 ? _EVAL_3144 : _EVAL_2998;
  assign _EVAL_0 = _EVAL_5994 ? _EVAL_685 : _EVAL_2343;
  assign _EVAL_99 = _EVAL_1226 ? _EVAL_5955 : _EVAL_724;
  assign _EVAL_62 = _EVAL_5994 ? _EVAL_804 : _EVAL_5642;
  assign _EVAL_84 = _EVAL_5994 ? _EVAL_5045 : _EVAL_75;
  assign _EVAL_82 = _EVAL_5994 ? _EVAL_3314 : _EVAL_152;
  assign _EVAL_3 = _EVAL_1226 ? _EVAL_3452 : _EVAL_2377;
  assign _EVAL_10 = _EVAL_43;
  assign _EVAL_153 = _EVAL_1226 ? _EVAL_611 : _EVAL_605;
  assign _EVAL_115 = _EVAL_5994 ? _EVAL_1447 : _EVAL_2080;
  assign _EVAL_148 = _EVAL_5994 ? _EVAL_3249 : _EVAL_200;
  assign _EVAL_119 = _EVAL_532 + _EVAL_5722;
  assign _EVAL_128 = _EVAL_1226 ? _EVAL_3698 : _EVAL_5666;
  assign _EVAL_45 = _EVAL_5994 ? _EVAL_4033 : _EVAL_1;
  assign _EVAL_93 = _EVAL_108;
  assign _EVAL_133 = _EVAL_95;
  assign _EVAL_150 = _EVAL_1226 ? _EVAL_1456 : _EVAL_2575;
  assign _EVAL_63 = _EVAL_1226 ? _EVAL_5308 : _EVAL_748;
  assign _EVAL_123 = _EVAL_5994 ? _EVAL_970 : _EVAL_1190;
  assign _EVAL_65 = _EVAL_5994 ? _EVAL_2008 : _EVAL_127;
  assign _EVAL_34 = _EVAL_5437;
  assign _EVAL_74 = _EVAL_1226 ? _EVAL_1740 : _EVAL_3073;
  assign _EVAL_59 = _EVAL_5994 ? _EVAL_6102 : _EVAL_8;
  assign _EVAL_22 = _EVAL_122;
  assign _EVAL_35 = _EVAL_5994 ? _EVAL_3359 : 1'h0;
  assign _EVAL_40 = _EVAL_29;
  assign _EVAL_106 = _EVAL_5994 ? _EVAL_2004 : _EVAL_122;
  assign _EVAL_11 = _EVAL_5994 ? _EVAL_4356 : _EVAL_1711;
  assign _EVAL_5 = _EVAL_5994 ? _EVAL_3801 : _EVAL_1351;
  assign _EVAL_41 = _EVAL_1226 ? _EVAL_2141 : _EVAL_5368;
  assign _EVAL_149 = _EVAL_1;
  assign _EVAL_50 = _EVAL_3266 != 4'h0;
  assign _EVAL_112 = _EVAL_1226 ? _EVAL_4588 : _EVAL_2199;
  assign _EVAL_158 = _EVAL_1226 ? _EVAL_5607 : _EVAL_2037;
  assign _EVAL_125 = _EVAL_5994 ? _EVAL_1530 : _EVAL_117;
  assign _EVAL_54 = _EVAL_4099 | _EVAL_3918;
  assign _EVAL_38 = _EVAL_1226 ? _EVAL_3456 : _EVAL_5237;
  assign _EVAL_81 = _EVAL_3771 != 4'h0;
  assign _EVAL_14 = _EVAL_1226 ? _EVAL_4203 : _EVAL_3998;
  assign _EVAL_70 = _EVAL_5994 ? _EVAL_1813 : _EVAL_13;
  assign _EVAL_69 = _EVAL_5994 ? _EVAL_2567 : _EVAL_1750;
  assign _EVAL_28 = _EVAL_5994 ? _EVAL_796 : _EVAL_47;
  assign _EVAL_113 = _EVAL_5052 & _EVAL_4675;
  assign _EVAL_120 = _EVAL_61;
  assign _EVAL_130 = _EVAL_5994 ? _EVAL_4664 : _EVAL_4533;
  assign _EVAL_71 = _EVAL_5994 ? _EVAL_3433 : _EVAL_12;
  assign _EVAL_86 = _EVAL_42;
  assign _EVAL_37 = _EVAL_1226 ? _EVAL_1867 : _EVAL_1896;
  assign _EVAL_83 = _EVAL_5994 ? _EVAL_4097 : _EVAL_245;
  assign _EVAL_16 = _EVAL_110;
  assign _EVAL_121 = _EVAL_5994 ? _EVAL_5951 : _EVAL_143;
  assign _EVAL_155 = _EVAL_47;
  assign _EVAL_141 = _EVAL_5994 ? _EVAL_1694 : _EVAL_4378;
  assign _EVAL_137 = _EVAL_1226 ? _EVAL_4455 : _EVAL_1363;
  assign _EVAL_15 = _EVAL_92;
  assign _EVAL_146 = _EVAL_152;
  assign _EVAL_46 = _EVAL_26 & _EVAL_1959;
  assign _EVAL_131 = _EVAL_5994 ? _EVAL_5552 : _EVAL_43;
  assign _EVAL_135 = _EVAL_2167 != 4'h0;
  assign _EVAL_17 = _EVAL_12;
  assign _EVAL_88 = _EVAL_5994 ? _EVAL_3240 : _EVAL_5765;
  assign _EVAL_76 = _EVAL_5994 ? _EVAL_2447 : _EVAL_4006;
  assign _EVAL_2 = _EVAL_117;
  assign _EVAL_134 = _EVAL_127;
  assign _EVAL_4 = _EVAL_5994 ? _EVAL_4849 : _EVAL_2721;
  assign _EVAL_55 = _EVAL_1226 ? _EVAL_6050 : _EVAL_5328;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_372 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_701 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_717 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_718 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_788 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_815 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_1171 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_1563 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_1726 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_2135 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_2202 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_2241 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_2281 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {4{`RANDOM}};
  _EVAL_2740 = _RAND_13[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_3403 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_3526 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_3907 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_4123 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_4261 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_4273 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_4664 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_4774 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_4793 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_5094 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_5165 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_5225 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_5335 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_5437 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_5648 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_5701 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_5994 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_6019 = _RAND_31[14:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_51) begin
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_372 <= _EVAL_143;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_701 <= _EVAL_43;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_717 <= _EVAL_127;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_718 <= _EVAL_12;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_788 <= _EVAL_42;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_815 <= _EVAL_29;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        if (_EVAL_1365) begin
          _EVAL_1171 <= 1'h1;
        end else begin
          if (_EVAL_314) begin
            _EVAL_1171 <= 1'h1;
          end else begin
            _EVAL_1171 <= _EVAL_5852;
          end
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_1563 <= _EVAL_13;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_1726 <= _EVAL_73;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_2135 <= _EVAL_75;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_2202 <= _EVAL_110;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        if (_EVAL_1660) begin
          _EVAL_2241 <= 1'h1;
        end else begin
          if (_EVAL_4736) begin
            _EVAL_2241 <= 1'h1;
          end else begin
            _EVAL_2241 <= _EVAL_5518;
          end
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_2281 <= _EVAL_8;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_2740 <= _EVAL_117;
      end
    end
    _EVAL_3403 <= _EVAL_5212[1:0];
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        if (_EVAL_3955) begin
          _EVAL_3526 <= _EVAL_2086;
        end else begin
          if (_EVAL_1365) begin
            _EVAL_3526 <= _EVAL_5417;
          end else begin
            if (_EVAL_1660) begin
              _EVAL_3526 <= _EVAL_1015;
            end else begin
              if (_EVAL_5472) begin
                _EVAL_3526 <= _EVAL_5787;
              end else begin
                _EVAL_3526 <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_3907 <= _EVAL_47;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_4123 <= _EVAL_122;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_4261 <= _EVAL_61;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_4273 <= _EVAL_92;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_4664 <= _EVAL_6115;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_4774 <= _EVAL_95;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        if (_EVAL_5472) begin
          _EVAL_4793 <= 1'h1;
        end else begin
          if (_EVAL_5748) begin
            _EVAL_4793 <= 1'h1;
          end else begin
            _EVAL_4793 <= _EVAL_6011;
          end
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_5094 <= _EVAL_2666;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        if (_EVAL_3955) begin
          _EVAL_5165 <= _EVAL_2357;
        end else begin
          if (_EVAL_1365) begin
            _EVAL_5165 <= _EVAL_527;
          end else begin
            if (_EVAL_1660) begin
              _EVAL_5165 <= _EVAL_3758;
            end else begin
              if (_EVAL_5472) begin
                _EVAL_5165 <= _EVAL_1048;
              end else begin
                _EVAL_5165 <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_5225 <= _EVAL_152;
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        if (_EVAL_3955) begin
          _EVAL_5335 <= 1'h1;
        end else begin
          if (_EVAL_661) begin
            _EVAL_5335 <= 1'h1;
          end else begin
            _EVAL_5335 <= _EVAL_4700;
          end
        end
      end
    end
    _EVAL_5437 <= _EVAL_52 & _EVAL_5957;
    if (_EVAL_66) begin
      _EVAL_5648 <= 1'h0;
    end else begin
      if (_EVAL_5414) begin
        _EVAL_5648 <= 1'h0;
      end else begin
        if (_EVAL_113) begin
          _EVAL_5648 <= 1'h1;
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_5701 <= _EVAL_1;
      end
    end
    if (_EVAL_66) begin
      _EVAL_5994 <= 1'h0;
    end else begin
      if (_EVAL_5414) begin
        _EVAL_5994 <= _EVAL_3810;
      end else begin
        if (_EVAL_113) begin
          _EVAL_5994 <= 1'h0;
        end
      end
    end
    if (_EVAL_5414) begin
      if (_EVAL_3810) begin
        _EVAL_6019 <= _EVAL_108;
      end
    end
  end
endmodule
