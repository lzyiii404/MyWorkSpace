//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_320(
  input  [63:0] _EVAL,
  input         _EVAL_0,
  output [31:0] _EVAL_1,
  output [6:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  output        _EVAL_5,
  output [2:0]  _EVAL_6,
  input  [63:0] _EVAL_7,
  input  [31:0] _EVAL_8,
  output [8:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  output [2:0]  _EVAL_14,
  output [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [6:0]  _EVAL_21,
  input         _EVAL_22,
  input  [2:0]  _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output [1:0]  _EVAL_26,
  output [63:0] _EVAL_27,
  input  [63:0] _EVAL_28,
  output        _EVAL_29,
  input  [2:0]  _EVAL_30,
  output [31:0] _EVAL_31,
  input  [8:0]  _EVAL_32,
  input         _EVAL_33,
  output        _EVAL_34,
  output [2:0]  _EVAL_35,
  output [7:0]  _EVAL_36,
  input  [2:0]  _EVAL_37,
  output        _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  output        _EVAL_43,
  output [1:0]  _EVAL_44,
  output        _EVAL_45,
  input  [6:0]  _EVAL_46,
  input         _EVAL_47,
  output [2:0]  _EVAL_48,
  input  [7:0]  _EVAL_49,
  output [63:0] _EVAL_50,
  input  [31:0] _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53
);
  wire  TLBroadcastTracker_1__EVAL;
  wire  TLBroadcastTracker_1__EVAL_0;
  wire  TLBroadcastTracker_1__EVAL_1;
  wire  TLBroadcastTracker_1__EVAL_2;
  wire  TLBroadcastTracker_1__EVAL_3;
  wire [6:0] TLBroadcastTracker_1__EVAL_4;
  wire  TLBroadcastTracker_1__EVAL_5;
  wire  TLBroadcastTracker_1__EVAL_6;
  wire [7:0] TLBroadcastTracker_1__EVAL_7;
  wire  TLBroadcastTracker_1__EVAL_8;
  wire [63:0] TLBroadcastTracker_1__EVAL_9;
  wire [2:0] TLBroadcastTracker_1__EVAL_10;
  wire [2:0] TLBroadcastTracker_1__EVAL_11;
  wire  TLBroadcastTracker_1__EVAL_12;
  wire  TLBroadcastTracker_1__EVAL_13;
  wire [31:0] TLBroadcastTracker_1__EVAL_14;
  wire [31:0] TLBroadcastTracker_1__EVAL_15;
  wire [2:0] TLBroadcastTracker_1__EVAL_16;
  wire [2:0] TLBroadcastTracker_1__EVAL_17;
  wire [8:0] TLBroadcastTracker_1__EVAL_18;
  wire [25:0] TLBroadcastTracker_1__EVAL_19;
  wire [6:0] TLBroadcastTracker_1__EVAL_20;
  wire [7:0] TLBroadcastTracker_1__EVAL_21;
  wire  TLBroadcastTracker_1__EVAL_22;
  wire  TLBroadcastTracker_1__EVAL_23;
  wire [2:0] TLBroadcastTracker_1__EVAL_24;
  wire  TLBroadcastTracker_1__EVAL_25;
  wire  TLBroadcastTracker_1__EVAL_26;
  wire [63:0] TLBroadcastTracker_1__EVAL_27;
  wire [2:0] TLBroadcastTracker_1__EVAL_28;
  wire  TLBroadcastTracker_1__EVAL_29;
  wire [7:0] TLBroadcastTracker__EVAL;
  wire  TLBroadcastTracker__EVAL_0;
  wire  TLBroadcastTracker__EVAL_1;
  wire [8:0] TLBroadcastTracker__EVAL_2;
  wire  TLBroadcastTracker__EVAL_3;
  wire  TLBroadcastTracker__EVAL_4;
  wire  TLBroadcastTracker__EVAL_5;
  wire [31:0] TLBroadcastTracker__EVAL_6;
  wire  TLBroadcastTracker__EVAL_7;
  wire [2:0] TLBroadcastTracker__EVAL_8;
  wire  TLBroadcastTracker__EVAL_9;
  wire [2:0] TLBroadcastTracker__EVAL_10;
  wire [63:0] TLBroadcastTracker__EVAL_11;
  wire  TLBroadcastTracker__EVAL_12;
  wire [2:0] TLBroadcastTracker__EVAL_13;
  wire  TLBroadcastTracker__EVAL_14;
  wire [2:0] TLBroadcastTracker__EVAL_15;
  wire [63:0] TLBroadcastTracker__EVAL_16;
  wire [25:0] TLBroadcastTracker__EVAL_17;
  wire [2:0] TLBroadcastTracker__EVAL_18;
  wire [31:0] TLBroadcastTracker__EVAL_19;
  wire  TLBroadcastTracker__EVAL_20;
  wire [7:0] TLBroadcastTracker__EVAL_21;
  wire  TLBroadcastTracker__EVAL_22;
  wire [6:0] TLBroadcastTracker__EVAL_23;
  wire  TLBroadcastTracker__EVAL_24;
  wire [2:0] TLBroadcastTracker__EVAL_25;
  wire  TLBroadcastTracker__EVAL_26;
  wire [6:0] TLBroadcastTracker__EVAL_27;
  wire  TLBroadcastTracker__EVAL_28;
  wire  TLBroadcastTracker__EVAL_29;
  reg [25:0] _EVAL_69;
  reg [31:0] _RAND_0;
  reg  _EVAL_81;
  reg [31:0] _RAND_1;
  reg  _EVAL_101;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_135;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_158;
  reg [31:0] _RAND_4;
  reg  _EVAL_197;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_267;
  reg [31:0] _RAND_6;
  reg  _EVAL_272;
  reg [31:0] _RAND_7;
  reg  _EVAL_276;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_322;
  reg [31:0] _RAND_9;
  reg  _EVAL_337;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_384;
  reg [31:0] _RAND_11;
  wire  _EVAL_140;
  wire  _EVAL_76;
  wire  _EVAL_260;
  wire  _EVAL_415;
  wire  _EVAL_116;
  wire [2:0] _EVAL_106;
  wire [3:0] _EVAL_145;
  wire [2:0] _EVAL_70;
  wire [2:0] _EVAL_354;
  wire [4:0] _EVAL_84;
  wire [2:0] _EVAL_356;
  wire [2:0] _EVAL_54;
  wire [3:0] _EVAL_144;
  wire [2:0] _EVAL_329;
  wire [2:0] _EVAL_175;
  wire  _EVAL_172;
  wire  _EVAL_194;
  wire  _EVAL_126;
  wire [122:0] _EVAL_151;
  wire [122:0] _EVAL_64;
  wire  _EVAL_321;
  wire [1:0] _EVAL_318;
  wire  _EVAL_401;
  wire  _EVAL_74;
  wire [2:0] _EVAL_269;
  wire [2:0] _EVAL_231;
  wire  _EVAL_315;
  wire [12:0] _EVAL_320;
  wire [5:0] _EVAL_300;
  wire [5:0] _EVAL_233;
  wire [2:0] _EVAL_195;
  wire [2:0] _EVAL_306;
  wire  _EVAL_271;
  wire  _EVAL_311;
  wire [1:0] _EVAL_188;
  wire [3:0] _EVAL_235;
  wire [2:0] _EVAL_313;
  wire [2:0] _EVAL_211;
  wire  _EVAL_292;
  wire  _EVAL_136;
  wire  _EVAL_56;
  wire  _EVAL_257;
  wire  _EVAL_153;
  wire  _EVAL_192;
  wire  _EVAL_103;
  wire  _EVAL_95;
  wire  _EVAL_208;
  wire  _EVAL_371;
  wire  _EVAL_281;
  wire  _EVAL_78;
  wire  _EVAL_73;
  wire  _EVAL_131;
  wire  _EVAL_123;
  wire  _EVAL_288;
  wire  _EVAL_277;
  wire  _EVAL_382;
  wire  _EVAL_83;
  wire [2:0] _EVAL_254;
  wire  _EVAL_308;
  wire  _EVAL_65;
  wire  _EVAL_183;
  wire  _EVAL_59;
  wire  _EVAL_380;
  wire  _EVAL_206;
  wire  _EVAL_273;
  wire  _EVAL_307;
  wire [1:0] _EVAL_407;
  wire [2:0] _EVAL_331;
  wire [25:0] _EVAL_379;
  wire  _EVAL_255;
  wire  _EVAL_268;
  wire [1:0] _EVAL_262;
  wire  _EVAL_349;
  wire [2:0] _EVAL_79;
  wire [1:0] _EVAL_137;
  wire [1:0] _EVAL_325;
  wire [2:0] _EVAL_339;
  wire [2:0] _EVAL_159;
  wire [2:0] _EVAL_166;
  wire [2:0] _EVAL_215;
  wire  _EVAL_187;
  wire  _EVAL_399;
  wire  _EVAL_146;
  wire  _EVAL_370;
  wire  _EVAL_242;
  wire  _EVAL_124;
  wire [6:0] _EVAL_212;
  wire  _EVAL_147;
  wire  _EVAL_238;
  wire  _EVAL_222;
  wire  _EVAL_330;
  wire [1:0] _EVAL_250;
  wire  _EVAL_310;
  wire  _EVAL_75;
  wire  _EVAL_412;
  wire  _EVAL_89;
  wire  _EVAL_378;
  wire  _EVAL_243;
  wire  _EVAL_148;
  wire [1:0] _EVAL_229;
  wire [2:0] _EVAL_237;
  wire [1:0] _EVAL_191;
  wire [1:0] _EVAL_309;
  wire [2:0] _EVAL_130;
  wire [1:0] _EVAL_284;
  wire [1:0] _EVAL_275;
  wire  _EVAL_246;
  wire  _EVAL_164;
  wire  _EVAL_174;
  wire  _EVAL_293;
  wire  _EVAL_248;
  wire  _EVAL_94;
  wire  _EVAL_280;
  wire  _EVAL_141;
  wire [1:0] _EVAL_305;
  wire  _EVAL_156;
  wire  _EVAL_125;
  wire  _EVAL_189;
  wire [12:0] _EVAL_150;
  wire  _EVAL_184;
  wire  _EVAL_118;
  wire  _EVAL_154;
  wire  _EVAL_204;
  wire  _EVAL_361;
  wire  _EVAL_114;
  wire  _EVAL_63;
  wire  _EVAL_294;
  wire  _EVAL_120;
  wire  _EVAL_253;
  wire [1:0] _EVAL_352;
  wire [2:0] _EVAL_408;
  wire [2:0] _EVAL_397;
  wire  _EVAL_402;
  wire  _EVAL_227;
  wire  _EVAL_87;
  wire  _EVAL_152;
  wire  _EVAL_261;
  wire  _EVAL_369;
  wire  _EVAL_179;
  wire [1:0] _EVAL_143;
  wire [1:0] _EVAL_80;
  wire [1:0] _EVAL_247;
  wire [1:0] _EVAL_400;
  wire [1:0] _EVAL_224;
  wire [1:0] _EVAL_102;
  wire [1:0] _EVAL_113;
  wire [1:0] _EVAL_216;
  wire  _EVAL_139;
  wire  _EVAL_85;
  wire  _EVAL_180;
  wire  _EVAL_385;
  wire [5:0] _EVAL_341;
  wire  _EVAL_77;
  wire  _EVAL_57;
  wire  _EVAL_373;
  wire  _EVAL_377;
  wire [81:0] _EVAL_169;
  wire [81:0] _EVAL_335;
  wire  _EVAL_72;
  wire  _EVAL_171;
  wire  _EVAL_279;
  wire  _EVAL_357;
  wire [12:0] _EVAL_117;
  wire [5:0] _EVAL_282;
  wire [5:0] _EVAL_323;
  wire [2:0] _EVAL_223;
  wire [2:0] _EVAL_67;
  wire  _EVAL_342;
  wire  _EVAL_386;
  wire [12:0] _EVAL_362;
  wire [5:0] _EVAL_291;
  wire [5:0] _EVAL_176;
  wire [2:0] _EVAL_58;
  wire [2:0] _EVAL_111;
  wire [2:0] _EVAL_193;
  wire  _EVAL_326;
  wire  _EVAL_201;
  wire  _EVAL_96;
  wire  _EVAL_413;
  wire  _EVAL_91;
  wire  _EVAL_367;
  wire  _EVAL_363;
  wire [25:0] _EVAL_61;
  wire  _EVAL_417;
  wire  _EVAL_68;
  wire  _EVAL_336;
  wire  _EVAL_266;
  wire [12:0] _EVAL_207;
  wire [5:0] _EVAL_345;
  wire [5:0] _EVAL_162;
  wire [2:0] _EVAL_366;
  wire [2:0] _EVAL_395;
  wire [2:0] _EVAL_82;
  wire  _EVAL_383;
  wire [5:0] _EVAL_360;
  wire [2:0] _EVAL_332;
  wire [2:0] _EVAL_240;
  wire [2:0] _EVAL_286;
  wire [2:0] _EVAL_301;
  wire [2:0] _EVAL_365;
  wire  _EVAL_202;
  wire  _EVAL_259;
  wire  _EVAL_163;
  wire  _EVAL_219;
  wire  _EVAL_133;
  wire  _EVAL_119;
  wire  _EVAL_107;
  wire  _EVAL_66;
  wire  _EVAL_220;
  wire  _EVAL_350;
  wire  _EVAL_90;
  wire  _EVAL_388;
  wire  _EVAL_328;
  wire  _EVAL_285;
  wire [1:0] _EVAL_319;
  wire [1:0] _EVAL_62;
  wire [1:0] _EVAL_161;
  wire  _EVAL_358;
  wire [81:0] _EVAL_278;
  wire  _EVAL_346;
  wire  _EVAL_122;
  wire  _EVAL_92;
  wire  _EVAL_289;
  wire  _EVAL_128;
  wire  _EVAL_376;
  wire  _EVAL_115;
  wire [6:0] _EVAL_213;
  wire  _EVAL_344;
  wire  _EVAL_302;
  wire  _EVAL_105;
  wire  _EVAL_97;
  wire  _EVAL_263;
  wire  _EVAL_93;
  wire  _EVAL_416;
  wire  _EVAL_312;
  wire  _EVAL_340;
  wire  _EVAL_112;
  wire  _EVAL_177;
  wire  _EVAL_167;
  wire  _EVAL_108;
  wire  _EVAL_200;
  wire  _EVAL_299;
  wire  _EVAL_199;
  wire  _EVAL_387;
  wire  _EVAL_198;
  wire  _EVAL_99;
  wire  _EVAL_409;
  wire  _EVAL_88;
  wire  _EVAL_304;
  wire  _EVAL_60;
  wire  _EVAL_127;
  wire  _EVAL_410;
  wire [64:0] _EVAL_104;
  wire [104:0] _EVAL_316;
  wire  _EVAL_351;
  wire  _EVAL_155;
  wire [2:0] _EVAL_368;
  wire  _EVAL_186;
  wire  _EVAL_391;
  wire  _EVAL_334;
  wire [1:0] _EVAL_160;
  wire  _EVAL_264;
  wire  _EVAL_375;
  wire  _EVAL_374;
  wire [6:0] _EVAL_190;
  wire [6:0] _EVAL_182;
  wire [6:0] _EVAL_251;
  wire [122:0] _EVAL_347;
  wire [122:0] _EVAL_157;
  wire [2:0] _EVAL_178;
  wire  _EVAL_181;
  wire  _EVAL_55;
  wire  _EVAL_228;
  wire  _EVAL_218;
  wire  _EVAL_100;
  wire [122:0] _EVAL_209;
  wire [122:0] _EVAL_98;
  wire [122:0] _EVAL_245;
  wire  _EVAL_394;
  wire  _EVAL_142;
  wire [122:0] _EVAL_297;
  wire [81:0] _EVAL_405;
  wire  _EVAL_355;
  wire [2:0] _EVAL_324;
  wire  _EVAL_230;
  wire [81:0] _EVAL_225;
  wire  _EVAL_270;
  wire  _EVAL_256;
  wire  _EVAL_372;
  SiFive__EVAL_319 TLBroadcastTracker_1 (
    ._EVAL(TLBroadcastTracker_1__EVAL),
    ._EVAL_0(TLBroadcastTracker_1__EVAL_0),
    ._EVAL_1(TLBroadcastTracker_1__EVAL_1),
    ._EVAL_2(TLBroadcastTracker_1__EVAL_2),
    ._EVAL_3(TLBroadcastTracker_1__EVAL_3),
    ._EVAL_4(TLBroadcastTracker_1__EVAL_4),
    ._EVAL_5(TLBroadcastTracker_1__EVAL_5),
    ._EVAL_6(TLBroadcastTracker_1__EVAL_6),
    ._EVAL_7(TLBroadcastTracker_1__EVAL_7),
    ._EVAL_8(TLBroadcastTracker_1__EVAL_8),
    ._EVAL_9(TLBroadcastTracker_1__EVAL_9),
    ._EVAL_10(TLBroadcastTracker_1__EVAL_10),
    ._EVAL_11(TLBroadcastTracker_1__EVAL_11),
    ._EVAL_12(TLBroadcastTracker_1__EVAL_12),
    ._EVAL_13(TLBroadcastTracker_1__EVAL_13),
    ._EVAL_14(TLBroadcastTracker_1__EVAL_14),
    ._EVAL_15(TLBroadcastTracker_1__EVAL_15),
    ._EVAL_16(TLBroadcastTracker_1__EVAL_16),
    ._EVAL_17(TLBroadcastTracker_1__EVAL_17),
    ._EVAL_18(TLBroadcastTracker_1__EVAL_18),
    ._EVAL_19(TLBroadcastTracker_1__EVAL_19),
    ._EVAL_20(TLBroadcastTracker_1__EVAL_20),
    ._EVAL_21(TLBroadcastTracker_1__EVAL_21),
    ._EVAL_22(TLBroadcastTracker_1__EVAL_22),
    ._EVAL_23(TLBroadcastTracker_1__EVAL_23),
    ._EVAL_24(TLBroadcastTracker_1__EVAL_24),
    ._EVAL_25(TLBroadcastTracker_1__EVAL_25),
    ._EVAL_26(TLBroadcastTracker_1__EVAL_26),
    ._EVAL_27(TLBroadcastTracker_1__EVAL_27),
    ._EVAL_28(TLBroadcastTracker_1__EVAL_28),
    ._EVAL_29(TLBroadcastTracker_1__EVAL_29)
  );
  SiFive__EVAL_318 TLBroadcastTracker (
    ._EVAL(TLBroadcastTracker__EVAL),
    ._EVAL_0(TLBroadcastTracker__EVAL_0),
    ._EVAL_1(TLBroadcastTracker__EVAL_1),
    ._EVAL_2(TLBroadcastTracker__EVAL_2),
    ._EVAL_3(TLBroadcastTracker__EVAL_3),
    ._EVAL_4(TLBroadcastTracker__EVAL_4),
    ._EVAL_5(TLBroadcastTracker__EVAL_5),
    ._EVAL_6(TLBroadcastTracker__EVAL_6),
    ._EVAL_7(TLBroadcastTracker__EVAL_7),
    ._EVAL_8(TLBroadcastTracker__EVAL_8),
    ._EVAL_9(TLBroadcastTracker__EVAL_9),
    ._EVAL_10(TLBroadcastTracker__EVAL_10),
    ._EVAL_11(TLBroadcastTracker__EVAL_11),
    ._EVAL_12(TLBroadcastTracker__EVAL_12),
    ._EVAL_13(TLBroadcastTracker__EVAL_13),
    ._EVAL_14(TLBroadcastTracker__EVAL_14),
    ._EVAL_15(TLBroadcastTracker__EVAL_15),
    ._EVAL_16(TLBroadcastTracker__EVAL_16),
    ._EVAL_17(TLBroadcastTracker__EVAL_17),
    ._EVAL_18(TLBroadcastTracker__EVAL_18),
    ._EVAL_19(TLBroadcastTracker__EVAL_19),
    ._EVAL_20(TLBroadcastTracker__EVAL_20),
    ._EVAL_21(TLBroadcastTracker__EVAL_21),
    ._EVAL_22(TLBroadcastTracker__EVAL_22),
    ._EVAL_23(TLBroadcastTracker__EVAL_23),
    ._EVAL_24(TLBroadcastTracker__EVAL_24),
    ._EVAL_25(TLBroadcastTracker__EVAL_25),
    ._EVAL_26(TLBroadcastTracker__EVAL_26),
    ._EVAL_27(TLBroadcastTracker__EVAL_27),
    ._EVAL_28(TLBroadcastTracker__EVAL_28),
    ._EVAL_29(TLBroadcastTracker__EVAL_29)
  );
  assign _EVAL_140 = _EVAL_322 == 3'h0;
  assign _EVAL_76 = _EVAL_20 == 3'h5;
  assign _EVAL_260 = _EVAL_20 == 3'h7;
  assign _EVAL_415 = _EVAL_76 | _EVAL_260;
  assign _EVAL_116 = _EVAL_3 & _EVAL_415;
  assign _EVAL_106 = {TLBroadcastTracker_1__EVAL_25,TLBroadcastTracker__EVAL_29,_EVAL_116};
  assign _EVAL_145 = {_EVAL_106, 1'h0};
  assign _EVAL_70 = _EVAL_145[2:0];
  assign _EVAL_354 = _EVAL_106 | _EVAL_70;
  assign _EVAL_84 = {_EVAL_354, 2'h0};
  assign _EVAL_356 = _EVAL_84[2:0];
  assign _EVAL_54 = _EVAL_354 | _EVAL_356;
  assign _EVAL_144 = {_EVAL_54, 1'h0};
  assign _EVAL_329 = _EVAL_144[2:0];
  assign _EVAL_175 = ~ _EVAL_329;
  assign _EVAL_172 = _EVAL_175[2];
  assign _EVAL_194 = _EVAL_172 & TLBroadcastTracker_1__EVAL_25;
  assign _EVAL_126 = _EVAL_140 ? _EVAL_194 : _EVAL_337;
  assign _EVAL_151 = {TLBroadcastTracker_1__EVAL_24,TLBroadcastTracker_1__EVAL_17,TLBroadcastTracker_1__EVAL_28,TLBroadcastTracker_1__EVAL_18,TLBroadcastTracker_1__EVAL_14,TLBroadcastTracker_1__EVAL_21,TLBroadcastTracker_1__EVAL_27,1'h0};
  assign _EVAL_64 = _EVAL_126 ? _EVAL_151 : 123'h0;
  assign _EVAL_321 = _EVAL_135 == 3'h1;
  assign _EVAL_318 = _EVAL_32[8:7];
  assign _EVAL_401 = _EVAL_318[1];
  assign _EVAL_74 = _EVAL_11[0];
  assign _EVAL_269 = _EVAL_74 ? 3'h5 : 3'h6;
  assign _EVAL_231 = _EVAL_401 ? _EVAL_269 : _EVAL_11;
  assign _EVAL_315 = _EVAL_231[0];
  assign _EVAL_320 = 13'h3f << _EVAL_4;
  assign _EVAL_300 = _EVAL_320[5:0];
  assign _EVAL_233 = ~ _EVAL_300;
  assign _EVAL_195 = _EVAL_233[5:3];
  assign _EVAL_306 = _EVAL_315 ? _EVAL_195 : 3'h0;
  assign _EVAL_271 = _EVAL_306 == 3'h0;
  assign _EVAL_311 = _EVAL_321 | _EVAL_271;
  assign _EVAL_188 = _EVAL_23[1:0];
  assign _EVAL_235 = 4'h1 << _EVAL_188;
  assign _EVAL_313 = _EVAL_235[2:0];
  assign _EVAL_211 = _EVAL_313 | 3'h1;
  assign _EVAL_292 = _EVAL_211[0];
  assign _EVAL_136 = _EVAL_51[2];
  assign _EVAL_56 = _EVAL_136 == 1'h0;
  assign _EVAL_257 = _EVAL_51[1];
  assign _EVAL_153 = _EVAL_257 == 1'h0;
  assign _EVAL_192 = _EVAL_56 & _EVAL_153;
  assign _EVAL_103 = _EVAL_51[0];
  assign _EVAL_95 = _EVAL_103 == 1'h0;
  assign _EVAL_208 = _EVAL_192 & _EVAL_95;
  assign _EVAL_371 = _EVAL_292 & _EVAL_208;
  assign _EVAL_281 = _EVAL_116 | TLBroadcastTracker__EVAL_29;
  assign _EVAL_78 = _EVAL_281 | TLBroadcastTracker_1__EVAL_25;
  assign _EVAL_73 = _EVAL_276 ? _EVAL_116 : 1'h0;
  assign _EVAL_131 = _EVAL_272 ? TLBroadcastTracker__EVAL_29 : 1'h0;
  assign _EVAL_123 = _EVAL_73 | _EVAL_131;
  assign _EVAL_288 = _EVAL_337 ? TLBroadcastTracker_1__EVAL_25 : 1'h0;
  assign _EVAL_277 = _EVAL_123 | _EVAL_288;
  assign _EVAL_382 = _EVAL_140 ? _EVAL_78 : _EVAL_277;
  assign _EVAL_83 = _EVAL_13 & _EVAL_382;
  assign _EVAL_254 = {{2'd0}, _EVAL_83};
  assign _EVAL_308 = _EVAL_175[0];
  assign _EVAL_65 = _EVAL_308 & _EVAL_116;
  assign _EVAL_183 = _EVAL_175[1];
  assign _EVAL_59 = _EVAL_183 & TLBroadcastTracker__EVAL_29;
  assign _EVAL_380 = TLBroadcastTracker_1__EVAL_24[2];
  assign _EVAL_206 = _EVAL_380 == 1'h0;
  assign _EVAL_273 = TLBroadcastTracker_1__EVAL_29;
  assign _EVAL_307 = TLBroadcastTracker__EVAL_3;
  assign _EVAL_407 = {_EVAL_273,_EVAL_307};
  assign _EVAL_331 = {{1'd0}, _EVAL_407};
  assign _EVAL_379 = _EVAL_8[31:6];
  assign _EVAL_255 = TLBroadcastTracker_1__EVAL_19 == _EVAL_379;
  assign _EVAL_268 = TLBroadcastTracker__EVAL_17 == _EVAL_379;
  assign _EVAL_262 = {_EVAL_255,_EVAL_268};
  assign _EVAL_349 = _EVAL_262 != 2'h0;
  assign _EVAL_79 = {_EVAL_407, 1'h0};
  assign _EVAL_137 = _EVAL_79[1:0];
  assign _EVAL_325 = _EVAL_407 | _EVAL_137;
  assign _EVAL_339 = {_EVAL_325, 1'h0};
  assign _EVAL_159 = ~ _EVAL_339;
  assign _EVAL_166 = _EVAL_331 & _EVAL_159;
  assign _EVAL_215 = _EVAL_349 ? {{1'd0}, _EVAL_262} : _EVAL_166;
  assign _EVAL_187 = _EVAL_215[0];
  assign _EVAL_399 = _EVAL_215[1];
  assign _EVAL_146 = _EVAL_23 >= 3'h3;
  assign _EVAL_370 = _EVAL_211[2];
  assign _EVAL_242 = _EVAL_370 & _EVAL_56;
  assign _EVAL_124 = _EVAL_146 | _EVAL_242;
  assign _EVAL_212 = _EVAL_32[6:0];
  assign _EVAL_147 = TLBroadcastTracker_1__EVAL_20 == _EVAL_212;
  assign _EVAL_238 = TLBroadcastTracker_1__EVAL_6 & _EVAL_147;
  assign _EVAL_222 = TLBroadcastTracker__EVAL_23 == _EVAL_212;
  assign _EVAL_330 = TLBroadcastTracker__EVAL_22 & _EVAL_222;
  assign _EVAL_250 = {_EVAL_238,_EVAL_330};
  assign _EVAL_310 = _EVAL_250[0];
  assign _EVAL_75 = _EVAL_267 == 3'h0;
  assign _EVAL_412 = _EVAL_318 == 2'h1;
  assign _EVAL_89 = _EVAL_412 == 1'h0;
  assign _EVAL_378 = _EVAL_22 & _EVAL_89;
  assign _EVAL_243 = _EVAL_20 == 3'h6;
  assign _EVAL_148 = _EVAL_3 & _EVAL_243;
  assign _EVAL_229 = {_EVAL_378,_EVAL_148};
  assign _EVAL_237 = {_EVAL_229, 1'h0};
  assign _EVAL_191 = _EVAL_237[1:0];
  assign _EVAL_309 = _EVAL_229 | _EVAL_191;
  assign _EVAL_130 = {_EVAL_309, 1'h0};
  assign _EVAL_284 = _EVAL_130[1:0];
  assign _EVAL_275 = ~ _EVAL_284;
  assign _EVAL_246 = _EVAL_275[1];
  assign _EVAL_164 = _EVAL_75 ? _EVAL_246 : _EVAL_197;
  assign _EVAL_174 = _EVAL_10 & _EVAL_164;
  assign _EVAL_293 = _EVAL_174 & _EVAL_378;
  assign _EVAL_248 = _EVAL_310 & _EVAL_293;
  assign _EVAL_94 = _EVAL_401 == 1'h0;
  assign _EVAL_280 = _EVAL_74 | _EVAL_94;
  assign _EVAL_141 = _EVAL_248 & _EVAL_280;
  assign _EVAL_305 = _EVAL_260 ? 2'h2 : 2'h1;
  assign _EVAL_156 = _EVAL_136 & _EVAL_257;
  assign _EVAL_125 = _EVAL_156 & _EVAL_95;
  assign _EVAL_189 = _EVAL_292 & _EVAL_125;
  assign _EVAL_150 = 13'h3f << TLBroadcastTracker_1__EVAL_28;
  assign _EVAL_184 = _EVAL_370 & _EVAL_136;
  assign _EVAL_118 = _EVAL_246 & _EVAL_378;
  assign _EVAL_154 = _EVAL_275[0];
  assign _EVAL_204 = _EVAL_75 ? _EVAL_154 : _EVAL_81;
  assign _EVAL_361 = _EVAL_158 == 3'h0;
  assign _EVAL_114 = _EVAL_361 == 1'h0;
  assign _EVAL_63 = _EVAL_101 == 1'h0;
  assign _EVAL_294 = _EVAL_114 | _EVAL_63;
  assign _EVAL_120 = TLBroadcastTracker_1__EVAL_8;
  assign _EVAL_253 = TLBroadcastTracker__EVAL_20;
  assign _EVAL_352 = {_EVAL_120,_EVAL_253};
  assign _EVAL_408 = {{1'd0}, _EVAL_352};
  assign _EVAL_397 = _EVAL_215 & _EVAL_408;
  assign _EVAL_402 = _EVAL_397 != 3'h0;
  assign _EVAL_227 = _EVAL_294 & _EVAL_402;
  assign _EVAL_87 = _EVAL_227 & _EVAL_39;
  assign _EVAL_152 = _EVAL_87 & _EVAL_361;
  assign _EVAL_261 = _EVAL_21 == 7'h40;
  assign _EVAL_369 = ~ _EVAL_261;
  assign _EVAL_179 = _EVAL_24 & _EVAL_101;
  assign _EVAL_143 = {{1'd0}, _EVAL_101};
  assign _EVAL_80 = {_EVAL_101, 1'h0};
  assign _EVAL_247 = ~ _EVAL_80;
  assign _EVAL_400 = _EVAL_143 & _EVAL_247;
  assign _EVAL_224 = ~ _EVAL_400;
  assign _EVAL_102 = _EVAL_143 & _EVAL_224;
  assign _EVAL_113 = _EVAL_179 ? _EVAL_102 : {{1'd0}, _EVAL_101};
  assign _EVAL_216 = _EVAL_152 ? {{1'd0}, _EVAL_369} : _EVAL_113;
  assign _EVAL_139 = _EVAL_174 | _EVAL_412;
  assign _EVAL_85 = _EVAL_30 == 3'h4;
  assign _EVAL_180 = _EVAL_156 & _EVAL_103;
  assign _EVAL_385 = _EVAL_292 & _EVAL_180;
  assign _EVAL_341 = _EVAL_150[5:0];
  assign _EVAL_77 = _EVAL_211[1];
  assign _EVAL_57 = 3'h2 == _EVAL_17;
  assign _EVAL_373 = _EVAL_154 & _EVAL_148;
  assign _EVAL_377 = _EVAL_75 ? _EVAL_373 : _EVAL_81;
  assign _EVAL_169 = {5'h18,_EVAL_23,_EVAL_46,67'h0};
  assign _EVAL_335 = _EVAL_377 ? _EVAL_169 : 82'h0;
  assign _EVAL_72 = 3'h2 == _EVAL_12;
  assign _EVAL_171 = 3'h1 == _EVAL_12;
  assign _EVAL_279 = _EVAL_17[2];
  assign _EVAL_357 = _EVAL_279 == 1'h0;
  assign _EVAL_117 = 13'h3f << _EVAL_37;
  assign _EVAL_282 = _EVAL_117[5:0];
  assign _EVAL_323 = ~ _EVAL_282;
  assign _EVAL_223 = _EVAL_323[5:3];
  assign _EVAL_67 = _EVAL_158 - 3'h1;
  assign _EVAL_342 = TLBroadcastTracker__EVAL_13[2];
  assign _EVAL_386 = _EVAL_342 == 1'h0;
  assign _EVAL_362 = 13'h3f << TLBroadcastTracker__EVAL_25;
  assign _EVAL_291 = _EVAL_362[5:0];
  assign _EVAL_176 = ~ _EVAL_291;
  assign _EVAL_58 = _EVAL_176[5:3];
  assign _EVAL_111 = _EVAL_386 ? _EVAL_58 : 3'h0;
  assign _EVAL_193 = _EVAL_59 ? _EVAL_111 : 3'h0;
  assign _EVAL_326 = _EVAL_20 == 3'h4;
  assign _EVAL_201 = _EVAL_10 & _EVAL_204;
  assign _EVAL_96 = _EVAL_140 ? _EVAL_308 : _EVAL_276;
  assign _EVAL_413 = _EVAL_13 & _EVAL_96;
  assign _EVAL_91 = _EVAL_243 ? _EVAL_201 : _EVAL_413;
  assign _EVAL_367 = _EVAL_326 | _EVAL_91;
  assign _EVAL_363 = _EVAL_367 & _EVAL_3;
  assign _EVAL_61 = _EVAL_51[31:6];
  assign _EVAL_417 = TLBroadcastTracker_1__EVAL_19 == _EVAL_61;
  assign _EVAL_68 = _EVAL_363 & _EVAL_417;
  assign _EVAL_336 = _EVAL_326 | _EVAL_76;
  assign _EVAL_266 = _EVAL_68 & _EVAL_336;
  assign _EVAL_207 = 13'h3f << _EVAL_23;
  assign _EVAL_345 = _EVAL_207[5:0];
  assign _EVAL_162 = ~ _EVAL_345;
  assign _EVAL_366 = _EVAL_162[5:3];
  assign _EVAL_395 = _EVAL_65 ? _EVAL_366 : 3'h0;
  assign _EVAL_82 = _EVAL_395 | _EVAL_193;
  assign _EVAL_383 = _EVAL_140 & _EVAL_13;
  assign _EVAL_360 = ~ _EVAL_341;
  assign _EVAL_332 = _EVAL_360[5:3];
  assign _EVAL_240 = _EVAL_206 ? _EVAL_332 : 3'h0;
  assign _EVAL_286 = _EVAL_194 ? _EVAL_240 : 3'h0;
  assign _EVAL_301 = _EVAL_82 | _EVAL_286;
  assign _EVAL_365 = _EVAL_322 - _EVAL_254;
  assign _EVAL_202 = _EVAL_146 | _EVAL_184;
  assign _EVAL_259 = _EVAL_77 & _EVAL_156;
  assign _EVAL_163 = _EVAL_202 | _EVAL_259;
  assign _EVAL_219 = _EVAL_163 | _EVAL_189;
  assign _EVAL_133 = 3'h5 == _EVAL_17;
  assign _EVAL_119 = TLBroadcastTracker__EVAL_17 == _EVAL_61;
  assign _EVAL_107 = _EVAL_363 & _EVAL_119;
  assign _EVAL_66 = _EVAL_107 & _EVAL_336;
  assign _EVAL_220 = 3'h3 == _EVAL_17;
  assign _EVAL_350 = 3'h4 == _EVAL_17;
  assign _EVAL_90 = 3'h0 == _EVAL_12;
  assign _EVAL_388 = 3'h6 == _EVAL_17;
  assign _EVAL_328 = 3'h7 == _EVAL_17;
  assign _EVAL_285 = _EVAL_318[0];
  assign _EVAL_319 = _EVAL_285 ? 2'h0 : 2'h1;
  assign _EVAL_62 = _EVAL_74 ? _EVAL_319 : 2'h0;
  assign _EVAL_161 = _EVAL_401 ? _EVAL_62 : 2'h0;
  assign _EVAL_358 = _EVAL_250[1];
  assign _EVAL_278 = {_EVAL_231,_EVAL_161,_EVAL_4,_EVAL_212,_EVAL_358,_EVAL_40,_EVAL_7,_EVAL_16};
  assign _EVAL_346 = _EVAL_39 & _EVAL_187;
  assign _EVAL_122 = _EVAL_75 ? _EVAL_118 : _EVAL_197;
  assign _EVAL_92 = _EVAL_148 | _EVAL_378;
  assign _EVAL_289 = _EVAL_81 ? _EVAL_148 : 1'h0;
  assign _EVAL_128 = _EVAL_197 ? _EVAL_378 : 1'h0;
  assign _EVAL_376 = _EVAL_289 | _EVAL_128;
  assign _EVAL_115 = _EVAL_75 ? _EVAL_92 : _EVAL_376;
  assign _EVAL_213 = _EVAL_119 ? TLBroadcastTracker__EVAL_23 : 7'h0;
  assign _EVAL_344 = _EVAL_163 | _EVAL_385;
  assign _EVAL_302 = _EVAL_136 & _EVAL_153;
  assign _EVAL_105 = _EVAL_77 & _EVAL_302;
  assign _EVAL_97 = _EVAL_202 | _EVAL_105;
  assign _EVAL_263 = _EVAL_302 & _EVAL_103;
  assign _EVAL_93 = _EVAL_292 & _EVAL_263;
  assign _EVAL_416 = _EVAL_97 | _EVAL_93;
  assign _EVAL_312 = _EVAL_302 & _EVAL_95;
  assign _EVAL_340 = _EVAL_292 & _EVAL_312;
  assign _EVAL_112 = _EVAL_97 | _EVAL_340;
  assign _EVAL_177 = _EVAL_56 & _EVAL_257;
  assign _EVAL_167 = _EVAL_77 & _EVAL_177;
  assign _EVAL_108 = _EVAL_124 | _EVAL_167;
  assign _EVAL_200 = _EVAL_177 & _EVAL_103;
  assign _EVAL_299 = _EVAL_292 & _EVAL_200;
  assign _EVAL_199 = _EVAL_108 | _EVAL_299;
  assign _EVAL_387 = _EVAL_177 & _EVAL_95;
  assign _EVAL_198 = _EVAL_292 & _EVAL_387;
  assign _EVAL_99 = _EVAL_108 | _EVAL_198;
  assign _EVAL_409 = _EVAL_77 & _EVAL_192;
  assign _EVAL_88 = _EVAL_124 | _EVAL_409;
  assign _EVAL_304 = _EVAL_192 & _EVAL_103;
  assign _EVAL_60 = _EVAL_292 & _EVAL_304;
  assign _EVAL_127 = _EVAL_88 | _EVAL_60;
  assign _EVAL_410 = _EVAL_88 | _EVAL_371;
  assign _EVAL_104 = {_EVAL,1'h0};
  assign _EVAL_316 = {_EVAL_51,_EVAL_344,_EVAL_219,_EVAL_416,_EVAL_112,_EVAL_199,_EVAL_99,_EVAL_127,_EVAL_410,_EVAL_104};
  assign _EVAL_351 = _EVAL_363 & _EVAL_326;
  assign _EVAL_155 = _EVAL_10 & _EVAL_115;
  assign _EVAL_368 = {{2'd0}, _EVAL_155};
  assign _EVAL_186 = _EVAL_75 & _EVAL_10;
  assign _EVAL_391 = _EVAL_139 & _EVAL_22;
  assign _EVAL_334 = _EVAL_135 == 3'h0;
  assign _EVAL_160 = 2'h1 << _EVAL_53;
  assign _EVAL_264 = _EVAL_160[1];
  assign _EVAL_375 = 3'h0 == _EVAL_17;
  assign _EVAL_374 = _EVAL_140 ? _EVAL_65 : _EVAL_276;
  assign _EVAL_190 = _EVAL_417 ? TLBroadcastTracker_1__EVAL_20 : 7'h0;
  assign _EVAL_182 = _EVAL_213 | _EVAL_190;
  assign _EVAL_251 = _EVAL_260 ? _EVAL_46 : _EVAL_182;
  assign _EVAL_347 = {6'h0,_EVAL_23,_EVAL_305,_EVAL_251,_EVAL_316};
  assign _EVAL_157 = _EVAL_374 ? _EVAL_347 : 123'h0;
  assign _EVAL_178 = _EVAL_135 - 3'h1;
  assign _EVAL_181 = _EVAL_310 & _EVAL_391;
  assign _EVAL_55 = 3'h1 == _EVAL_17;
  assign _EVAL_228 = _EVAL_30 == 3'h0;
  assign _EVAL_218 = _EVAL_140 ? _EVAL_183 : _EVAL_272;
  assign _EVAL_100 = _EVAL_140 ? _EVAL_59 : _EVAL_272;
  assign _EVAL_209 = {TLBroadcastTracker__EVAL_13,TLBroadcastTracker__EVAL_8,TLBroadcastTracker__EVAL_25,TLBroadcastTracker__EVAL_2,TLBroadcastTracker__EVAL_19,TLBroadcastTracker__EVAL,TLBroadcastTracker__EVAL_11,1'h0};
  assign _EVAL_98 = _EVAL_100 ? _EVAL_209 : 123'h0;
  assign _EVAL_245 = _EVAL_157 | _EVAL_98;
  assign _EVAL_394 = _EVAL_358 & _EVAL_293;
  assign _EVAL_142 = _EVAL_394 & _EVAL_280;
  assign _EVAL_297 = _EVAL_245 | _EVAL_64;
  assign _EVAL_405 = _EVAL_122 ? _EVAL_278 : 82'h0;
  assign _EVAL_355 = _EVAL_140 ? _EVAL_172 : _EVAL_337;
  assign _EVAL_324 = _EVAL_267 - _EVAL_368;
  assign _EVAL_230 = _EVAL_39 & _EVAL_399;
  assign _EVAL_225 = _EVAL_335 | _EVAL_405;
  assign _EVAL_270 = _EVAL_228 | _EVAL_85;
  assign _EVAL_256 = _EVAL_160[0];
  assign _EVAL_372 = _EVAL_358 & _EVAL_391;
  assign _EVAL_15 = _EVAL_297[116:114];
  assign _EVAL_27 = _EVAL_225[64:1];
  assign _EVAL_6 = _EVAL_225[81:79];
  assign _EVAL_36 = _EVAL_297[72:65];
  assign TLBroadcastTracker_1__EVAL_11 = _EVAL_37;
  assign _EVAL_25 = _EVAL_225[65];
  assign _EVAL_9 = _EVAL_297[113:105];
  assign _EVAL_44 = _EVAL_384;
  assign TLBroadcastTracker_1__EVAL_15 = _EVAL_8;
  assign _EVAL_5 = _EVAL_101;
  assign TLBroadcastTracker__EVAL_4 = _EVAL_158 == 3'h0;
  assign _EVAL_43 = _EVAL_174 | _EVAL_412;
  assign _EVAL_45 = _EVAL_140 ? _EVAL_78 : _EVAL_277;
  assign TLBroadcastTracker__EVAL_15 = _EVAL_37;
  assign TLBroadcastTracker__EVAL_27 = _EVAL_21;
  assign _EVAL_42 = _EVAL_326 | _EVAL_91;
  assign _EVAL_26 = _EVAL_225[78:77];
  assign TLBroadcastTracker_1__EVAL_12 = _EVAL_19;
  assign _EVAL_35 = _EVAL_225[76:74];
  assign _EVAL_29 = _EVAL_225[66];
  assign TLBroadcastTracker__EVAL_12 = _EVAL_256 & _EVAL_0;
  assign TLBroadcastTracker__EVAL_28 = _EVAL_66 & _EVAL_270;
  assign TLBroadcastTracker_1__EVAL_26 = _EVAL_33;
  assign TLBroadcastTracker_1__EVAL_13 = _EVAL_351 & _EVAL_417;
  assign TLBroadcastTracker_1__EVAL_22 = _EVAL_13 & _EVAL_355;
  assign TLBroadcastTracker_1__EVAL_1 = _EVAL_261 ? 1'h0 : 1'h1;
  assign TLBroadcastTracker__EVAL_18 = _EVAL_17;
  assign _EVAL_2 = _EVAL_225[73:67];
  assign _EVAL_41 = _EVAL_225[0];
  assign _EVAL_50 = _EVAL_297[64:1];
  assign _EVAL_14 = _EVAL_297[122:120];
  assign TLBroadcastTracker_1__EVAL_16 = _EVAL_17;
  assign TLBroadcastTracker__EVAL_7 = _EVAL_346 & _EVAL_294;
  assign TLBroadcastTracker_1__EVAL_5 = _EVAL_142 & _EVAL_311;
  assign _EVAL_34 = _EVAL_75 ? _EVAL_92 : _EVAL_376;
  assign TLBroadcastTracker_1__EVAL_9 = _EVAL_28;
  assign _EVAL_18 = _EVAL_297[0];
  assign TLBroadcastTracker_1__EVAL_2 = _EVAL_266 & _EVAL_270;
  assign TLBroadcastTracker__EVAL_0 = _EVAL_13 & _EVAL_218;
  assign TLBroadcastTracker__EVAL_9 = _EVAL_141 & _EVAL_311;
  assign TLBroadcastTracker_1__EVAL_10 = _EVAL_12;
  assign TLBroadcastTracker_1__EVAL_3 = _EVAL_158 == 3'h0;
  assign TLBroadcastTracker__EVAL_6 = _EVAL_8;
  assign TLBroadcastTracker_1__EVAL_0 = _EVAL_264 & _EVAL_0;
  assign TLBroadcastTracker__EVAL_14 = _EVAL_261 ? 1'h0 : 1'h1;
  assign _EVAL_31 = {_EVAL_69, 6'h0};
  assign _EVAL_1 = _EVAL_297[104:73];
  assign TLBroadcastTracker__EVAL_16 = _EVAL_28;
  assign TLBroadcastTracker__EVAL_1 = _EVAL_181 & _EVAL_412;
  assign TLBroadcastTracker__EVAL_21 = _EVAL_49;
  assign TLBroadcastTracker_1__EVAL_23 = _EVAL_230 & _EVAL_294;
  assign TLBroadcastTracker__EVAL_5 = _EVAL_19;
  assign _EVAL_38 = _EVAL_294 & _EVAL_402;
  assign TLBroadcastTracker_1__EVAL_4 = _EVAL_21;
  assign TLBroadcastTracker__EVAL_24 = _EVAL_351 & _EVAL_119;
  assign TLBroadcastTracker_1__EVAL = _EVAL_372 & _EVAL_412;
  assign _EVAL_48 = _EVAL_297[119:117];
  assign TLBroadcastTracker__EVAL_10 = _EVAL_12;
  assign TLBroadcastTracker__EVAL_26 = _EVAL_33;
  assign TLBroadcastTracker_1__EVAL_7 = _EVAL_49;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_69 = _RAND_0[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_81 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_101 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_135 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_158 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_197 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_267 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_272 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_276 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_322 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_337 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_384 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_33) begin
    if (_EVAL_152) begin
      _EVAL_69 <= _EVAL_379;
    end
    if (_EVAL_19) begin
      _EVAL_81 <= 1'h0;
    end else begin
      if (_EVAL_75) begin
        _EVAL_81 <= _EVAL_373;
      end
    end
    if (_EVAL_19) begin
      _EVAL_101 <= 1'h0;
    end else begin
      _EVAL_101 <= _EVAL_216[0];
    end
    if (_EVAL_19) begin
      _EVAL_135 <= 3'h0;
    end else begin
      if (_EVAL_293) begin
        if (_EVAL_334) begin
          if (_EVAL_315) begin
            _EVAL_135 <= _EVAL_195;
          end else begin
            _EVAL_135 <= 3'h0;
          end
        end else begin
          _EVAL_135 <= _EVAL_178;
        end
      end
    end
    if (_EVAL_19) begin
      _EVAL_158 <= 3'h0;
    end else begin
      if (_EVAL_87) begin
        if (_EVAL_361) begin
          if (_EVAL_357) begin
            _EVAL_158 <= _EVAL_223;
          end else begin
            _EVAL_158 <= 3'h0;
          end
        end else begin
          _EVAL_158 <= _EVAL_67;
        end
      end
    end
    if (_EVAL_19) begin
      _EVAL_197 <= 1'h0;
    end else begin
      if (_EVAL_75) begin
        _EVAL_197 <= _EVAL_118;
      end
    end
    if (_EVAL_19) begin
      _EVAL_267 <= 3'h0;
    end else begin
      if (_EVAL_186) begin
        if (_EVAL_118) begin
          if (_EVAL_315) begin
            _EVAL_267 <= _EVAL_195;
          end else begin
            _EVAL_267 <= 3'h0;
          end
        end else begin
          _EVAL_267 <= 3'h0;
        end
      end else begin
        _EVAL_267 <= _EVAL_324;
      end
    end
    if (_EVAL_19) begin
      _EVAL_272 <= 1'h0;
    end else begin
      if (_EVAL_140) begin
        _EVAL_272 <= _EVAL_59;
      end
    end
    if (_EVAL_19) begin
      _EVAL_276 <= 1'h0;
    end else begin
      if (_EVAL_140) begin
        _EVAL_276 <= _EVAL_65;
      end
    end
    if (_EVAL_19) begin
      _EVAL_322 <= 3'h0;
    end else begin
      if (_EVAL_383) begin
        _EVAL_322 <= _EVAL_301;
      end else begin
        _EVAL_322 <= _EVAL_365;
      end
    end
    if (_EVAL_19) begin
      _EVAL_337 <= 1'h0;
    end else begin
      if (_EVAL_140) begin
        _EVAL_337 <= _EVAL_194;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_375) begin
        _EVAL_384 <= 2'h2;
      end else begin
        if (_EVAL_55) begin
          _EVAL_384 <= 2'h2;
        end else begin
          if (_EVAL_57) begin
            _EVAL_384 <= 2'h2;
          end else begin
            if (_EVAL_220) begin
              _EVAL_384 <= 2'h2;
            end else begin
              if (_EVAL_350) begin
                _EVAL_384 <= 2'h1;
              end else begin
                if (_EVAL_133) begin
                  if (_EVAL_90) begin
                    _EVAL_384 <= 2'h1;
                  end else begin
                    if (_EVAL_171) begin
                      _EVAL_384 <= 2'h2;
                    end else begin
                      _EVAL_384 <= 2'h0;
                    end
                  end
                end else begin
                  if (_EVAL_388) begin
                    if (_EVAL_90) begin
                      _EVAL_384 <= 2'h1;
                    end else begin
                      if (_EVAL_171) begin
                        _EVAL_384 <= 2'h2;
                      end else begin
                        if (_EVAL_72) begin
                          _EVAL_384 <= 2'h2;
                        end else begin
                          _EVAL_384 <= 2'h0;
                        end
                      end
                    end
                  end else begin
                    if (_EVAL_328) begin
                      if (_EVAL_90) begin
                        _EVAL_384 <= 2'h1;
                      end else begin
                        if (_EVAL_171) begin
                          _EVAL_384 <= 2'h2;
                        end else begin
                          if (_EVAL_72) begin
                            _EVAL_384 <= 2'h2;
                          end else begin
                            _EVAL_384 <= 2'h0;
                          end
                        end
                      end
                    end else begin
                      _EVAL_384 <= 2'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
