//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_36_assert(
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_7,
  input  [6:0]  _EVAL_8,
  input  [7:0]  _EVAL_9,
  input  [6:0]  _EVAL_10,
  input  [30:0] _EVAL_13,
  input         _EVAL_16,
  input         _EVAL_18,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  input  [2:0]  _EVAL_32,
  input  [2:0]  _EVAL_34,
  input         _EVAL_45,
  input         _EVAL_80,
  input         Repeater__EVAL_6
);
  wire  TLMonitor__EVAL;
  wire [2:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire [2:0] TLMonitor__EVAL_4;
  wire [7:0] TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire [30:0] TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire  TLMonitor__EVAL_12;
  wire [6:0] TLMonitor__EVAL_13;
  wire [2:0] TLMonitor__EVAL_14;
  wire [6:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  SiFive__EVAL_34_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16)
  );
  assign TLMonitor__EVAL_4 = _EVAL_32;
  assign TLMonitor__EVAL_5 = _EVAL_9;
  assign TLMonitor__EVAL_10 = _EVAL_18;
  assign TLMonitor__EVAL_16 = _EVAL_0 | _EVAL_45;
  assign TLMonitor__EVAL_7 = _EVAL_2 & _EVAL_80;
  assign TLMonitor__EVAL_3 = _EVAL_25;
  assign TLMonitor__EVAL_9 = _EVAL_13;
  assign TLMonitor__EVAL_15 = _EVAL_8;
  assign TLMonitor__EVAL_1 = _EVAL_16;
  assign TLMonitor__EVAL_8 = _EVAL_7;
  assign TLMonitor__EVAL_2 = _EVAL_1;
  assign TLMonitor__EVAL_13 = _EVAL_10;
  assign TLMonitor__EVAL_6 = _EVAL_26;
  assign TLMonitor__EVAL_12 = _EVAL_27;
  assign TLMonitor__EVAL_11 = _EVAL_34;
  assign TLMonitor__EVAL = Repeater__EVAL_6;
  assign TLMonitor__EVAL_0 = _EVAL_29;
  assign TLMonitor__EVAL_14 = _EVAL_28;

endmodule
