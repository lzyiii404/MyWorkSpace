//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_181_assert(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [27:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [11:0] _EVAL_13,
  input  [11:0] _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2335:0] _EVAL_33;
  reg [2335:0] _RAND_0;
  reg  _EVAL_51;
  reg [31:0] _RAND_1;
  reg [11:0] _EVAL_64;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_79;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_127;
  reg [31:0] _RAND_4;
  reg [27:0] _EVAL_138;
  reg [31:0] _RAND_5;
  reg [31:0] _EVAL_143;
  reg [31:0] _RAND_6;
  reg  _EVAL_145;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_166;
  reg [31:0] _RAND_8;
  reg [1:0] _EVAL_171;
  reg [31:0] _RAND_9;
  reg [11:0] _EVAL_177;
  reg [31:0] _RAND_10;
  reg  _EVAL_200;
  reg [31:0] _RAND_11;
  reg  _EVAL_215;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_235;
  reg [31:0] _RAND_13;
  wire  _EVAL_112;
  wire  _EVAL_44;
  wire  _EVAL_18;
  wire  _EVAL_163;
  wire  _EVAL_39;
  wire  _EVAL_80;
  wire  _EVAL_181;
  wire  _EVAL_37;
  wire  _EVAL_147;
  wire [4095:0] _EVAL_161;
  wire [4095:0] _EVAL_175;
  wire [2335:0] _EVAL_35;
  wire  _EVAL_155;
  wire  _EVAL_128;
  wire  _EVAL_136;
  wire  _EVAL_69;
  wire  _EVAL_186;
  wire  _EVAL_211;
  wire [4095:0] _EVAL_150;
  wire [4095:0] _EVAL_108;
  wire [2335:0] _EVAL_220;
  wire  _EVAL_205;
  wire  _EVAL_125;
  wire  _EVAL_99;
  wire  _EVAL_121;
  wire  _EVAL_47;
  wire  _EVAL_105;
  wire  _EVAL_78;
  wire  _EVAL_137;
  wire  _EVAL_231;
  wire  _EVAL_89;
  wire  _EVAL_229;
  wire  _EVAL_16;
  wire  _EVAL_90;
  wire  _EVAL_189;
  wire [4:0] _EVAL_216;
  wire  _EVAL_29;
  wire  _EVAL_170;
  wire [1:0] _EVAL_173;
  wire [1:0] _EVAL_180;
  wire  _EVAL_106;
  wire  _EVAL_116;
  wire  _EVAL_144;
  wire  _EVAL_135;
  wire  _EVAL_72;
  wire  _EVAL_146;
  wire  _EVAL_42;
  wire  _EVAL_76;
  wire  _EVAL_139;
  wire  _EVAL_226;
  wire  _EVAL_195;
  wire  _EVAL_178;
  wire  _EVAL_208;
  wire  _EVAL_201;
  wire [2335:0] _EVAL_191;
  wire [2335:0] _EVAL_36;
  wire  _EVAL_65;
  wire  _EVAL_55;
  wire  _EVAL_228;
  wire [1:0] _EVAL_190;
  wire [1:0] _EVAL_27;
  wire [27:0] _EVAL_221;
  wire [28:0] _EVAL_57;
  wire [28:0] _EVAL_50;
  wire [28:0] _EVAL_101;
  wire  _EVAL_210;
  wire  _EVAL_169;
  wire  _EVAL_62;
  wire  _EVAL_162;
  wire  _EVAL_87;
  wire  _EVAL_193;
  wire  _EVAL_113;
  wire  _EVAL_56;
  wire  _EVAL_202;
  wire  _EVAL_151;
  wire  _EVAL_213;
  wire  _EVAL_95;
  wire  _EVAL_46;
  wire  _EVAL_179;
  wire  _EVAL_227;
  wire  _EVAL_88;
  wire  _EVAL_98;
  wire  _EVAL_49;
  wire  _EVAL_74;
  wire  _EVAL_126;
  wire [2335:0] _EVAL_168;
  wire  _EVAL_96;
  wire  _EVAL_70;
  wire  _EVAL_160;
  wire  _EVAL_114;
  wire  _EVAL_140;
  wire  _EVAL_153;
  wire  _EVAL_148;
  wire  _EVAL_223;
  wire  _EVAL_104;
  wire  _EVAL_154;
  wire  _EVAL_100;
  wire  _EVAL_52;
  wire  _EVAL_34;
  wire  _EVAL_230;
  wire [27:0] _EVAL_182;
  wire [27:0] _EVAL_59;
  wire  _EVAL_86;
  wire  _EVAL_183;
  wire  _EVAL_73;
  wire  _EVAL_85;
  wire  _EVAL_54;
  wire  _EVAL_233;
  wire  _EVAL_167;
  wire  _EVAL_26;
  wire  _EVAL_156;
  wire  _EVAL_184;
  wire  _EVAL_129;
  wire  _EVAL_30;
  wire  _EVAL_24;
  wire  _EVAL_31;
  wire  _EVAL_60;
  wire  _EVAL_48;
  wire  _EVAL_84;
  wire  _EVAL_25;
  wire  _EVAL_174;
  wire  _EVAL_40;
  wire  _EVAL_23;
  wire  _EVAL_124;
  wire [3:0] _EVAL_238;
  wire  _EVAL_117;
  wire  _EVAL_157;
  wire [3:0] _EVAL_225;
  wire  _EVAL_93;
  wire  _EVAL_159;
  wire  _EVAL_199;
  wire  _EVAL_17;
  wire  _EVAL_91;
  wire [2335:0] _EVAL_134;
  wire  _EVAL_152;
  wire  _EVAL_217;
  wire  _EVAL_103;
  wire  _EVAL_236;
  wire  _EVAL_119;
  wire  _EVAL_58;
  wire  _EVAL_110;
  wire  _EVAL_75;
  wire  _EVAL_71;
  wire  _EVAL_123;
  wire  _EVAL_218;
  wire  _EVAL_53;
  wire [3:0] _EVAL_15;
  wire [3:0] _EVAL_224;
  wire  _EVAL_219;
  wire  _EVAL_63;
  wire  _EVAL_83;
  wire  _EVAL_118;
  wire  _EVAL_207;
  wire  _EVAL_77;
  wire  _EVAL_131;
  wire  _EVAL_43;
  wire  _EVAL_67;
  wire  _EVAL_102;
  wire  _EVAL_41;
  wire  _EVAL_149;
  wire  _EVAL_198;
  wire  _EVAL_192;
  wire  _EVAL_21;
  wire  _EVAL_212;
  wire  _EVAL_158;
  wire [31:0] _EVAL_222;
  wire  _EVAL_32;
  wire  _EVAL_107;
  wire  _EVAL_66;
  wire  _EVAL_92;
  wire  _EVAL_197;
  wire  _EVAL_172;
  wire  _EVAL_141;
  wire  _EVAL_22;
  wire  _EVAL_68;
  wire  _EVAL_185;
  wire  _EVAL_203;
  wire  _EVAL_122;
  wire  _EVAL_204;
  wire  _EVAL_188;
  wire  _EVAL_232;
  wire  _EVAL_115;
  wire  _EVAL_164;
  wire  _EVAL_19;
  wire [2335:0] _EVAL_38;
  wire  _EVAL_61;
  wire  _EVAL_234;
  wire  _EVAL_111;
  wire  _EVAL_130;
  wire  _EVAL_133;
  wire  _EVAL_20;
  wire  _EVAL_97;
  wire  _EVAL_109;
  wire [2335:0] _EVAL_132;
  wire  _EVAL_176;
  wire  _EVAL_187;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_112 = _EVAL_200 == 1'h0;
  assign _EVAL_44 = _EVAL_200 - 1'h1;
  assign _EVAL_18 = _EVAL_0 == 3'h5;
  assign _EVAL_163 = _EVAL_7 & _EVAL_18;
  assign _EVAL_39 = _EVAL_6 == _EVAL_127;
  assign _EVAL_80 = _EVAL_39 | _EVAL_3;
  assign _EVAL_181 = _EVAL_11 & _EVAL_7;
  assign _EVAL_37 = _EVAL_51 == 1'h0;
  assign _EVAL_147 = _EVAL_181 & _EVAL_37;
  assign _EVAL_161 = 4096'h1 << _EVAL_13;
  assign _EVAL_175 = _EVAL_147 ? _EVAL_161 : 4096'h0;
  assign _EVAL_35 = _EVAL_175[2335:0];
  assign _EVAL_155 = _EVAL_5 & _EVAL_9;
  assign _EVAL_128 = _EVAL_215 == 1'h0;
  assign _EVAL_136 = _EVAL_155 & _EVAL_128;
  assign _EVAL_69 = _EVAL_6 == 3'h6;
  assign _EVAL_186 = _EVAL_69 == 1'h0;
  assign _EVAL_211 = _EVAL_136 & _EVAL_186;
  assign _EVAL_150 = 4096'h1 << _EVAL_14;
  assign _EVAL_108 = _EVAL_211 ? _EVAL_150 : 4096'h0;
  assign _EVAL_220 = _EVAL_108[2335:0];
  assign _EVAL_205 = _EVAL_35 != _EVAL_220;
  assign _EVAL_125 = _EVAL_35 != 2336'h0;
  assign _EVAL_99 = _EVAL_125 == 1'h0;
  assign _EVAL_121 = _EVAL_205 | _EVAL_99;
  assign _EVAL_47 = _EVAL_121 | _EVAL_3;
  assign _EVAL_105 = _EVAL_47 == 1'h0;
  assign _EVAL_78 = _EVAL_13 == _EVAL_177;
  assign _EVAL_137 = _EVAL != 3'h0;
  assign _EVAL_231 = _EVAL_137 | _EVAL_3;
  assign _EVAL_89 = _EVAL_231 == 1'h0;
  assign _EVAL_229 = _EVAL_9 & _EVAL_69;
  assign _EVAL_16 = _EVAL_51 - 1'h1;
  assign _EVAL_90 = _EVAL_6 == 3'h4;
  assign _EVAL_189 = _EVAL_9 & _EVAL_90;
  assign _EVAL_216 = 5'h3 << _EVAL_8;
  assign _EVAL_29 = _EVAL_8 >= 2'h2;
  assign _EVAL_170 = _EVAL_8[0];
  assign _EVAL_173 = 2'h1 << _EVAL_170;
  assign _EVAL_180 = _EVAL_173 | 2'h1;
  assign _EVAL_106 = _EVAL_180[1];
  assign _EVAL_116 = _EVAL_2[1];
  assign _EVAL_144 = _EVAL_116 == 1'h0;
  assign _EVAL_135 = _EVAL_106 & _EVAL_144;
  assign _EVAL_72 = _EVAL_29 | _EVAL_135;
  assign _EVAL_146 = _EVAL_180[0];
  assign _EVAL_42 = _EVAL_2[0];
  assign _EVAL_76 = _EVAL_42 == 1'h0;
  assign _EVAL_139 = _EVAL_144 & _EVAL_76;
  assign _EVAL_226 = _EVAL_146 & _EVAL_139;
  assign _EVAL_195 = _EVAL_72 | _EVAL_226;
  assign _EVAL_178 = _EVAL_0 == 3'h1;
  assign _EVAL_208 = _EVAL_7 & _EVAL_178;
  assign _EVAL_201 = plusarg_reader_out == 32'h0;
  assign _EVAL_191 = _EVAL_35 | _EVAL_33;
  assign _EVAL_36 = _EVAL_191 >> _EVAL_14;
  assign _EVAL_65 = _EVAL_36[0];
  assign _EVAL_55 = _EVAL_65 | _EVAL_3;
  assign _EVAL_228 = _EVAL_55 == 1'h0;
  assign _EVAL_190 = _EVAL_216[1:0];
  assign _EVAL_27 = ~ _EVAL_190;
  assign _EVAL_221 = _EVAL_2 ^ 28'hc000000;
  assign _EVAL_57 = {1'b0,$signed(_EVAL_221)};
  assign _EVAL_50 = $signed(_EVAL_57) & $signed(-29'sh4000000);
  assign _EVAL_101 = $signed(_EVAL_50);
  assign _EVAL_210 = _EVAL_2 == _EVAL_138;
  assign _EVAL_169 = _EVAL_210 | _EVAL_3;
  assign _EVAL_62 = _EVAL_169 == 1'h0;
  assign _EVAL_162 = _EVAL_8 <= 2'h2;
  assign _EVAL_87 = $signed(_EVAL_101) == $signed(29'sh0);
  assign _EVAL_193 = _EVAL_162 & _EVAL_87;
  assign _EVAL_113 = _EVAL <= 3'h3;
  assign _EVAL_56 = _EVAL_113 | _EVAL_3;
  assign _EVAL_202 = _EVAL_56 == 1'h0;
  assign _EVAL_151 = _EVAL_1 == 1'h0;
  assign _EVAL_213 = _EVAL_33 != 2336'h0;
  assign _EVAL_95 = _EVAL_213 == 1'h0;
  assign _EVAL_46 = _EVAL_95 | _EVAL_201;
  assign _EVAL_179 = _EVAL_143 < plusarg_reader_out;
  assign _EVAL_227 = _EVAL_46 | _EVAL_179;
  assign _EVAL_88 = _EVAL_227 | _EVAL_3;
  assign _EVAL_98 = _EVAL_88 == 1'h0;
  assign _EVAL_49 = _EVAL_0 == 3'h3;
  assign _EVAL_74 = _EVAL == _EVAL_166;
  assign _EVAL_126 = _EVAL_151 | _EVAL_3;
  assign _EVAL_168 = ~ _EVAL_220;
  assign _EVAL_96 = _EVAL == 3'h0;
  assign _EVAL_70 = _EVAL_96 | _EVAL_3;
  assign _EVAL_160 = _EVAL_116 & _EVAL_42;
  assign _EVAL_114 = _EVAL_145 == 1'h0;
  assign _EVAL_140 = _EVAL_145 - 1'h1;
  assign _EVAL_153 = _EVAL_0 == 3'h6;
  assign _EVAL_148 = _EVAL_112 == 1'h0;
  assign _EVAL_223 = _EVAL_9 & _EVAL_148;
  assign _EVAL_104 = _EVAL_0 == 3'h2;
  assign _EVAL_154 = _EVAL_14 <= 12'h91f;
  assign _EVAL_100 = _EVAL_154 | _EVAL_3;
  assign _EVAL_52 = _EVAL_100 == 1'h0;
  assign _EVAL_34 = _EVAL <= 3'h2;
  assign _EVAL_230 = _EVAL_34 | _EVAL_3;
  assign _EVAL_182 = {{26'd0}, _EVAL_27};
  assign _EVAL_59 = _EVAL_2 & _EVAL_182;
  assign _EVAL_86 = _EVAL_59 == 28'h0;
  assign _EVAL_183 = _EVAL_86 | _EVAL_3;
  assign _EVAL_73 = _EVAL_6 == 3'h2;
  assign _EVAL_85 = _EVAL_181 | _EVAL_155;
  assign _EVAL_54 = _EVAL_106 & _EVAL_116;
  assign _EVAL_233 = _EVAL_29 | _EVAL_54;
  assign _EVAL_167 = _EVAL_146 & _EVAL_160;
  assign _EVAL_26 = _EVAL_233 | _EVAL_167;
  assign _EVAL_156 = _EVAL_13 <= 12'h91f;
  assign _EVAL_184 = _EVAL_126 == 1'h0;
  assign _EVAL_129 = _EVAL <= 3'h4;
  assign _EVAL_30 = _EVAL_129 | _EVAL_3;
  assign _EVAL_24 = _EVAL_30 == 1'h0;
  assign _EVAL_31 = _EVAL_144 & _EVAL_42;
  assign _EVAL_60 = _EVAL_6 <= 3'h6;
  assign _EVAL_48 = _EVAL_60 | _EVAL_3;
  assign _EVAL_84 = _EVAL_48 == 1'h0;
  assign _EVAL_25 = _EVAL_116 & _EVAL_76;
  assign _EVAL_174 = _EVAL_146 & _EVAL_25;
  assign _EVAL_40 = _EVAL_233 | _EVAL_174;
  assign _EVAL_23 = _EVAL_146 & _EVAL_31;
  assign _EVAL_124 = _EVAL_72 | _EVAL_23;
  assign _EVAL_238 = {_EVAL_26,_EVAL_40,_EVAL_124,_EVAL_195};
  assign _EVAL_117 = _EVAL_12 == _EVAL_238;
  assign _EVAL_157 = _EVAL_117 | _EVAL_3;
  assign _EVAL_225 = ~ _EVAL_12;
  assign _EVAL_93 = _EVAL_225 == 4'h0;
  assign _EVAL_159 = _EVAL_93 | _EVAL_3;
  assign _EVAL_199 = _EVAL_159 == 1'h0;
  assign _EVAL_17 = _EVAL_0 == _EVAL_79;
  assign _EVAL_91 = _EVAL_17 | _EVAL_3;
  assign _EVAL_134 = _EVAL_33 >> _EVAL_13;
  assign _EVAL_152 = _EVAL_134[0];
  assign _EVAL_217 = _EVAL_152 == 1'h0;
  assign _EVAL_103 = _EVAL_217 | _EVAL_3;
  assign _EVAL_236 = _EVAL_10 >= 2'h2;
  assign _EVAL_119 = _EVAL_236 | _EVAL_3;
  assign _EVAL_58 = _EVAL_10 == _EVAL_235;
  assign _EVAL_110 = _EVAL_74 | _EVAL_3;
  assign _EVAL_75 = _EVAL_110 == 1'h0;
  assign _EVAL_71 = _EVAL_114 == 1'h0;
  assign _EVAL_123 = _EVAL_9 & _EVAL_73;
  assign _EVAL_218 = _EVAL_215 - 1'h1;
  assign _EVAL_53 = _EVAL_0 == 3'h4;
  assign _EVAL_15 = ~ _EVAL_238;
  assign _EVAL_224 = _EVAL_12 & _EVAL_15;
  assign _EVAL_219 = _EVAL_224 == 4'h0;
  assign _EVAL_63 = _EVAL_219 | _EVAL_3;
  assign _EVAL_83 = _EVAL_6 == 3'h0;
  assign _EVAL_118 = _EVAL_91 == 1'h0;
  assign _EVAL_207 = _EVAL_7 & _EVAL_53;
  assign _EVAL_77 = _EVAL_58 | _EVAL_3;
  assign _EVAL_131 = _EVAL_77 == 1'h0;
  assign _EVAL_43 = _EVAL_8 == _EVAL_171;
  assign _EVAL_67 = _EVAL_43 | _EVAL_3;
  assign _EVAL_102 = _EVAL_6 == 3'h5;
  assign _EVAL_41 = _EVAL_14 == _EVAL_64;
  assign _EVAL_149 = _EVAL_41 | _EVAL_3;
  assign _EVAL_198 = _EVAL_149 == 1'h0;
  assign _EVAL_192 = _EVAL_3 == 1'h0;
  assign _EVAL_21 = _EVAL_7 & _EVAL_153;
  assign _EVAL_212 = _EVAL_155 & _EVAL_112;
  assign _EVAL_158 = _EVAL_80 == 1'h0;
  assign _EVAL_222 = _EVAL_143 + 32'h1;
  assign _EVAL_32 = _EVAL_67 == 1'h0;
  assign _EVAL_107 = _EVAL_181 & _EVAL_114;
  assign _EVAL_66 = _EVAL_0 == 3'h7;
  assign _EVAL_92 = _EVAL_0 == 3'h0;
  assign _EVAL_197 = _EVAL_78 | _EVAL_3;
  assign _EVAL_172 = _EVAL_197 == 1'h0;
  assign _EVAL_141 = _EVAL_70 == 1'h0;
  assign _EVAL_22 = _EVAL_9 & _EVAL_102;
  assign _EVAL_68 = _EVAL_119 == 1'h0;
  assign _EVAL_185 = _EVAL_6 == 3'h1;
  assign _EVAL_203 = _EVAL_9 & _EVAL_185;
  assign _EVAL_122 = _EVAL_157 == 1'h0;
  assign _EVAL_204 = _EVAL_63 == 1'h0;
  assign _EVAL_188 = _EVAL_9 & _EVAL_83;
  assign _EVAL_232 = _EVAL_156 | _EVAL_3;
  assign _EVAL_115 = _EVAL_29 | _EVAL_3;
  assign _EVAL_164 = _EVAL_115 == 1'h0;
  assign _EVAL_19 = _EVAL_183 == 1'h0;
  assign _EVAL_38 = _EVAL_33 | _EVAL_35;
  assign _EVAL_61 = _EVAL_7 & _EVAL_49;
  assign _EVAL_234 = _EVAL_7 & _EVAL_66;
  assign _EVAL_111 = _EVAL_7 & _EVAL_104;
  assign _EVAL_130 = _EVAL_230 == 1'h0;
  assign _EVAL_133 = _EVAL_193 | _EVAL_3;
  assign _EVAL_20 = _EVAL_133 == 1'h0;
  assign _EVAL_97 = _EVAL_103 == 1'h0;
  assign _EVAL_109 = _EVAL_232 == 1'h0;
  assign _EVAL_132 = _EVAL_38 & _EVAL_168;
  assign _EVAL_176 = _EVAL_7 & _EVAL_71;
  assign _EVAL_187 = _EVAL_7 & _EVAL_92;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {73{`RANDOM}};
  _EVAL_33 = _RAND_0[2335:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_51 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_79 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_127 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_138 = _RAND_5[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_143 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_145 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_166 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_171 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_177 = _RAND_10[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_200 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_215 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_235 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_3) begin
      _EVAL_33 <= 2336'h0;
    end else begin
      _EVAL_33 <= _EVAL_132;
    end
    if (_EVAL_3) begin
      _EVAL_51 <= 1'h0;
    end else begin
      if (_EVAL_181) begin
        if (_EVAL_37) begin
          _EVAL_51 <= 1'h0;
        end else begin
          _EVAL_51 <= _EVAL_16;
        end
      end
    end
    if (_EVAL_212) begin
      _EVAL_64 <= _EVAL_14;
    end
    if (_EVAL_107) begin
      _EVAL_79 <= _EVAL_0;
    end
    if (_EVAL_212) begin
      _EVAL_127 <= _EVAL_6;
    end
    if (_EVAL_107) begin
      _EVAL_138 <= _EVAL_2;
    end
    if (_EVAL_3) begin
      _EVAL_143 <= 32'h0;
    end else begin
      if (_EVAL_85) begin
        _EVAL_143 <= 32'h0;
      end else begin
        _EVAL_143 <= _EVAL_222;
      end
    end
    if (_EVAL_3) begin
      _EVAL_145 <= 1'h0;
    end else begin
      if (_EVAL_181) begin
        if (_EVAL_114) begin
          _EVAL_145 <= 1'h0;
        end else begin
          _EVAL_145 <= _EVAL_140;
        end
      end
    end
    if (_EVAL_107) begin
      _EVAL_166 <= _EVAL;
    end
    if (_EVAL_107) begin
      _EVAL_171 <= _EVAL_8;
    end
    if (_EVAL_107) begin
      _EVAL_177 <= _EVAL_13;
    end
    if (_EVAL_3) begin
      _EVAL_200 <= 1'h0;
    end else begin
      if (_EVAL_155) begin
        if (_EVAL_112) begin
          _EVAL_200 <= 1'h0;
        end else begin
          _EVAL_200 <= _EVAL_44;
        end
      end
    end
    if (_EVAL_3) begin
      _EVAL_215 <= 1'h0;
    end else begin
      if (_EVAL_155) begin
        if (_EVAL_128) begin
          _EVAL_215 <= 1'h0;
        end else begin
          _EVAL_215 <= _EVAL_218;
        end
      end
    end
    if (_EVAL_212) begin
      _EVAL_235 <= _EVAL_10;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adb9543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41af69c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97ce01ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24c0342e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5428059c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c7ebd80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aa4f0cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf6b1da4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30e8d4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72c2439c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfea87eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a3fe56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d85715b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35d7dda2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f507a900)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76a23f77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a907b8cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(871ff20f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(518932e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac84c543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf33a86c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a96f94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfc9e3d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42dbdc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6eff4b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6e467e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b77c82a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(669c9ff8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb56a9a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9b55191)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8fd4096)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a580767f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ad753ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90af529c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(532b2800)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6243b8b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de5157e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(626f625d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7bf0c2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0b536ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1088ab9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aa7c129)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9af1f6c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c415586)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bfa26cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1febaaad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531cca50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa23acb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fdd68f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(420b21da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afadcc49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed32d2ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(202c6f5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c1284a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a951f6f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c923bd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cea28ba8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f366654)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33031838)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa205140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e5ed9a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72820793)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39e85a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(209714a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(172c12d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c43ab094)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d934160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a4f762d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14088283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d02f7301)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8356124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f274c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
