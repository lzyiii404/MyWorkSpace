//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_180(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  output [1:0]  _EVAL_2,
  output [2:0]  _EVAL_3,
  output [3:0]  _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  output [27:0] _EVAL_9,
  output [1:0]  _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  output [1:0]  _EVAL_14,
  input  [31:0] _EVAL_15,
  output [6:0]  _EVAL_16,
  output [31:0] _EVAL_17,
  output [29:0] _EVAL_18,
  output [31:0] _EVAL_19,
  input  [2:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  output        _EVAL_22,
  input  [29:0] _EVAL_23,
  output [1:0]  _EVAL_24,
  input         _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [1:0]  _EVAL_27,
  output [6:0]  _EVAL_28,
  input  [6:0]  _EVAL_29,
  input         _EVAL_30,
  input  [2:0]  _EVAL_31,
  output [3:0]  _EVAL_32,
  input  [1:0]  _EVAL_33,
  output [3:0]  _EVAL_34,
  output [2:0]  _EVAL_35,
  output        _EVAL_36,
  output [3:0]  _EVAL_37,
  output        _EVAL_38,
  output [1:0]  _EVAL_39,
  output [2:0]  _EVAL_40,
  input  [1:0]  _EVAL_41,
  input  [31:0] _EVAL_42,
  output        _EVAL_43,
  input         _EVAL_44,
  input  [2:0]  _EVAL_45,
  output [31:0] _EVAL_46,
  output [7:0]  _EVAL_47,
  output        _EVAL_48,
  output [31:0] _EVAL_49,
  input  [2:0]  _EVAL_50,
  input         _EVAL_51,
  input  [1:0]  _EVAL_52,
  input         _EVAL_53,
  input  [31:0] _EVAL_54,
  output [2:0]  _EVAL_55,
  output [3:0]  _EVAL_56,
  input  [31:0] _EVAL_57,
  input         _EVAL_58,
  output [31:0] _EVAL_59,
  output [1:0]  _EVAL_60,
  output [1:0]  _EVAL_61,
  input  [1:0]  _EVAL_62,
  input         _EVAL_63,
  output [2:0]  _EVAL_64,
  output        _EVAL_65,
  output [2:0]  _EVAL_66,
  input  [2:0]  _EVAL_67,
  output [2:0]  _EVAL_68,
  output        _EVAL_69,
  output [24:0] _EVAL_70,
  output        _EVAL_71,
  input  [11:0] _EVAL_72,
  output [1:0]  _EVAL_73,
  output [2:0]  _EVAL_74,
  output [11:0] _EVAL_75,
  output [3:0]  _EVAL_76,
  input  [2:0]  _EVAL_77,
  output [14:0] _EVAL_78,
  output [7:0]  _EVAL_79,
  input  [2:0]  _EVAL_80,
  output [11:0] _EVAL_81,
  input         _EVAL_82,
  input  [11:0] _EVAL_83,
  input         _EVAL_84,
  input         _EVAL_85,
  input         _EVAL_86,
  output [31:0] _EVAL_87,
  output        _EVAL_88,
  input  [6:0]  _EVAL_89,
  input         _EVAL_90,
  output [25:0] _EVAL_91,
  output        _EVAL_92,
  output [2:0]  _EVAL_93,
  input  [2:0]  _EVAL_94,
  output        _EVAL_95,
  output        _EVAL_96,
  output [11:0] _EVAL_97,
  input         _EVAL_98,
  output [3:0]  _EVAL_99,
  output [29:0] _EVAL_100,
  output [2:0]  _EVAL_101,
  input  [2:0]  _EVAL_102,
  output        _EVAL_103,
  input         _EVAL_104,
  input  [1:0]  _EVAL_105,
  output        _EVAL_106,
  input         _EVAL_107,
  output [24:0] _EVAL_108,
  input  [1:0]  _EVAL_109,
  output        _EVAL_110,
  output        _EVAL_111,
  output [3:0]  _EVAL_112,
  output [11:0] _EVAL_113,
  output [2:0]  _EVAL_114,
  output [6:0]  _EVAL_115,
  input         _EVAL_116,
  input         _EVAL_117,
  output [3:0]  _EVAL_118,
  output        _EVAL_119,
  output [31:0] _EVAL_120,
  input         _EVAL_121,
  input         _EVAL_122,
  output [3:0]  _EVAL_123,
  input         _EVAL_124,
  output [2:0]  _EVAL_125,
  output [2:0]  _EVAL_126,
  input  [1:0]  _EVAL_127,
  input         _EVAL_128,
  output        _EVAL_129,
  input         _EVAL_130,
  input         _EVAL_131,
  output [2:0]  _EVAL_132,
  output [31:0] _EVAL_133,
  output [11:0] _EVAL_134,
  output        _EVAL_135,
  output        _EVAL_136,
  input  [31:0] _EVAL_137,
  input  [11:0] _EVAL_138,
  output        _EVAL_139,
  input  [6:0]  _EVAL_140,
  input  [11:0] _EVAL_141,
  output        _EVAL_142,
  output        _EVAL_143,
  input  [3:0]  _EVAL_144,
  input  [1:0]  _EVAL_145,
  input         _EVAL_146,
  input  [31:0] _EVAL_147,
  output [3:0]  _EVAL_148,
  output        _EVAL_149,
  output        _EVAL_150,
  output        _EVAL_151,
  output [1:0]  _EVAL_152,
  input         _EVAL_153,
  output        _EVAL_154,
  output [2:0]  _EVAL_155,
  output [2:0]  _EVAL_156,
  output [3:0]  _EVAL_157,
  output        _EVAL_158,
  input  [2:0]  _EVAL_159
);
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_0;
  wire [7:0] coupler_to_port_named_axi4_periph_port__EVAL_1;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_2;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_3;
  wire [1:0] coupler_to_port_named_axi4_periph_port__EVAL_4;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_5;
  wire [1:0] coupler_to_port_named_axi4_periph_port__EVAL_6;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_7;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_8;
  wire [29:0] coupler_to_port_named_axi4_periph_port__EVAL_9;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_10;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_11;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_12;
  wire [3:0] coupler_to_port_named_axi4_periph_port__EVAL_13;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_14;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_15;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_16;
  wire [6:0] coupler_to_port_named_axi4_periph_port__EVAL_17;
  wire [3:0] coupler_to_port_named_axi4_periph_port__EVAL_18;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_19;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_20;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_21;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_22;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_23;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_24;
  wire [3:0] coupler_to_port_named_axi4_periph_port__EVAL_25;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_26;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_27;
  wire [6:0] coupler_to_port_named_axi4_periph_port__EVAL_28;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_29;
  wire [31:0] coupler_to_port_named_axi4_periph_port__EVAL_30;
  wire [3:0] coupler_to_port_named_axi4_periph_port__EVAL_31;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_32;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_33;
  wire [31:0] coupler_to_port_named_axi4_periph_port__EVAL_34;
  wire [7:0] coupler_to_port_named_axi4_periph_port__EVAL_35;
  wire [3:0] coupler_to_port_named_axi4_periph_port__EVAL_36;
  wire [29:0] coupler_to_port_named_axi4_periph_port__EVAL_37;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_38;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_39;
  wire [1:0] coupler_to_port_named_axi4_periph_port__EVAL_40;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_41;
  wire [31:0] coupler_to_port_named_axi4_periph_port__EVAL_42;
  wire [3:0] coupler_to_port_named_axi4_periph_port__EVAL_43;
  wire [29:0] coupler_to_port_named_axi4_periph_port__EVAL_44;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_45;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_46;
  wire [31:0] coupler_to_port_named_axi4_periph_port__EVAL_47;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_48;
  wire [2:0] coupler_to_port_named_axi4_periph_port__EVAL_49;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_50;
  wire [1:0] coupler_to_port_named_axi4_periph_port__EVAL_51;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_52;
  wire  coupler_to_port_named_axi4_periph_port__EVAL_53;
  wire [27:0] out_xbar__EVAL;
  wire  out_xbar__EVAL_0;
  wire [31:0] out_xbar__EVAL_1;
  wire [2:0] out_xbar__EVAL_2;
  wire  out_xbar__EVAL_3;
  wire [2:0] out_xbar__EVAL_4;
  wire [6:0] out_xbar__EVAL_5;
  wire [3:0] out_xbar__EVAL_6;
  wire  out_xbar__EVAL_7;
  wire [2:0] out_xbar__EVAL_8;
  wire [2:0] out_xbar__EVAL_9;
  wire [29:0] out_xbar__EVAL_10;
  wire [2:0] out_xbar__EVAL_11;
  wire [3:0] out_xbar__EVAL_12;
  wire  out_xbar__EVAL_13;
  wire  out_xbar__EVAL_14;
  wire [6:0] out_xbar__EVAL_15;
  wire  out_xbar__EVAL_16;
  wire  out_xbar__EVAL_17;
  wire [2:0] out_xbar__EVAL_18;
  wire [2:0] out_xbar__EVAL_19;
  wire [6:0] out_xbar__EVAL_20;
  wire [2:0] out_xbar__EVAL_21;
  wire [2:0] out_xbar__EVAL_22;
  wire [13:0] out_xbar__EVAL_23;
  wire  out_xbar__EVAL_24;
  wire  out_xbar__EVAL_25;
  wire [6:0] out_xbar__EVAL_26;
  wire [2:0] out_xbar__EVAL_27;
  wire [2:0] out_xbar__EVAL_28;
  wire  out_xbar__EVAL_29;
  wire [2:0] out_xbar__EVAL_30;
  wire  out_xbar__EVAL_31;
  wire [2:0] out_xbar__EVAL_32;
  wire  out_xbar__EVAL_33;
  wire [3:0] out_xbar__EVAL_34;
  wire [6:0] out_xbar__EVAL_35;
  wire [6:0] out_xbar__EVAL_36;
  wire  out_xbar__EVAL_37;
  wire [29:0] out_xbar__EVAL_38;
  wire  out_xbar__EVAL_39;
  wire [31:0] out_xbar__EVAL_40;
  wire  out_xbar__EVAL_41;
  wire [2:0] out_xbar__EVAL_42;
  wire [2:0] out_xbar__EVAL_43;
  wire [31:0] out_xbar__EVAL_44;
  wire  out_xbar__EVAL_45;
  wire [6:0] out_xbar__EVAL_46;
  wire [2:0] out_xbar__EVAL_47;
  wire [6:0] out_xbar__EVAL_48;
  wire  out_xbar__EVAL_49;
  wire [6:0] out_xbar__EVAL_50;
  wire [2:0] out_xbar__EVAL_51;
  wire [31:0] out_xbar__EVAL_52;
  wire [6:0] out_xbar__EVAL_53;
  wire [6:0] out_xbar__EVAL_54;
  wire [14:0] out_xbar__EVAL_55;
  wire [3:0] out_xbar__EVAL_56;
  wire  out_xbar__EVAL_57;
  wire [2:0] out_xbar__EVAL_58;
  wire [3:0] out_xbar__EVAL_59;
  wire  out_xbar__EVAL_60;
  wire  out_xbar__EVAL_61;
  wire [2:0] out_xbar__EVAL_62;
  wire  out_xbar__EVAL_63;
  wire  out_xbar__EVAL_64;
  wire [31:0] out_xbar__EVAL_65;
  wire  out_xbar__EVAL_66;
  wire  out_xbar__EVAL_67;
  wire [3:0] out_xbar__EVAL_68;
  wire [3:0] out_xbar__EVAL_69;
  wire  out_xbar__EVAL_70;
  wire [3:0] out_xbar__EVAL_71;
  wire  out_xbar__EVAL_72;
  wire  out_xbar__EVAL_73;
  wire [31:0] out_xbar__EVAL_74;
  wire [6:0] out_xbar__EVAL_75;
  wire  out_xbar__EVAL_76;
  wire  out_xbar__EVAL_77;
  wire  out_xbar__EVAL_78;
  wire  out_xbar__EVAL_79;
  wire  out_xbar__EVAL_80;
  wire [31:0] out_xbar__EVAL_81;
  wire  out_xbar__EVAL_82;
  wire [24:0] out_xbar__EVAL_83;
  wire  out_xbar__EVAL_84;
  wire [2:0] out_xbar__EVAL_85;
  wire [6:0] out_xbar__EVAL_86;
  wire  out_xbar__EVAL_87;
  wire  out_xbar__EVAL_88;
  wire [1:0] out_xbar__EVAL_89;
  wire [6:0] out_xbar__EVAL_90;
  wire [2:0] out_xbar__EVAL_91;
  wire  out_xbar__EVAL_92;
  wire [31:0] out_xbar__EVAL_93;
  wire [3:0] out_xbar__EVAL_94;
  wire [2:0] out_xbar__EVAL_95;
  wire [31:0] out_xbar__EVAL_96;
  wire  out_xbar__EVAL_97;
  wire [25:0] out_xbar__EVAL_98;
  wire [3:0] out_xbar__EVAL_99;
  wire  out_xbar__EVAL_100;
  wire  out_xbar__EVAL_101;
  wire [2:0] out_xbar__EVAL_102;
  wire  out_xbar__EVAL_103;
  wire [2:0] out_xbar__EVAL_104;
  wire [2:0] out_xbar__EVAL_105;
  wire [31:0] out_xbar__EVAL_106;
  wire [2:0] out_xbar__EVAL_107;
  wire [6:0] out_xbar__EVAL_108;
  wire  out_xbar__EVAL_109;
  wire [31:0] out_xbar__EVAL_110;
  wire [2:0] out_xbar__EVAL_111;
  wire  out_xbar__EVAL_112;
  wire [3:0] out_xbar__EVAL_113;
  wire [6:0] out_xbar__EVAL_114;
  wire [11:0] out_xbar__EVAL_115;
  wire [2:0] out_xbar__EVAL_116;
  wire [2:0] out_xbar__EVAL_117;
  wire  out_xbar__EVAL_118;
  wire [31:0] out_xbar__EVAL_119;
  wire [31:0] out_xbar__EVAL_120;
  wire [2:0] out_xbar__EVAL_121;
  wire  out_xbar__EVAL_122;
  wire  out_xbar__EVAL_123;
  wire  out_xbar__EVAL_124;
  wire [2:0] out_xbar__EVAL_125;
  wire [2:0] out_xbar__EVAL_126;
  wire [3:0] out_xbar__EVAL_127;
  wire  out_xbar__EVAL_128;
  wire  out_xbar__EVAL_129;
  wire  out_xbar__EVAL_130;
  wire  out_xbar__EVAL_131;
  wire [1:0] out_xbar__EVAL_132;
  wire [2:0] out_xbar__EVAL_133;
  wire  out_xbar__EVAL_134;
  wire [1:0] out_xbar__EVAL_135;
  wire [2:0] out_xbar__EVAL_136;
  wire  out_xbar__EVAL_137;
  wire [31:0] out_xbar__EVAL_138;
  wire [2:0] out_xbar__EVAL_139;
  wire [31:0] out_xbar__EVAL_140;
  wire [2:0] out_xbar__EVAL_141;
  wire  coupler_to_debug__EVAL;
  wire  coupler_to_debug__EVAL_0;
  wire [11:0] coupler_to_debug__EVAL_1;
  wire [31:0] coupler_to_debug__EVAL_2;
  wire [2:0] coupler_to_debug__EVAL_3;
  wire [3:0] coupler_to_debug__EVAL_4;
  wire [11:0] coupler_to_debug__EVAL_5;
  wire  coupler_to_debug__EVAL_6;
  wire  coupler_to_debug__EVAL_7;
  wire [31:0] coupler_to_debug__EVAL_8;
  wire  coupler_to_debug__EVAL_9;
  wire  coupler_to_debug__EVAL_10;
  wire [11:0] coupler_to_debug__EVAL_11;
  wire [6:0] coupler_to_debug__EVAL_12;
  wire [2:0] coupler_to_debug__EVAL_13;
  wire [11:0] coupler_to_debug__EVAL_14;
  wire [6:0] coupler_to_debug__EVAL_15;
  wire [2:0] coupler_to_debug__EVAL_16;
  wire [1:0] coupler_to_debug__EVAL_17;
  wire [3:0] coupler_to_debug__EVAL_18;
  wire [2:0] coupler_to_debug__EVAL_19;
  wire [2:0] coupler_to_debug__EVAL_20;
  wire [31:0] coupler_to_debug__EVAL_21;
  wire [2:0] coupler_to_debug__EVAL_22;
  wire [31:0] coupler_to_debug__EVAL_23;
  wire  coupler_to_debug__EVAL_24;
  wire  coupler_to_debug__EVAL_25;
  wire  coupler_to_debug__EVAL_26;
  wire  coupler_to_debug__EVAL_27;
  wire [1:0] coupler_to_debug__EVAL_28;
  wire  coupler_to_debug__EVAL_29;
  wire [2:0] coupler_to_debug__EVAL_30;
  wire [2:0] coupler_to_debug__EVAL_31;
  wire  coupler_to_debug__EVAL_32;
  wire [31:0] in_xbar__EVAL;
  wire  in_xbar__EVAL_0;
  wire [1:0] in_xbar__EVAL_1;
  wire [3:0] in_xbar__EVAL_2;
  wire [31:0] in_xbar__EVAL_3;
  wire [29:0] in_xbar__EVAL_4;
  wire [31:0] in_xbar__EVAL_5;
  wire [3:0] in_xbar__EVAL_6;
  wire  in_xbar__EVAL_7;
  wire  in_xbar__EVAL_8;
  wire [31:0] in_xbar__EVAL_9;
  wire  in_xbar__EVAL_10;
  wire [6:0] in_xbar__EVAL_11;
  wire  in_xbar__EVAL_12;
  wire  in_xbar__EVAL_13;
  wire  in_xbar__EVAL_14;
  wire [2:0] in_xbar__EVAL_15;
  wire [29:0] in_xbar__EVAL_16;
  wire [2:0] in_xbar__EVAL_17;
  wire [6:0] in_xbar__EVAL_18;
  wire [3:0] in_xbar__EVAL_19;
  wire [3:0] in_xbar__EVAL_20;
  wire [6:0] in_xbar__EVAL_21;
  wire  in_xbar__EVAL_22;
  wire [6:0] in_xbar__EVAL_23;
  wire  in_xbar__EVAL_24;
  wire  in_xbar__EVAL_25;
  wire  in_xbar__EVAL_26;
  wire [2:0] in_xbar__EVAL_27;
  wire [3:0] in_xbar__EVAL_28;
  wire  in_xbar__EVAL_29;
  wire [2:0] in_xbar__EVAL_30;
  wire [1:0] in_xbar__EVAL_31;
  wire  in_xbar__EVAL_32;
  wire  in_xbar__EVAL_33;
  wire  in_xbar__EVAL_34;
  wire [3:0] in_xbar__EVAL_35;
  wire  in_xbar__EVAL_36;
  wire  in_xbar__EVAL_37;
  wire [2:0] in_xbar__EVAL_38;
  wire [2:0] in_xbar__EVAL_39;
  wire  in_xbar__EVAL_40;
  wire  buffer__EVAL;
  wire [6:0] buffer__EVAL_0;
  wire [6:0] buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire [3:0] buffer__EVAL_3;
  wire [2:0] buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [31:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [3:0] buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [2:0] buffer__EVAL_10;
  wire [6:0] buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire [31:0] buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire [2:0] buffer__EVAL_16;
  wire [29:0] buffer__EVAL_17;
  wire [6:0] buffer__EVAL_18;
  wire [2:0] buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire [31:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire [31:0] buffer__EVAL_25;
  wire [1:0] buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [29:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [3:0] buffer__EVAL_33;
  wire [3:0] buffer__EVAL_34;
  wire [2:0] buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [3:0] buffer__EVAL_37;
  wire [2:0] buffer__EVAL_38;
  wire [1:0] buffer__EVAL_39;
  wire [3:0] buffer__EVAL_40;
  wire [2:0] buffer_1__EVAL;
  wire  buffer_1__EVAL_0;
  wire  buffer_1__EVAL_1;
  wire [1:0] buffer_1__EVAL_2;
  wire [3:0] buffer_1__EVAL_3;
  wire [1:0] buffer_1__EVAL_4;
  wire  buffer_1__EVAL_5;
  wire  buffer_1__EVAL_6;
  wire [3:0] buffer_1__EVAL_7;
  wire  buffer_1__EVAL_8;
  wire [3:0] buffer_1__EVAL_9;
  wire [6:0] buffer_1__EVAL_10;
  wire [2:0] buffer_1__EVAL_11;
  wire  buffer_1__EVAL_12;
  wire [31:0] buffer_1__EVAL_13;
  wire  buffer_1__EVAL_14;
  wire  buffer_1__EVAL_15;
  wire  buffer_1__EVAL_16;
  wire [29:0] buffer_1__EVAL_17;
  wire  buffer_1__EVAL_18;
  wire [2:0] buffer_1__EVAL_19;
  wire [3:0] buffer_1__EVAL_20;
  wire [6:0] buffer_1__EVAL_21;
  wire  buffer_1__EVAL_22;
  wire [3:0] buffer_1__EVAL_23;
  wire  buffer_1__EVAL_24;
  wire [6:0] buffer_1__EVAL_25;
  wire  buffer_1__EVAL_26;
  wire  buffer_1__EVAL_27;
  wire [31:0] buffer_1__EVAL_28;
  wire [31:0] buffer_1__EVAL_29;
  wire [6:0] buffer_1__EVAL_30;
  wire [29:0] buffer_1__EVAL_31;
  wire [31:0] buffer_1__EVAL_32;
  wire  buffer_1__EVAL_33;
  wire [3:0] buffer_1__EVAL_34;
  wire [2:0] buffer_1__EVAL_35;
  wire  buffer_1__EVAL_36;
  wire [2:0] buffer_1__EVAL_37;
  wire [2:0] buffer_1__EVAL_38;
  wire  buffer_1__EVAL_39;
  wire  buffer_1__EVAL_40;
  wire [2:0] coupler_to_tile_with_no_name__EVAL;
  wire  coupler_to_tile_with_no_name__EVAL_0;
  wire  coupler_to_tile_with_no_name__EVAL_1;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_2;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_3;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_4;
  wire [6:0] coupler_to_tile_with_no_name__EVAL_5;
  wire  coupler_to_tile_with_no_name__EVAL_6;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_7;
  wire [6:0] coupler_to_tile_with_no_name__EVAL_8;
  wire  coupler_to_tile_with_no_name__EVAL_9;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_10;
  wire [31:0] coupler_to_tile_with_no_name__EVAL_11;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_12;
  wire [6:0] coupler_to_tile_with_no_name__EVAL_13;
  wire  coupler_to_tile_with_no_name__EVAL_14;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_15;
  wire  coupler_to_tile_with_no_name__EVAL_16;
  wire  coupler_to_tile_with_no_name__EVAL_17;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_18;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_19;
  wire  coupler_to_tile_with_no_name__EVAL_20;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_21;
  wire  coupler_to_tile_with_no_name__EVAL_22;
  wire  coupler_to_tile_with_no_name__EVAL_23;
  wire [6:0] coupler_to_tile_with_no_name__EVAL_24;
  wire [3:0] coupler_to_tile_with_no_name__EVAL_25;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_26;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_27;
  wire  coupler_to_tile_with_no_name__EVAL_28;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_29;
  wire  coupler_to_tile_with_no_name__EVAL_30;
  wire [3:0] coupler_to_tile_with_no_name__EVAL_31;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_32;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_33;
  wire  coupler_to_tile_with_no_name__EVAL_34;
  wire [24:0] coupler_to_tile_with_no_name__EVAL_35;
  wire [6:0] coupler_to_tile_with_no_name__EVAL_36;
  wire  coupler_to_tile_with_no_name__EVAL_37;
  wire [24:0] coupler_to_tile_with_no_name__EVAL_38;
  wire  coupler_to_tile_with_no_name__EVAL_39;
  wire [6:0] coupler_to_tile_with_no_name__EVAL_40;
  wire  coupler_to_tile_with_no_name__EVAL_41;
  wire [31:0] coupler_to_tile_with_no_name__EVAL_42;
  wire  coupler_to_tile_with_no_name__EVAL_43;
  wire [24:0] coupler_to_tile_with_no_name__EVAL_44;
  wire [31:0] coupler_to_tile_with_no_name__EVAL_45;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_46;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_47;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_48;
  wire  coupler_to_tile_with_no_name__EVAL_49;
  wire [1:0] coupler_to_tile_with_no_name__EVAL_50;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_51;
  wire [2:0] coupler_to_tile_with_no_name__EVAL_52;
  wire  coupler_to_tile_with_no_name__EVAL_53;
  wire [3:0] coupler_to_tile_with_no_name__EVAL_54;
  wire  coupler_to_tile_with_no_name__EVAL_55;
  wire  coupler_to_tile_with_no_name__EVAL_56;
  wire [31:0] coupler_to_tile_with_no_name__EVAL_57;
  wire [31:0] coupler_to_tile_with_no_name__EVAL_58;
  wire [31:0] coupler_to_tile_with_no_name__EVAL_59;
  wire  coupler_to_tile_with_no_name__EVAL_60;
  wire [2:0] wrapped_error_device__EVAL;
  wire  wrapped_error_device__EVAL_0;
  wire [31:0] wrapped_error_device__EVAL_1;
  wire [13:0] wrapped_error_device__EVAL_2;
  wire  wrapped_error_device__EVAL_3;
  wire  wrapped_error_device__EVAL_4;
  wire [3:0] wrapped_error_device__EVAL_5;
  wire  wrapped_error_device__EVAL_6;
  wire  wrapped_error_device__EVAL_7;
  wire  wrapped_error_device__EVAL_8;
  wire  wrapped_error_device__EVAL_9;
  wire  wrapped_error_device__EVAL_10;
  wire [2:0] wrapped_error_device__EVAL_11;
  wire  wrapped_error_device__EVAL_12;
  wire [2:0] wrapped_error_device__EVAL_13;
  wire [6:0] wrapped_error_device__EVAL_14;
  wire [3:0] wrapped_error_device__EVAL_15;
  wire [3:0] wrapped_error_device__EVAL_16;
  wire  wrapped_error_device__EVAL_17;
  wire [1:0] wrapped_error_device__EVAL_18;
  wire [6:0] wrapped_error_device__EVAL_19;
  wire [2:0] fixer__EVAL;
  wire  fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire [2:0] fixer__EVAL_2;
  wire [3:0] fixer__EVAL_3;
  wire  fixer__EVAL_4;
  wire  fixer__EVAL_5;
  wire [31:0] fixer__EVAL_6;
  wire [29:0] fixer__EVAL_7;
  wire [31:0] fixer__EVAL_8;
  wire  fixer__EVAL_9;
  wire  fixer__EVAL_10;
  wire  fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire [2:0] fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire [1:0] fixer__EVAL_15;
  wire [29:0] fixer__EVAL_16;
  wire [6:0] fixer__EVAL_17;
  wire [3:0] fixer__EVAL_18;
  wire [2:0] fixer__EVAL_19;
  wire  fixer__EVAL_20;
  wire [6:0] fixer__EVAL_21;
  wire [2:0] fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire  fixer__EVAL_24;
  wire [31:0] fixer__EVAL_25;
  wire [3:0] fixer__EVAL_26;
  wire  fixer__EVAL_27;
  wire [3:0] fixer__EVAL_28;
  wire [31:0] fixer__EVAL_29;
  wire [6:0] fixer__EVAL_30;
  wire [3:0] fixer__EVAL_31;
  wire  fixer__EVAL_32;
  wire  fixer__EVAL_33;
  wire [6:0] fixer__EVAL_34;
  wire [1:0] fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire [2:0] fixer__EVAL_37;
  wire  fixer__EVAL_38;
  wire  fixer__EVAL_39;
  wire [3:0] fixer__EVAL_40;
  wire  coupler_to_testindicator__EVAL;
  wire [2:0] coupler_to_testindicator__EVAL_0;
  wire [2:0] coupler_to_testindicator__EVAL_1;
  wire  coupler_to_testindicator__EVAL_2;
  wire  coupler_to_testindicator__EVAL_3;
  wire  coupler_to_testindicator__EVAL_4;
  wire [1:0] coupler_to_testindicator__EVAL_5;
  wire [11:0] coupler_to_testindicator__EVAL_6;
  wire [3:0] coupler_to_testindicator__EVAL_7;
  wire [2:0] coupler_to_testindicator__EVAL_8;
  wire [2:0] coupler_to_testindicator__EVAL_9;
  wire [14:0] coupler_to_testindicator__EVAL_10;
  wire [11:0] coupler_to_testindicator__EVAL_11;
  wire [3:0] coupler_to_testindicator__EVAL_12;
  wire  coupler_to_testindicator__EVAL_13;
  wire [6:0] coupler_to_testindicator__EVAL_14;
  wire [2:0] coupler_to_testindicator__EVAL_15;
  wire [14:0] coupler_to_testindicator__EVAL_16;
  wire  coupler_to_testindicator__EVAL_17;
  wire [31:0] coupler_to_testindicator__EVAL_18;
  wire  coupler_to_testindicator__EVAL_19;
  wire [31:0] coupler_to_testindicator__EVAL_20;
  wire  coupler_to_testindicator__EVAL_21;
  wire  coupler_to_testindicator__EVAL_22;
  wire  coupler_to_testindicator__EVAL_23;
  wire [2:0] coupler_to_testindicator__EVAL_24;
  wire [2:0] coupler_to_testindicator__EVAL_25;
  wire  coupler_to_testindicator__EVAL_26;
  wire [6:0] coupler_to_testindicator__EVAL_27;
  wire [31:0] coupler_to_testindicator__EVAL_28;
  wire [31:0] coupler_to_testindicator__EVAL_29;
  wire  coupler_to_testindicator__EVAL_30;
  wire [1:0] coupler_to_testindicator__EVAL_31;
  wire [2:0] coupler_to_testindicator__EVAL_32;
  wire [2:0] coupler_to_clint__EVAL;
  wire [25:0] coupler_to_clint__EVAL_0;
  wire [2:0] coupler_to_clint__EVAL_1;
  wire [31:0] coupler_to_clint__EVAL_2;
  wire  coupler_to_clint__EVAL_3;
  wire [1:0] coupler_to_clint__EVAL_4;
  wire [1:0] coupler_to_clint__EVAL_5;
  wire  coupler_to_clint__EVAL_6;
  wire [2:0] coupler_to_clint__EVAL_7;
  wire  coupler_to_clint__EVAL_8;
  wire [11:0] coupler_to_clint__EVAL_9;
  wire [11:0] coupler_to_clint__EVAL_10;
  wire  coupler_to_clint__EVAL_11;
  wire  coupler_to_clint__EVAL_12;
  wire [25:0] coupler_to_clint__EVAL_13;
  wire [2:0] coupler_to_clint__EVAL_14;
  wire [2:0] coupler_to_clint__EVAL_15;
  wire [6:0] coupler_to_clint__EVAL_16;
  wire [2:0] coupler_to_clint__EVAL_17;
  wire [6:0] coupler_to_clint__EVAL_18;
  wire  coupler_to_clint__EVAL_19;
  wire [31:0] coupler_to_clint__EVAL_20;
  wire [31:0] coupler_to_clint__EVAL_21;
  wire  coupler_to_clint__EVAL_22;
  wire [3:0] coupler_to_clint__EVAL_23;
  wire  coupler_to_clint__EVAL_24;
  wire  coupler_to_clint__EVAL_25;
  wire  coupler_to_clint__EVAL_26;
  wire  coupler_to_clint__EVAL_27;
  wire [31:0] coupler_to_clint__EVAL_28;
  wire [2:0] coupler_to_clint__EVAL_29;
  wire  coupler_to_clint__EVAL_30;
  wire [3:0] coupler_to_clint__EVAL_31;
  wire [2:0] coupler_to_clint__EVAL_32;
  wire [2:0] coupler_to_plic__EVAL;
  wire  coupler_to_plic__EVAL_0;
  wire  coupler_to_plic__EVAL_1;
  wire [31:0] coupler_to_plic__EVAL_2;
  wire [11:0] coupler_to_plic__EVAL_3;
  wire  coupler_to_plic__EVAL_4;
  wire  coupler_to_plic__EVAL_5;
  wire [11:0] coupler_to_plic__EVAL_6;
  wire [2:0] coupler_to_plic__EVAL_7;
  wire [1:0] coupler_to_plic__EVAL_8;
  wire  coupler_to_plic__EVAL_9;
  wire [2:0] coupler_to_plic__EVAL_10;
  wire [27:0] coupler_to_plic__EVAL_11;
  wire [2:0] coupler_to_plic__EVAL_12;
  wire  coupler_to_plic__EVAL_13;
  wire [3:0] coupler_to_plic__EVAL_14;
  wire [2:0] coupler_to_plic__EVAL_15;
  wire  coupler_to_plic__EVAL_16;
  wire  coupler_to_plic__EVAL_17;
  wire [2:0] coupler_to_plic__EVAL_18;
  wire [6:0] coupler_to_plic__EVAL_19;
  wire [2:0] coupler_to_plic__EVAL_20;
  wire [31:0] coupler_to_plic__EVAL_21;
  wire  coupler_to_plic__EVAL_22;
  wire [27:0] coupler_to_plic__EVAL_23;
  wire [3:0] coupler_to_plic__EVAL_24;
  wire  coupler_to_plic__EVAL_25;
  wire [2:0] coupler_to_plic__EVAL_26;
  wire [31:0] coupler_to_plic__EVAL_27;
  wire [31:0] coupler_to_plic__EVAL_28;
  wire  coupler_to_plic__EVAL_29;
  wire  coupler_to_plic__EVAL_30;
  wire [6:0] coupler_to_plic__EVAL_31;
  wire [1:0] coupler_to_plic__EVAL_32;
  wire  atomics__EVAL;
  wire [31:0] atomics__EVAL_0;
  wire  atomics__EVAL_1;
  wire  atomics__EVAL_2;
  wire [1:0] atomics__EVAL_3;
  wire  atomics__EVAL_4;
  wire [1:0] atomics__EVAL_5;
  wire [6:0] atomics__EVAL_6;
  wire  atomics__EVAL_7;
  wire  atomics__EVAL_8;
  wire  atomics__EVAL_9;
  wire  atomics__EVAL_10;
  wire [29:0] atomics__EVAL_11;
  wire [2:0] atomics__EVAL_12;
  wire [3:0] atomics__EVAL_13;
  wire [2:0] atomics__EVAL_14;
  wire [3:0] atomics__EVAL_15;
  wire [2:0] atomics__EVAL_16;
  wire  atomics__EVAL_17;
  wire [2:0] atomics__EVAL_18;
  wire [31:0] atomics__EVAL_19;
  wire  atomics__EVAL_20;
  wire [6:0] atomics__EVAL_21;
  wire [6:0] atomics__EVAL_22;
  wire  atomics__EVAL_23;
  wire  atomics__EVAL_24;
  wire [3:0] atomics__EVAL_25;
  wire  atomics__EVAL_26;
  wire [29:0] atomics__EVAL_27;
  wire [31:0] atomics__EVAL_28;
  wire [3:0] atomics__EVAL_29;
  wire  atomics__EVAL_30;
  wire  atomics__EVAL_31;
  wire  atomics__EVAL_32;
  wire [6:0] atomics__EVAL_33;
  wire  atomics__EVAL_34;
  wire [3:0] atomics__EVAL_35;
  wire [2:0] atomics__EVAL_36;
  wire [3:0] atomics__EVAL_37;
  wire  atomics__EVAL_38;
  wire [31:0] atomics__EVAL_39;
  wire [2:0] atomics__EVAL_40;
  SiFive__EVAL_177 coupler_to_port_named_axi4_periph_port (
    ._EVAL(coupler_to_port_named_axi4_periph_port__EVAL),
    ._EVAL_0(coupler_to_port_named_axi4_periph_port__EVAL_0),
    ._EVAL_1(coupler_to_port_named_axi4_periph_port__EVAL_1),
    ._EVAL_2(coupler_to_port_named_axi4_periph_port__EVAL_2),
    ._EVAL_3(coupler_to_port_named_axi4_periph_port__EVAL_3),
    ._EVAL_4(coupler_to_port_named_axi4_periph_port__EVAL_4),
    ._EVAL_5(coupler_to_port_named_axi4_periph_port__EVAL_5),
    ._EVAL_6(coupler_to_port_named_axi4_periph_port__EVAL_6),
    ._EVAL_7(coupler_to_port_named_axi4_periph_port__EVAL_7),
    ._EVAL_8(coupler_to_port_named_axi4_periph_port__EVAL_8),
    ._EVAL_9(coupler_to_port_named_axi4_periph_port__EVAL_9),
    ._EVAL_10(coupler_to_port_named_axi4_periph_port__EVAL_10),
    ._EVAL_11(coupler_to_port_named_axi4_periph_port__EVAL_11),
    ._EVAL_12(coupler_to_port_named_axi4_periph_port__EVAL_12),
    ._EVAL_13(coupler_to_port_named_axi4_periph_port__EVAL_13),
    ._EVAL_14(coupler_to_port_named_axi4_periph_port__EVAL_14),
    ._EVAL_15(coupler_to_port_named_axi4_periph_port__EVAL_15),
    ._EVAL_16(coupler_to_port_named_axi4_periph_port__EVAL_16),
    ._EVAL_17(coupler_to_port_named_axi4_periph_port__EVAL_17),
    ._EVAL_18(coupler_to_port_named_axi4_periph_port__EVAL_18),
    ._EVAL_19(coupler_to_port_named_axi4_periph_port__EVAL_19),
    ._EVAL_20(coupler_to_port_named_axi4_periph_port__EVAL_20),
    ._EVAL_21(coupler_to_port_named_axi4_periph_port__EVAL_21),
    ._EVAL_22(coupler_to_port_named_axi4_periph_port__EVAL_22),
    ._EVAL_23(coupler_to_port_named_axi4_periph_port__EVAL_23),
    ._EVAL_24(coupler_to_port_named_axi4_periph_port__EVAL_24),
    ._EVAL_25(coupler_to_port_named_axi4_periph_port__EVAL_25),
    ._EVAL_26(coupler_to_port_named_axi4_periph_port__EVAL_26),
    ._EVAL_27(coupler_to_port_named_axi4_periph_port__EVAL_27),
    ._EVAL_28(coupler_to_port_named_axi4_periph_port__EVAL_28),
    ._EVAL_29(coupler_to_port_named_axi4_periph_port__EVAL_29),
    ._EVAL_30(coupler_to_port_named_axi4_periph_port__EVAL_30),
    ._EVAL_31(coupler_to_port_named_axi4_periph_port__EVAL_31),
    ._EVAL_32(coupler_to_port_named_axi4_periph_port__EVAL_32),
    ._EVAL_33(coupler_to_port_named_axi4_periph_port__EVAL_33),
    ._EVAL_34(coupler_to_port_named_axi4_periph_port__EVAL_34),
    ._EVAL_35(coupler_to_port_named_axi4_periph_port__EVAL_35),
    ._EVAL_36(coupler_to_port_named_axi4_periph_port__EVAL_36),
    ._EVAL_37(coupler_to_port_named_axi4_periph_port__EVAL_37),
    ._EVAL_38(coupler_to_port_named_axi4_periph_port__EVAL_38),
    ._EVAL_39(coupler_to_port_named_axi4_periph_port__EVAL_39),
    ._EVAL_40(coupler_to_port_named_axi4_periph_port__EVAL_40),
    ._EVAL_41(coupler_to_port_named_axi4_periph_port__EVAL_41),
    ._EVAL_42(coupler_to_port_named_axi4_periph_port__EVAL_42),
    ._EVAL_43(coupler_to_port_named_axi4_periph_port__EVAL_43),
    ._EVAL_44(coupler_to_port_named_axi4_periph_port__EVAL_44),
    ._EVAL_45(coupler_to_port_named_axi4_periph_port__EVAL_45),
    ._EVAL_46(coupler_to_port_named_axi4_periph_port__EVAL_46),
    ._EVAL_47(coupler_to_port_named_axi4_periph_port__EVAL_47),
    ._EVAL_48(coupler_to_port_named_axi4_periph_port__EVAL_48),
    ._EVAL_49(coupler_to_port_named_axi4_periph_port__EVAL_49),
    ._EVAL_50(coupler_to_port_named_axi4_periph_port__EVAL_50),
    ._EVAL_51(coupler_to_port_named_axi4_periph_port__EVAL_51),
    ._EVAL_52(coupler_to_port_named_axi4_periph_port__EVAL_52),
    ._EVAL_53(coupler_to_port_named_axi4_periph_port__EVAL_53)
  );
  SiFive__EVAL_116 out_xbar (
    ._EVAL(out_xbar__EVAL),
    ._EVAL_0(out_xbar__EVAL_0),
    ._EVAL_1(out_xbar__EVAL_1),
    ._EVAL_2(out_xbar__EVAL_2),
    ._EVAL_3(out_xbar__EVAL_3),
    ._EVAL_4(out_xbar__EVAL_4),
    ._EVAL_5(out_xbar__EVAL_5),
    ._EVAL_6(out_xbar__EVAL_6),
    ._EVAL_7(out_xbar__EVAL_7),
    ._EVAL_8(out_xbar__EVAL_8),
    ._EVAL_9(out_xbar__EVAL_9),
    ._EVAL_10(out_xbar__EVAL_10),
    ._EVAL_11(out_xbar__EVAL_11),
    ._EVAL_12(out_xbar__EVAL_12),
    ._EVAL_13(out_xbar__EVAL_13),
    ._EVAL_14(out_xbar__EVAL_14),
    ._EVAL_15(out_xbar__EVAL_15),
    ._EVAL_16(out_xbar__EVAL_16),
    ._EVAL_17(out_xbar__EVAL_17),
    ._EVAL_18(out_xbar__EVAL_18),
    ._EVAL_19(out_xbar__EVAL_19),
    ._EVAL_20(out_xbar__EVAL_20),
    ._EVAL_21(out_xbar__EVAL_21),
    ._EVAL_22(out_xbar__EVAL_22),
    ._EVAL_23(out_xbar__EVAL_23),
    ._EVAL_24(out_xbar__EVAL_24),
    ._EVAL_25(out_xbar__EVAL_25),
    ._EVAL_26(out_xbar__EVAL_26),
    ._EVAL_27(out_xbar__EVAL_27),
    ._EVAL_28(out_xbar__EVAL_28),
    ._EVAL_29(out_xbar__EVAL_29),
    ._EVAL_30(out_xbar__EVAL_30),
    ._EVAL_31(out_xbar__EVAL_31),
    ._EVAL_32(out_xbar__EVAL_32),
    ._EVAL_33(out_xbar__EVAL_33),
    ._EVAL_34(out_xbar__EVAL_34),
    ._EVAL_35(out_xbar__EVAL_35),
    ._EVAL_36(out_xbar__EVAL_36),
    ._EVAL_37(out_xbar__EVAL_37),
    ._EVAL_38(out_xbar__EVAL_38),
    ._EVAL_39(out_xbar__EVAL_39),
    ._EVAL_40(out_xbar__EVAL_40),
    ._EVAL_41(out_xbar__EVAL_41),
    ._EVAL_42(out_xbar__EVAL_42),
    ._EVAL_43(out_xbar__EVAL_43),
    ._EVAL_44(out_xbar__EVAL_44),
    ._EVAL_45(out_xbar__EVAL_45),
    ._EVAL_46(out_xbar__EVAL_46),
    ._EVAL_47(out_xbar__EVAL_47),
    ._EVAL_48(out_xbar__EVAL_48),
    ._EVAL_49(out_xbar__EVAL_49),
    ._EVAL_50(out_xbar__EVAL_50),
    ._EVAL_51(out_xbar__EVAL_51),
    ._EVAL_52(out_xbar__EVAL_52),
    ._EVAL_53(out_xbar__EVAL_53),
    ._EVAL_54(out_xbar__EVAL_54),
    ._EVAL_55(out_xbar__EVAL_55),
    ._EVAL_56(out_xbar__EVAL_56),
    ._EVAL_57(out_xbar__EVAL_57),
    ._EVAL_58(out_xbar__EVAL_58),
    ._EVAL_59(out_xbar__EVAL_59),
    ._EVAL_60(out_xbar__EVAL_60),
    ._EVAL_61(out_xbar__EVAL_61),
    ._EVAL_62(out_xbar__EVAL_62),
    ._EVAL_63(out_xbar__EVAL_63),
    ._EVAL_64(out_xbar__EVAL_64),
    ._EVAL_65(out_xbar__EVAL_65),
    ._EVAL_66(out_xbar__EVAL_66),
    ._EVAL_67(out_xbar__EVAL_67),
    ._EVAL_68(out_xbar__EVAL_68),
    ._EVAL_69(out_xbar__EVAL_69),
    ._EVAL_70(out_xbar__EVAL_70),
    ._EVAL_71(out_xbar__EVAL_71),
    ._EVAL_72(out_xbar__EVAL_72),
    ._EVAL_73(out_xbar__EVAL_73),
    ._EVAL_74(out_xbar__EVAL_74),
    ._EVAL_75(out_xbar__EVAL_75),
    ._EVAL_76(out_xbar__EVAL_76),
    ._EVAL_77(out_xbar__EVAL_77),
    ._EVAL_78(out_xbar__EVAL_78),
    ._EVAL_79(out_xbar__EVAL_79),
    ._EVAL_80(out_xbar__EVAL_80),
    ._EVAL_81(out_xbar__EVAL_81),
    ._EVAL_82(out_xbar__EVAL_82),
    ._EVAL_83(out_xbar__EVAL_83),
    ._EVAL_84(out_xbar__EVAL_84),
    ._EVAL_85(out_xbar__EVAL_85),
    ._EVAL_86(out_xbar__EVAL_86),
    ._EVAL_87(out_xbar__EVAL_87),
    ._EVAL_88(out_xbar__EVAL_88),
    ._EVAL_89(out_xbar__EVAL_89),
    ._EVAL_90(out_xbar__EVAL_90),
    ._EVAL_91(out_xbar__EVAL_91),
    ._EVAL_92(out_xbar__EVAL_92),
    ._EVAL_93(out_xbar__EVAL_93),
    ._EVAL_94(out_xbar__EVAL_94),
    ._EVAL_95(out_xbar__EVAL_95),
    ._EVAL_96(out_xbar__EVAL_96),
    ._EVAL_97(out_xbar__EVAL_97),
    ._EVAL_98(out_xbar__EVAL_98),
    ._EVAL_99(out_xbar__EVAL_99),
    ._EVAL_100(out_xbar__EVAL_100),
    ._EVAL_101(out_xbar__EVAL_101),
    ._EVAL_102(out_xbar__EVAL_102),
    ._EVAL_103(out_xbar__EVAL_103),
    ._EVAL_104(out_xbar__EVAL_104),
    ._EVAL_105(out_xbar__EVAL_105),
    ._EVAL_106(out_xbar__EVAL_106),
    ._EVAL_107(out_xbar__EVAL_107),
    ._EVAL_108(out_xbar__EVAL_108),
    ._EVAL_109(out_xbar__EVAL_109),
    ._EVAL_110(out_xbar__EVAL_110),
    ._EVAL_111(out_xbar__EVAL_111),
    ._EVAL_112(out_xbar__EVAL_112),
    ._EVAL_113(out_xbar__EVAL_113),
    ._EVAL_114(out_xbar__EVAL_114),
    ._EVAL_115(out_xbar__EVAL_115),
    ._EVAL_116(out_xbar__EVAL_116),
    ._EVAL_117(out_xbar__EVAL_117),
    ._EVAL_118(out_xbar__EVAL_118),
    ._EVAL_119(out_xbar__EVAL_119),
    ._EVAL_120(out_xbar__EVAL_120),
    ._EVAL_121(out_xbar__EVAL_121),
    ._EVAL_122(out_xbar__EVAL_122),
    ._EVAL_123(out_xbar__EVAL_123),
    ._EVAL_124(out_xbar__EVAL_124),
    ._EVAL_125(out_xbar__EVAL_125),
    ._EVAL_126(out_xbar__EVAL_126),
    ._EVAL_127(out_xbar__EVAL_127),
    ._EVAL_128(out_xbar__EVAL_128),
    ._EVAL_129(out_xbar__EVAL_129),
    ._EVAL_130(out_xbar__EVAL_130),
    ._EVAL_131(out_xbar__EVAL_131),
    ._EVAL_132(out_xbar__EVAL_132),
    ._EVAL_133(out_xbar__EVAL_133),
    ._EVAL_134(out_xbar__EVAL_134),
    ._EVAL_135(out_xbar__EVAL_135),
    ._EVAL_136(out_xbar__EVAL_136),
    ._EVAL_137(out_xbar__EVAL_137),
    ._EVAL_138(out_xbar__EVAL_138),
    ._EVAL_139(out_xbar__EVAL_139),
    ._EVAL_140(out_xbar__EVAL_140),
    ._EVAL_141(out_xbar__EVAL_141)
  );
  SiFive__EVAL_141 coupler_to_debug (
    ._EVAL(coupler_to_debug__EVAL),
    ._EVAL_0(coupler_to_debug__EVAL_0),
    ._EVAL_1(coupler_to_debug__EVAL_1),
    ._EVAL_2(coupler_to_debug__EVAL_2),
    ._EVAL_3(coupler_to_debug__EVAL_3),
    ._EVAL_4(coupler_to_debug__EVAL_4),
    ._EVAL_5(coupler_to_debug__EVAL_5),
    ._EVAL_6(coupler_to_debug__EVAL_6),
    ._EVAL_7(coupler_to_debug__EVAL_7),
    ._EVAL_8(coupler_to_debug__EVAL_8),
    ._EVAL_9(coupler_to_debug__EVAL_9),
    ._EVAL_10(coupler_to_debug__EVAL_10),
    ._EVAL_11(coupler_to_debug__EVAL_11),
    ._EVAL_12(coupler_to_debug__EVAL_12),
    ._EVAL_13(coupler_to_debug__EVAL_13),
    ._EVAL_14(coupler_to_debug__EVAL_14),
    ._EVAL_15(coupler_to_debug__EVAL_15),
    ._EVAL_16(coupler_to_debug__EVAL_16),
    ._EVAL_17(coupler_to_debug__EVAL_17),
    ._EVAL_18(coupler_to_debug__EVAL_18),
    ._EVAL_19(coupler_to_debug__EVAL_19),
    ._EVAL_20(coupler_to_debug__EVAL_20),
    ._EVAL_21(coupler_to_debug__EVAL_21),
    ._EVAL_22(coupler_to_debug__EVAL_22),
    ._EVAL_23(coupler_to_debug__EVAL_23),
    ._EVAL_24(coupler_to_debug__EVAL_24),
    ._EVAL_25(coupler_to_debug__EVAL_25),
    ._EVAL_26(coupler_to_debug__EVAL_26),
    ._EVAL_27(coupler_to_debug__EVAL_27),
    ._EVAL_28(coupler_to_debug__EVAL_28),
    ._EVAL_29(coupler_to_debug__EVAL_29),
    ._EVAL_30(coupler_to_debug__EVAL_30),
    ._EVAL_31(coupler_to_debug__EVAL_31),
    ._EVAL_32(coupler_to_debug__EVAL_32)
  );
  SiFive__EVAL_114 in_xbar (
    ._EVAL(in_xbar__EVAL),
    ._EVAL_0(in_xbar__EVAL_0),
    ._EVAL_1(in_xbar__EVAL_1),
    ._EVAL_2(in_xbar__EVAL_2),
    ._EVAL_3(in_xbar__EVAL_3),
    ._EVAL_4(in_xbar__EVAL_4),
    ._EVAL_5(in_xbar__EVAL_5),
    ._EVAL_6(in_xbar__EVAL_6),
    ._EVAL_7(in_xbar__EVAL_7),
    ._EVAL_8(in_xbar__EVAL_8),
    ._EVAL_9(in_xbar__EVAL_9),
    ._EVAL_10(in_xbar__EVAL_10),
    ._EVAL_11(in_xbar__EVAL_11),
    ._EVAL_12(in_xbar__EVAL_12),
    ._EVAL_13(in_xbar__EVAL_13),
    ._EVAL_14(in_xbar__EVAL_14),
    ._EVAL_15(in_xbar__EVAL_15),
    ._EVAL_16(in_xbar__EVAL_16),
    ._EVAL_17(in_xbar__EVAL_17),
    ._EVAL_18(in_xbar__EVAL_18),
    ._EVAL_19(in_xbar__EVAL_19),
    ._EVAL_20(in_xbar__EVAL_20),
    ._EVAL_21(in_xbar__EVAL_21),
    ._EVAL_22(in_xbar__EVAL_22),
    ._EVAL_23(in_xbar__EVAL_23),
    ._EVAL_24(in_xbar__EVAL_24),
    ._EVAL_25(in_xbar__EVAL_25),
    ._EVAL_26(in_xbar__EVAL_26),
    ._EVAL_27(in_xbar__EVAL_27),
    ._EVAL_28(in_xbar__EVAL_28),
    ._EVAL_29(in_xbar__EVAL_29),
    ._EVAL_30(in_xbar__EVAL_30),
    ._EVAL_31(in_xbar__EVAL_31),
    ._EVAL_32(in_xbar__EVAL_32),
    ._EVAL_33(in_xbar__EVAL_33),
    ._EVAL_34(in_xbar__EVAL_34),
    ._EVAL_35(in_xbar__EVAL_35),
    ._EVAL_36(in_xbar__EVAL_36),
    ._EVAL_37(in_xbar__EVAL_37),
    ._EVAL_38(in_xbar__EVAL_38),
    ._EVAL_39(in_xbar__EVAL_39),
    ._EVAL_40(in_xbar__EVAL_40)
  );
  SiFive__EVAL_120 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40)
  );
  SiFive__EVAL_179 buffer_1 (
    ._EVAL(buffer_1__EVAL),
    ._EVAL_0(buffer_1__EVAL_0),
    ._EVAL_1(buffer_1__EVAL_1),
    ._EVAL_2(buffer_1__EVAL_2),
    ._EVAL_3(buffer_1__EVAL_3),
    ._EVAL_4(buffer_1__EVAL_4),
    ._EVAL_5(buffer_1__EVAL_5),
    ._EVAL_6(buffer_1__EVAL_6),
    ._EVAL_7(buffer_1__EVAL_7),
    ._EVAL_8(buffer_1__EVAL_8),
    ._EVAL_9(buffer_1__EVAL_9),
    ._EVAL_10(buffer_1__EVAL_10),
    ._EVAL_11(buffer_1__EVAL_11),
    ._EVAL_12(buffer_1__EVAL_12),
    ._EVAL_13(buffer_1__EVAL_13),
    ._EVAL_14(buffer_1__EVAL_14),
    ._EVAL_15(buffer_1__EVAL_15),
    ._EVAL_16(buffer_1__EVAL_16),
    ._EVAL_17(buffer_1__EVAL_17),
    ._EVAL_18(buffer_1__EVAL_18),
    ._EVAL_19(buffer_1__EVAL_19),
    ._EVAL_20(buffer_1__EVAL_20),
    ._EVAL_21(buffer_1__EVAL_21),
    ._EVAL_22(buffer_1__EVAL_22),
    ._EVAL_23(buffer_1__EVAL_23),
    ._EVAL_24(buffer_1__EVAL_24),
    ._EVAL_25(buffer_1__EVAL_25),
    ._EVAL_26(buffer_1__EVAL_26),
    ._EVAL_27(buffer_1__EVAL_27),
    ._EVAL_28(buffer_1__EVAL_28),
    ._EVAL_29(buffer_1__EVAL_29),
    ._EVAL_30(buffer_1__EVAL_30),
    ._EVAL_31(buffer_1__EVAL_31),
    ._EVAL_32(buffer_1__EVAL_32),
    ._EVAL_33(buffer_1__EVAL_33),
    ._EVAL_34(buffer_1__EVAL_34),
    ._EVAL_35(buffer_1__EVAL_35),
    ._EVAL_36(buffer_1__EVAL_36),
    ._EVAL_37(buffer_1__EVAL_37),
    ._EVAL_38(buffer_1__EVAL_38),
    ._EVAL_39(buffer_1__EVAL_39),
    ._EVAL_40(buffer_1__EVAL_40)
  );
  SiFive__EVAL_152 coupler_to_tile_with_no_name (
    ._EVAL(coupler_to_tile_with_no_name__EVAL),
    ._EVAL_0(coupler_to_tile_with_no_name__EVAL_0),
    ._EVAL_1(coupler_to_tile_with_no_name__EVAL_1),
    ._EVAL_2(coupler_to_tile_with_no_name__EVAL_2),
    ._EVAL_3(coupler_to_tile_with_no_name__EVAL_3),
    ._EVAL_4(coupler_to_tile_with_no_name__EVAL_4),
    ._EVAL_5(coupler_to_tile_with_no_name__EVAL_5),
    ._EVAL_6(coupler_to_tile_with_no_name__EVAL_6),
    ._EVAL_7(coupler_to_tile_with_no_name__EVAL_7),
    ._EVAL_8(coupler_to_tile_with_no_name__EVAL_8),
    ._EVAL_9(coupler_to_tile_with_no_name__EVAL_9),
    ._EVAL_10(coupler_to_tile_with_no_name__EVAL_10),
    ._EVAL_11(coupler_to_tile_with_no_name__EVAL_11),
    ._EVAL_12(coupler_to_tile_with_no_name__EVAL_12),
    ._EVAL_13(coupler_to_tile_with_no_name__EVAL_13),
    ._EVAL_14(coupler_to_tile_with_no_name__EVAL_14),
    ._EVAL_15(coupler_to_tile_with_no_name__EVAL_15),
    ._EVAL_16(coupler_to_tile_with_no_name__EVAL_16),
    ._EVAL_17(coupler_to_tile_with_no_name__EVAL_17),
    ._EVAL_18(coupler_to_tile_with_no_name__EVAL_18),
    ._EVAL_19(coupler_to_tile_with_no_name__EVAL_19),
    ._EVAL_20(coupler_to_tile_with_no_name__EVAL_20),
    ._EVAL_21(coupler_to_tile_with_no_name__EVAL_21),
    ._EVAL_22(coupler_to_tile_with_no_name__EVAL_22),
    ._EVAL_23(coupler_to_tile_with_no_name__EVAL_23),
    ._EVAL_24(coupler_to_tile_with_no_name__EVAL_24),
    ._EVAL_25(coupler_to_tile_with_no_name__EVAL_25),
    ._EVAL_26(coupler_to_tile_with_no_name__EVAL_26),
    ._EVAL_27(coupler_to_tile_with_no_name__EVAL_27),
    ._EVAL_28(coupler_to_tile_with_no_name__EVAL_28),
    ._EVAL_29(coupler_to_tile_with_no_name__EVAL_29),
    ._EVAL_30(coupler_to_tile_with_no_name__EVAL_30),
    ._EVAL_31(coupler_to_tile_with_no_name__EVAL_31),
    ._EVAL_32(coupler_to_tile_with_no_name__EVAL_32),
    ._EVAL_33(coupler_to_tile_with_no_name__EVAL_33),
    ._EVAL_34(coupler_to_tile_with_no_name__EVAL_34),
    ._EVAL_35(coupler_to_tile_with_no_name__EVAL_35),
    ._EVAL_36(coupler_to_tile_with_no_name__EVAL_36),
    ._EVAL_37(coupler_to_tile_with_no_name__EVAL_37),
    ._EVAL_38(coupler_to_tile_with_no_name__EVAL_38),
    ._EVAL_39(coupler_to_tile_with_no_name__EVAL_39),
    ._EVAL_40(coupler_to_tile_with_no_name__EVAL_40),
    ._EVAL_41(coupler_to_tile_with_no_name__EVAL_41),
    ._EVAL_42(coupler_to_tile_with_no_name__EVAL_42),
    ._EVAL_43(coupler_to_tile_with_no_name__EVAL_43),
    ._EVAL_44(coupler_to_tile_with_no_name__EVAL_44),
    ._EVAL_45(coupler_to_tile_with_no_name__EVAL_45),
    ._EVAL_46(coupler_to_tile_with_no_name__EVAL_46),
    ._EVAL_47(coupler_to_tile_with_no_name__EVAL_47),
    ._EVAL_48(coupler_to_tile_with_no_name__EVAL_48),
    ._EVAL_49(coupler_to_tile_with_no_name__EVAL_49),
    ._EVAL_50(coupler_to_tile_with_no_name__EVAL_50),
    ._EVAL_51(coupler_to_tile_with_no_name__EVAL_51),
    ._EVAL_52(coupler_to_tile_with_no_name__EVAL_52),
    ._EVAL_53(coupler_to_tile_with_no_name__EVAL_53),
    ._EVAL_54(coupler_to_tile_with_no_name__EVAL_54),
    ._EVAL_55(coupler_to_tile_with_no_name__EVAL_55),
    ._EVAL_56(coupler_to_tile_with_no_name__EVAL_56),
    ._EVAL_57(coupler_to_tile_with_no_name__EVAL_57),
    ._EVAL_58(coupler_to_tile_with_no_name__EVAL_58),
    ._EVAL_59(coupler_to_tile_with_no_name__EVAL_59),
    ._EVAL_60(coupler_to_tile_with_no_name__EVAL_60)
  );
  SiFive__EVAL_129 wrapped_error_device (
    ._EVAL(wrapped_error_device__EVAL),
    ._EVAL_0(wrapped_error_device__EVAL_0),
    ._EVAL_1(wrapped_error_device__EVAL_1),
    ._EVAL_2(wrapped_error_device__EVAL_2),
    ._EVAL_3(wrapped_error_device__EVAL_3),
    ._EVAL_4(wrapped_error_device__EVAL_4),
    ._EVAL_5(wrapped_error_device__EVAL_5),
    ._EVAL_6(wrapped_error_device__EVAL_6),
    ._EVAL_7(wrapped_error_device__EVAL_7),
    ._EVAL_8(wrapped_error_device__EVAL_8),
    ._EVAL_9(wrapped_error_device__EVAL_9),
    ._EVAL_10(wrapped_error_device__EVAL_10),
    ._EVAL_11(wrapped_error_device__EVAL_11),
    ._EVAL_12(wrapped_error_device__EVAL_12),
    ._EVAL_13(wrapped_error_device__EVAL_13),
    ._EVAL_14(wrapped_error_device__EVAL_14),
    ._EVAL_15(wrapped_error_device__EVAL_15),
    ._EVAL_16(wrapped_error_device__EVAL_16),
    ._EVAL_17(wrapped_error_device__EVAL_17),
    ._EVAL_18(wrapped_error_device__EVAL_18),
    ._EVAL_19(wrapped_error_device__EVAL_19)
  );
  SiFive__EVAL_112 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40)
  );
  SiFive__EVAL_158 coupler_to_testindicator (
    ._EVAL(coupler_to_testindicator__EVAL),
    ._EVAL_0(coupler_to_testindicator__EVAL_0),
    ._EVAL_1(coupler_to_testindicator__EVAL_1),
    ._EVAL_2(coupler_to_testindicator__EVAL_2),
    ._EVAL_3(coupler_to_testindicator__EVAL_3),
    ._EVAL_4(coupler_to_testindicator__EVAL_4),
    ._EVAL_5(coupler_to_testindicator__EVAL_5),
    ._EVAL_6(coupler_to_testindicator__EVAL_6),
    ._EVAL_7(coupler_to_testindicator__EVAL_7),
    ._EVAL_8(coupler_to_testindicator__EVAL_8),
    ._EVAL_9(coupler_to_testindicator__EVAL_9),
    ._EVAL_10(coupler_to_testindicator__EVAL_10),
    ._EVAL_11(coupler_to_testindicator__EVAL_11),
    ._EVAL_12(coupler_to_testindicator__EVAL_12),
    ._EVAL_13(coupler_to_testindicator__EVAL_13),
    ._EVAL_14(coupler_to_testindicator__EVAL_14),
    ._EVAL_15(coupler_to_testindicator__EVAL_15),
    ._EVAL_16(coupler_to_testindicator__EVAL_16),
    ._EVAL_17(coupler_to_testindicator__EVAL_17),
    ._EVAL_18(coupler_to_testindicator__EVAL_18),
    ._EVAL_19(coupler_to_testindicator__EVAL_19),
    ._EVAL_20(coupler_to_testindicator__EVAL_20),
    ._EVAL_21(coupler_to_testindicator__EVAL_21),
    ._EVAL_22(coupler_to_testindicator__EVAL_22),
    ._EVAL_23(coupler_to_testindicator__EVAL_23),
    ._EVAL_24(coupler_to_testindicator__EVAL_24),
    ._EVAL_25(coupler_to_testindicator__EVAL_25),
    ._EVAL_26(coupler_to_testindicator__EVAL_26),
    ._EVAL_27(coupler_to_testindicator__EVAL_27),
    ._EVAL_28(coupler_to_testindicator__EVAL_28),
    ._EVAL_29(coupler_to_testindicator__EVAL_29),
    ._EVAL_30(coupler_to_testindicator__EVAL_30),
    ._EVAL_31(coupler_to_testindicator__EVAL_31),
    ._EVAL_32(coupler_to_testindicator__EVAL_32)
  );
  SiFive__EVAL_137 coupler_to_clint (
    ._EVAL(coupler_to_clint__EVAL),
    ._EVAL_0(coupler_to_clint__EVAL_0),
    ._EVAL_1(coupler_to_clint__EVAL_1),
    ._EVAL_2(coupler_to_clint__EVAL_2),
    ._EVAL_3(coupler_to_clint__EVAL_3),
    ._EVAL_4(coupler_to_clint__EVAL_4),
    ._EVAL_5(coupler_to_clint__EVAL_5),
    ._EVAL_6(coupler_to_clint__EVAL_6),
    ._EVAL_7(coupler_to_clint__EVAL_7),
    ._EVAL_8(coupler_to_clint__EVAL_8),
    ._EVAL_9(coupler_to_clint__EVAL_9),
    ._EVAL_10(coupler_to_clint__EVAL_10),
    ._EVAL_11(coupler_to_clint__EVAL_11),
    ._EVAL_12(coupler_to_clint__EVAL_12),
    ._EVAL_13(coupler_to_clint__EVAL_13),
    ._EVAL_14(coupler_to_clint__EVAL_14),
    ._EVAL_15(coupler_to_clint__EVAL_15),
    ._EVAL_16(coupler_to_clint__EVAL_16),
    ._EVAL_17(coupler_to_clint__EVAL_17),
    ._EVAL_18(coupler_to_clint__EVAL_18),
    ._EVAL_19(coupler_to_clint__EVAL_19),
    ._EVAL_20(coupler_to_clint__EVAL_20),
    ._EVAL_21(coupler_to_clint__EVAL_21),
    ._EVAL_22(coupler_to_clint__EVAL_22),
    ._EVAL_23(coupler_to_clint__EVAL_23),
    ._EVAL_24(coupler_to_clint__EVAL_24),
    ._EVAL_25(coupler_to_clint__EVAL_25),
    ._EVAL_26(coupler_to_clint__EVAL_26),
    ._EVAL_27(coupler_to_clint__EVAL_27),
    ._EVAL_28(coupler_to_clint__EVAL_28),
    ._EVAL_29(coupler_to_clint__EVAL_29),
    ._EVAL_30(coupler_to_clint__EVAL_30),
    ._EVAL_31(coupler_to_clint__EVAL_31),
    ._EVAL_32(coupler_to_clint__EVAL_32)
  );
  SiFive__EVAL_133 coupler_to_plic (
    ._EVAL(coupler_to_plic__EVAL),
    ._EVAL_0(coupler_to_plic__EVAL_0),
    ._EVAL_1(coupler_to_plic__EVAL_1),
    ._EVAL_2(coupler_to_plic__EVAL_2),
    ._EVAL_3(coupler_to_plic__EVAL_3),
    ._EVAL_4(coupler_to_plic__EVAL_4),
    ._EVAL_5(coupler_to_plic__EVAL_5),
    ._EVAL_6(coupler_to_plic__EVAL_6),
    ._EVAL_7(coupler_to_plic__EVAL_7),
    ._EVAL_8(coupler_to_plic__EVAL_8),
    ._EVAL_9(coupler_to_plic__EVAL_9),
    ._EVAL_10(coupler_to_plic__EVAL_10),
    ._EVAL_11(coupler_to_plic__EVAL_11),
    ._EVAL_12(coupler_to_plic__EVAL_12),
    ._EVAL_13(coupler_to_plic__EVAL_13),
    ._EVAL_14(coupler_to_plic__EVAL_14),
    ._EVAL_15(coupler_to_plic__EVAL_15),
    ._EVAL_16(coupler_to_plic__EVAL_16),
    ._EVAL_17(coupler_to_plic__EVAL_17),
    ._EVAL_18(coupler_to_plic__EVAL_18),
    ._EVAL_19(coupler_to_plic__EVAL_19),
    ._EVAL_20(coupler_to_plic__EVAL_20),
    ._EVAL_21(coupler_to_plic__EVAL_21),
    ._EVAL_22(coupler_to_plic__EVAL_22),
    ._EVAL_23(coupler_to_plic__EVAL_23),
    ._EVAL_24(coupler_to_plic__EVAL_24),
    ._EVAL_25(coupler_to_plic__EVAL_25),
    ._EVAL_26(coupler_to_plic__EVAL_26),
    ._EVAL_27(coupler_to_plic__EVAL_27),
    ._EVAL_28(coupler_to_plic__EVAL_28),
    ._EVAL_29(coupler_to_plic__EVAL_29),
    ._EVAL_30(coupler_to_plic__EVAL_30),
    ._EVAL_31(coupler_to_plic__EVAL_31),
    ._EVAL_32(coupler_to_plic__EVAL_32)
  );
  SiFive__EVAL_122 atomics (
    ._EVAL(atomics__EVAL),
    ._EVAL_0(atomics__EVAL_0),
    ._EVAL_1(atomics__EVAL_1),
    ._EVAL_2(atomics__EVAL_2),
    ._EVAL_3(atomics__EVAL_3),
    ._EVAL_4(atomics__EVAL_4),
    ._EVAL_5(atomics__EVAL_5),
    ._EVAL_6(atomics__EVAL_6),
    ._EVAL_7(atomics__EVAL_7),
    ._EVAL_8(atomics__EVAL_8),
    ._EVAL_9(atomics__EVAL_9),
    ._EVAL_10(atomics__EVAL_10),
    ._EVAL_11(atomics__EVAL_11),
    ._EVAL_12(atomics__EVAL_12),
    ._EVAL_13(atomics__EVAL_13),
    ._EVAL_14(atomics__EVAL_14),
    ._EVAL_15(atomics__EVAL_15),
    ._EVAL_16(atomics__EVAL_16),
    ._EVAL_17(atomics__EVAL_17),
    ._EVAL_18(atomics__EVAL_18),
    ._EVAL_19(atomics__EVAL_19),
    ._EVAL_20(atomics__EVAL_20),
    ._EVAL_21(atomics__EVAL_21),
    ._EVAL_22(atomics__EVAL_22),
    ._EVAL_23(atomics__EVAL_23),
    ._EVAL_24(atomics__EVAL_24),
    ._EVAL_25(atomics__EVAL_25),
    ._EVAL_26(atomics__EVAL_26),
    ._EVAL_27(atomics__EVAL_27),
    ._EVAL_28(atomics__EVAL_28),
    ._EVAL_29(atomics__EVAL_29),
    ._EVAL_30(atomics__EVAL_30),
    ._EVAL_31(atomics__EVAL_31),
    ._EVAL_32(atomics__EVAL_32),
    ._EVAL_33(atomics__EVAL_33),
    ._EVAL_34(atomics__EVAL_34),
    ._EVAL_35(atomics__EVAL_35),
    ._EVAL_36(atomics__EVAL_36),
    ._EVAL_37(atomics__EVAL_37),
    ._EVAL_38(atomics__EVAL_38),
    ._EVAL_39(atomics__EVAL_39),
    ._EVAL_40(atomics__EVAL_40)
  );
  assign coupler_to_tile_with_no_name__EVAL_37 = _EVAL_25;
  assign buffer__EVAL_38 = atomics__EVAL_18;
  assign _EVAL_118 = buffer_1__EVAL_3;
  assign out_xbar__EVAL_127 = fixer__EVAL_28;
  assign coupler_to_port_named_axi4_periph_port__EVAL_29 = _EVAL_82;
  assign _EVAL_112 = coupler_to_debug__EVAL_18;
  assign _EVAL_39 = coupler_to_testindicator__EVAL_31;
  assign _EVAL_81 = coupler_to_debug__EVAL_5;
  assign _EVAL_43 = coupler_to_port_named_axi4_periph_port__EVAL_14;
  assign in_xbar__EVAL_19 = buffer_1__EVAL_9;
  assign _EVAL_74 = coupler_to_tile_with_no_name__EVAL_48;
  assign out_xbar__EVAL_81 = coupler_to_plic__EVAL_27;
  assign _EVAL_48 = buffer_1__EVAL_5;
  assign buffer__EVAL_5 = fixer__EVAL_38;
  assign _EVAL_34 = coupler_to_port_named_axi4_periph_port__EVAL_43;
  assign in_xbar__EVAL_36 = buffer_1__EVAL_40;
  assign fixer__EVAL_9 = buffer__EVAL_2;
  assign coupler_to_port_named_axi4_periph_port__EVAL_53 = _EVAL_116;
  assign coupler_to_plic__EVAL_23 = out_xbar__EVAL;
  assign coupler_to_debug__EVAL_7 = out_xbar__EVAL_112;
  assign _EVAL_93 = coupler_to_port_named_axi4_periph_port__EVAL_11;
  assign fixer__EVAL_31 = buffer__EVAL_37;
  assign _EVAL_111 = coupler_to_tile_with_no_name__EVAL_20;
  assign out_xbar__EVAL_70 = coupler_to_testindicator__EVAL_23;
  assign coupler_to_testindicator__EVAL_16 = out_xbar__EVAL_55;
  assign atomics__EVAL_23 = in_xbar__EVAL_24;
  assign _EVAL_151 = coupler_to_plic__EVAL_9;
  assign _EVAL_87 = coupler_to_tile_with_no_name__EVAL_58;
  assign coupler_to_port_named_axi4_periph_port__EVAL_26 = _EVAL_12;
  assign _EVAL_10 = buffer_1__EVAL_4;
  assign _EVAL_135 = coupler_to_clint__EVAL_12;
  assign coupler_to_plic__EVAL_0 = _EVAL_90;
  assign _EVAL_148 = coupler_to_port_named_axi4_periph_port__EVAL_13;
  assign buffer_1__EVAL_35 = _EVAL_102;
  assign coupler_to_tile_with_no_name__EVAL_18 = _EVAL_105;
  assign _EVAL_114 = coupler_to_clint__EVAL;
  assign out_xbar__EVAL_116 = coupler_to_port_named_axi4_periph_port__EVAL_24;
  assign _EVAL_26 = coupler_to_tile_with_no_name__EVAL;
  assign buffer_1__EVAL_18 = in_xbar__EVAL_7;
  assign out_xbar__EVAL_133 = fixer__EVAL_19;
  assign buffer__EVAL_15 = atomics__EVAL_10;
  assign _EVAL_70 = coupler_to_tile_with_no_name__EVAL_44;
  assign _EVAL_71 = buffer_1__EVAL_24;
  assign coupler_to_clint__EVAL_20 = out_xbar__EVAL_93;
  assign fixer__EVAL_1 = out_xbar__EVAL_88;
  assign coupler_to_debug__EVAL_14 = _EVAL_141;
  assign coupler_to_tile_with_no_name__EVAL_35 = out_xbar__EVAL_83;
  assign coupler_to_tile_with_no_name__EVAL_22 = _EVAL_82;
  assign fixer__EVAL_14 = buffer__EVAL_12;
  assign coupler_to_plic__EVAL = out_xbar__EVAL_43;
  assign coupler_to_tile_with_no_name__EVAL_45 = _EVAL_42;
  assign out_xbar__EVAL_33 = coupler_to_debug__EVAL_9;
  assign out_xbar__EVAL_102 = coupler_to_plic__EVAL_20;
  assign buffer_1__EVAL_25 = in_xbar__EVAL_21;
  assign fixer__EVAL_5 = out_xbar__EVAL_14;
  assign _EVAL_56 = coupler_to_port_named_axi4_periph_port__EVAL_36;
  assign coupler_to_port_named_axi4_periph_port__EVAL_34 = _EVAL_57;
  assign _EVAL_119 = buffer_1__EVAL_12;
  assign _EVAL_79 = coupler_to_port_named_axi4_periph_port__EVAL_35;
  assign coupler_to_tile_with_no_name__EVAL_6 = _EVAL_30;
  assign out_xbar__EVAL_92 = coupler_to_port_named_axi4_periph_port__EVAL_20;
  assign out_xbar__EVAL_129 = coupler_to_plic__EVAL_29;
  assign buffer_1__EVAL_7 = in_xbar__EVAL_35;
  assign coupler_to_plic__EVAL_2 = _EVAL_54;
  assign coupler_to_port_named_axi4_periph_port__EVAL_17 = out_xbar__EVAL_50;
  assign coupler_to_testindicator__EVAL_4 = _EVAL_90;
  assign in_xbar__EVAL_12 = atomics__EVAL_24;
  assign coupler_to_debug__EVAL_8 = _EVAL_8;
  assign _EVAL_154 = coupler_to_debug__EVAL_29;
  assign _EVAL_97 = coupler_to_plic__EVAL_6;
  assign _EVAL_115 = buffer_1__EVAL_30;
  assign coupler_to_testindicator__EVAL_20 = _EVAL_147;
  assign coupler_to_debug__EVAL_26 = out_xbar__EVAL_130;
  assign _EVAL_99 = coupler_to_port_named_axi4_periph_port__EVAL_18;
  assign atomics__EVAL_21 = in_xbar__EVAL_18;
  assign in_xbar__EVAL_15 = buffer_1__EVAL_19;
  assign coupler_to_tile_with_no_name__EVAL_3 = _EVAL_31;
  assign coupler_to_plic__EVAL_28 = out_xbar__EVAL_119;
  assign coupler_to_clint__EVAL_32 = out_xbar__EVAL_104;
  assign coupler_to_clint__EVAL_16 = out_xbar__EVAL_54;
  assign _EVAL_4 = coupler_to_plic__EVAL_14;
  assign coupler_to_plic__EVAL_7 = out_xbar__EVAL_111;
  assign coupler_to_tile_with_no_name__EVAL_24 = _EVAL_29;
  assign in_xbar__EVAL_5 = buffer_1__EVAL_28;
  assign _EVAL_36 = coupler_to_port_named_axi4_periph_port__EVAL_16;
  assign coupler_to_port_named_axi4_periph_port__EVAL_37 = out_xbar__EVAL_38;
  assign wrapped_error_device__EVAL_19 = out_xbar__EVAL_114;
  assign buffer_1__EVAL_8 = in_xbar__EVAL_25;
  assign coupler_to_clint__EVAL_29 = _EVAL_77;
  assign buffer_1__EVAL = _EVAL_45;
  assign _EVAL_40 = coupler_to_tile_with_no_name__EVAL_51;
  assign coupler_to_port_named_axi4_periph_port__EVAL = out_xbar__EVAL_95;
  assign in_xbar__EVAL_29 = atomics__EVAL_9;
  assign wrapped_error_device__EVAL_10 = _EVAL_90;
  assign in_xbar__EVAL_10 = atomics__EVAL_31;
  assign coupler_to_port_named_axi4_periph_port__EVAL_42 = out_xbar__EVAL_140;
  assign buffer__EVAL_29 = fixer__EVAL_36;
  assign buffer__EVAL_3 = atomics__EVAL_15;
  assign in_xbar__EVAL_3 = atomics__EVAL_19;
  assign out_xbar__EVAL_73 = coupler_to_port_named_axi4_periph_port__EVAL_0;
  assign buffer_1__EVAL_2 = in_xbar__EVAL_31;
  assign atomics__EVAL_1 = _EVAL_90;
  assign _EVAL_2 = coupler_to_tile_with_no_name__EVAL_19;
  assign coupler_to_tile_with_no_name__EVAL_2 = _EVAL_67;
  assign atomics__EVAL_2 = in_xbar__EVAL_33;
  assign in_xbar__EVAL_34 = atomics__EVAL_34;
  assign _EVAL_47 = coupler_to_port_named_axi4_periph_port__EVAL_1;
  assign in_xbar__EVAL_40 = atomics__EVAL_30;
  assign _EVAL_143 = coupler_to_port_named_axi4_periph_port__EVAL_19;
  assign _EVAL_152 = coupler_to_plic__EVAL_32;
  assign _EVAL_14 = coupler_to_tile_with_no_name__EVAL_26;
  assign _EVAL_60 = coupler_to_debug__EVAL_17;
  assign fixer__EVAL_4 = buffer__EVAL_9;
  assign buffer__EVAL_1 = fixer__EVAL_30;
  assign atomics__EVAL_14 = in_xbar__EVAL_27;
  assign coupler_to_testindicator__EVAL_14 = out_xbar__EVAL_86;
  assign out_xbar__EVAL_66 = wrapped_error_device__EVAL_6;
  assign in_xbar__EVAL_22 = _EVAL_90;
  assign coupler_to_tile_with_no_name__EVAL_10 = _EVAL_52;
  assign in_xbar__EVAL_37 = buffer_1__EVAL_22;
  assign out_xbar__EVAL_138 = coupler_to_testindicator__EVAL_18;
  assign in_xbar__EVAL_30 = buffer_1__EVAL_37;
  assign buffer_1__EVAL_36 = _EVAL_117;
  assign _EVAL_156 = coupler_to_tile_with_no_name__EVAL_27;
  assign _EVAL_55 = coupler_to_clint__EVAL_7;
  assign coupler_to_testindicator__EVAL_28 = out_xbar__EVAL_120;
  assign coupler_to_tile_with_no_name__EVAL_13 = _EVAL_89;
  assign fixer__EVAL_23 = out_xbar__EVAL_100;
  assign out_xbar__EVAL_72 = coupler_to_tile_with_no_name__EVAL_23;
  assign _EVAL_101 = coupler_to_tile_with_no_name__EVAL_21;
  assign atomics__EVAL_12 = buffer__EVAL_16;
  assign _EVAL_76 = coupler_to_port_named_axi4_periph_port__EVAL_25;
  assign coupler_to_plic__EVAL_1 = out_xbar__EVAL_78;
  assign atomics__EVAL_17 = buffer__EVAL_14;
  assign atomics__EVAL_27 = in_xbar__EVAL_4;
  assign buffer__EVAL_31 = _EVAL_90;
  assign out_xbar__EVAL_17 = coupler_to_clint__EVAL_6;
  assign buffer__EVAL_7 = atomics__EVAL;
  assign _EVAL_158 = coupler_to_port_named_axi4_periph_port__EVAL_22;
  assign in_xbar__EVAL_39 = atomics__EVAL_16;
  assign wrapped_error_device__EVAL_5 = out_xbar__EVAL_71;
  assign out_xbar__EVAL_49 = _EVAL_82;
  assign _EVAL_123 = coupler_to_testindicator__EVAL_12;
  assign _EVAL_65 = coupler_to_debug__EVAL_27;
  assign coupler_to_debug__EVAL_10 = _EVAL_86;
  assign coupler_to_testindicator__EVAL_11 = _EVAL_138;
  assign _EVAL_100 = coupler_to_port_named_axi4_periph_port__EVAL_44;
  assign in_xbar__EVAL_14 = _EVAL_82;
  assign out_xbar__EVAL_11 = coupler_to_debug__EVAL_20;
  assign fixer__EVAL_39 = out_xbar__EVAL_57;
  assign coupler_to_testindicator__EVAL_22 = _EVAL_122;
  assign coupler_to_testindicator__EVAL_3 = out_xbar__EVAL_97;
  assign _EVAL_126 = coupler_to_testindicator__EVAL_15;
  assign in_xbar__EVAL_11 = buffer_1__EVAL_21;
  assign buffer__EVAL_24 = atomics__EVAL_4;
  assign out_xbar__EVAL_3 = coupler_to_plic__EVAL_17;
  assign buffer__EVAL_17 = atomics__EVAL_11;
  assign _EVAL_6 = coupler_to_testindicator__EVAL_19;
  assign _EVAL_5 = coupler_to_testindicator__EVAL_26;
  assign coupler_to_testindicator__EVAL_7 = out_xbar__EVAL_59;
  assign coupler_to_port_named_axi4_periph_port__EVAL_3 = _EVAL_44;
  assign out_xbar__EVAL_60 = wrapped_error_device__EVAL_12;
  assign out_xbar__EVAL_106 = coupler_to_debug__EVAL_2;
  assign atomics__EVAL_3 = buffer__EVAL_39;
  assign out_xbar__EVAL_31 = coupler_to_tile_with_no_name__EVAL_1;
  assign coupler_to_tile_with_no_name__EVAL_9 = _EVAL_0;
  assign coupler_to_plic__EVAL_24 = out_xbar__EVAL_69;
  assign coupler_to_debug__EVAL_28 = _EVAL_145;
  assign _EVAL_9 = coupler_to_plic__EVAL_11;
  assign _EVAL = coupler_to_debug__EVAL_13;
  assign _EVAL_38 = coupler_to_testindicator__EVAL;
  assign out_xbar__EVAL_15 = wrapped_error_device__EVAL_14;
  assign fixer__EVAL_2 = out_xbar__EVAL_105;
  assign out_xbar__EVAL_27 = coupler_to_tile_with_no_name__EVAL_29;
  assign atomics__EVAL_13 = in_xbar__EVAL_2;
  assign _EVAL_22 = coupler_to_debug__EVAL_6;
  assign in_xbar__EVAL_1 = atomics__EVAL_5;
  assign _EVAL_46 = coupler_to_debug__EVAL_21;
  assign coupler_to_tile_with_no_name__EVAL_46 = _EVAL_62;
  assign coupler_to_testindicator__EVAL_32 = out_xbar__EVAL_125;
  assign coupler_to_tile_with_no_name__EVAL_43 = _EVAL_51;
  assign coupler_to_plic__EVAL_4 = _EVAL_85;
  assign buffer_1__EVAL_29 = _EVAL_15;
  assign out_xbar__EVAL_123 = coupler_to_tile_with_no_name__EVAL_30;
  assign _EVAL_17 = coupler_to_plic__EVAL_21;
  assign coupler_to_port_named_axi4_periph_port__EVAL_41 = out_xbar__EVAL_118;
  assign coupler_to_testindicator__EVAL_17 = out_xbar__EVAL_41;
  assign wrapped_error_device__EVAL_16 = out_xbar__EVAL_68;
  assign buffer_1__EVAL_1 = in_xbar__EVAL_8;
  assign buffer__EVAL_25 = fixer__EVAL_25;
  assign atomics__EVAL_0 = buffer__EVAL_13;
  assign coupler_to_debug__EVAL_4 = out_xbar__EVAL_99;
  assign coupler_to_port_named_axi4_periph_port__EVAL_31 = out_xbar__EVAL_94;
  assign _EVAL_136 = coupler_to_clint__EVAL_11;
  assign out_xbar__EVAL_132 = coupler_to_tile_with_no_name__EVAL_32;
  assign _EVAL_78 = coupler_to_testindicator__EVAL_10;
  assign buffer__EVAL = fixer__EVAL_12;
  assign fixer__EVAL_22 = buffer__EVAL_19;
  assign coupler_to_tile_with_no_name__EVAL_53 = out_xbar__EVAL_37;
  assign coupler_to_plic__EVAL_15 = _EVAL_50;
  assign wrapped_error_device__EVAL_0 = out_xbar__EVAL_134;
  assign coupler_to_debug__EVAL_30 = out_xbar__EVAL_30;
  assign coupler_to_clint__EVAL_8 = _EVAL_82;
  assign wrapped_error_device__EVAL_17 = _EVAL_82;
  assign coupler_to_tile_with_no_name__EVAL_56 = _EVAL_90;
  assign atomics__EVAL_8 = _EVAL_82;
  assign out_xbar__EVAL_1 = coupler_to_tile_with_no_name__EVAL_59;
  assign coupler_to_port_named_axi4_periph_port__EVAL_45 = _EVAL_128;
  assign _EVAL_150 = coupler_to_port_named_axi4_periph_port__EVAL_50;
  assign out_xbar__EVAL_63 = coupler_to_port_named_axi4_periph_port__EVAL_52;
  assign _EVAL_75 = coupler_to_debug__EVAL_1;
  assign out_xbar__EVAL_108 = coupler_to_debug__EVAL_12;
  assign atomics__EVAL_20 = buffer__EVAL_36;
  assign out_xbar__EVAL_46 = coupler_to_tile_with_no_name__EVAL_5;
  assign coupler_to_tile_with_no_name__EVAL_33 = out_xbar__EVAL_136;
  assign buffer__EVAL_26 = fixer__EVAL_35;
  assign coupler_to_debug__EVAL_23 = out_xbar__EVAL_65;
  assign fixer__EVAL_15 = out_xbar__EVAL_89;
  assign _EVAL_108 = coupler_to_tile_with_no_name__EVAL_38;
  assign out_xbar__EVAL_44 = wrapped_error_device__EVAL_1;
  assign coupler_to_tile_with_no_name__EVAL_41 = out_xbar__EVAL_109;
  assign buffer_1__EVAL_10 = _EVAL_140;
  assign coupler_to_clint__EVAL_24 = out_xbar__EVAL_124;
  assign out_xbar__EVAL_19 = wrapped_error_device__EVAL;
  assign _EVAL_61 = coupler_to_clint__EVAL_5;
  assign out_xbar__EVAL_82 = coupler_to_tile_with_no_name__EVAL_49;
  assign coupler_to_tile_with_no_name__EVAL_16 = _EVAL_153;
  assign coupler_to_tile_with_no_name__EVAL_40 = out_xbar__EVAL_36;
  assign fixer__EVAL_3 = buffer__EVAL_8;
  assign coupler_to_plic__EVAL_13 = out_xbar__EVAL_103;
  assign fixer__EVAL_11 = _EVAL_90;
  assign coupler_to_debug__EVAL_3 = out_xbar__EVAL_126;
  assign coupler_to_clint__EVAL_4 = _EVAL_33;
  assign coupler_to_clint__EVAL_13 = out_xbar__EVAL_98;
  assign out_xbar__EVAL_139 = coupler_to_port_named_axi4_periph_port__EVAL_39;
  assign coupler_to_testindicator__EVAL_13 = _EVAL_146;
  assign out_xbar__EVAL_5 = coupler_to_plic__EVAL_19;
  assign fixer__EVAL_0 = _EVAL_82;
  assign coupler_to_tile_with_no_name__EVAL_60 = _EVAL_121;
  assign out_xbar__EVAL_107 = coupler_to_debug__EVAL_31;
  assign buffer_1__EVAL_31 = _EVAL_23;
  assign out_xbar__EVAL_76 = coupler_to_tile_with_no_name__EVAL_55;
  assign out_xbar__EVAL_45 = coupler_to_clint__EVAL_19;
  assign in_xbar__EVAL_6 = atomics__EVAL_35;
  assign coupler_to_plic__EVAL_31 = out_xbar__EVAL_26;
  assign fixer__EVAL = buffer__EVAL_10;
  assign out_xbar__EVAL_113 = fixer__EVAL_26;
  assign buffer__EVAL_33 = atomics__EVAL_25;
  assign _EVAL_95 = coupler_to_port_named_axi4_periph_port__EVAL_10;
  assign coupler_to_clint__EVAL_31 = out_xbar__EVAL_12;
  assign _EVAL_133 = coupler_to_tile_with_no_name__EVAL_42;
  assign coupler_to_debug__EVAL_11 = out_xbar__EVAL_115;
  assign buffer_1__EVAL_20 = _EVAL_7;
  assign out_xbar__EVAL_48 = coupler_to_clint__EVAL_18;
  assign coupler_to_port_named_axi4_periph_port__EVAL_12 = out_xbar__EVAL_0;
  assign coupler_to_debug__EVAL_15 = out_xbar__EVAL_35;
  assign coupler_to_testindicator__EVAL_5 = _EVAL_1;
  assign coupler_to_clint__EVAL_25 = out_xbar__EVAL_79;
  assign _EVAL_24 = coupler_to_port_named_axi4_periph_port__EVAL_4;
  assign _EVAL_19 = coupler_to_clint__EVAL_28;
  assign _EVAL_11 = coupler_to_port_named_axi4_periph_port__EVAL_33;
  assign _EVAL_149 = coupler_to_tile_with_no_name__EVAL_28;
  assign out_xbar__EVAL_101 = coupler_to_debug__EVAL_25;
  assign out_xbar__EVAL_9 = coupler_to_plic__EVAL_12;
  assign buffer_1__EVAL_27 = _EVAL_82;
  assign buffer__EVAL_27 = fixer__EVAL_27;
  assign _EVAL_129 = buffer_1__EVAL_16;
  assign _EVAL_32 = coupler_to_tile_with_no_name__EVAL_54;
  assign buffer_1__EVAL_23 = _EVAL_144;
  assign out_xbar__EVAL_16 = _EVAL_90;
  assign _EVAL_28 = coupler_to_tile_with_no_name__EVAL_8;
  assign coupler_to_port_named_axi4_periph_port__EVAL_38 = out_xbar__EVAL_80;
  assign coupler_to_clint__EVAL_26 = _EVAL_90;
  assign _EVAL_125 = coupler_to_port_named_axi4_periph_port__EVAL_48;
  assign coupler_to_clint__EVAL_1 = out_xbar__EVAL_21;
  assign coupler_to_port_named_axi4_periph_port__EVAL_2 = _EVAL_84;
  assign wrapped_error_device__EVAL_13 = out_xbar__EVAL_117;
  assign coupler_to_port_named_axi4_periph_port__EVAL_40 = _EVAL_109;
  assign out_xbar__EVAL_20 = coupler_to_port_named_axi4_periph_port__EVAL_28;
  assign coupler_to_port_named_axi4_periph_port__EVAL_27 = out_xbar__EVAL_18;
  assign out_xbar__EVAL_4 = coupler_to_testindicator__EVAL_25;
  assign coupler_to_plic__EVAL_8 = _EVAL_127;
  assign out_xbar__EVAL_40 = coupler_to_port_named_axi4_periph_port__EVAL_47;
  assign _EVAL_157 = coupler_to_clint__EVAL_23;
  assign out_xbar__EVAL_96 = fixer__EVAL_8;
  assign coupler_to_tile_with_no_name__EVAL_47 = out_xbar__EVAL_8;
  assign buffer__EVAL_35 = fixer__EVAL_37;
  assign out_xbar__EVAL_61 = fixer__EVAL_32;
  assign _EVAL_92 = coupler_to_clint__EVAL_22;
  assign fixer__EVAL_21 = out_xbar__EVAL_90;
  assign buffer__EVAL_21 = atomics__EVAL_28;
  assign coupler_to_plic__EVAL_26 = out_xbar__EVAL_32;
  assign _EVAL_120 = buffer_1__EVAL_32;
  assign _EVAL_3 = coupler_to_tile_with_no_name__EVAL_52;
  assign out_xbar__EVAL_84 = wrapped_error_device__EVAL_7;
  assign buffer__EVAL_40 = fixer__EVAL_18;
  assign out_xbar__EVAL_91 = coupler_to_clint__EVAL_14;
  assign coupler_to_tile_with_no_name__EVAL_17 = _EVAL_104;
  assign buffer__EVAL_0 = atomics__EVAL_33;
  assign _EVAL_139 = coupler_to_tile_with_no_name__EVAL_34;
  assign _EVAL_113 = coupler_to_testindicator__EVAL_6;
  assign coupler_to_clint__EVAL_15 = out_xbar__EVAL_51;
  assign wrapped_error_device__EVAL_3 = out_xbar__EVAL_39;
  assign coupler_to_port_named_axi4_periph_port__EVAL_8 = _EVAL_130;
  assign coupler_to_plic__EVAL_5 = out_xbar__EVAL_67;
  assign coupler_to_tile_with_no_name__EVAL_50 = _EVAL_27;
  assign coupler_to_debug__EVAL_19 = out_xbar__EVAL_42;
  assign coupler_to_tile_with_no_name__EVAL_11 = _EVAL_137;
  assign out_xbar__EVAL_64 = fixer__EVAL_20;
  assign buffer__EVAL_22 = fixer__EVAL_33;
  assign coupler_to_debug__EVAL_24 = _EVAL_82;
  assign _EVAL_68 = buffer_1__EVAL_38;
  assign coupler_to_debug__EVAL_16 = _EVAL_20;
  assign coupler_to_tile_with_no_name__EVAL_12 = _EVAL_159;
  assign _EVAL_16 = coupler_to_tile_with_no_name__EVAL_36;
  assign coupler_to_clint__EVAL_27 = _EVAL_124;
  assign atomics__EVAL_38 = buffer__EVAL_23;
  assign buffer_1__EVAL_39 = _EVAL_98;
  assign coupler_to_clint__EVAL_3 = _EVAL_58;
  assign _EVAL_106 = coupler_to_port_named_axi4_periph_port__EVAL_32;
  assign atomics__EVAL_6 = buffer__EVAL_18;
  assign coupler_to_tile_with_no_name__EVAL_31 = out_xbar__EVAL_6;
  assign atomics__EVAL_29 = in_xbar__EVAL_28;
  assign coupler_to_clint__EVAL_30 = out_xbar__EVAL_7;
  assign _EVAL_142 = coupler_to_port_named_axi4_periph_port__EVAL_23;
  assign _EVAL_134 = coupler_to_clint__EVAL_10;
  assign coupler_to_debug__EVAL_32 = out_xbar__EVAL_87;
  assign buffer_1__EVAL_11 = in_xbar__EVAL_17;
  assign out_xbar__EVAL_24 = coupler_to_port_named_axi4_periph_port__EVAL_5;
  assign _EVAL_91 = coupler_to_clint__EVAL_0;
  assign buffer_1__EVAL_13 = in_xbar__EVAL;
  assign wrapped_error_device__EVAL_11 = out_xbar__EVAL_47;
  assign buffer__EVAL_20 = _EVAL_82;
  assign coupler_to_plic__EVAL_16 = _EVAL_131;
  assign coupler_to_clint__EVAL_9 = _EVAL_72;
  assign atomics__EVAL_26 = buffer__EVAL_28;
  assign coupler_to_debug__EVAL = _EVAL_107;
  assign fixer__EVAL_6 = buffer__EVAL_6;
  assign out_xbar__EVAL_29 = wrapped_error_device__EVAL_4;
  assign fixer__EVAL_40 = out_xbar__EVAL_34;
  assign coupler_to_plic__EVAL_3 = _EVAL_83;
  assign fixer__EVAL_24 = out_xbar__EVAL_13;
  assign coupler_to_testindicator__EVAL_30 = out_xbar__EVAL_122;
  assign buffer_1__EVAL_6 = in_xbar__EVAL_13;
  assign atomics__EVAL_40 = in_xbar__EVAL_38;
  assign in_xbar__EVAL_20 = buffer_1__EVAL_34;
  assign coupler_to_testindicator__EVAL_1 = _EVAL_80;
  assign coupler_to_tile_with_no_name__EVAL_39 = out_xbar__EVAL_137;
  assign out_xbar__EVAL_2 = coupler_to_clint__EVAL_17;
  assign out_xbar__EVAL_75 = coupler_to_testindicator__EVAL_27;
  assign out_xbar__EVAL_53 = fixer__EVAL_17;
  assign _EVAL_21 = coupler_to_plic__EVAL_10;
  assign atomics__EVAL_7 = buffer__EVAL_32;
  assign coupler_to_tile_with_no_name__EVAL_15 = _EVAL_94;
  assign coupler_to_port_named_axi4_periph_port__EVAL_51 = _EVAL_41;
  assign coupler_to_testindicator__EVAL_0 = out_xbar__EVAL_85;
  assign coupler_to_clint__EVAL_2 = _EVAL_13;
  assign out_xbar__EVAL_25 = fixer__EVAL_10;
  assign wrapped_error_device__EVAL_9 = out_xbar__EVAL_131;
  assign _EVAL_88 = coupler_to_plic__EVAL_30;
  assign coupler_to_plic__EVAL_22 = _EVAL_82;
  assign buffer_1__EVAL_15 = _EVAL_90;
  assign in_xbar__EVAL_0 = buffer_1__EVAL_26;
  assign coupler_to_port_named_axi4_periph_port__EVAL_21 = _EVAL_90;
  assign out_xbar__EVAL_121 = fixer__EVAL_13;
  assign fixer__EVAL_34 = buffer__EVAL_11;
  assign out_xbar__EVAL_128 = wrapped_error_device__EVAL_8;
  assign _EVAL_59 = coupler_to_port_named_axi4_periph_port__EVAL_30;
  assign coupler_to_tile_with_no_name__EVAL_7 = out_xbar__EVAL_28;
  assign fixer__EVAL_16 = buffer__EVAL_30;
  assign _EVAL_155 = coupler_to_testindicator__EVAL_9;
  assign out_xbar__EVAL_10 = fixer__EVAL_7;
  assign atomics__EVAL_32 = in_xbar__EVAL_32;
  assign out_xbar__EVAL_135 = wrapped_error_device__EVAL_18;
  assign out_xbar__EVAL_22 = coupler_to_testindicator__EVAL_8;
  assign atomics__EVAL_39 = in_xbar__EVAL_9;
  assign coupler_to_debug__EVAL_0 = _EVAL_90;
  assign coupler_to_port_named_axi4_periph_port__EVAL_46 = out_xbar__EVAL_62;
  assign _EVAL_103 = buffer_1__EVAL_33;
  assign buffer_1__EVAL_14 = in_xbar__EVAL_26;
  assign buffer__EVAL_4 = atomics__EVAL_36;
  assign _EVAL_73 = coupler_to_port_named_axi4_periph_port__EVAL_6;
  assign _EVAL_49 = coupler_to_testindicator__EVAL_29;
  assign coupler_to_testindicator__EVAL_24 = out_xbar__EVAL_141;
  assign buffer_1__EVAL_0 = _EVAL_53;
  assign in_xbar__EVAL_16 = buffer_1__EVAL_17;
  assign coupler_to_tile_with_no_name__EVAL_0 = _EVAL_63;
  assign in_xbar__EVAL_23 = atomics__EVAL_22;
  assign coupler_to_testindicator__EVAL_21 = _EVAL_82;
  assign _EVAL_18 = coupler_to_port_named_axi4_periph_port__EVAL_9;
  assign _EVAL_69 = coupler_to_tile_with_no_name__EVAL_14;
  assign _EVAL_66 = coupler_to_plic__EVAL_18;
  assign _EVAL_64 = coupler_to_port_named_axi4_periph_port__EVAL_7;
  assign _EVAL_132 = coupler_to_debug__EVAL_22;
  assign out_xbar__EVAL_56 = wrapped_error_device__EVAL_15;
  assign _EVAL_96 = coupler_to_plic__EVAL_25;
  assign atomics__EVAL_37 = buffer__EVAL_34;
  assign _EVAL_35 = coupler_to_port_named_axi4_periph_port__EVAL_49;
  assign fixer__EVAL_29 = out_xbar__EVAL_74;
  assign out_xbar__EVAL_52 = coupler_to_clint__EVAL_21;
  assign _EVAL_37 = coupler_to_tile_with_no_name__EVAL_25;
  assign _EVAL_110 = coupler_to_port_named_axi4_periph_port__EVAL_15;
  assign wrapped_error_device__EVAL_2 = out_xbar__EVAL_23;
  assign out_xbar__EVAL_77 = coupler_to_testindicator__EVAL_2;
  assign coupler_to_tile_with_no_name__EVAL_57 = out_xbar__EVAL_110;
  assign out_xbar__EVAL_58 = coupler_to_tile_with_no_name__EVAL_4;
endmodule
