//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_73(
  output        _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  output [31:0] _EVAL_2,
  output [6:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [5:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [1:0]  _EVAL_9,
  output [6:0]  _EVAL_10,
  input  [7:0]  _EVAL_11,
  output [7:0]  _EVAL_12,
  output [1:0]  _EVAL_13,
  output [1:0]  _EVAL_14,
  output [1:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  input  [2:0]  _EVAL_20,
  output [31:0] _EVAL_21,
  input  [2:0]  _EVAL_22,
  output        _EVAL_23,
  input  [1:0]  _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input  [5:0]  _EVAL_27,
  input         _EVAL_28,
  output        _EVAL_29,
  input  [3:0]  _EVAL_30,
  input  [31:0] _EVAL_31,
  output        _EVAL_32,
  output [1:0]  _EVAL_33,
  output [3:0]  _EVAL_34,
  output        _EVAL_35,
  input         _EVAL_36,
  output [1:0]  _EVAL_37,
  input  [1:0]  _EVAL_38,
  input  [6:0]  _EVAL_39,
  output [2:0]  _EVAL_40,
  output [5:0]  _EVAL_41,
  output [7:0]  _EVAL_42,
  input  [31:0] _EVAL_43,
  output        _EVAL_44,
  input  [31:0] _EVAL_45,
  output [5:0]  _EVAL_46,
  input  [1:0]  _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  output        _EVAL_50,
  input  [1:0]  _EVAL_51,
  output [1:0]  _EVAL_52,
  input         _EVAL_53,
  input  [1:0]  _EVAL_54,
  output        _EVAL_55,
  output [31:0] _EVAL_56,
  input         _EVAL_57,
  input  [1:0]  _EVAL_58,
  input  [1:0]  _EVAL_59,
  input         _EVAL_60,
  output        _EVAL_61,
  input  [31:0] _EVAL_62,
  input  [6:0]  _EVAL_63,
  input  [7:0]  _EVAL_64
);
  wire [1:0] Queue_1__EVAL;
  wire [1:0] Queue_1__EVAL_0;
  wire [2:0] Queue_1__EVAL_1;
  wire [5:0] Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire [5:0] Queue_1__EVAL_4;
  wire [2:0] Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire [31:0] Queue_1__EVAL_7;
  wire [7:0] Queue_1__EVAL_8;
  wire [1:0] Queue_1__EVAL_9;
  wire  Queue_1__EVAL_10;
  wire  Queue_1__EVAL_11;
  wire [1:0] Queue_1__EVAL_12;
  wire  Queue_1__EVAL_13;
  wire [31:0] Queue_1__EVAL_14;
  wire [7:0] Queue_1__EVAL_15;
  wire  Queue_1__EVAL_16;
  wire  Queue_2__EVAL;
  wire  Queue_2__EVAL_0;
  wire [3:0] Queue_2__EVAL_1;
  wire  Queue_2__EVAL_2;
  wire [31:0] Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire  Queue_2__EVAL_5;
  wire  Queue_2__EVAL_6;
  wire  Queue_2__EVAL_7;
  wire [3:0] Queue_2__EVAL_8;
  wire  Queue_2__EVAL_9;
  wire [31:0] Queue_2__EVAL_10;
  wire [1:0] Queue__EVAL;
  wire [1:0] Queue__EVAL_0;
  wire [2:0] Queue__EVAL_1;
  wire [5:0] Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire [5:0] Queue__EVAL_4;
  wire [2:0] Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire [31:0] Queue__EVAL_7;
  wire [7:0] Queue__EVAL_8;
  wire [1:0] Queue__EVAL_9;
  wire  Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire [1:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire [31:0] Queue__EVAL_14;
  wire [7:0] Queue__EVAL_15;
  wire  Queue__EVAL_16;
  reg [31:0] _EVAL_71;
  reg [31:0] _RAND_0;
  reg [1:0] _EVAL_101;
  reg [31:0] _RAND_1;
  reg  _EVAL_112;
  reg [31:0] _RAND_2;
  reg [7:0] _EVAL_132;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_136;
  reg [31:0] _RAND_4;
  reg [7:0] _EVAL_172;
  reg [31:0] _RAND_5;
  reg  _EVAL_182;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_213;
  reg [31:0] _RAND_7;
  reg  _EVAL_229;
  reg [31:0] _RAND_8;
  reg [1:0] _EVAL_296;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_356;
  reg [31:0] _RAND_10;
  reg [8:0] _EVAL_407;
  reg [31:0] _RAND_11;
  wire  _EVAL_170;
  wire [1:0] _EVAL_252;
  wire [31:0] _EVAL_267;
  wire [31:0] _EVAL_211;
  wire [31:0] _EVAL_287;
  wire [32:0] _EVAL_305;
  wire [32:0] _EVAL_323;
  wire [32:0] _EVAL_271;
  wire  _EVAL_362;
  wire [1:0] _EVAL_238;
  wire  _EVAL_134;
  wire [2:0] _EVAL_227;
  wire  _EVAL_180;
  wire  _EVAL_177;
  wire [8:0] _EVAL_131;
  wire [1:0] _EVAL_232;
  wire [7:0] _EVAL_338;
  wire [7:0] _EVAL_73;
  wire [6:0] _EVAL_206;
  wire [7:0] _EVAL_249;
  wire [7:0] _EVAL_282;
  wire [5:0] _EVAL_266;
  wire [7:0] _EVAL_233;
  wire [7:0] _EVAL_390;
  wire [3:0] _EVAL_87;
  wire [7:0] _EVAL_294;
  wire [32:0] _EVAL_121;
  wire [32:0] _EVAL_216;
  wire [32:0] _EVAL_273;
  wire  _EVAL_185;
  wire [1:0] _EVAL_191;
  wire [8:0] _EVAL_212;
  wire [7:0] _EVAL_226;
  wire [6:0] _EVAL_283;
  wire [7:0] _EVAL_124;
  wire [7:0] _EVAL_375;
  wire [8:0] _EVAL_354;
  wire [7:0] _EVAL_263;
  wire [7:0] _EVAL_243;
  wire [9:0] _EVAL_393;
  wire [7:0] _EVAL_334;
  wire [7:0] _EVAL_149;
  wire [11:0] _EVAL_348;
  wire [7:0] _EVAL_158;
  wire [7:0] _EVAL_187;
  wire [7:0] _EVAL_106;
  wire [7:0] _EVAL_329;
  wire [31:0] _EVAL_69;
  wire [31:0] _EVAL_74;
  wire [7:0] _EVAL_368;
  wire [8:0] _EVAL_76;
  wire [7:0] _EVAL_278;
  wire [7:0] _EVAL_404;
  wire [9:0] _EVAL_95;
  wire [7:0] _EVAL_199;
  wire [7:0] _EVAL_167;
  wire [11:0] _EVAL_246;
  wire [7:0] _EVAL_275;
  wire [7:0] _EVAL_358;
  wire [7:0] _EVAL_388;
  wire [7:0] _EVAL_234;
  wire [31:0] _EVAL_302;
  wire [32:0] _EVAL_270;
  wire [32:0] _EVAL_82;
  wire [32:0] _EVAL_204;
  wire  _EVAL_406;
  wire [5:0] _EVAL_276;
  wire [31:0] _EVAL_222;
  wire [32:0] _EVAL_85;
  wire [32:0] _EVAL_139;
  wire [32:0] _EVAL_118;
  wire  _EVAL_308;
  wire [31:0] _EVAL_290;
  wire [32:0] _EVAL_79;
  wire [32:0] _EVAL_190;
  wire [32:0] _EVAL_321;
  wire  _EVAL_160;
  wire  _EVAL_72;
  wire [31:0] _EVAL_144;
  wire [32:0] _EVAL_186;
  wire [32:0] _EVAL_269;
  wire [32:0] _EVAL_104;
  wire  _EVAL_310;
  wire  _EVAL_174;
  wire [31:0] _EVAL_319;
  wire [32:0] _EVAL_382;
  wire [32:0] _EVAL_391;
  wire [32:0] _EVAL_350;
  wire  _EVAL_197;
  wire  _EVAL_242;
  wire [32:0] _EVAL_357;
  wire [32:0] _EVAL_162;
  wire [32:0] _EVAL_231;
  wire  _EVAL_311;
  wire  _EVAL_352;
  wire [31:0] _EVAL_395;
  wire [32:0] _EVAL_111;
  wire [32:0] _EVAL_389;
  wire [32:0] _EVAL_207;
  wire  _EVAL_285;
  wire  _EVAL_108;
  wire [31:0] _EVAL_145;
  wire [32:0] _EVAL_397;
  wire [32:0] _EVAL_360;
  wire [32:0] _EVAL_373;
  wire  _EVAL_257;
  wire  _EVAL_353;
  wire [3:0] _EVAL_123;
  wire [5:0] _EVAL_154;
  wire [5:0] _EVAL_91;
  wire [7:0] _EVAL_307;
  wire [7:0] _EVAL_183;
  wire [7:0] _EVAL_126;
  wire [8:0] _EVAL_392;
  wire [8:0] _EVAL_102;
  wire [8:0] _EVAL_284;
  wire [8:0] _EVAL_90;
  wire [8:0] _EVAL_208;
  wire [15:0] _EVAL_117;
  wire [22:0] _EVAL_94;
  wire [22:0] _EVAL_140;
  wire [14:0] _EVAL_66;
  wire [31:0] _EVAL_255;
  wire [1:0] _EVAL_259;
  wire [31:0] _EVAL_214;
  wire [31:0] _EVAL_309;
  wire  _EVAL_219;
  wire  _EVAL_274;
  wire  _EVAL_262;
  wire  _EVAL_398;
  wire  _EVAL_103;
  wire  _EVAL_83;
  wire  _EVAL_394;
  wire  _EVAL_135;
  wire  _EVAL_75;
  wire [15:0] _EVAL_235;
  wire [15:0] _EVAL_344;
  wire [1:0] _EVAL_194;
  wire  _EVAL_381;
  wire [2:0] _EVAL_221;
  wire  _EVAL_288;
  wire  _EVAL_408;
  wire [7:0] _EVAL_340;
  wire [7:0] _EVAL_272;
  wire [6:0] _EVAL_68;
  wire [7:0] _EVAL_156;
  wire [7:0] _EVAL_120;
  wire [5:0] _EVAL_295;
  wire [7:0] _EVAL_320;
  wire [7:0] _EVAL_279;
  wire [3:0] _EVAL_220;
  wire [7:0] _EVAL_250;
  wire [7:0] _EVAL_372;
  wire [6:0] _EVAL_176;
  wire [7:0] _EVAL_343;
  wire [7:0] _EVAL_210;
  wire [8:0] _EVAL_384;
  wire [7:0] _EVAL_330;
  wire [7:0] _EVAL_96;
  wire [9:0] _EVAL_258;
  wire [7:0] _EVAL_128;
  wire [7:0] _EVAL_223;
  wire [11:0] _EVAL_322;
  wire [7:0] _EVAL_301;
  wire [7:0] _EVAL_138;
  wire [7:0] _EVAL_317;
  wire [7:0] _EVAL_77;
  wire [7:0] _EVAL_159;
  wire [8:0] _EVAL_146;
  wire [7:0] _EVAL_286;
  wire [7:0] _EVAL_163;
  wire [9:0] _EVAL_92;
  wire [7:0] _EVAL_218;
  wire [7:0] _EVAL_304;
  wire [11:0] _EVAL_240;
  wire [7:0] _EVAL_299;
  wire [7:0] _EVAL_105;
  wire [7:0] _EVAL_402;
  wire [7:0] _EVAL_386;
  wire [31:0] _EVAL_253;
  wire [32:0] _EVAL_173;
  wire [32:0] _EVAL_327;
  wire [32:0] _EVAL_316;
  wire  _EVAL_268;
  wire [5:0] _EVAL_336;
  wire [31:0] _EVAL_333;
  wire [32:0] _EVAL_178;
  wire [32:0] _EVAL_157;
  wire [32:0] _EVAL_261;
  wire  _EVAL_193;
  wire  _EVAL_109;
  wire [31:0] _EVAL_318;
  wire [32:0] _EVAL_260;
  wire [32:0] _EVAL_209;
  wire [32:0] _EVAL_378;
  wire  _EVAL_127;
  wire  _EVAL_217;
  wire [31:0] _EVAL_385;
  wire [32:0] _EVAL_335;
  wire [32:0] _EVAL_143;
  wire [32:0] _EVAL_148;
  wire  _EVAL_251;
  wire  _EVAL_86;
  wire  _EVAL_150;
  wire [31:0] _EVAL_341;
  wire [32:0] _EVAL_277;
  wire [32:0] _EVAL_97;
  wire [32:0] _EVAL_324;
  wire  _EVAL_351;
  wire  _EVAL_137;
  wire [31:0] _EVAL_200;
  wire [32:0] _EVAL_151;
  wire [32:0] _EVAL_241;
  wire [32:0] _EVAL_228;
  wire  _EVAL_129;
  wire  _EVAL_169;
  wire [3:0] _EVAL_401;
  wire [5:0] _EVAL_289;
  wire [5:0] _EVAL_300;
  wire [7:0] _EVAL_326;
  wire [7:0] _EVAL_332;
  wire [7:0] _EVAL_347;
  wire [8:0] _EVAL_215;
  wire  _EVAL_107;
  wire  _EVAL_181;
  wire [8:0] _EVAL_363;
  wire [8:0] _EVAL_265;
  wire [8:0] _EVAL_331;
  wire [8:0] _EVAL_203;
  wire [31:0] _EVAL_387;
  wire [8:0] _EVAL_161;
  wire [8:0] _EVAL_369;
  wire [8:0] _EVAL_248;
  wire [8:0] _EVAL_339;
  wire [8:0] _EVAL_88;
  wire [8:0] _EVAL_244;
  wire [8:0] _EVAL_230;
  wire [1:0] _EVAL_78;
  wire [31:0] _EVAL_141;
  wire [31:0] _EVAL_130;
  wire [31:0] _EVAL_312;
  wire [31:0] _EVAL_205;
  wire [31:0] _EVAL_361;
  wire [31:0] _EVAL_93;
  wire [31:0] _EVAL_379;
  wire  _EVAL_113;
  wire  _EVAL_89;
  wire  _EVAL_291;
  wire [8:0] _EVAL_298;
  wire [1:0] _EVAL_349;
  wire [15:0] _EVAL_224;
  wire [15:0] _EVAL_147;
  wire [31:0] _EVAL_325;
  wire [31:0] _EVAL_119;
  wire [15:0] _EVAL_346;
  wire [22:0] _EVAL_247;
  wire [22:0] _EVAL_281;
  wire [14:0] _EVAL_399;
  wire [31:0] _EVAL_125;
  wire [31:0] _EVAL_202;
  wire [3:0] _EVAL_355;
  wire  _EVAL_225;
  wire  _EVAL_345;
  wire  _EVAL_188;
  wire  _EVAL_264;
  wire  _EVAL_192;
  wire  _EVAL_81;
  wire  _EVAL_116;
  wire [31:0] _EVAL_198;
  wire  _EVAL_110;
  wire  _EVAL_237;
  wire [1:0] _EVAL_256;
  wire [1:0] _EVAL_396;
  wire [31:0] _EVAL_366;
  wire [1:0] _EVAL_403;
  wire [1:0] _EVAL_337;
  wire [31:0] _EVAL_342;
  wire [31:0] _EVAL_155;
  wire  _EVAL_377;
  wire [31:0] _EVAL_313;
  wire [31:0] _EVAL_364;
  wire  _EVAL_239;
  wire  _EVAL_114;
  wire  _EVAL_236;
  wire [31:0] _EVAL_189;
  wire [1:0] _EVAL_245;
  wire  _EVAL_115;
  wire  _EVAL_65;
  wire  _EVAL_153;
  wire  _EVAL_166;
  wire [8:0] _EVAL_371;
  wire [8:0] _EVAL_142;
  wire [5:0] _EVAL_171;
  wire  _EVAL_164;
  wire [5:0] _EVAL_168;
  wire  _EVAL_328;
  wire  _EVAL_67;
  wire  _EVAL_280;
  SiFive__EVAL_72 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14),
    ._EVAL_15(Queue_1__EVAL_15),
    ._EVAL_16(Queue_1__EVAL_16)
  );
  SiFive__EVAL_31 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6),
    ._EVAL_7(Queue_2__EVAL_7),
    ._EVAL_8(Queue_2__EVAL_8),
    ._EVAL_9(Queue_2__EVAL_9),
    ._EVAL_10(Queue_2__EVAL_10)
  );
  SiFive__EVAL_72 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16)
  );
  assign _EVAL_170 = _EVAL_39[0];
  assign _EVAL_252 = _EVAL_101 | _EVAL_38;
  assign _EVAL_267 = Queue__EVAL_7;
  assign _EVAL_211 = _EVAL_182 ? _EVAL_71 : _EVAL_267;
  assign _EVAL_287 = _EVAL_211 ^ 32'h40000000;
  assign _EVAL_305 = {1'b0,$signed(_EVAL_287)};
  assign _EVAL_323 = $signed(_EVAL_305) & $signed(33'sheb000000);
  assign _EVAL_271 = $signed(_EVAL_323);
  assign _EVAL_362 = $signed(_EVAL_271) == $signed(33'sh0);
  assign _EVAL_238 = Queue_1__EVAL_12;
  assign _EVAL_134 = _EVAL_238 == 2'h0;
  assign _EVAL_227 = Queue_1__EVAL_5;
  assign _EVAL_180 = _EVAL_227 != 3'h2;
  assign _EVAL_177 = _EVAL_134 | _EVAL_180;
  assign _EVAL_131 = 9'h3 << _EVAL_227;
  assign _EVAL_232 = _EVAL_131[1:0];
  assign _EVAL_338 = Queue_1__EVAL_8;
  assign _EVAL_73 = _EVAL_229 ? _EVAL_132 : _EVAL_338;
  assign _EVAL_206 = _EVAL_73[7:1];
  assign _EVAL_249 = {{1'd0}, _EVAL_206};
  assign _EVAL_282 = _EVAL_73 | _EVAL_249;
  assign _EVAL_266 = _EVAL_282[7:2];
  assign _EVAL_233 = {{2'd0}, _EVAL_266};
  assign _EVAL_390 = _EVAL_282 | _EVAL_233;
  assign _EVAL_87 = _EVAL_390[7:4];
  assign _EVAL_294 = {{4'd0}, _EVAL_87};
  assign _EVAL_121 = {1'b0,$signed(_EVAL_211)};
  assign _EVAL_216 = $signed(_EVAL_121) & $signed(33'sheb001000);
  assign _EVAL_273 = $signed(_EVAL_216);
  assign _EVAL_185 = $signed(_EVAL_273) == $signed(33'sh0);
  assign _EVAL_191 = _EVAL_296 | _EVAL_38;
  assign _EVAL_212 = {{1'd0}, _EVAL_73};
  assign _EVAL_226 = _EVAL_390 | _EVAL_294;
  assign _EVAL_283 = _EVAL_226[7:1];
  assign _EVAL_124 = {{1'd0}, _EVAL_283};
  assign _EVAL_375 = ~ _EVAL_73;
  assign _EVAL_354 = {_EVAL_375, 1'h0};
  assign _EVAL_263 = _EVAL_354[7:0];
  assign _EVAL_243 = _EVAL_375 | _EVAL_263;
  assign _EVAL_393 = {_EVAL_243, 2'h0};
  assign _EVAL_334 = _EVAL_393[7:0];
  assign _EVAL_149 = _EVAL_243 | _EVAL_334;
  assign _EVAL_348 = {_EVAL_149, 4'h0};
  assign _EVAL_158 = _EVAL_348[7:0];
  assign _EVAL_187 = _EVAL_149 | _EVAL_158;
  assign _EVAL_106 = ~ _EVAL_187;
  assign _EVAL_329 = _EVAL_124 | _EVAL_106;
  assign _EVAL_69 = Queue_1__EVAL_7;
  assign _EVAL_74 = _EVAL_229 ? _EVAL_213 : _EVAL_69;
  assign _EVAL_368 = _EVAL_74[9:2];
  assign _EVAL_76 = {_EVAL_368, 1'h0};
  assign _EVAL_278 = _EVAL_76[7:0];
  assign _EVAL_404 = _EVAL_368 | _EVAL_278;
  assign _EVAL_95 = {_EVAL_404, 2'h0};
  assign _EVAL_199 = _EVAL_95[7:0];
  assign _EVAL_167 = _EVAL_404 | _EVAL_199;
  assign _EVAL_246 = {_EVAL_167, 4'h0};
  assign _EVAL_275 = _EVAL_246[7:0];
  assign _EVAL_358 = _EVAL_167 | _EVAL_275;
  assign _EVAL_388 = ~ _EVAL_358;
  assign _EVAL_234 = _EVAL_329 & _EVAL_388;
  assign _EVAL_302 = _EVAL_74 ^ 32'h1000;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_302)};
  assign _EVAL_82 = $signed(_EVAL_270) & $signed(33'sheb001000);
  assign _EVAL_204 = $signed(_EVAL_82);
  assign _EVAL_406 = $signed(_EVAL_204) == $signed(33'sh0);
  assign _EVAL_276 = _EVAL_406 ? 6'h3f : 6'h0;
  assign _EVAL_222 = _EVAL_74 ^ 32'h40000000;
  assign _EVAL_85 = {1'b0,$signed(_EVAL_222)};
  assign _EVAL_139 = $signed(_EVAL_85) & $signed(33'sheb000000);
  assign _EVAL_118 = $signed(_EVAL_139);
  assign _EVAL_308 = $signed(_EVAL_118) == $signed(33'sh0);
  assign _EVAL_290 = _EVAL_74 ^ 32'h80000000;
  assign _EVAL_79 = {1'b0,$signed(_EVAL_290)};
  assign _EVAL_190 = $signed(_EVAL_79) & $signed(33'sheb000000);
  assign _EVAL_321 = $signed(_EVAL_190);
  assign _EVAL_160 = $signed(_EVAL_321) == $signed(33'sh0);
  assign _EVAL_72 = _EVAL_308 | _EVAL_160;
  assign _EVAL_144 = _EVAL_74 ^ 32'h8000000;
  assign _EVAL_186 = {1'b0,$signed(_EVAL_144)};
  assign _EVAL_269 = $signed(_EVAL_186) & $signed(33'she8000000);
  assign _EVAL_104 = $signed(_EVAL_269);
  assign _EVAL_310 = $signed(_EVAL_104) == $signed(33'sh0);
  assign _EVAL_174 = _EVAL_72 | _EVAL_310;
  assign _EVAL_319 = _EVAL_74 ^ 32'h2000000;
  assign _EVAL_382 = {1'b0,$signed(_EVAL_319)};
  assign _EVAL_391 = $signed(_EVAL_382) & $signed(33'sheb000000);
  assign _EVAL_350 = $signed(_EVAL_391);
  assign _EVAL_197 = $signed(_EVAL_350) == $signed(33'sh0);
  assign _EVAL_242 = _EVAL_174 | _EVAL_197;
  assign _EVAL_357 = {1'b0,$signed(_EVAL_74)};
  assign _EVAL_162 = $signed(_EVAL_357) & $signed(33'sheb001000);
  assign _EVAL_231 = $signed(_EVAL_162);
  assign _EVAL_311 = $signed(_EVAL_231) == $signed(33'sh0);
  assign _EVAL_352 = _EVAL_242 | _EVAL_311;
  assign _EVAL_395 = _EVAL_74 ^ 32'h1000000;
  assign _EVAL_111 = {1'b0,$signed(_EVAL_395)};
  assign _EVAL_389 = $signed(_EVAL_111) & $signed(33'sheb000000);
  assign _EVAL_207 = $signed(_EVAL_389);
  assign _EVAL_285 = $signed(_EVAL_207) == $signed(33'sh0);
  assign _EVAL_108 = _EVAL_352 | _EVAL_285;
  assign _EVAL_145 = _EVAL_74 ^ 32'h20000000;
  assign _EVAL_397 = {1'b0,$signed(_EVAL_145)};
  assign _EVAL_360 = $signed(_EVAL_397) & $signed(33'sheb000000);
  assign _EVAL_373 = $signed(_EVAL_360);
  assign _EVAL_257 = $signed(_EVAL_373) == $signed(33'sh0);
  assign _EVAL_353 = _EVAL_108 | _EVAL_257;
  assign _EVAL_123 = _EVAL_353 ? 4'hf : 4'h0;
  assign _EVAL_154 = {{2'd0}, _EVAL_123};
  assign _EVAL_91 = _EVAL_276 | _EVAL_154;
  assign _EVAL_307 = {{2'd0}, _EVAL_91};
  assign _EVAL_183 = _EVAL_234 & _EVAL_307;
  assign _EVAL_126 = _EVAL_177 ? 8'h0 : _EVAL_183;
  assign _EVAL_392 = {_EVAL_126, 1'h0};
  assign _EVAL_102 = _EVAL_392 | 9'h1;
  assign _EVAL_284 = {1'h0,_EVAL_126};
  assign _EVAL_90 = ~ _EVAL_284;
  assign _EVAL_208 = _EVAL_102 & _EVAL_90;
  assign _EVAL_117 = {_EVAL_338,8'hff};
  assign _EVAL_94 = {{7'd0}, _EVAL_117};
  assign _EVAL_140 = _EVAL_94 << _EVAL_227;
  assign _EVAL_66 = _EVAL_140[22:8];
  assign _EVAL_255 = ~ _EVAL_74;
  assign _EVAL_259 = ~ _EVAL_232;
  assign _EVAL_214 = {{30'd0}, _EVAL_259};
  assign _EVAL_309 = _EVAL_255 | _EVAL_214;
  assign _EVAL_219 = Queue_2__EVAL;
  assign _EVAL_274 = _EVAL_407 == 9'h0;
  assign _EVAL_262 = _EVAL_274 == 1'h0;
  assign _EVAL_398 = Queue_1__EVAL_3;
  assign _EVAL_103 = _EVAL_112 == 1'h0;
  assign _EVAL_83 = _EVAL_398 & _EVAL_103;
  assign _EVAL_394 = _EVAL_262 | _EVAL_83;
  assign _EVAL_135 = _EVAL_219 & _EVAL_394;
  assign _EVAL_75 = _EVAL_60 & _EVAL_135;
  assign _EVAL_235 = {{7'd0}, _EVAL_208};
  assign _EVAL_344 = _EVAL_235 << _EVAL_227;
  assign _EVAL_194 = Queue__EVAL_12;
  assign _EVAL_381 = _EVAL_194 == 2'h0;
  assign _EVAL_221 = Queue__EVAL_5;
  assign _EVAL_288 = _EVAL_221 != 3'h2;
  assign _EVAL_408 = _EVAL_381 | _EVAL_288;
  assign _EVAL_340 = Queue__EVAL_8;
  assign _EVAL_272 = _EVAL_182 ? _EVAL_172 : _EVAL_340;
  assign _EVAL_68 = _EVAL_272[7:1];
  assign _EVAL_156 = {{1'd0}, _EVAL_68};
  assign _EVAL_120 = _EVAL_272 | _EVAL_156;
  assign _EVAL_295 = _EVAL_120[7:2];
  assign _EVAL_320 = {{2'd0}, _EVAL_295};
  assign _EVAL_279 = _EVAL_120 | _EVAL_320;
  assign _EVAL_220 = _EVAL_279[7:4];
  assign _EVAL_250 = {{4'd0}, _EVAL_220};
  assign _EVAL_372 = _EVAL_279 | _EVAL_250;
  assign _EVAL_176 = _EVAL_372[7:1];
  assign _EVAL_343 = {{1'd0}, _EVAL_176};
  assign _EVAL_210 = ~ _EVAL_272;
  assign _EVAL_384 = {_EVAL_210, 1'h0};
  assign _EVAL_330 = _EVAL_384[7:0];
  assign _EVAL_96 = _EVAL_210 | _EVAL_330;
  assign _EVAL_258 = {_EVAL_96, 2'h0};
  assign _EVAL_128 = _EVAL_258[7:0];
  assign _EVAL_223 = _EVAL_96 | _EVAL_128;
  assign _EVAL_322 = {_EVAL_223, 4'h0};
  assign _EVAL_301 = _EVAL_322[7:0];
  assign _EVAL_138 = _EVAL_223 | _EVAL_301;
  assign _EVAL_317 = ~ _EVAL_138;
  assign _EVAL_77 = _EVAL_343 | _EVAL_317;
  assign _EVAL_159 = _EVAL_211[9:2];
  assign _EVAL_146 = {_EVAL_159, 1'h0};
  assign _EVAL_286 = _EVAL_146[7:0];
  assign _EVAL_163 = _EVAL_159 | _EVAL_286;
  assign _EVAL_92 = {_EVAL_163, 2'h0};
  assign _EVAL_218 = _EVAL_92[7:0];
  assign _EVAL_304 = _EVAL_163 | _EVAL_218;
  assign _EVAL_240 = {_EVAL_304, 4'h0};
  assign _EVAL_299 = _EVAL_240[7:0];
  assign _EVAL_105 = _EVAL_304 | _EVAL_299;
  assign _EVAL_402 = ~ _EVAL_105;
  assign _EVAL_386 = _EVAL_77 & _EVAL_402;
  assign _EVAL_253 = _EVAL_211 ^ 32'h1000;
  assign _EVAL_173 = {1'b0,$signed(_EVAL_253)};
  assign _EVAL_327 = $signed(_EVAL_173) & $signed(33'sheb001000);
  assign _EVAL_316 = $signed(_EVAL_327);
  assign _EVAL_268 = $signed(_EVAL_316) == $signed(33'sh0);
  assign _EVAL_336 = _EVAL_268 ? 6'h3f : 6'h0;
  assign _EVAL_333 = _EVAL_211 ^ 32'h80000000;
  assign _EVAL_178 = {1'b0,$signed(_EVAL_333)};
  assign _EVAL_157 = $signed(_EVAL_178) & $signed(33'sheb000000);
  assign _EVAL_261 = $signed(_EVAL_157);
  assign _EVAL_193 = $signed(_EVAL_261) == $signed(33'sh0);
  assign _EVAL_109 = _EVAL_362 | _EVAL_193;
  assign _EVAL_318 = _EVAL_211 ^ 32'h8000000;
  assign _EVAL_260 = {1'b0,$signed(_EVAL_318)};
  assign _EVAL_209 = $signed(_EVAL_260) & $signed(33'she8000000);
  assign _EVAL_378 = $signed(_EVAL_209);
  assign _EVAL_127 = $signed(_EVAL_378) == $signed(33'sh0);
  assign _EVAL_217 = _EVAL_109 | _EVAL_127;
  assign _EVAL_385 = _EVAL_211 ^ 32'h2000000;
  assign _EVAL_335 = {1'b0,$signed(_EVAL_385)};
  assign _EVAL_143 = $signed(_EVAL_335) & $signed(33'sheb000000);
  assign _EVAL_148 = $signed(_EVAL_143);
  assign _EVAL_251 = $signed(_EVAL_148) == $signed(33'sh0);
  assign _EVAL_86 = _EVAL_217 | _EVAL_251;
  assign _EVAL_150 = _EVAL_86 | _EVAL_185;
  assign _EVAL_341 = _EVAL_211 ^ 32'h1000000;
  assign _EVAL_277 = {1'b0,$signed(_EVAL_341)};
  assign _EVAL_97 = $signed(_EVAL_277) & $signed(33'sheb000000);
  assign _EVAL_324 = $signed(_EVAL_97);
  assign _EVAL_351 = $signed(_EVAL_324) == $signed(33'sh0);
  assign _EVAL_137 = _EVAL_150 | _EVAL_351;
  assign _EVAL_200 = _EVAL_211 ^ 32'h20000000;
  assign _EVAL_151 = {1'b0,$signed(_EVAL_200)};
  assign _EVAL_241 = $signed(_EVAL_151) & $signed(33'sheb000000);
  assign _EVAL_228 = $signed(_EVAL_241);
  assign _EVAL_129 = $signed(_EVAL_228) == $signed(33'sh0);
  assign _EVAL_169 = _EVAL_137 | _EVAL_129;
  assign _EVAL_401 = _EVAL_169 ? 4'hf : 4'h0;
  assign _EVAL_289 = {{2'd0}, _EVAL_401};
  assign _EVAL_300 = _EVAL_336 | _EVAL_289;
  assign _EVAL_326 = {{2'd0}, _EVAL_300};
  assign _EVAL_332 = _EVAL_386 & _EVAL_326;
  assign _EVAL_347 = _EVAL_408 ? 8'h0 : _EVAL_332;
  assign _EVAL_215 = {_EVAL_347, 1'h0};
  assign _EVAL_107 = Queue__EVAL_3;
  assign _EVAL_181 = _EVAL_49 & _EVAL_107;
  assign _EVAL_363 = _EVAL_83 ? _EVAL_208 : 9'h0;
  assign _EVAL_265 = _EVAL_274 ? _EVAL_363 : _EVAL_407;
  assign _EVAL_331 = {{8'd0}, _EVAL_75};
  assign _EVAL_203 = _EVAL_265 - _EVAL_331;
  assign _EVAL_387 = {{16'd0}, _EVAL_344};
  assign _EVAL_161 = {{1'd0}, _EVAL_272};
  assign _EVAL_369 = _EVAL_215 | 9'h1;
  assign _EVAL_248 = {1'h0,_EVAL_347};
  assign _EVAL_339 = ~ _EVAL_248;
  assign _EVAL_88 = _EVAL_369 & _EVAL_339;
  assign _EVAL_244 = _EVAL_161 - _EVAL_88;
  assign _EVAL_230 = _EVAL_181 ? _EVAL_244 : {{1'd0}, _EVAL_172};
  assign _EVAL_78 = _EVAL_136 | _EVAL_38;
  assign _EVAL_141 = _EVAL_74 + _EVAL_387;
  assign _EVAL_130 = {{17'd0}, _EVAL_66};
  assign _EVAL_312 = _EVAL_141 & _EVAL_130;
  assign _EVAL_205 = ~ _EVAL_69;
  assign _EVAL_361 = _EVAL_205 | _EVAL_130;
  assign _EVAL_93 = ~ _EVAL_361;
  assign _EVAL_379 = _EVAL_312 | _EVAL_93;
  assign _EVAL_113 = _EVAL_274 | _EVAL_112;
  assign _EVAL_89 = _EVAL_398 & _EVAL_113;
  assign _EVAL_291 = _EVAL_28 & _EVAL_89;
  assign _EVAL_298 = 9'h3 << _EVAL_221;
  assign _EVAL_349 = _EVAL_298[1:0];
  assign _EVAL_224 = {{7'd0}, _EVAL_88};
  assign _EVAL_147 = _EVAL_224 << _EVAL_221;
  assign _EVAL_325 = {{16'd0}, _EVAL_147};
  assign _EVAL_119 = _EVAL_211 + _EVAL_325;
  assign _EVAL_346 = {_EVAL_340,8'hff};
  assign _EVAL_247 = {{7'd0}, _EVAL_346};
  assign _EVAL_281 = _EVAL_247 << _EVAL_221;
  assign _EVAL_399 = _EVAL_281[22:8];
  assign _EVAL_125 = {{17'd0}, _EVAL_399};
  assign _EVAL_202 = _EVAL_119 & _EVAL_125;
  assign _EVAL_355 = 4'h1 << _EVAL_54;
  assign _EVAL_225 = _EVAL_355[3];
  assign _EVAL_345 = _EVAL_170 == 1'h0;
  assign _EVAL_188 = _EVAL_18 | _EVAL_345;
  assign _EVAL_264 = _EVAL_188 & _EVAL_36;
  assign _EVAL_192 = _EVAL_225 & _EVAL_264;
  assign _EVAL_81 = _EVAL_355[2];
  assign _EVAL_116 = _EVAL_81 & _EVAL_264;
  assign _EVAL_198 = ~ _EVAL_211;
  assign _EVAL_110 = _EVAL_355[1];
  assign _EVAL_237 = _EVAL_110 & _EVAL_264;
  assign _EVAL_256 = _EVAL_356 | _EVAL_38;
  assign _EVAL_396 = ~ _EVAL_349;
  assign _EVAL_366 = {{30'd0}, _EVAL_396};
  assign _EVAL_403 = 2'h1 == _EVAL_54 ? _EVAL_356 : _EVAL_296;
  assign _EVAL_337 = 2'h2 == _EVAL_54 ? _EVAL_136 : _EVAL_403;
  assign _EVAL_342 = ~ _EVAL_267;
  assign _EVAL_155 = _EVAL_342 | _EVAL_125;
  assign _EVAL_377 = _EVAL_194 == 2'h2;
  assign _EVAL_313 = ~ _EVAL_155;
  assign _EVAL_364 = _EVAL_202 | _EVAL_313;
  assign _EVAL_239 = _EVAL_347 == _EVAL_272;
  assign _EVAL_114 = _EVAL_239 == 1'h0;
  assign _EVAL_236 = _EVAL_83 & _EVAL_274;
  assign _EVAL_189 = _EVAL_198 | _EVAL_366;
  assign _EVAL_245 = 2'h3 == _EVAL_54 ? _EVAL_101 : _EVAL_337;
  assign _EVAL_115 = _EVAL_238 == 2'h2;
  assign _EVAL_65 = _EVAL_355[0];
  assign _EVAL_153 = _EVAL_28 & _EVAL_113;
  assign _EVAL_166 = _EVAL_153 & _EVAL_398;
  assign _EVAL_371 = _EVAL_212 - _EVAL_208;
  assign _EVAL_142 = _EVAL_166 ? _EVAL_371 : {{1'd0}, _EVAL_132};
  assign _EVAL_171 = Queue_1__EVAL_2;
  assign _EVAL_164 = _EVAL_65 & _EVAL_264;
  assign _EVAL_168 = Queue__EVAL_2;
  assign _EVAL_328 = _EVAL_126 == _EVAL_73;
  assign _EVAL_67 = _EVAL_328 == 1'h0;
  assign _EVAL_280 = _EVAL_63[0];
  assign Queue_1__EVAL_13 = _EVAL_153 & _EVAL_328;
  assign Queue_1__EVAL_1 = _EVAL_22;
  assign Queue_2__EVAL_9 = _EVAL_26;
  assign _EVAL_44 = _EVAL_18 | _EVAL_345;
  assign _EVAL_16 = _EVAL_43;
  assign _EVAL_0 = _EVAL_219 & _EVAL_394;
  assign Queue__EVAL_11 = _EVAL_57;
  assign Queue__EVAL_0 = _EVAL_24;
  assign Queue_1__EVAL_0 = _EVAL_59;
  assign _EVAL_23 = Queue__EVAL_6;
  assign _EVAL_32 = _EVAL_265 == 9'h1;
  assign _EVAL_21 = ~ _EVAL_189;
  assign _EVAL_61 = _EVAL_5 & _EVAL_280;
  assign Queue_1__EVAL_4 = _EVAL_6;
  assign Queue_1__EVAL_10 = _EVAL_1;
  assign Queue__EVAL_13 = _EVAL_49 & _EVAL_239;
  assign Queue__EVAL_14 = _EVAL_45;
  assign _EVAL_48 = _EVAL_398 & _EVAL_113;
  assign _EVAL_35 = _EVAL_8;
  assign _EVAL_29 = Queue_2__EVAL_6;
  assign Queue_2__EVAL_0 = _EVAL_7;
  assign _EVAL_14 = Queue__EVAL;
  assign _EVAL_33 = _EVAL_47;
  assign _EVAL_15 = _EVAL_54;
  assign _EVAL_56 = Queue_2__EVAL_10;
  assign Queue__EVAL_15 = _EVAL_11;
  assign _EVAL_55 = Queue_1__EVAL_6;
  assign Queue_2__EVAL_4 = _EVAL_60 & _EVAL_394;
  assign Queue_2__EVAL_3 = _EVAL_31;
  assign Queue_1__EVAL_14 = _EVAL_62;
  assign _EVAL_19 = _EVAL_17;
  assign _EVAL_41 = _EVAL_63[6:1];
  assign _EVAL_4 = Queue_1__EVAL_5;
  assign _EVAL_40 = Queue__EVAL_5;
  assign Queue_2__EVAL_5 = _EVAL_1;
  assign _EVAL_46 = _EVAL_39[6:1];
  assign _EVAL_13 = _EVAL_38 | _EVAL_245;
  assign Queue_2__EVAL_8 = _EVAL_30;
  assign _EVAL_37 = Queue_1__EVAL;
  assign Queue__EVAL_4 = _EVAL_27;
  assign _EVAL_10 = {_EVAL_171,_EVAL_328};
  assign Queue_1__EVAL_11 = _EVAL_53;
  assign Queue_2__EVAL_2 = _EVAL_25;
  assign Queue_1__EVAL_15 = _EVAL_64;
  assign _EVAL_34 = Queue_2__EVAL_1;
  assign Queue__EVAL_1 = _EVAL_20;
  assign _EVAL_2 = ~ _EVAL_309;
  assign _EVAL_3 = {_EVAL_168,_EVAL_239};
  assign _EVAL_50 = Queue__EVAL_3;
  assign Queue__EVAL_16 = _EVAL_26;
  assign _EVAL_12 = _EVAL_408 ? 8'h0 : _EVAL_332;
  assign Queue_1__EVAL_9 = _EVAL_58;
  assign Queue__EVAL_9 = _EVAL_9;
  assign Queue_1__EVAL_16 = _EVAL_26;
  assign Queue__EVAL_10 = _EVAL_1;
  assign _EVAL = _EVAL_36 & _EVAL_170;
  assign _EVAL_52 = _EVAL_51;
  assign _EVAL_42 = _EVAL_177 ? 8'h0 : _EVAL_183;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_71 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_101 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_112 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_132 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_136 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_172 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_182 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_213 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_229 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_296 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_356 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_407 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_1) begin
    if (_EVAL_181) begin
      if (_EVAL_381) begin
        _EVAL_71 <= _EVAL_267;
      end else begin
        if (_EVAL_377) begin
          _EVAL_71 <= _EVAL_364;
        end else begin
          _EVAL_71 <= _EVAL_119;
        end
      end
    end
    if (_EVAL_26) begin
      _EVAL_101 <= 2'h0;
    end else begin
      if (_EVAL_192) begin
        if (_EVAL_170) begin
          _EVAL_101 <= 2'h0;
        end else begin
          _EVAL_101 <= _EVAL_252;
        end
      end
    end
    if (_EVAL_26) begin
      _EVAL_112 <= 1'h0;
    end else begin
      if (_EVAL_291) begin
        _EVAL_112 <= 1'h0;
      end else begin
        if (_EVAL_236) begin
          _EVAL_112 <= 1'h1;
        end
      end
    end
    _EVAL_132 <= _EVAL_142[7:0];
    if (_EVAL_26) begin
      _EVAL_136 <= 2'h0;
    end else begin
      if (_EVAL_116) begin
        if (_EVAL_170) begin
          _EVAL_136 <= 2'h0;
        end else begin
          _EVAL_136 <= _EVAL_78;
        end
      end
    end
    _EVAL_172 <= _EVAL_230[7:0];
    if (_EVAL_26) begin
      _EVAL_182 <= 1'h0;
    end else begin
      if (_EVAL_181) begin
        _EVAL_182 <= _EVAL_114;
      end
    end
    if (_EVAL_166) begin
      if (_EVAL_134) begin
        _EVAL_213 <= _EVAL_69;
      end else begin
        if (_EVAL_115) begin
          _EVAL_213 <= _EVAL_379;
        end else begin
          _EVAL_213 <= _EVAL_141;
        end
      end
    end
    if (_EVAL_26) begin
      _EVAL_229 <= 1'h0;
    end else begin
      if (_EVAL_166) begin
        _EVAL_229 <= _EVAL_67;
      end
    end
    if (_EVAL_26) begin
      _EVAL_296 <= 2'h0;
    end else begin
      if (_EVAL_164) begin
        if (_EVAL_170) begin
          _EVAL_296 <= 2'h0;
        end else begin
          _EVAL_296 <= _EVAL_191;
        end
      end
    end
    if (_EVAL_26) begin
      _EVAL_356 <= 2'h0;
    end else begin
      if (_EVAL_237) begin
        if (_EVAL_170) begin
          _EVAL_356 <= 2'h0;
        end else begin
          _EVAL_356 <= _EVAL_256;
        end
      end
    end
    if (_EVAL_26) begin
      _EVAL_407 <= 9'h0;
    end else begin
      _EVAL_407 <= _EVAL_203;
    end
  end
endmodule
