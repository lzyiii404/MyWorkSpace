//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_102_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [7:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_19;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_41;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_82;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_90;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_98;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_103;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_131;
  reg [31:0] _RAND_6;
  reg  _EVAL_158;
  reg [31:0] _RAND_7;
  reg  _EVAL_181;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_195;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_205;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_225;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_249;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_269;
  reg [31:0] _RAND_13;
  reg  _EVAL_283;
  reg [31:0] _RAND_14;
  wire  _EVAL_266;
  wire [1:0] _EVAL_245;
  wire [3:0] _EVAL_244;
  wire [2:0] _EVAL_85;
  wire [2:0] _EVAL_128;
  wire  _EVAL_233;
  wire  _EVAL_65;
  wire  _EVAL_118;
  wire  _EVAL_25;
  wire  _EVAL_216;
  wire  _EVAL_93;
  wire  _EVAL_68;
  wire  _EVAL_262;
  wire  _EVAL_36;
  wire  _EVAL_276;
  wire  _EVAL_72;
  wire  _EVAL_282;
  wire  _EVAL_28;
  wire  _EVAL_213;
  wire  _EVAL_175;
  wire  _EVAL_220;
  wire  _EVAL_212;
  wire  _EVAL_60;
  wire  _EVAL_201;
  wire  _EVAL_214;
  wire  _EVAL_58;
  wire  _EVAL_134;
  wire  _EVAL_116;
  wire  _EVAL_44;
  wire  _EVAL_176;
  wire  _EVAL_112;
  wire  _EVAL_243;
  wire  _EVAL_239;
  wire  _EVAL_187;
  wire  _EVAL_32;
  wire  _EVAL_259;
  wire  _EVAL_241;
  wire  _EVAL_53;
  wire  _EVAL_240;
  wire  _EVAL_135;
  wire  _EVAL_235;
  wire  _EVAL_149;
  wire [1:0] _EVAL_101;
  wire [1:0] _EVAL_22;
  wire [1:0] _EVAL_86;
  wire [1:0] _EVAL_96;
  wire  _EVAL_224;
  wire  _EVAL_57;
  wire  _EVAL_219;
  wire  _EVAL_33;
  wire [12:0] _EVAL_236;
  wire [5:0] _EVAL_207;
  wire [5:0] _EVAL_43;
  wire [31:0] _EVAL_199;
  wire [31:0] _EVAL_66;
  wire  _EVAL_150;
  wire  _EVAL_141;
  wire  _EVAL_48;
  wire  _EVAL_156;
  wire  _EVAL_268;
  wire  _EVAL_143;
  wire [1:0] _EVAL_162;
  wire [1:0] _EVAL_61;
  wire  _EVAL_140;
  wire  _EVAL_67;
  wire  _EVAL_153;
  wire  _EVAL_121;
  wire  _EVAL_280;
  wire  _EVAL_94;
  wire  _EVAL_49;
  wire  _EVAL_200;
  wire  _EVAL_139;
  wire [31:0] _EVAL_281;
  wire  _EVAL_229;
  wire [12:0] _EVAL_27;
  wire [5:0] _EVAL_70;
  wire [5:0] _EVAL_79;
  wire [2:0] _EVAL_26;
  wire [2:0] _EVAL_73;
  wire  _EVAL_104;
  wire  _EVAL_186;
  wire  _EVAL_91;
  wire  _EVAL_29;
  wire  _EVAL_109;
  wire  _EVAL_211;
  wire  _EVAL_50;
  wire  _EVAL_238;
  wire [2:0] _EVAL_267;
  wire [2:0] _EVAL_237;
  wire  _EVAL_100;
  wire  _EVAL_260;
  wire  _EVAL_127;
  wire  _EVAL_88;
  wire  _EVAL_144;
  wire  _EVAL_102;
  wire  _EVAL_51;
  wire  _EVAL_136;
  wire  _EVAL_166;
  wire  _EVAL_20;
  wire  _EVAL_167;
  wire  _EVAL_59;
  wire  _EVAL_228;
  wire  _EVAL_99;
  wire  _EVAL_80;
  wire  _EVAL_274;
  wire  _EVAL_23;
  wire  _EVAL_163;
  wire  _EVAL_115;
  wire  _EVAL_246;
  wire  _EVAL_35;
  wire  _EVAL_114;
  wire  _EVAL_89;
  wire  _EVAL_75;
  wire  _EVAL_34;
  wire  _EVAL_168;
  wire [7:0] _EVAL_226;
  wire [7:0] _EVAL_189;
  wire [7:0] _EVAL_203;
  wire [1:0] _EVAL_137;
  wire  _EVAL_180;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_151;
  wire  _EVAL_173;
  wire  _EVAL_210;
  wire  _EVAL_160;
  wire  _EVAL_227;
  wire  _EVAL_170;
  wire  _EVAL_263;
  wire  _EVAL_230;
  wire  _EVAL_64;
  wire  _EVAL_184;
  wire  _EVAL_258;
  wire  _EVAL_106;
  wire  _EVAL_159;
  wire  _EVAL_47;
  wire  _EVAL_146;
  wire  _EVAL_87;
  wire  _EVAL_39;
  wire  _EVAL_161;
  wire  _EVAL_275;
  wire  _EVAL_196;
  wire  _EVAL_279;
  wire  _EVAL_261;
  wire  _EVAL_97;
  wire  _EVAL_74;
  wire  _EVAL_251;
  wire  _EVAL_172;
  wire [7:0] _EVAL_54;
  wire  _EVAL_253;
  wire  _EVAL_217;
  wire  _EVAL_209;
  wire  _EVAL_24;
  wire  _EVAL_111;
  wire  _EVAL_171;
  wire  _EVAL_18;
  wire  _EVAL_174;
  wire  _EVAL_63;
  wire  _EVAL_133;
  wire  _EVAL_117;
  wire  _EVAL_154;
  wire  _EVAL_165;
  wire [31:0] _EVAL_31;
  wire [32:0] _EVAL_108;
  wire [32:0] _EVAL_105;
  wire [32:0] _EVAL_130;
  wire  _EVAL_126;
  wire  _EVAL_92;
  wire  _EVAL_157;
  wire [2:0] _EVAL_257;
  wire  _EVAL_232;
  wire  _EVAL_84;
  wire  _EVAL_129;
  wire  _EVAL_147;
  wire  _EVAL_37;
  wire  _EVAL_271;
  wire  _EVAL_190;
  wire  _EVAL_152;
  wire  _EVAL_132;
  wire  _EVAL_142;
  wire  _EVAL_204;
  wire  _EVAL_215;
  wire  _EVAL_234;
  wire  _EVAL_198;
  wire  _EVAL_38;
  wire  _EVAL_193;
  wire  _EVAL_17;
  wire  _EVAL_145;
  wire  _EVAL_202;
  wire  _EVAL_81;
  wire  _EVAL_247;
  wire  _EVAL_265;
  wire  _EVAL_78;
  wire  _EVAL_69;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_188;
  wire [1:0] _EVAL_191;
  wire  _EVAL_273;
  wire  _EVAL_148;
  wire  _EVAL_113;
  wire  _EVAL_223;
  wire  _EVAL_192;
  wire  _EVAL_155;
  wire  _EVAL_264;
  wire  _EVAL_250;
  wire  _EVAL_242;
  wire [1:0] _EVAL_208;
  wire  _EVAL_83;
  wire  _EVAL_123;
  wire  _EVAL_177;
  wire  _EVAL_71;
  wire [1:0] _EVAL_52;
  wire  _EVAL_179;
  wire  _EVAL_30;
  wire  _EVAL_272;
  wire  _EVAL_46;
  wire  _EVAL_182;
  wire  _EVAL_231;
  wire [2:0] _EVAL_252;
  wire  _EVAL_164;
  wire  _EVAL_62;
  wire  _EVAL_56;
  wire  _EVAL_194;
  wire  _EVAL_40;
  wire  _EVAL_277;
  wire  _EVAL_21;
  wire  _EVAL_76;
  wire  _EVAL_124;
  wire  _EVAL_42;
  wire  _EVAL_95;
  wire  _EVAL_248;
  wire  _EVAL_77;
  wire  _EVAL_221;
  wire  _EVAL_278;
  wire  _EVAL_178;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_266 = _EVAL_11 >= 3'h3;
  assign _EVAL_245 = _EVAL_11[1:0];
  assign _EVAL_244 = 4'h1 << _EVAL_245;
  assign _EVAL_85 = _EVAL_244[2:0];
  assign _EVAL_128 = _EVAL_85 | 3'h1;
  assign _EVAL_233 = _EVAL_128[2];
  assign _EVAL_65 = _EVAL_7[2];
  assign _EVAL_118 = _EVAL_65 == 1'h0;
  assign _EVAL_25 = _EVAL_233 & _EVAL_118;
  assign _EVAL_216 = _EVAL_266 | _EVAL_25;
  assign _EVAL_93 = _EVAL_128[1];
  assign _EVAL_68 = _EVAL_7[1];
  assign _EVAL_262 = _EVAL_118 & _EVAL_68;
  assign _EVAL_36 = _EVAL_93 & _EVAL_262;
  assign _EVAL_276 = _EVAL_216 | _EVAL_36;
  assign _EVAL_72 = _EVAL_128[0];
  assign _EVAL_282 = _EVAL_7[0];
  assign _EVAL_28 = _EVAL_282 == 1'h0;
  assign _EVAL_213 = _EVAL_262 & _EVAL_28;
  assign _EVAL_175 = _EVAL_72 & _EVAL_213;
  assign _EVAL_220 = _EVAL_276 | _EVAL_175;
  assign _EVAL_212 = _EVAL_15 == 3'h2;
  assign _EVAL_60 = _EVAL_3 == 3'h5;
  assign _EVAL_201 = _EVAL_65 & _EVAL_68;
  assign _EVAL_214 = _EVAL_201 & _EVAL_28;
  assign _EVAL_58 = _EVAL_3 == 3'h2;
  assign _EVAL_134 = _EVAL_6 & _EVAL_58;
  assign _EVAL_116 = _EVAL_98 != 2'h0;
  assign _EVAL_44 = _EVAL_116 == 1'h0;
  assign _EVAL_176 = plusarg_reader_out == 32'h0;
  assign _EVAL_112 = _EVAL_44 | _EVAL_176;
  assign _EVAL_243 = _EVAL_225 < plusarg_reader_out;
  assign _EVAL_239 = _EVAL_112 | _EVAL_243;
  assign _EVAL_187 = _EVAL_239 | _EVAL_9;
  assign _EVAL_32 = _EVAL_187 == 1'h0;
  assign _EVAL_259 = _EVAL_68 == 1'h0;
  assign _EVAL_241 = _EVAL_65 & _EVAL_259;
  assign _EVAL_53 = _EVAL_16 == 1'h0;
  assign _EVAL_240 = _EVAL_53 | _EVAL_9;
  assign _EVAL_135 = _EVAL_13 & _EVAL_6;
  assign _EVAL_235 = _EVAL_269 == 3'h0;
  assign _EVAL_149 = _EVAL_135 & _EVAL_235;
  assign _EVAL_101 = 2'h1 << _EVAL_4;
  assign _EVAL_22 = _EVAL_149 ? _EVAL_101 : 2'h0;
  assign _EVAL_86 = _EVAL_22 | _EVAL_98;
  assign _EVAL_96 = _EVAL_86 >> _EVAL_0;
  assign _EVAL_224 = _EVAL_96[0];
  assign _EVAL_57 = _EVAL_224 | _EVAL_9;
  assign _EVAL_219 = _EVAL_3 == 3'h6;
  assign _EVAL_33 = _EVAL_6 & _EVAL_219;
  assign _EVAL_236 = 13'h3f << _EVAL_11;
  assign _EVAL_207 = _EVAL_236[5:0];
  assign _EVAL_43 = ~ _EVAL_207;
  assign _EVAL_199 = {{26'd0}, _EVAL_43};
  assign _EVAL_66 = _EVAL_7 & _EVAL_199;
  assign _EVAL_150 = _EVAL_8 & _EVAL_5;
  assign _EVAL_141 = _EVAL_205 == 3'h0;
  assign _EVAL_48 = _EVAL_150 & _EVAL_141;
  assign _EVAL_156 = _EVAL_15 == 3'h6;
  assign _EVAL_268 = _EVAL_156 == 1'h0;
  assign _EVAL_143 = _EVAL_48 & _EVAL_268;
  assign _EVAL_162 = 2'h1 << _EVAL_0;
  assign _EVAL_61 = _EVAL_143 ? _EVAL_162 : 2'h0;
  assign _EVAL_140 = _EVAL_241 & _EVAL_282;
  assign _EVAL_67 = _EVAL_72 & _EVAL_140;
  assign _EVAL_153 = _EVAL_15 == _EVAL_82;
  assign _EVAL_121 = _EVAL_153 | _EVAL_9;
  assign _EVAL_280 = _EVAL_121 == 1'h0;
  assign _EVAL_94 = _EVAL_1 <= 3'h2;
  assign _EVAL_49 = _EVAL_94 | _EVAL_9;
  assign _EVAL_200 = _EVAL_49 == 1'h0;
  assign _EVAL_139 = _EVAL_135 | _EVAL_150;
  assign _EVAL_281 = _EVAL_225 + 32'h1;
  assign _EVAL_229 = _EVAL_15[0];
  assign _EVAL_27 = 13'h3f << _EVAL_10;
  assign _EVAL_70 = _EVAL_27[5:0];
  assign _EVAL_79 = ~ _EVAL_70;
  assign _EVAL_26 = _EVAL_79[5:3];
  assign _EVAL_73 = _EVAL_205 - 3'h1;
  assign _EVAL_104 = _EVAL_12 == _EVAL_283;
  assign _EVAL_186 = _EVAL_104 | _EVAL_9;
  assign _EVAL_91 = _EVAL_118 & _EVAL_259;
  assign _EVAL_29 = _EVAL_91 & _EVAL_28;
  assign _EVAL_109 = _EVAL_72 & _EVAL_29;
  assign _EVAL_211 = _EVAL_15 == 3'h5;
  assign _EVAL_50 = _EVAL_3[2];
  assign _EVAL_238 = _EVAL_50 == 1'h0;
  assign _EVAL_267 = _EVAL_43[5:3];
  assign _EVAL_237 = _EVAL_269 - 3'h1;
  assign _EVAL_100 = _EVAL_266 | _EVAL_9;
  assign _EVAL_260 = _EVAL_100 == 1'h0;
  assign _EVAL_127 = _EVAL_233 & _EVAL_65;
  assign _EVAL_88 = _EVAL_266 | _EVAL_127;
  assign _EVAL_144 = _EVAL_93 & _EVAL_201;
  assign _EVAL_102 = _EVAL_88 | _EVAL_144;
  assign _EVAL_51 = _EVAL_201 & _EVAL_282;
  assign _EVAL_136 = _EVAL_72 & _EVAL_51;
  assign _EVAL_166 = _EVAL_102 | _EVAL_136;
  assign _EVAL_20 = _EVAL_72 & _EVAL_214;
  assign _EVAL_167 = _EVAL_102 | _EVAL_20;
  assign _EVAL_59 = _EVAL_93 & _EVAL_241;
  assign _EVAL_228 = _EVAL_88 | _EVAL_59;
  assign _EVAL_99 = _EVAL_228 | _EVAL_67;
  assign _EVAL_80 = _EVAL_241 & _EVAL_28;
  assign _EVAL_274 = _EVAL_72 & _EVAL_80;
  assign _EVAL_23 = _EVAL_228 | _EVAL_274;
  assign _EVAL_163 = _EVAL_262 & _EVAL_282;
  assign _EVAL_115 = _EVAL_72 & _EVAL_163;
  assign _EVAL_246 = _EVAL_276 | _EVAL_115;
  assign _EVAL_35 = _EVAL_93 & _EVAL_91;
  assign _EVAL_114 = _EVAL_216 | _EVAL_35;
  assign _EVAL_89 = _EVAL_91 & _EVAL_282;
  assign _EVAL_75 = _EVAL_72 & _EVAL_89;
  assign _EVAL_34 = _EVAL_114 | _EVAL_75;
  assign _EVAL_168 = _EVAL_114 | _EVAL_109;
  assign _EVAL_226 = {_EVAL_166,_EVAL_167,_EVAL_99,_EVAL_23,_EVAL_246,_EVAL_220,_EVAL_34,_EVAL_168};
  assign _EVAL_189 = ~ _EVAL_226;
  assign _EVAL_203 = _EVAL_14 & _EVAL_189;
  assign _EVAL_137 = _EVAL_98 >> _EVAL_4;
  assign _EVAL_180 = _EVAL_7 == _EVAL_19;
  assign _EVAL_255 = _EVAL_180 | _EVAL_9;
  assign _EVAL_256 = _EVAL_15 == 3'h0;
  assign _EVAL_151 = _EVAL_5 & _EVAL_256;
  assign _EVAL_173 = _EVAL_10 == _EVAL_131;
  assign _EVAL_210 = _EVAL_173 | _EVAL_9;
  assign _EVAL_160 = _EVAL_210 == 1'h0;
  assign _EVAL_227 = _EVAL_15 == 3'h4;
  assign _EVAL_170 = _EVAL_3 == 3'h4;
  assign _EVAL_263 = _EVAL_0 == _EVAL_181;
  assign _EVAL_230 = _EVAL_263 | _EVAL_9;
  assign _EVAL_64 = _EVAL_230 == 1'h0;
  assign _EVAL_184 = _EVAL_4 == _EVAL_158;
  assign _EVAL_258 = _EVAL_184 | _EVAL_9;
  assign _EVAL_106 = _EVAL_258 == 1'h0;
  assign _EVAL_159 = _EVAL == 1'h0;
  assign _EVAL_47 = _EVAL_1 == _EVAL_41;
  assign _EVAL_146 = _EVAL_11 <= 3'h6;
  assign _EVAL_87 = _EVAL_1 <= 3'h3;
  assign _EVAL_39 = _EVAL_87 | _EVAL_9;
  assign _EVAL_161 = _EVAL_39 == 1'h0;
  assign _EVAL_275 = _EVAL_22 != _EVAL_61;
  assign _EVAL_196 = _EVAL_22 != 2'h0;
  assign _EVAL_279 = _EVAL_196 == 1'h0;
  assign _EVAL_261 = _EVAL_275 | _EVAL_279;
  assign _EVAL_97 = _EVAL_261 | _EVAL_9;
  assign _EVAL_74 = _EVAL_11 == _EVAL_249;
  assign _EVAL_251 = _EVAL_137[0];
  assign _EVAL_172 = _EVAL_251 == 1'h0;
  assign _EVAL_54 = ~ _EVAL_14;
  assign _EVAL_253 = _EVAL_54 == 8'h0;
  assign _EVAL_217 = _EVAL_253 | _EVAL_9;
  assign _EVAL_209 = _EVAL_5 & _EVAL_227;
  assign _EVAL_24 = _EVAL_97 == 1'h0;
  assign _EVAL_111 = _EVAL_1 != 3'h0;
  assign _EVAL_171 = _EVAL_111 | _EVAL_9;
  assign _EVAL_18 = _EVAL_171 == 1'h0;
  assign _EVAL_174 = _EVAL_57 == 1'h0;
  assign _EVAL_63 = _EVAL_3 == _EVAL_103;
  assign _EVAL_133 = _EVAL_90 == 3'h0;
  assign _EVAL_117 = _EVAL_203 == 8'h0;
  assign _EVAL_154 = _EVAL_1 <= 3'h4;
  assign _EVAL_165 = _EVAL_5 & _EVAL_212;
  assign _EVAL_31 = _EVAL_7 ^ 32'h80000000;
  assign _EVAL_108 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_105 = $signed(_EVAL_108) & $signed(-33'sh20000);
  assign _EVAL_130 = $signed(_EVAL_105);
  assign _EVAL_126 = $signed(_EVAL_130) == $signed(33'sh0);
  assign _EVAL_92 = _EVAL_3 == 3'h3;
  assign _EVAL_157 = _EVAL_195 == 3'h0;
  assign _EVAL_257 = _EVAL_195 - 3'h1;
  assign _EVAL_232 = _EVAL_15 <= 3'h6;
  assign _EVAL_84 = _EVAL_232 | _EVAL_9;
  assign _EVAL_129 = _EVAL_217 == 1'h0;
  assign _EVAL_147 = _EVAL_5 & _EVAL_156;
  assign _EVAL_37 = _EVAL_3 == 3'h1;
  assign _EVAL_271 = _EVAL_6 & _EVAL_37;
  assign _EVAL_190 = _EVAL_146 & _EVAL_126;
  assign _EVAL_152 = _EVAL_190 | _EVAL_9;
  assign _EVAL_132 = _EVAL_152 == 1'h0;
  assign _EVAL_142 = _EVAL_63 | _EVAL_9;
  assign _EVAL_204 = _EVAL_142 == 1'h0;
  assign _EVAL_215 = _EVAL_66 == 32'h0;
  assign _EVAL_234 = _EVAL_84 == 1'h0;
  assign _EVAL_198 = _EVAL_255 == 1'h0;
  assign _EVAL_38 = _EVAL_154 | _EVAL_9;
  assign _EVAL_193 = _EVAL_157 == 1'h0;
  assign _EVAL_17 = _EVAL_6 & _EVAL_193;
  assign _EVAL_145 = _EVAL_14 == _EVAL_226;
  assign _EVAL_202 = _EVAL_3 == 3'h0;
  assign _EVAL_81 = _EVAL_6 & _EVAL_202;
  assign _EVAL_247 = _EVAL_9 == 1'h0;
  assign _EVAL_265 = _EVAL_6 & _EVAL_60;
  assign _EVAL_78 = _EVAL_1 == 3'h0;
  assign _EVAL_69 = _EVAL_10 >= 3'h3;
  assign _EVAL_119 = _EVAL_69 | _EVAL_9;
  assign _EVAL_120 = _EVAL_119 == 1'h0;
  assign _EVAL_188 = _EVAL_5 & _EVAL_211;
  assign _EVAL_191 = ~ _EVAL_61;
  assign _EVAL_273 = _EVAL_3 == 3'h7;
  assign _EVAL_148 = _EVAL_47 | _EVAL_9;
  assign _EVAL_113 = _EVAL_148 == 1'h0;
  assign _EVAL_223 = _EVAL_12 == 1'h0;
  assign _EVAL_192 = _EVAL_223 | _EVAL_9;
  assign _EVAL_155 = _EVAL_192 == 1'h0;
  assign _EVAL_264 = _EVAL_223 | _EVAL_16;
  assign _EVAL_250 = _EVAL_117 | _EVAL_9;
  assign _EVAL_242 = _EVAL_250 == 1'h0;
  assign _EVAL_208 = _EVAL_98 | _EVAL_22;
  assign _EVAL_83 = _EVAL_264 | _EVAL_9;
  assign _EVAL_123 = _EVAL_83 == 1'h0;
  assign _EVAL_177 = _EVAL_150 & _EVAL_133;
  assign _EVAL_71 = _EVAL_159 | _EVAL_9;
  assign _EVAL_52 = _EVAL_208 & _EVAL_191;
  assign _EVAL_179 = _EVAL_6 & _EVAL_170;
  assign _EVAL_30 = _EVAL_71 == 1'h0;
  assign _EVAL_272 = _EVAL_15 == 3'h1;
  assign _EVAL_46 = _EVAL_172 | _EVAL_9;
  assign _EVAL_182 = _EVAL_46 == 1'h0;
  assign _EVAL_231 = _EVAL_135 & _EVAL_157;
  assign _EVAL_252 = _EVAL_90 - 3'h1;
  assign _EVAL_164 = _EVAL_78 | _EVAL_9;
  assign _EVAL_62 = _EVAL_164 == 1'h0;
  assign _EVAL_56 = _EVAL_6 & _EVAL_92;
  assign _EVAL_194 = _EVAL_133 == 1'h0;
  assign _EVAL_40 = _EVAL_5 & _EVAL_194;
  assign _EVAL_277 = _EVAL_240 == 1'h0;
  assign _EVAL_21 = _EVAL_6 & _EVAL_273;
  assign _EVAL_76 = _EVAL_74 | _EVAL_9;
  assign _EVAL_124 = _EVAL_76 == 1'h0;
  assign _EVAL_42 = _EVAL_186 == 1'h0;
  assign _EVAL_95 = _EVAL_215 | _EVAL_9;
  assign _EVAL_248 = _EVAL_95 == 1'h0;
  assign _EVAL_77 = _EVAL_5 & _EVAL_272;
  assign _EVAL_221 = _EVAL_38 == 1'h0;
  assign _EVAL_278 = _EVAL_145 | _EVAL_9;
  assign _EVAL_178 = _EVAL_278 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_19 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_41 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_82 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_90 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_98 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_103 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_131 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_158 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_181 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_195 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_205 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_225 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_249 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_269 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_283 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_231) begin
      _EVAL_19 <= _EVAL_7;
    end
    if (_EVAL_231) begin
      _EVAL_41 <= _EVAL_1;
    end
    if (_EVAL_177) begin
      _EVAL_82 <= _EVAL_15;
    end
    if (_EVAL_9) begin
      _EVAL_90 <= 3'h0;
    end else begin
      if (_EVAL_150) begin
        if (_EVAL_133) begin
          if (_EVAL_229) begin
            _EVAL_90 <= _EVAL_26;
          end else begin
            _EVAL_90 <= 3'h0;
          end
        end else begin
          _EVAL_90 <= _EVAL_252;
        end
      end
    end
    if (_EVAL_9) begin
      _EVAL_98 <= 2'h0;
    end else begin
      _EVAL_98 <= _EVAL_52;
    end
    if (_EVAL_231) begin
      _EVAL_103 <= _EVAL_3;
    end
    if (_EVAL_177) begin
      _EVAL_131 <= _EVAL_10;
    end
    if (_EVAL_231) begin
      _EVAL_158 <= _EVAL_4;
    end
    if (_EVAL_177) begin
      _EVAL_181 <= _EVAL_0;
    end
    if (_EVAL_9) begin
      _EVAL_195 <= 3'h0;
    end else begin
      if (_EVAL_135) begin
        if (_EVAL_157) begin
          if (_EVAL_238) begin
            _EVAL_195 <= _EVAL_267;
          end else begin
            _EVAL_195 <= 3'h0;
          end
        end else begin
          _EVAL_195 <= _EVAL_257;
        end
      end
    end
    if (_EVAL_9) begin
      _EVAL_205 <= 3'h0;
    end else begin
      if (_EVAL_150) begin
        if (_EVAL_141) begin
          if (_EVAL_229) begin
            _EVAL_205 <= _EVAL_26;
          end else begin
            _EVAL_205 <= 3'h0;
          end
        end else begin
          _EVAL_205 <= _EVAL_73;
        end
      end
    end
    if (_EVAL_9) begin
      _EVAL_225 <= 32'h0;
    end else begin
      if (_EVAL_139) begin
        _EVAL_225 <= 32'h0;
      end else begin
        _EVAL_225 <= _EVAL_281;
      end
    end
    if (_EVAL_231) begin
      _EVAL_249 <= _EVAL_11;
    end
    if (_EVAL_9) begin
      _EVAL_269 <= 3'h0;
    end else begin
      if (_EVAL_135) begin
        if (_EVAL_235) begin
          if (_EVAL_238) begin
            _EVAL_269 <= _EVAL_267;
          end else begin
            _EVAL_269 <= 3'h0;
          end
        end else begin
          _EVAL_269 <= _EVAL_237;
        end
      end
    end
    if (_EVAL_177) begin
      _EVAL_283 <= _EVAL_12;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17b82870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a31061ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d5aceaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cee40c88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c7a12ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84b04a5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa756c83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a9ec047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc052cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6230477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60ace749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b26d2f75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8ba476)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e475088)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41fe89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff63c5a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c448c8d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7338ad5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16a47fae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce79cc75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac3e0bde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93bb9d07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7d30f33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28d6351e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edcf9636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e9842b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51495ccb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ce811f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d81781d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73dd17e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90c6b80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c089d00e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e5a55ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2d7195e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70f68c1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4500353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cb4b93d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cc69ae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a15576)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(156be40b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(166be2cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b85c6f47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e9fcdab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8923a66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cf0fe99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49344fc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6081fc4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b05c5fd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(535b8b89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e2b970e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db61aeb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff7d121f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2474456c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41c11a0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdf90d22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a40acacc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(368a79c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86758aa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f664afb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5dd2ad0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52186f06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa88c781)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(729c9205)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6ca1bff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df91ed32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65dfb62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
