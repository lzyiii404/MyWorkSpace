//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_273_assert(
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_7,
  input  [3:0]  _EVAL_12,
  input         _EVAL_17,
  input  [3:0]  _EVAL_22,
  input         _EVAL_23,
  input  [3:0]  _EVAL_26,
  input         _EVAL_29,
  input         _EVAL_42,
  input  [2:0]  _EVAL_56,
  input  [31:0] _EVAL_62,
  input         _EVAL_67,
  input  [2:0]  _EVAL_69,
  input  [31:0] _EVAL_71,
  input  [2:0]  _EVAL_74,
  input  [2:0]  _EVAL_82,
  input         _EVAL_96,
  input  [7:0]  _EVAL_100,
  input         _EVAL_104,
  input  [3:0]  _EVAL_106,
  input         RationalCrossingSource_2__EVAL_3,
  input         RationalCrossingSource_1__EVAL_1,
  input  [1:0]  RationalCrossingSink__EVAL_21,
  input         RationalCrossingSink__EVAL_3,
  input         RationalCrossingSink_1__EVAL_4,
  input  [31:0] RationalCrossingSink_1__EVAL_9,
  input  [3:0]  RationalCrossingSink__EVAL_27,
  input  [1:0]  RationalCrossingSink_1__EVAL_2,
  input         RationalCrossingSink__EVAL_9,
  input  [2:0]  RationalCrossingSink__EVAL_8,
  input         RationalCrossingSink__EVAL_28,
  input  [3:0]  RationalCrossingSink__EVAL_17,
  input         RationalCrossingSource__EVAL_12,
  input         RationalCrossingSink__EVAL_19
);
  wire [2:0] TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire [3:0] TLMonitor__EVAL_5;
  wire [31:0] TLMonitor__EVAL_6;
  wire [7:0] TLMonitor__EVAL_7;
  wire [1:0] TLMonitor__EVAL_8;
  wire [2:0] TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire [31:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [2:0] TLMonitor__EVAL_14;
  wire [31:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire  TLMonitor__EVAL_17;
  wire  TLMonitor__EVAL_18;
  wire [3:0] TLMonitor__EVAL_19;
  wire  TLMonitor__EVAL_20;
  wire [3:0] TLMonitor__EVAL_21;
  wire  TLMonitor__EVAL_22;
  wire [1:0] TLMonitor__EVAL_23;
  wire  TLMonitor__EVAL_24;
  wire [2:0] TLMonitor__EVAL_25;
  wire  TLMonitor__EVAL_26;
  wire [3:0] TLMonitor__EVAL_27;
  wire  TLMonitor__EVAL_28;
  wire  TLMonitor__EVAL_29;
  wire  TLMonitor__EVAL_30;
  wire [3:0] TLMonitor__EVAL_31;
  wire [3:0] TLMonitor__EVAL_32;
  wire  TLMonitor__EVAL_33;
  SiFive__EVAL_267_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18),
    ._EVAL_19(TLMonitor__EVAL_19),
    ._EVAL_20(TLMonitor__EVAL_20),
    ._EVAL_21(TLMonitor__EVAL_21),
    ._EVAL_22(TLMonitor__EVAL_22),
    ._EVAL_23(TLMonitor__EVAL_23),
    ._EVAL_24(TLMonitor__EVAL_24),
    ._EVAL_25(TLMonitor__EVAL_25),
    ._EVAL_26(TLMonitor__EVAL_26),
    ._EVAL_27(TLMonitor__EVAL_27),
    ._EVAL_28(TLMonitor__EVAL_28),
    ._EVAL_29(TLMonitor__EVAL_29),
    ._EVAL_30(TLMonitor__EVAL_30),
    ._EVAL_31(TLMonitor__EVAL_31),
    ._EVAL_32(TLMonitor__EVAL_32),
    ._EVAL_33(TLMonitor__EVAL_33)
  );
  assign TLMonitor__EVAL_12 = _EVAL_71;
  assign TLMonitor__EVAL_10 = RationalCrossingSource_2__EVAL_3;
  assign TLMonitor__EVAL_27 = _EVAL_22;
  assign TLMonitor__EVAL_3 = RationalCrossingSource_1__EVAL_1;
  assign TLMonitor__EVAL_8 = RationalCrossingSink__EVAL_21;
  assign TLMonitor__EVAL_9 = _EVAL_74;
  assign TLMonitor__EVAL_6 = _EVAL_62;
  assign TLMonitor__EVAL_2 = _EVAL_67;
  assign TLMonitor__EVAL_26 = _EVAL_104;
  assign TLMonitor__EVAL_7 = _EVAL_100;
  assign TLMonitor__EVAL_11 = _EVAL_82;
  assign TLMonitor__EVAL_30 = _EVAL_3;
  assign TLMonitor__EVAL_1 = RationalCrossingSink__EVAL_3;
  assign TLMonitor__EVAL_17 = _EVAL_4;
  assign TLMonitor__EVAL = _EVAL_56;
  assign TLMonitor__EVAL_18 = _EVAL_23;
  assign TLMonitor__EVAL_4 = RationalCrossingSink_1__EVAL_4;
  assign TLMonitor__EVAL_24 = _EVAL_17;
  assign TLMonitor__EVAL_15 = RationalCrossingSink_1__EVAL_9;
  assign TLMonitor__EVAL_19 = RationalCrossingSink__EVAL_27;
  assign TLMonitor__EVAL_21 = _EVAL_106;
  assign TLMonitor__EVAL_23 = RationalCrossingSink_1__EVAL_2;
  assign TLMonitor__EVAL_25 = _EVAL_69;
  assign TLMonitor__EVAL_31 = _EVAL_26;
  assign TLMonitor__EVAL_5 = _EVAL_12;
  assign TLMonitor__EVAL_13 = RationalCrossingSink__EVAL_9;
  assign TLMonitor__EVAL_20 = _EVAL_96;
  assign TLMonitor__EVAL_0 = _EVAL_7;
  assign TLMonitor__EVAL_14 = RationalCrossingSink__EVAL_8;
  assign TLMonitor__EVAL_22 = RationalCrossingSink__EVAL_28;
  assign TLMonitor__EVAL_32 = RationalCrossingSink__EVAL_17;
  assign TLMonitor__EVAL_16 = RationalCrossingSource__EVAL_12;
  assign TLMonitor__EVAL_29 = RationalCrossingSink__EVAL_19;
  assign TLMonitor__EVAL_28 = _EVAL_42;
  assign TLMonitor__EVAL_33 = _EVAL_29;

endmodule
