//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_211_assert(
  input        _EVAL,
  input  [2:0] _EVAL_0,
  input        _EVAL_1,
  input  [2:0] _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input        _EVAL_5,
  input        _EVAL_6,
  input  [2:0] _EVAL_7,
  input        _EVAL_8,
  input  [3:0] _EVAL_9,
  input  [1:0] _EVAL_10,
  input  [8:0] _EVAL_11,
  input  [1:0] _EVAL_12,
  input        _EVAL_13,
  input        _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [1:0] _EVAL_37;
  reg [31:0] _RAND_0;
  reg [1:0] _EVAL_50;
  reg [31:0] _RAND_1;
  reg  _EVAL_117;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_123;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_127;
  reg [31:0] _RAND_4;
  reg  _EVAL_134;
  reg [31:0] _RAND_5;
  reg  _EVAL_135;
  reg [31:0] _RAND_6;
  reg  _EVAL_157;
  reg [31:0] _RAND_7;
  reg  _EVAL_174;
  reg [31:0] _RAND_8;
  reg [8:0] _EVAL_184;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_203;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_212;
  reg [31:0] _RAND_11;
  reg  _EVAL_221;
  reg [31:0] _RAND_12;
  reg  _EVAL_233;
  reg [31:0] _RAND_13;
  wire  _EVAL_63;
  wire [8:0] _EVAL_54;
  wire  _EVAL_109;
  wire [8:0] _EVAL_176;
  wire [9:0] _EVAL_26;
  wire [9:0] _EVAL_172;
  wire [9:0] _EVAL_144;
  wire  _EVAL_17;
  wire  _EVAL_160;
  wire  _EVAL_68;
  wire  _EVAL_121;
  wire [9:0] _EVAL_83;
  wire [9:0] _EVAL_153;
  wire [9:0] _EVAL_146;
  wire  _EVAL_138;
  wire  _EVAL_226;
  wire  _EVAL_31;
  wire  _EVAL_209;
  wire  _EVAL_53;
  wire [1:0] _EVAL_178;
  wire [1:0] _EVAL_238;
  wire  _EVAL_230;
  wire  _EVAL_98;
  wire  _EVAL_139;
  wire  _EVAL_122;
  wire  _EVAL_245;
  wire  _EVAL_234;
  wire [31:0] _EVAL_220;
  wire [4:0] _EVAL_130;
  wire [1:0] _EVAL_177;
  wire  _EVAL_106;
  wire  _EVAL_110;
  wire [8:0] _EVAL_70;
  wire [9:0] _EVAL_142;
  wire [9:0] _EVAL_152;
  wire [9:0] _EVAL_161;
  wire  _EVAL_81;
  wire  _EVAL_188;
  wire [8:0] _EVAL_143;
  wire [9:0] _EVAL_87;
  wire [9:0] _EVAL_90;
  wire [9:0] _EVAL_133;
  wire  _EVAL_148;
  wire  _EVAL_242;
  wire  _EVAL_249;
  wire [9:0] _EVAL_171;
  wire [9:0] _EVAL_61;
  wire [9:0] _EVAL_246;
  wire  _EVAL_187;
  wire  _EVAL_251;
  wire [8:0] _EVAL_119;
  wire [9:0] _EVAL_118;
  wire [9:0] _EVAL_40;
  wire [9:0] _EVAL_215;
  wire  _EVAL_207;
  wire  _EVAL_96;
  wire  _EVAL_225;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_257;
  wire  _EVAL_29;
  wire  _EVAL_155;
  wire [1:0] _EVAL_84;
  wire [1:0] _EVAL_197;
  wire  _EVAL_49;
  wire  _EVAL_79;
  wire  _EVAL_125;
  wire  _EVAL_217;
  wire  _EVAL_101;
  wire  _EVAL_73;
  wire  _EVAL_204;
  wire  _EVAL_193;
  wire  _EVAL_115;
  wire  _EVAL_169;
  wire  _EVAL_64;
  wire  _EVAL_56;
  wire  _EVAL_45;
  wire  _EVAL_182;
  wire  _EVAL_74;
  wire  _EVAL_38;
  wire  _EVAL_202;
  wire  _EVAL_94;
  wire  _EVAL_131;
  wire  _EVAL_16;
  wire  _EVAL_241;
  wire  _EVAL_191;
  wire  _EVAL_65;
  wire  _EVAL_82;
  wire  _EVAL_206;
  wire  _EVAL_108;
  wire  _EVAL_99;
  wire  _EVAL_243;
  wire  _EVAL_231;
  wire  _EVAL_165;
  wire  _EVAL_114;
  wire  _EVAL_210;
  wire [1:0] _EVAL_77;
  wire [1:0] _EVAL_48;
  wire  _EVAL_158;
  wire  _EVAL_71;
  wire  _EVAL_104;
  wire  _EVAL_58;
  wire  _EVAL_67;
  wire [3:0] _EVAL_126;
  wire  _EVAL_173;
  wire  _EVAL_44;
  wire  _EVAL_72;
  wire  _EVAL_192;
  wire  _EVAL_156;
  wire  _EVAL_69;
  wire  _EVAL_147;
  wire  _EVAL_78;
  wire  _EVAL_132;
  wire  _EVAL_227;
  wire  _EVAL_137;
  wire  _EVAL_247;
  wire  _EVAL_52;
  wire  _EVAL_189;
  wire  _EVAL_180;
  wire  _EVAL_240;
  wire  _EVAL_30;
  wire [3:0] _EVAL_229;
  wire [3:0] _EVAL_116;
  wire [3:0] _EVAL_103;
  wire  _EVAL_35;
  wire  _EVAL_256;
  wire  _EVAL_23;
  wire  _EVAL_55;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_97;
  wire  _EVAL_162;
  wire  _EVAL_124;
  wire  _EVAL_51;
  wire  _EVAL_25;
  wire  _EVAL_32;
  wire  _EVAL_255;
  wire  _EVAL_15;
  wire  _EVAL_92;
  wire  _EVAL_236;
  wire  _EVAL_105;
  wire  _EVAL_34;
  wire  _EVAL_232;
  wire  _EVAL_21;
  wire  _EVAL_183;
  wire  _EVAL_89;
  wire  _EVAL_167;
  wire  _EVAL_166;
  wire  _EVAL_258;
  wire  _EVAL_95;
  wire  _EVAL_46;
  wire  _EVAL_223;
  wire  _EVAL_113;
  wire  _EVAL_244;
  wire  _EVAL_235;
  wire  _EVAL_100;
  wire  _EVAL_239;
  wire  _EVAL_211;
  wire [1:0] _EVAL_200;
  wire  _EVAL_175;
  wire  _EVAL_91;
  wire  _EVAL_250;
  wire  _EVAL_219;
  wire  _EVAL_195;
  wire  _EVAL_28;
  wire  _EVAL_185;
  wire  _EVAL_218;
  wire  _EVAL_66;
  wire  _EVAL_102;
  wire  _EVAL_60;
  wire  _EVAL_93;
  wire  _EVAL_140;
  wire  _EVAL_112;
  wire  _EVAL_141;
  wire  _EVAL_248;
  wire  _EVAL_88;
  wire  _EVAL_205;
  wire  _EVAL_76;
  wire [8:0] _EVAL_136;
  wire [8:0] _EVAL_208;
  wire  _EVAL_80;
  wire  _EVAL_47;
  wire  _EVAL_42;
  wire  _EVAL_24;
  wire  _EVAL_43;
  wire  _EVAL_159;
  wire  _EVAL_168;
  wire  _EVAL_201;
  wire  _EVAL_170;
  wire  _EVAL_75;
  wire  _EVAL_196;
  wire  _EVAL_149;
  wire  _EVAL_20;
  wire  _EVAL_128;
  wire  _EVAL_254;
  wire  _EVAL_120;
  wire  _EVAL_19;
  wire  _EVAL_190;
  wire  _EVAL_163;
  wire  _EVAL_33;
  wire  _EVAL_107;
  wire  _EVAL_111;
  wire  _EVAL_27;
  wire  _EVAL_39;
  wire  _EVAL_199;
  wire  _EVAL_154;
  wire  _EVAL_186;
  wire  _EVAL_224;
  wire  _EVAL_228;
  wire  _EVAL_18;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_36;
  wire  _EVAL_85;
  wire  _EVAL_194;
  wire  _EVAL_198;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_63 = _EVAL_2 == 3'h0;
  assign _EVAL_54 = _EVAL_11 ^ 9'h80;
  assign _EVAL_109 = _EVAL_123 < plusarg_reader_out;
  assign _EVAL_176 = _EVAL_11 ^ 9'h60;
  assign _EVAL_26 = {1'b0,$signed(_EVAL_176)};
  assign _EVAL_172 = $signed(_EVAL_26) & $signed(-10'sh20);
  assign _EVAL_144 = $signed(_EVAL_172);
  assign _EVAL_17 = $signed(_EVAL_144) == $signed(10'sh0);
  assign _EVAL_160 = _EVAL_7 == 3'h0;
  assign _EVAL_68 = _EVAL_160 | _EVAL_14;
  assign _EVAL_121 = _EVAL_68 == 1'h0;
  assign _EVAL_83 = {1'b0,$signed(_EVAL_11)};
  assign _EVAL_153 = $signed(_EVAL_83) & $signed(-10'sh40);
  assign _EVAL_146 = $signed(_EVAL_153);
  assign _EVAL_138 = _EVAL_134 == 1'h0;
  assign _EVAL_226 = _EVAL_138 == 1'h0;
  assign _EVAL_31 = _EVAL_4 & _EVAL_8;
  assign _EVAL_209 = _EVAL_135 == 1'h0;
  assign _EVAL_53 = _EVAL_31 & _EVAL_209;
  assign _EVAL_178 = 2'h1 << _EVAL_6;
  assign _EVAL_238 = _EVAL_53 ? _EVAL_178 : 2'h0;
  assign _EVAL_230 = _EVAL_238[0];
  assign _EVAL_98 = _EVAL_230 | _EVAL_117;
  assign _EVAL_139 = _EVAL_98 >> _EVAL_3;
  assign _EVAL_122 = _EVAL_139 | _EVAL_14;
  assign _EVAL_245 = _EVAL_13 & _EVAL_1;
  assign _EVAL_234 = _EVAL_31 | _EVAL_245;
  assign _EVAL_220 = _EVAL_123 + 32'h1;
  assign _EVAL_130 = 5'h3 << _EVAL_10;
  assign _EVAL_177 = _EVAL_130[1:0];
  assign _EVAL_106 = _EVAL_10 <= 2'h2;
  assign _EVAL_110 = $signed(_EVAL_146) == $signed(10'sh0);
  assign _EVAL_70 = _EVAL_11 ^ 9'h44;
  assign _EVAL_142 = {1'b0,$signed(_EVAL_70)};
  assign _EVAL_152 = $signed(_EVAL_142) & $signed(-10'sh4);
  assign _EVAL_161 = $signed(_EVAL_152);
  assign _EVAL_81 = $signed(_EVAL_161) == $signed(10'sh0);
  assign _EVAL_188 = _EVAL_110 | _EVAL_81;
  assign _EVAL_143 = _EVAL_11 ^ 9'h48;
  assign _EVAL_87 = {1'b0,$signed(_EVAL_143)};
  assign _EVAL_90 = $signed(_EVAL_87) & $signed(-10'sh18);
  assign _EVAL_133 = $signed(_EVAL_90);
  assign _EVAL_148 = $signed(_EVAL_133) == $signed(10'sh0);
  assign _EVAL_242 = _EVAL_188 | _EVAL_148;
  assign _EVAL_249 = _EVAL_242 | _EVAL_17;
  assign _EVAL_171 = {1'b0,$signed(_EVAL_54)};
  assign _EVAL_61 = $signed(_EVAL_171) & $signed(-10'sh80);
  assign _EVAL_246 = $signed(_EVAL_61);
  assign _EVAL_187 = $signed(_EVAL_246) == $signed(10'sh0);
  assign _EVAL_251 = _EVAL_249 | _EVAL_187;
  assign _EVAL_119 = _EVAL_11 ^ 9'h100;
  assign _EVAL_118 = {1'b0,$signed(_EVAL_119)};
  assign _EVAL_40 = $signed(_EVAL_118) & $signed(-10'sh100);
  assign _EVAL_215 = $signed(_EVAL_40);
  assign _EVAL_207 = $signed(_EVAL_215) == $signed(10'sh0);
  assign _EVAL_96 = _EVAL_251 | _EVAL_207;
  assign _EVAL_225 = _EVAL_106 & _EVAL_96;
  assign _EVAL_213 = _EVAL_157 == 1'h0;
  assign _EVAL_214 = _EVAL_213 == 1'h0;
  assign _EVAL_257 = _EVAL_1 & _EVAL_214;
  assign _EVAL_29 = _EVAL_10 >= 2'h2;
  assign _EVAL_155 = _EVAL_10[0];
  assign _EVAL_84 = 2'h1 << _EVAL_155;
  assign _EVAL_197 = _EVAL_84 | 2'h1;
  assign _EVAL_49 = _EVAL_197[1];
  assign _EVAL_79 = _EVAL_11[1];
  assign _EVAL_125 = _EVAL_49 & _EVAL_79;
  assign _EVAL_217 = _EVAL_29 | _EVAL_125;
  assign _EVAL_101 = _EVAL_197[0];
  assign _EVAL_73 = _EVAL_11[0];
  assign _EVAL_204 = _EVAL_79 & _EVAL_73;
  assign _EVAL_193 = _EVAL_101 & _EVAL_204;
  assign _EVAL_115 = _EVAL_217 | _EVAL_193;
  assign _EVAL_169 = _EVAL_79 == 1'h0;
  assign _EVAL_64 = _EVAL_49 & _EVAL_169;
  assign _EVAL_56 = _EVAL_29 | _EVAL_64;
  assign _EVAL_45 = _EVAL_12 == _EVAL_37;
  assign _EVAL_182 = _EVAL_45 | _EVAL_14;
  assign _EVAL_74 = _EVAL_2 == 3'h3;
  assign _EVAL_38 = _EVAL_8 & _EVAL_74;
  assign _EVAL_202 = _EVAL_134 - 1'h1;
  assign _EVAL_94 = _EVAL_117 == 1'h0;
  assign _EVAL_131 = plusarg_reader_out == 32'h0;
  assign _EVAL_16 = _EVAL_94 | _EVAL_131;
  assign _EVAL_241 = _EVAL_16 | _EVAL_109;
  assign _EVAL_191 = _EVAL_241 | _EVAL_14;
  assign _EVAL_65 = _EVAL_0 == 3'h6;
  assign _EVAL_82 = _EVAL_0 == 3'h2;
  assign _EVAL_206 = _EVAL_1 & _EVAL_82;
  assign _EVAL_108 = _EVAL_1 & _EVAL_65;
  assign _EVAL_99 = _EVAL_12 >= 2'h2;
  assign _EVAL_243 = _EVAL_117 | _EVAL_230;
  assign _EVAL_231 = _EVAL_233 == 1'h0;
  assign _EVAL_165 = _EVAL_245 & _EVAL_231;
  assign _EVAL_114 = _EVAL_65 == 1'h0;
  assign _EVAL_210 = _EVAL_165 & _EVAL_114;
  assign _EVAL_77 = 2'h1 << _EVAL_3;
  assign _EVAL_48 = _EVAL_210 ? _EVAL_77 : 2'h0;
  assign _EVAL_158 = _EVAL_48[0];
  assign _EVAL_71 = ~ _EVAL_158;
  assign _EVAL_104 = _EVAL_243 & _EVAL_71;
  assign _EVAL_58 = _EVAL_0 == 3'h5;
  assign _EVAL_67 = _EVAL_1 & _EVAL_58;
  assign _EVAL_126 = ~ _EVAL_9;
  assign _EVAL_173 = _EVAL_5 == 1'h0;
  assign _EVAL_44 = _EVAL_173 | _EVAL_14;
  assign _EVAL_72 = _EVAL_7 <= 3'h2;
  assign _EVAL_192 = _EVAL_2 == 3'h7;
  assign _EVAL_156 = _EVAL_8 & _EVAL_192;
  assign _EVAL_69 = _EVAL_0 == _EVAL_203;
  assign _EVAL_147 = _EVAL_69 | _EVAL_14;
  assign _EVAL_78 = _EVAL_73 == 1'h0;
  assign _EVAL_132 = _EVAL_79 & _EVAL_78;
  assign _EVAL_227 = _EVAL_101 & _EVAL_132;
  assign _EVAL_137 = _EVAL_217 | _EVAL_227;
  assign _EVAL_247 = _EVAL_169 & _EVAL_73;
  assign _EVAL_52 = _EVAL_101 & _EVAL_247;
  assign _EVAL_189 = _EVAL_56 | _EVAL_52;
  assign _EVAL_180 = _EVAL_169 & _EVAL_78;
  assign _EVAL_240 = _EVAL_101 & _EVAL_180;
  assign _EVAL_30 = _EVAL_56 | _EVAL_240;
  assign _EVAL_229 = {_EVAL_115,_EVAL_137,_EVAL_189,_EVAL_30};
  assign _EVAL_116 = ~ _EVAL_229;
  assign _EVAL_103 = _EVAL_9 & _EVAL_116;
  assign _EVAL_35 = _EVAL_103 == 4'h0;
  assign _EVAL_256 = _EVAL_35 | _EVAL_14;
  assign _EVAL_23 = _EVAL_256 == 1'h0;
  assign _EVAL_55 = _EVAL_0 <= 3'h6;
  assign _EVAL_179 = _EVAL_55 | _EVAL_14;
  assign _EVAL_181 = _EVAL_0 == 3'h1;
  assign _EVAL_97 = _EVAL_1 & _EVAL_181;
  assign _EVAL_162 = _EVAL_117 >> _EVAL_6;
  assign _EVAL_124 = _EVAL_162 == 1'h0;
  assign _EVAL_51 = _EVAL_124 | _EVAL_14;
  assign _EVAL_25 = _EVAL_0 == 3'h0;
  assign _EVAL_32 = _EVAL_1 & _EVAL_25;
  assign _EVAL_255 = _EVAL_6 == 1'h0;
  assign _EVAL_15 = _EVAL_255 | _EVAL_14;
  assign _EVAL_92 = _EVAL_15 == 1'h0;
  assign _EVAL_236 = _EVAL_233 - 1'h1;
  assign _EVAL_105 = _EVAL_29 | _EVAL_14;
  assign _EVAL_34 = _EVAL_2 == _EVAL_212;
  assign _EVAL_232 = _EVAL_3 == _EVAL_221;
  assign _EVAL_21 = _EVAL_232 | _EVAL_14;
  assign _EVAL_183 = _EVAL_21 == 1'h0;
  assign _EVAL_89 = _EVAL_10 == _EVAL_50;
  assign _EVAL_167 = _EVAL_225 | _EVAL_14;
  assign _EVAL_166 = _EVAL_167 == 1'h0;
  assign _EVAL_258 = _EVAL_2 == 3'h2;
  assign _EVAL_95 = _EVAL_34 | _EVAL_14;
  assign _EVAL_46 = _EVAL_6 == _EVAL_174;
  assign _EVAL_223 = _EVAL_46 | _EVAL_14;
  assign _EVAL_113 = _EVAL_3 == 1'h0;
  assign _EVAL_244 = _EVAL_7 <= 3'h3;
  assign _EVAL_235 = _EVAL_7 != 3'h0;
  assign _EVAL_100 = _EVAL_235 | _EVAL_14;
  assign _EVAL_239 = _EVAL_135 - 1'h1;
  assign _EVAL_211 = _EVAL_89 | _EVAL_14;
  assign _EVAL_200 = ~ _EVAL_177;
  assign _EVAL_175 = _EVAL_105 == 1'h0;
  assign _EVAL_91 = _EVAL_8 & _EVAL_226;
  assign _EVAL_250 = _EVAL_2 == 3'h4;
  assign _EVAL_219 = _EVAL_8 & _EVAL_250;
  assign _EVAL_195 = _EVAL_44 == 1'h0;
  assign _EVAL_28 = _EVAL_244 | _EVAL_14;
  assign _EVAL_185 = _EVAL_2 == 3'h6;
  assign _EVAL_218 = _EVAL_147 == 1'h0;
  assign _EVAL_66 = _EVAL_11 == _EVAL_184;
  assign _EVAL_102 = _EVAL_66 | _EVAL_14;
  assign _EVAL_60 = _EVAL_102 == 1'h0;
  assign _EVAL_93 = _EVAL_51 == 1'h0;
  assign _EVAL_140 = _EVAL_157 - 1'h1;
  assign _EVAL_112 = _EVAL_7 == _EVAL_127;
  assign _EVAL_141 = _EVAL_112 | _EVAL_14;
  assign _EVAL_248 = _EVAL_245 & _EVAL_213;
  assign _EVAL_88 = _EVAL_28 == 1'h0;
  assign _EVAL_205 = _EVAL_126 == 4'h0;
  assign _EVAL_76 = _EVAL_205 | _EVAL_14;
  assign _EVAL_136 = {{7'd0}, _EVAL_200};
  assign _EVAL_208 = _EVAL_11 & _EVAL_136;
  assign _EVAL_80 = _EVAL_122 == 1'h0;
  assign _EVAL_47 = _EVAL_211 == 1'h0;
  assign _EVAL_42 = _EVAL_113 | _EVAL_14;
  assign _EVAL_24 = _EVAL_99 | _EVAL_14;
  assign _EVAL_43 = _EVAL_191 == 1'h0;
  assign _EVAL_159 = _EVAL_95 == 1'h0;
  assign _EVAL_168 = _EVAL_100 == 1'h0;
  assign _EVAL_201 = _EVAL_7 <= 3'h4;
  assign _EVAL_170 = _EVAL_201 | _EVAL_14;
  assign _EVAL_75 = _EVAL_170 == 1'h0;
  assign _EVAL_196 = _EVAL_208 == 9'h0;
  assign _EVAL_149 = _EVAL_0 == 3'h4;
  assign _EVAL_20 = _EVAL_182 == 1'h0;
  assign _EVAL_128 = _EVAL_223 == 1'h0;
  assign _EVAL_254 = _EVAL_8 & _EVAL_258;
  assign _EVAL_120 = _EVAL_2 == 3'h5;
  assign _EVAL_19 = _EVAL_76 == 1'h0;
  assign _EVAL_190 = _EVAL_179 == 1'h0;
  assign _EVAL_163 = _EVAL_9 == _EVAL_229;
  assign _EVAL_33 = _EVAL_163 | _EVAL_14;
  assign _EVAL_107 = _EVAL_196 | _EVAL_14;
  assign _EVAL_111 = _EVAL_2 == 3'h1;
  assign _EVAL_27 = _EVAL_8 & _EVAL_111;
  assign _EVAL_39 = _EVAL_33 == 1'h0;
  assign _EVAL_199 = _EVAL_31 & _EVAL_138;
  assign _EVAL_154 = _EVAL_8 & _EVAL_63;
  assign _EVAL_186 = _EVAL_14 == 1'h0;
  assign _EVAL_224 = _EVAL_8 & _EVAL_120;
  assign _EVAL_228 = _EVAL_141 == 1'h0;
  assign _EVAL_18 = _EVAL_107 == 1'h0;
  assign _EVAL_150 = _EVAL_72 | _EVAL_14;
  assign _EVAL_151 = _EVAL_150 == 1'h0;
  assign _EVAL_36 = _EVAL_42 == 1'h0;
  assign _EVAL_85 = _EVAL_24 == 1'h0;
  assign _EVAL_194 = _EVAL_1 & _EVAL_149;
  assign _EVAL_198 = _EVAL_8 & _EVAL_185;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_37 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_50 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_117 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_123 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_127 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_134 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_135 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_157 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_174 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_184 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_203 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_212 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_221 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_233 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_248) begin
      _EVAL_37 <= _EVAL_12;
    end
    if (_EVAL_199) begin
      _EVAL_50 <= _EVAL_10;
    end
    if (_EVAL_14) begin
      _EVAL_117 <= 1'h0;
    end else begin
      _EVAL_117 <= _EVAL_104;
    end
    if (_EVAL_14) begin
      _EVAL_123 <= 32'h0;
    end else begin
      if (_EVAL_234) begin
        _EVAL_123 <= 32'h0;
      end else begin
        _EVAL_123 <= _EVAL_220;
      end
    end
    if (_EVAL_199) begin
      _EVAL_127 <= _EVAL_7;
    end
    if (_EVAL_14) begin
      _EVAL_134 <= 1'h0;
    end else begin
      if (_EVAL_31) begin
        if (_EVAL_138) begin
          _EVAL_134 <= 1'h0;
        end else begin
          _EVAL_134 <= _EVAL_202;
        end
      end
    end
    if (_EVAL_14) begin
      _EVAL_135 <= 1'h0;
    end else begin
      if (_EVAL_31) begin
        if (_EVAL_209) begin
          _EVAL_135 <= 1'h0;
        end else begin
          _EVAL_135 <= _EVAL_239;
        end
      end
    end
    if (_EVAL_14) begin
      _EVAL_157 <= 1'h0;
    end else begin
      if (_EVAL_245) begin
        if (_EVAL_213) begin
          _EVAL_157 <= 1'h0;
        end else begin
          _EVAL_157 <= _EVAL_140;
        end
      end
    end
    if (_EVAL_199) begin
      _EVAL_174 <= _EVAL_6;
    end
    if (_EVAL_199) begin
      _EVAL_184 <= _EVAL_11;
    end
    if (_EVAL_248) begin
      _EVAL_203 <= _EVAL_0;
    end
    if (_EVAL_199) begin
      _EVAL_212 <= _EVAL_2;
    end
    if (_EVAL_248) begin
      _EVAL_221 <= _EVAL_3;
    end
    if (_EVAL_14) begin
      _EVAL_233 <= 1'h0;
    end else begin
      if (_EVAL_245) begin
        if (_EVAL_231) begin
          _EVAL_233 <= 1'h0;
        end else begin
          _EVAL_233 <= _EVAL_236;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4f16e65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae8c647e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36aa1be4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ee2a07a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3477010)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8d32161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15e22ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f4037d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de8d6f77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c869348d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f412d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(581041ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(877132e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d42578fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34e08e9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5779b20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69021240)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f2e9ac9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8f782f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78102890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6475e9e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f3a0681)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd968690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d56dc4e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca6aa006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(575c089a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(946962ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38d67063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b98f097)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdda7bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3b99d71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3baa884b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bab7de1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de7ab9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7b77070)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50805480)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6d5d363)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(975d19e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6971d8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc52e753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56397583)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(886b9ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4550a444)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a439e59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c617f25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d11a4eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4de1ac38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18ee873c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d165f1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5541da04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88e8d444)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9167698e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aff83f68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d62c03a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8864732a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acfcfaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59a12a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efef4626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8d1c87e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(262adfd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dc099fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ad270d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9b20fd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c9908f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f6a822)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76a6b2fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ea6844b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da413053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13a9e7d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67eee3c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cdfabc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
