//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_133(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [11:0] _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output [11:0] _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  output        _EVAL_9,
  output [2:0]  _EVAL_10,
  output [27:0] _EVAL_11,
  output [2:0]  _EVAL_12,
  input         _EVAL_13,
  output [3:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  output [2:0]  _EVAL_18,
  output [6:0]  _EVAL_19,
  output [2:0]  _EVAL_20,
  output [31:0] _EVAL_21,
  input         _EVAL_22,
  input  [27:0] _EVAL_23,
  input  [3:0]  _EVAL_24,
  output        _EVAL_25,
  input  [2:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  input  [31:0] _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  input  [6:0]  _EVAL_31,
  output [1:0]  _EVAL_32
);
  wire [11:0] fragmenter__EVAL;
  wire [31:0] fragmenter__EVAL_0;
  wire  fragmenter__EVAL_1;
  wire [2:0] fragmenter__EVAL_2;
  wire [1:0] fragmenter__EVAL_3;
  wire  fragmenter__EVAL_4;
  wire  fragmenter__EVAL_5;
  wire [1:0] fragmenter__EVAL_6;
  wire [2:0] fragmenter__EVAL_7;
  wire [2:0] fragmenter__EVAL_8;
  wire  fragmenter__EVAL_9;
  wire [27:0] fragmenter__EVAL_10;
  wire [2:0] fragmenter__EVAL_11;
  wire [2:0] fragmenter__EVAL_12;
  wire [3:0] fragmenter__EVAL_13;
  wire [3:0] fragmenter__EVAL_14;
  wire [2:0] fragmenter__EVAL_15;
  wire [2:0] fragmenter__EVAL_16;
  wire  fragmenter__EVAL_17;
  wire [27:0] fragmenter__EVAL_18;
  wire [11:0] fragmenter__EVAL_19;
  wire  fragmenter__EVAL_20;
  wire [6:0] fragmenter__EVAL_21;
  wire [2:0] fragmenter__EVAL_22;
  wire [31:0] fragmenter__EVAL_23;
  wire  fragmenter__EVAL_24;
  wire [6:0] fragmenter__EVAL_25;
  wire  fragmenter__EVAL_26;
  wire  fragmenter__EVAL_27;
  wire [31:0] fragmenter__EVAL_28;
  wire  fragmenter__EVAL_29;
  wire [31:0] fragmenter__EVAL_30;
  wire  fragmenter__EVAL_31;
  wire  fragmenter__EVAL_32;
  SiFive__EVAL_132 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28),
    ._EVAL_29(fragmenter__EVAL_29),
    ._EVAL_30(fragmenter__EVAL_30),
    ._EVAL_31(fragmenter__EVAL_31),
    ._EVAL_32(fragmenter__EVAL_32)
  );
  assign fragmenter__EVAL_19 = _EVAL_3;
  assign fragmenter__EVAL_20 = _EVAL_22;
  assign _EVAL_32 = fragmenter__EVAL_3;
  assign _EVAL_27 = fragmenter__EVAL_23;
  assign fragmenter__EVAL_5 = _EVAL_13;
  assign _EVAL_25 = fragmenter__EVAL_17;
  assign fragmenter__EVAL_1 = _EVAL_1;
  assign _EVAL_21 = fragmenter__EVAL_0;
  assign _EVAL_12 = fragmenter__EVAL_22;
  assign _EVAL_10 = fragmenter__EVAL_16;
  assign fragmenter__EVAL_6 = _EVAL_8;
  assign fragmenter__EVAL_26 = _EVAL_0;
  assign fragmenter__EVAL_24 = _EVAL_4;
  assign _EVAL_29 = fragmenter__EVAL_4;
  assign fragmenter__EVAL_2 = _EVAL_15;
  assign fragmenter__EVAL_30 = _EVAL_28;
  assign _EVAL_17 = fragmenter__EVAL_31;
  assign _EVAL_6 = fragmenter__EVAL;
  assign _EVAL_14 = fragmenter__EVAL_14;
  assign fragmenter__EVAL_12 = _EVAL_7;
  assign fragmenter__EVAL_29 = _EVAL_16;
  assign fragmenter__EVAL_7 = _EVAL;
  assign _EVAL_30 = fragmenter__EVAL_9;
  assign fragmenter__EVAL_15 = _EVAL_26;
  assign fragmenter__EVAL_28 = _EVAL_2;
  assign _EVAL_9 = fragmenter__EVAL_27;
  assign fragmenter__EVAL_32 = _EVAL_5;
  assign fragmenter__EVAL_21 = _EVAL_31;
  assign _EVAL_11 = fragmenter__EVAL_18;
  assign fragmenter__EVAL_13 = _EVAL_24;
  assign _EVAL_20 = fragmenter__EVAL_8;
  assign fragmenter__EVAL_10 = _EVAL_23;
  assign _EVAL_18 = fragmenter__EVAL_11;
  assign _EVAL_19 = fragmenter__EVAL_25;
endmodule
