//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_66(
  input  [1:0]  _EVAL,
  output [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  output [2:0]  _EVAL_6,
  output [31:0] _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  output [31:0] _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [4:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input  [3:0]  _EVAL_21,
  output [4:0]  _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output [31:0] _EVAL_25,
  input         _EVAL_26,
  output        _EVAL_27,
  input  [3:0]  _EVAL_28,
  input  [31:0] _EVAL_29,
  output [4:0]  _EVAL_30,
  output [2:0]  _EVAL_31,
  output [2:0]  _EVAL_32,
  input         _EVAL_33,
  input  [31:0] _EVAL_34,
  input  [2:0]  _EVAL_35,
  input         _EVAL_36,
  output [3:0]  _EVAL_37,
  input  [4:0]  _EVAL_38
);
  assign _EVAL_16 = _EVAL_13;
  assign _EVAL_27 = _EVAL_10;
  assign _EVAL_19 = _EVAL_36;
  assign _EVAL_30 = _EVAL_38;
  assign _EVAL_18 = _EVAL_20;
  assign _EVAL_24 = _EVAL_26;
  assign _EVAL_3 = _EVAL_1;
  assign _EVAL_31 = _EVAL_15;
  assign _EVAL_6 = _EVAL_17;
  assign _EVAL_7 = _EVAL_8;
  assign _EVAL_22 = _EVAL_14;
  assign _EVAL_0 = _EVAL_28;
  assign _EVAL_5 = _EVAL_11;
  assign _EVAL_25 = _EVAL_34;
  assign _EVAL_23 = _EVAL_33;
  assign _EVAL_37 = _EVAL_21;
  assign _EVAL_32 = _EVAL_35;
  assign _EVAL_12 = _EVAL_29;
endmodule
