//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_325_assert(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [6:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [29:0] _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input  [6:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [7:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input  [2:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_21;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_45;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_83;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_97;
  reg [31:0] _RAND_3;
  reg [29:0] _EVAL_107;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_110;
  reg [31:0] _RAND_5;
  reg  _EVAL_151;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_176;
  reg [31:0] _RAND_7;
  reg [4:0] _EVAL_182;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_197;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_200;
  reg [31:0] _RAND_10;
  reg [72:0] _EVAL_223;
  reg [95:0] _RAND_11;
  reg [3:0] _EVAL_229;
  reg [31:0] _RAND_12;
  reg [6:0] _EVAL_292;
  reg [31:0] _RAND_13;
  reg  _EVAL_304;
  reg [31:0] _RAND_14;
  reg [1:0] _EVAL_340;
  reg [31:0] _RAND_15;
  reg [6:0] _EVAL_379;
  reg [31:0] _RAND_16;
  wire [3:0] _EVAL_224;
  wire  _EVAL_367;
  wire  _EVAL_361;
  wire  _EVAL_104;
  wire  _EVAL_342;
  wire  _EVAL_164;
  wire  _EVAL_333;
  wire [127:0] _EVAL_288;
  wire [127:0] _EVAL_234;
  wire [72:0] _EVAL_296;
  wire  _EVAL_370;
  wire  _EVAL_186;
  wire  _EVAL_237;
  wire  _EVAL_269;
  wire  _EVAL_308;
  wire [1:0] _EVAL_341;
  wire [3:0] _EVAL_317;
  wire [2:0] _EVAL_191;
  wire [2:0] _EVAL_158;
  wire  _EVAL_69;
  wire  _EVAL_218;
  wire  _EVAL_20;
  wire  _EVAL_313;
  wire  _EVAL_206;
  wire  _EVAL_26;
  wire  _EVAL_345;
  wire  _EVAL_295;
  wire  _EVAL_330;
  wire  _EVAL_306;
  wire  _EVAL_183;
  wire  _EVAL_321;
  wire  _EVAL_324;
  wire  _EVAL_173;
  wire  _EVAL_322;
  wire  _EVAL_172;
  wire  _EVAL_202;
  wire  _EVAL_184;
  wire  _EVAL_55;
  wire  _EVAL_246;
  wire  _EVAL_272;
  wire  _EVAL_96;
  wire  _EVAL_247;
  wire  _EVAL_133;
  wire  _EVAL_215;
  wire  _EVAL_90;
  wire  _EVAL_94;
  wire  _EVAL_35;
  wire  _EVAL_193;
  wire  _EVAL_323;
  wire  _EVAL_194;
  wire  _EVAL_353;
  wire  _EVAL_328;
  wire  _EVAL_301;
  wire  _EVAL_207;
  wire  _EVAL_39;
  wire  _EVAL_175;
  wire  _EVAL_219;
  wire  _EVAL_332;
  wire  _EVAL_111;
  wire  _EVAL_195;
  wire  _EVAL_369;
  wire  _EVAL_331;
  wire  _EVAL_67;
  wire  _EVAL_382;
  wire  _EVAL_144;
  wire  _EVAL_371;
  wire  _EVAL_249;
  wire  _EVAL_251;
  wire [7:0] _EVAL_320;
  wire  _EVAL_187;
  wire  _EVAL_362;
  wire  _EVAL_115;
  wire  _EVAL_227;
  wire  _EVAL_174;
  wire  _EVAL_145;
  wire  _EVAL_54;
  wire  _EVAL_244;
  wire [30:0] _EVAL_56;
  wire [30:0] _EVAL_278;
  wire [30:0] _EVAL_388;
  wire [72:0] _EVAL_266;
  wire  _EVAL_271;
  wire  _EVAL_360;
  wire  _EVAL_196;
  wire  _EVAL_72;
  wire  _EVAL_364;
  wire  _EVAL_78;
  wire  _EVAL_343;
  wire  _EVAL_126;
  wire  _EVAL_307;
  wire  _EVAL_138;
  wire  _EVAL_281;
  wire [29:0] _EVAL_316;
  wire [30:0] _EVAL_47;
  wire [30:0] _EVAL_89;
  wire [30:0] _EVAL_265;
  wire  _EVAL_276;
  wire [29:0] _EVAL_334;
  wire [30:0] _EVAL_282;
  wire [30:0] _EVAL_287;
  wire [30:0] _EVAL_49;
  wire  _EVAL_165;
  wire  _EVAL_178;
  wire [29:0] _EVAL_68;
  wire [30:0] _EVAL_291;
  wire [30:0] _EVAL_203;
  wire [30:0] _EVAL_142;
  wire  _EVAL_135;
  wire  _EVAL_357;
  wire  _EVAL_181;
  wire  _EVAL_318;
  wire  _EVAL_101;
  wire  _EVAL_392;
  wire  _EVAL_243;
  wire  _EVAL_254;
  wire  _EVAL_214;
  wire  _EVAL_88;
  wire  _EVAL_46;
  wire [127:0] _EVAL_192;
  wire [127:0] _EVAL_93;
  wire [72:0] _EVAL_24;
  wire  _EVAL_228;
  wire  _EVAL_31;
  wire  _EVAL_137;
  wire  _EVAL_60;
  wire  _EVAL_134;
  wire [29:0] _EVAL_87;
  wire [30:0] _EVAL_163;
  wire [30:0] _EVAL_239;
  wire [30:0] _EVAL_170;
  wire  _EVAL_118;
  wire [29:0] _EVAL_121;
  wire  _EVAL_255;
  wire  _EVAL_365;
  wire  _EVAL_216;
  wire [4:0] _EVAL_129;
  wire [7:0] _EVAL_381;
  wire  _EVAL_58;
  wire  _EVAL_319;
  wire [72:0] _EVAL_210;
  wire  _EVAL_190;
  wire  _EVAL_238;
  wire  _EVAL_347;
  wire  _EVAL_23;
  wire [22:0] _EVAL_275;
  wire [7:0] _EVAL_208;
  wire [7:0] _EVAL_245;
  wire [29:0] _EVAL_393;
  wire [29:0] _EVAL_153;
  wire  _EVAL_325;
  wire  _EVAL_314;
  wire  _EVAL_152;
  wire  _EVAL_368;
  wire  _EVAL_30;
  wire  _EVAL_285;
  wire  _EVAL_240;
  wire  _EVAL_236;
  wire  _EVAL_122;
  wire  _EVAL_298;
  wire  _EVAL_43;
  wire [22:0] _EVAL_50;
  wire [7:0] _EVAL_398;
  wire [7:0] _EVAL_310;
  wire  _EVAL_85;
  wire  _EVAL_312;
  wire  _EVAL_123;
  wire  _EVAL_394;
  wire  _EVAL_146;
  wire  _EVAL_171;
  wire  _EVAL_376;
  wire  _EVAL_286;
  wire  _EVAL_349;
  wire  _EVAL_179;
  wire  _EVAL_125;
  wire [2:0] _EVAL_81;
  wire  _EVAL_185;
  wire  _EVAL_222;
  wire  _EVAL_124;
  wire  _EVAL_262;
  wire  _EVAL_136;
  wire  _EVAL_366;
  wire  _EVAL_248;
  wire  _EVAL_252;
  wire  _EVAL_66;
  wire  _EVAL_150;
  wire  _EVAL_373;
  wire  _EVAL_225;
  wire  _EVAL_139;
  wire  _EVAL_102;
  wire  _EVAL_354;
  wire [3:0] _EVAL_387;
  wire  _EVAL_65;
  wire [2:0] _EVAL_267;
  wire  _EVAL_250;
  wire  _EVAL_231;
  wire  _EVAL_32;
  wire  _EVAL_108;
  wire  _EVAL_22;
  wire  _EVAL_338;
  wire  _EVAL_378;
  wire  _EVAL_395;
  wire  _EVAL_391;
  wire  _EVAL_209;
  wire  _EVAL_337;
  wire  _EVAL_63;
  wire [30:0] _EVAL_52;
  wire [30:0] _EVAL_257;
  wire [30:0] _EVAL_188;
  wire  _EVAL_315;
  wire  _EVAL_82;
  wire [29:0] _EVAL_44;
  wire [30:0] _EVAL_311;
  wire [30:0] _EVAL_106;
  wire [30:0] _EVAL_258;
  wire  _EVAL_36;
  wire  _EVAL_305;
  wire  _EVAL_213;
  wire  _EVAL_180;
  wire  _EVAL_168;
  wire  _EVAL_120;
  wire  _EVAL_149;
  wire  _EVAL_103;
  wire  _EVAL_162;
  wire  _EVAL_274;
  wire [4:0] _EVAL_399;
  wire [4:0] _EVAL_156;
  wire [4:0] _EVAL_348;
  wire  _EVAL_336;
  wire  _EVAL_160;
  wire  _EVAL_99;
  wire  _EVAL_157;
  wire  _EVAL_159;
  wire  _EVAL_212;
  wire  _EVAL_261;
  wire  _EVAL_41;
  wire  _EVAL_77;
  wire  _EVAL_350;
  wire  _EVAL_75;
  wire  _EVAL_84;
  wire  _EVAL_273;
  wire  _EVAL_300;
  wire  _EVAL_116;
  wire [7:0] _EVAL_242;
  wire [7:0] _EVAL_279;
  wire  _EVAL_53;
  wire  _EVAL_70;
  wire  _EVAL_268;
  wire  _EVAL_397;
  wire  _EVAL_25;
  wire  _EVAL_38;
  wire  _EVAL_199;
  wire  _EVAL_48;
  wire  _EVAL_344;
  wire  _EVAL_19;
  wire  _EVAL_309;
  wire  _EVAL_57;
  wire  _EVAL_389;
  wire  _EVAL_51;
  wire  _EVAL_375;
  wire  _EVAL_86;
  wire  _EVAL_339;
  wire  _EVAL_232;
  wire  _EVAL_299;
  wire  _EVAL_109;
  wire  _EVAL_64;
  wire  _EVAL_132;
  wire  _EVAL_28;
  wire  _EVAL_62;
  wire  _EVAL_117;
  wire [4:0] _EVAL_177;
  wire  _EVAL_130;
  wire  _EVAL_374;
  wire  _EVAL_112;
  wire  _EVAL_358;
  wire  _EVAL_167;
  wire  _EVAL_241;
  wire  _EVAL_127;
  wire [4:0] _EVAL_351;
  wire  _EVAL_264;
  wire  _EVAL_100;
  wire  _EVAL_147;
  wire  _EVAL_40;
  wire  _EVAL_198;
  wire  _EVAL_329;
  wire  _EVAL_293;
  wire  _EVAL_92;
  wire [72:0] _EVAL_235;
  wire  _EVAL_352;
  wire  _EVAL_105;
  wire  _EVAL_205;
  wire  _EVAL_383;
  wire  _EVAL_42;
  wire  _EVAL_226;
  wire  _EVAL_355;
  wire  _EVAL_384;
  wire  _EVAL_155;
  wire  _EVAL_98;
  wire  _EVAL_385;
  wire  _EVAL_27;
  wire [72:0] _EVAL_211;
  wire [72:0] _EVAL_302;
  wire [72:0] _EVAL_386;
  wire  _EVAL_377;
  wire  _EVAL_29;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_74;
  wire  _EVAL_263;
  wire  _EVAL_73;
  wire  _EVAL_189;
  wire  _EVAL_59;
  wire  _EVAL_148;
  wire  _EVAL_95;
  wire  _EVAL_113;
  wire  _EVAL_204;
  wire  _EVAL_201;
  wire  _EVAL_289;
  wire  _EVAL_335;
  wire  _EVAL_37;
  wire  _EVAL_359;
  wire  _EVAL_356;
  wire  _EVAL_61;
  wire  _EVAL_284;
  wire  _EVAL_230;
  wire  _EVAL_71;
  wire  _EVAL_346;
  wire [31:0] _EVAL_372;
  wire  _EVAL_233;
  wire  _EVAL_270;
  wire  _EVAL_143;
  wire  _EVAL_220;
  wire  _EVAL_119;
  wire  _EVAL_363;
  wire  _EVAL_290;
  wire  _EVAL_260;
  wire  _EVAL_76;
  wire  _EVAL_33;
  wire  _EVAL_80;
  wire  _EVAL_283;
  wire  _EVAL_326;
  wire  _EVAL_253;
  wire  _EVAL_169;
  wire  _EVAL_256;
  wire  _EVAL_259;
  wire  _EVAL_390;
  wire  _EVAL_221;
  wire  _EVAL_79;
  wire  _EVAL_217;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_224 = _EVAL_11[6:3];
  assign _EVAL_367 = _EVAL >= 4'h3;
  assign _EVAL_361 = _EVAL_367 | _EVAL_13;
  assign _EVAL_104 = _EVAL_361 == 1'h0;
  assign _EVAL_342 = _EVAL_10 & _EVAL_7;
  assign _EVAL_164 = _EVAL_110 == 5'h0;
  assign _EVAL_333 = _EVAL_342 & _EVAL_164;
  assign _EVAL_288 = 128'h1 << _EVAL_11;
  assign _EVAL_234 = _EVAL_333 ? _EVAL_288 : 128'h0;
  assign _EVAL_296 = _EVAL_234[72:0];
  assign _EVAL_370 = _EVAL_296 != 73'h0;
  assign _EVAL_186 = _EVAL_17 == _EVAL_340;
  assign _EVAL_237 = _EVAL_186 | _EVAL_13;
  assign _EVAL_269 = _EVAL_237 == 1'h0;
  assign _EVAL_308 = _EVAL_9 >= 4'h3;
  assign _EVAL_341 = _EVAL_9[1:0];
  assign _EVAL_317 = 4'h1 << _EVAL_341;
  assign _EVAL_191 = _EVAL_317[2:0];
  assign _EVAL_158 = _EVAL_191 | 3'h1;
  assign _EVAL_69 = _EVAL_158[2];
  assign _EVAL_218 = _EVAL_6[2];
  assign _EVAL_20 = _EVAL_69 & _EVAL_218;
  assign _EVAL_313 = _EVAL_308 | _EVAL_20;
  assign _EVAL_206 = _EVAL_158[1];
  assign _EVAL_26 = _EVAL_6[1];
  assign _EVAL_345 = _EVAL_218 & _EVAL_26;
  assign _EVAL_295 = _EVAL_206 & _EVAL_345;
  assign _EVAL_330 = _EVAL_313 | _EVAL_295;
  assign _EVAL_306 = _EVAL_158[0];
  assign _EVAL_183 = _EVAL_6[0];
  assign _EVAL_321 = _EVAL_345 & _EVAL_183;
  assign _EVAL_324 = _EVAL_306 & _EVAL_321;
  assign _EVAL_173 = _EVAL_330 | _EVAL_324;
  assign _EVAL_322 = _EVAL_183 == 1'h0;
  assign _EVAL_172 = _EVAL_345 & _EVAL_322;
  assign _EVAL_202 = _EVAL_306 & _EVAL_172;
  assign _EVAL_184 = _EVAL_330 | _EVAL_202;
  assign _EVAL_55 = _EVAL_26 == 1'h0;
  assign _EVAL_246 = _EVAL_218 & _EVAL_55;
  assign _EVAL_272 = _EVAL_206 & _EVAL_246;
  assign _EVAL_96 = _EVAL_313 | _EVAL_272;
  assign _EVAL_247 = _EVAL_246 & _EVAL_183;
  assign _EVAL_133 = _EVAL_306 & _EVAL_247;
  assign _EVAL_215 = _EVAL_96 | _EVAL_133;
  assign _EVAL_90 = _EVAL_246 & _EVAL_322;
  assign _EVAL_94 = _EVAL_306 & _EVAL_90;
  assign _EVAL_35 = _EVAL_96 | _EVAL_94;
  assign _EVAL_193 = _EVAL_218 == 1'h0;
  assign _EVAL_323 = _EVAL_69 & _EVAL_193;
  assign _EVAL_194 = _EVAL_308 | _EVAL_323;
  assign _EVAL_353 = _EVAL_193 & _EVAL_26;
  assign _EVAL_328 = _EVAL_206 & _EVAL_353;
  assign _EVAL_301 = _EVAL_194 | _EVAL_328;
  assign _EVAL_207 = _EVAL_353 & _EVAL_183;
  assign _EVAL_39 = _EVAL_306 & _EVAL_207;
  assign _EVAL_175 = _EVAL_301 | _EVAL_39;
  assign _EVAL_219 = _EVAL_353 & _EVAL_322;
  assign _EVAL_332 = _EVAL_306 & _EVAL_219;
  assign _EVAL_111 = _EVAL_301 | _EVAL_332;
  assign _EVAL_195 = _EVAL_193 & _EVAL_55;
  assign _EVAL_369 = _EVAL_206 & _EVAL_195;
  assign _EVAL_331 = _EVAL_194 | _EVAL_369;
  assign _EVAL_67 = _EVAL_195 & _EVAL_183;
  assign _EVAL_382 = _EVAL_306 & _EVAL_67;
  assign _EVAL_144 = _EVAL_331 | _EVAL_382;
  assign _EVAL_371 = _EVAL_195 & _EVAL_322;
  assign _EVAL_249 = _EVAL_306 & _EVAL_371;
  assign _EVAL_251 = _EVAL_331 | _EVAL_249;
  assign _EVAL_320 = {_EVAL_173,_EVAL_184,_EVAL_215,_EVAL_35,_EVAL_175,_EVAL_111,_EVAL_144,_EVAL_251};
  assign _EVAL_187 = _EVAL_14 == _EVAL_320;
  assign _EVAL_362 = _EVAL_308 | _EVAL_13;
  assign _EVAL_115 = _EVAL_12 == _EVAL_151;
  assign _EVAL_227 = _EVAL_115 | _EVAL_13;
  assign _EVAL_174 = _EVAL_227 == 1'h0;
  assign _EVAL_145 = _EVAL_1 <= 3'h3;
  assign _EVAL_54 = _EVAL_145 | _EVAL_13;
  assign _EVAL_244 = _EVAL_54 == 1'h0;
  assign _EVAL_56 = {1'b0,$signed(_EVAL_6)};
  assign _EVAL_278 = $signed(_EVAL_56) & $signed(-31'sh5000);
  assign _EVAL_388 = $signed(_EVAL_278);
  assign _EVAL_266 = _EVAL_296 | _EVAL_223;
  assign _EVAL_271 = _EVAL_2 <= 3'h6;
  assign _EVAL_360 = _EVAL_271 | _EVAL_13;
  assign _EVAL_196 = _EVAL_360 == 1'h0;
  assign _EVAL_72 = _EVAL_1 <= 3'h4;
  assign _EVAL_364 = _EVAL_72 | _EVAL_13;
  assign _EVAL_78 = _EVAL_1 == 3'h0;
  assign _EVAL_343 = _EVAL_78 | _EVAL_13;
  assign _EVAL_126 = _EVAL_343 == 1'h0;
  assign _EVAL_307 = _EVAL_83 == 5'h0;
  assign _EVAL_138 = _EVAL_307 == 1'h0;
  assign _EVAL_281 = _EVAL_3 == 7'h48;
  assign _EVAL_316 = _EVAL_6 ^ 30'h3000;
  assign _EVAL_47 = {1'b0,$signed(_EVAL_316)};
  assign _EVAL_89 = $signed(_EVAL_47) & $signed(-31'sh1000);
  assign _EVAL_265 = $signed(_EVAL_89);
  assign _EVAL_276 = $signed(_EVAL_265) == $signed(31'sh0);
  assign _EVAL_334 = _EVAL_6 ^ 30'hc000000;
  assign _EVAL_282 = {1'b0,$signed(_EVAL_334)};
  assign _EVAL_287 = $signed(_EVAL_282) & $signed(-31'sh4000000);
  assign _EVAL_49 = $signed(_EVAL_287);
  assign _EVAL_165 = $signed(_EVAL_49) == $signed(31'sh0);
  assign _EVAL_178 = _EVAL_276 | _EVAL_165;
  assign _EVAL_68 = _EVAL_6 ^ 30'h2000000;
  assign _EVAL_291 = {1'b0,$signed(_EVAL_68)};
  assign _EVAL_203 = $signed(_EVAL_291) & $signed(-31'sh10000);
  assign _EVAL_142 = $signed(_EVAL_203);
  assign _EVAL_135 = $signed(_EVAL_142) == $signed(31'sh0);
  assign _EVAL_357 = _EVAL_178 | _EVAL_135;
  assign _EVAL_181 = _EVAL_11 == 7'h40;
  assign _EVAL_318 = 4'h6 == _EVAL_9;
  assign _EVAL_101 = _EVAL_181 ? _EVAL_318 : 1'h0;
  assign _EVAL_392 = _EVAL_5 & _EVAL_4;
  assign _EVAL_243 = _EVAL_182 == 5'h0;
  assign _EVAL_254 = _EVAL_392 & _EVAL_243;
  assign _EVAL_214 = _EVAL_2 == 3'h6;
  assign _EVAL_88 = _EVAL_214 == 1'h0;
  assign _EVAL_46 = _EVAL_254 & _EVAL_88;
  assign _EVAL_192 = 128'h1 << _EVAL_3;
  assign _EVAL_93 = _EVAL_46 ? _EVAL_192 : 128'h0;
  assign _EVAL_24 = _EVAL_93[72:0];
  assign _EVAL_228 = _EVAL_296 != _EVAL_24;
  assign _EVAL_31 = _EVAL_370 == 1'h0;
  assign _EVAL_137 = _EVAL_228 | _EVAL_31;
  assign _EVAL_60 = _EVAL_137 | _EVAL_13;
  assign _EVAL_134 = _EVAL_101 | _EVAL_13;
  assign _EVAL_87 = _EVAL_6 ^ 30'h20000000;
  assign _EVAL_163 = {1'b0,$signed(_EVAL_87)};
  assign _EVAL_239 = $signed(_EVAL_163) & $signed(-31'sh2000);
  assign _EVAL_170 = $signed(_EVAL_239);
  assign _EVAL_118 = _EVAL_342 & _EVAL_307;
  assign _EVAL_121 = _EVAL_6 ^ 30'h1800000;
  assign _EVAL_255 = _EVAL_1 == _EVAL_21;
  assign _EVAL_365 = _EVAL_3 == 7'h40;
  assign _EVAL_216 = _EVAL_281 | _EVAL_365;
  assign _EVAL_129 = _EVAL_110 - 5'h1;
  assign _EVAL_381 = ~ _EVAL_14;
  assign _EVAL_58 = _EVAL_381 == 8'h0;
  assign _EVAL_319 = _EVAL_1 != 3'h0;
  assign _EVAL_210 = _EVAL_223 >> _EVAL_11;
  assign _EVAL_190 = _EVAL_210[0];
  assign _EVAL_238 = _EVAL_190 == 1'h0;
  assign _EVAL_347 = _EVAL_238 | _EVAL_13;
  assign _EVAL_23 = _EVAL_347 == 1'h0;
  assign _EVAL_275 = 23'hff << _EVAL_9;
  assign _EVAL_208 = _EVAL_275[7:0];
  assign _EVAL_245 = ~ _EVAL_208;
  assign _EVAL_393 = {{22'd0}, _EVAL_245};
  assign _EVAL_153 = _EVAL_6 & _EVAL_393;
  assign _EVAL_325 = _EVAL_153 == 30'h0;
  assign _EVAL_314 = _EVAL_325 | _EVAL_13;
  assign _EVAL_152 = _EVAL_2 == 3'h4;
  assign _EVAL_368 = _EVAL_4 & _EVAL_152;
  assign _EVAL_30 = _EVAL_223 != 73'h0;
  assign _EVAL_285 = _EVAL_30 == 1'h0;
  assign _EVAL_240 = plusarg_reader_out == 32'h0;
  assign _EVAL_236 = _EVAL_285 | _EVAL_240;
  assign _EVAL_122 = _EVAL_97 < plusarg_reader_out;
  assign _EVAL_298 = _EVAL_236 | _EVAL_122;
  assign _EVAL_43 = _EVAL_298 | _EVAL_13;
  assign _EVAL_50 = 23'hff << _EVAL;
  assign _EVAL_398 = _EVAL_50[7:0];
  assign _EVAL_310 = ~ _EVAL_398;
  assign _EVAL_85 = _EVAL_11 == _EVAL_292;
  assign _EVAL_312 = _EVAL_12 == 1'h0;
  assign _EVAL_123 = _EVAL_312 | _EVAL_13;
  assign _EVAL_394 = _EVAL_123 == 1'h0;
  assign _EVAL_146 = _EVAL_200 == 5'h0;
  assign _EVAL_171 = _EVAL_165 | _EVAL_135;
  assign _EVAL_376 = $signed(_EVAL_388) == $signed(31'sh0);
  assign _EVAL_286 = _EVAL_171 | _EVAL_376;
  assign _EVAL_349 = _EVAL_11 == 7'h48;
  assign _EVAL_179 = _EVAL_349 | _EVAL_181;
  assign _EVAL_125 = _EVAL_224 == 4'h8;
  assign _EVAL_81 = _EVAL_11[2:0];
  assign _EVAL_185 = 3'h1 <= _EVAL_81;
  assign _EVAL_222 = _EVAL_125 & _EVAL_185;
  assign _EVAL_124 = _EVAL_179 | _EVAL_222;
  assign _EVAL_262 = _EVAL_11 == 7'h20;
  assign _EVAL_136 = _EVAL_124 | _EVAL_262;
  assign _EVAL_366 = _EVAL_224 == 4'h0;
  assign _EVAL_248 = _EVAL_136 | _EVAL_366;
  assign _EVAL_252 = _EVAL_224 == 4'h1;
  assign _EVAL_66 = _EVAL_248 | _EVAL_252;
  assign _EVAL_150 = _EVAL_224 == 4'h2;
  assign _EVAL_373 = _EVAL_66 | _EVAL_150;
  assign _EVAL_225 = _EVAL_224 == 4'h3;
  assign _EVAL_139 = _EVAL_373 | _EVAL_225;
  assign _EVAL_102 = _EVAL_139 | _EVAL_13;
  assign _EVAL_354 = _EVAL_102 == 1'h0;
  assign _EVAL_387 = _EVAL_3[6:3];
  assign _EVAL_65 = _EVAL_387 == 4'h8;
  assign _EVAL_267 = _EVAL_3[2:0];
  assign _EVAL_250 = 3'h1 <= _EVAL_267;
  assign _EVAL_231 = _EVAL_65 & _EVAL_250;
  assign _EVAL_32 = _EVAL_216 | _EVAL_231;
  assign _EVAL_108 = _EVAL_3 == 7'h20;
  assign _EVAL_22 = _EVAL_32 | _EVAL_108;
  assign _EVAL_338 = _EVAL_387 == 4'h0;
  assign _EVAL_378 = _EVAL_22 | _EVAL_338;
  assign _EVAL_395 = _EVAL_387 == 4'h1;
  assign _EVAL_391 = _EVAL_378 | _EVAL_395;
  assign _EVAL_209 = _EVAL_9 <= 4'h8;
  assign _EVAL_337 = _EVAL_209 & _EVAL_276;
  assign _EVAL_63 = _EVAL_9 <= 4'h6;
  assign _EVAL_52 = {1'b0,$signed(_EVAL_121)};
  assign _EVAL_257 = $signed(_EVAL_52) & $signed(-31'sh8000);
  assign _EVAL_188 = $signed(_EVAL_257);
  assign _EVAL_315 = $signed(_EVAL_188) == $signed(31'sh0);
  assign _EVAL_82 = _EVAL_286 | _EVAL_315;
  assign _EVAL_44 = _EVAL_6 ^ 30'h1900000;
  assign _EVAL_311 = {1'b0,$signed(_EVAL_44)};
  assign _EVAL_106 = $signed(_EVAL_311) & $signed(-31'sh2000);
  assign _EVAL_258 = $signed(_EVAL_106);
  assign _EVAL_36 = $signed(_EVAL_258) == $signed(31'sh0);
  assign _EVAL_305 = _EVAL_82 | _EVAL_36;
  assign _EVAL_213 = $signed(_EVAL_170) == $signed(31'sh0);
  assign _EVAL_180 = _EVAL_305 | _EVAL_213;
  assign _EVAL_168 = _EVAL_63 & _EVAL_180;
  assign _EVAL_120 = _EVAL_337 | _EVAL_168;
  assign _EVAL_149 = _EVAL_16 == 1'h0;
  assign _EVAL_103 = _EVAL_149 | _EVAL_13;
  assign _EVAL_162 = _EVAL_103 == 1'h0;
  assign _EVAL_274 = _EVAL_2[0];
  assign _EVAL_399 = _EVAL_310[7:3];
  assign _EVAL_156 = _EVAL_200 - 5'h1;
  assign _EVAL_348 = _EVAL_245[7:3];
  assign _EVAL_336 = _EVAL_18 == _EVAL_45;
  assign _EVAL_160 = _EVAL_17 <= 2'h2;
  assign _EVAL_99 = _EVAL_160 | _EVAL_13;
  assign _EVAL_157 = _EVAL_99 == 1'h0;
  assign _EVAL_159 = _EVAL_146 == 1'h0;
  assign _EVAL_212 = _EVAL_4 & _EVAL_159;
  assign _EVAL_261 = _EVAL_2 == 3'h0;
  assign _EVAL_41 = _EVAL_4 & _EVAL_261;
  assign _EVAL_77 = _EVAL_0 == 1'h0;
  assign _EVAL_350 = _EVAL_77 | _EVAL_13;
  assign _EVAL_75 = _EVAL_350 == 1'h0;
  assign _EVAL_84 = _EVAL_18[2];
  assign _EVAL_273 = _EVAL_84 == 1'h0;
  assign _EVAL_300 = _EVAL_336 | _EVAL_13;
  assign _EVAL_116 = _EVAL_300 == 1'h0;
  assign _EVAL_242 = ~ _EVAL_320;
  assign _EVAL_279 = _EVAL_14 & _EVAL_242;
  assign _EVAL_53 = _EVAL_279 == 8'h0;
  assign _EVAL_70 = _EVAL_18 == 3'h1;
  assign _EVAL_268 = _EVAL_7 & _EVAL_70;
  assign _EVAL_397 = _EVAL_18 == 3'h5;
  assign _EVAL_25 = _EVAL_337 | _EVAL_13;
  assign _EVAL_38 = _EVAL_2 == 3'h2;
  assign _EVAL_199 = _EVAL_4 & _EVAL_214;
  assign _EVAL_48 = _EVAL_387 == 4'h2;
  assign _EVAL_344 = _EVAL_391 | _EVAL_48;
  assign _EVAL_19 = _EVAL_387 == 4'h3;
  assign _EVAL_309 = _EVAL_344 | _EVAL_19;
  assign _EVAL_57 = _EVAL_309 | _EVAL_13;
  assign _EVAL_389 = _EVAL_57 == 1'h0;
  assign _EVAL_51 = _EVAL_53 | _EVAL_13;
  assign _EVAL_375 = _EVAL_18 == 3'h6;
  assign _EVAL_86 = _EVAL_17 != 2'h2;
  assign _EVAL_339 = _EVAL_86 | _EVAL_13;
  assign _EVAL_232 = _EVAL_339 == 1'h0;
  assign _EVAL_299 = _EVAL_9 <= 4'h2;
  assign _EVAL_109 = _EVAL_357 | _EVAL_376;
  assign _EVAL_64 = _EVAL_109 | _EVAL_315;
  assign _EVAL_132 = _EVAL_64 | _EVAL_36;
  assign _EVAL_28 = _EVAL_132 | _EVAL_213;
  assign _EVAL_62 = _EVAL_299 & _EVAL_28;
  assign _EVAL_117 = _EVAL_62 | _EVAL_13;
  assign _EVAL_177 = _EVAL_83 - 5'h1;
  assign _EVAL_130 = _EVAL_17 == 2'h0;
  assign _EVAL_374 = _EVAL_319 | _EVAL_13;
  assign _EVAL_112 = _EVAL_374 == 1'h0;
  assign _EVAL_358 = _EVAL_6 == _EVAL_107;
  assign _EVAL_167 = _EVAL_358 | _EVAL_13;
  assign _EVAL_241 = _EVAL_85 | _EVAL_13;
  assign _EVAL_127 = _EVAL_241 == 1'h0;
  assign _EVAL_351 = _EVAL_182 - 5'h1;
  assign _EVAL_264 = _EVAL_3 == _EVAL_379;
  assign _EVAL_100 = _EVAL_264 | _EVAL_13;
  assign _EVAL_147 = _EVAL_100 == 1'h0;
  assign _EVAL_40 = _EVAL_18 == 3'h3;
  assign _EVAL_198 = _EVAL_7 & _EVAL_40;
  assign _EVAL_329 = _EVAL_25 == 1'h0;
  assign _EVAL_293 = _EVAL_58 | _EVAL_13;
  assign _EVAL_92 = _EVAL_187 | _EVAL_13;
  assign _EVAL_235 = _EVAL_266 >> _EVAL_3;
  assign _EVAL_352 = _EVAL_235[0];
  assign _EVAL_105 = _EVAL_352 | _EVAL_13;
  assign _EVAL_205 = _EVAL_1 <= 3'h2;
  assign _EVAL_383 = _EVAL_205 | _EVAL_13;
  assign _EVAL_42 = _EVAL_383 == 1'h0;
  assign _EVAL_226 = _EVAL_392 & _EVAL_146;
  assign _EVAL_355 = _EVAL_7 & _EVAL_397;
  assign _EVAL_384 = _EVAL_167 == 1'h0;
  assign _EVAL_155 = _EVAL_130 | _EVAL_13;
  assign _EVAL_98 = _EVAL_155 == 1'h0;
  assign _EVAL_385 = _EVAL_18 == 3'h2;
  assign _EVAL_27 = _EVAL_7 & _EVAL_385;
  assign _EVAL_211 = _EVAL_223 | _EVAL_296;
  assign _EVAL_302 = ~ _EVAL_24;
  assign _EVAL_386 = _EVAL_211 & _EVAL_302;
  assign _EVAL_377 = _EVAL_9 == _EVAL_197;
  assign _EVAL_29 = _EVAL_377 | _EVAL_13;
  assign _EVAL_140 = _EVAL_60 == 1'h0;
  assign _EVAL_141 = _EVAL_2 == 3'h5;
  assign _EVAL_74 = _EVAL_18 == 3'h7;
  assign _EVAL_263 = _EVAL_312 | _EVAL_0;
  assign _EVAL_73 = _EVAL_263 | _EVAL_13;
  assign _EVAL_189 = _EVAL_73 == 1'h0;
  assign _EVAL_59 = _EVAL_15 == _EVAL_304;
  assign _EVAL_148 = _EVAL_13 == 1'h0;
  assign _EVAL_95 = _EVAL_2 == _EVAL_176;
  assign _EVAL_113 = _EVAL_362 == 1'h0;
  assign _EVAL_204 = _EVAL_4 & _EVAL_141;
  assign _EVAL_201 = _EVAL_59 | _EVAL_13;
  assign _EVAL_289 = _EVAL_201 == 1'h0;
  assign _EVAL_335 = _EVAL == _EVAL_229;
  assign _EVAL_37 = _EVAL_335 | _EVAL_13;
  assign _EVAL_359 = _EVAL_37 == 1'h0;
  assign _EVAL_356 = _EVAL_51 == 1'h0;
  assign _EVAL_61 = _EVAL_7 & _EVAL_74;
  assign _EVAL_284 = _EVAL_342 | _EVAL_392;
  assign _EVAL_230 = _EVAL_364 == 1'h0;
  assign _EVAL_71 = _EVAL_255 | _EVAL_13;
  assign _EVAL_346 = _EVAL_71 == 1'h0;
  assign _EVAL_372 = _EVAL_97 + 32'h1;
  assign _EVAL_233 = _EVAL_120 | _EVAL_13;
  assign _EVAL_270 = _EVAL_7 & _EVAL_138;
  assign _EVAL_143 = _EVAL_314 == 1'h0;
  assign _EVAL_220 = _EVAL_29 == 1'h0;
  assign _EVAL_119 = _EVAL_134 == 1'h0;
  assign _EVAL_363 = _EVAL_2 == 3'h1;
  assign _EVAL_290 = _EVAL_4 & _EVAL_363;
  assign _EVAL_260 = _EVAL_95 | _EVAL_13;
  assign _EVAL_76 = _EVAL_4 & _EVAL_38;
  assign _EVAL_33 = _EVAL_233 == 1'h0;
  assign _EVAL_80 = _EVAL_117 == 1'h0;
  assign _EVAL_283 = _EVAL_18 == 3'h0;
  assign _EVAL_326 = _EVAL_7 & _EVAL_283;
  assign _EVAL_253 = _EVAL_18 == 3'h4;
  assign _EVAL_169 = _EVAL_7 & _EVAL_253;
  assign _EVAL_256 = _EVAL_260 == 1'h0;
  assign _EVAL_259 = _EVAL_105 == 1'h0;
  assign _EVAL_390 = _EVAL_7 & _EVAL_375;
  assign _EVAL_221 = _EVAL_43 == 1'h0;
  assign _EVAL_79 = _EVAL_92 == 1'h0;
  assign _EVAL_217 = _EVAL_293 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_21 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_45 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_83 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_97 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_107 = _RAND_4[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_110 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_151 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_176 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_182 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_197 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_200 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {3{`RANDOM}};
  _EVAL_223 = _RAND_11[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_229 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_292 = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_304 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_340 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_379 = _RAND_16[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_8) begin
    if (_EVAL_118) begin
      _EVAL_21 <= _EVAL_1;
    end
    if (_EVAL_118) begin
      _EVAL_45 <= _EVAL_18;
    end
    if (_EVAL_13) begin
      _EVAL_83 <= 5'h0;
    end else begin
      if (_EVAL_342) begin
        if (_EVAL_307) begin
          if (_EVAL_273) begin
            _EVAL_83 <= _EVAL_348;
          end else begin
            _EVAL_83 <= 5'h0;
          end
        end else begin
          _EVAL_83 <= _EVAL_177;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_97 <= 32'h0;
    end else begin
      if (_EVAL_284) begin
        _EVAL_97 <= 32'h0;
      end else begin
        _EVAL_97 <= _EVAL_372;
      end
    end
    if (_EVAL_118) begin
      _EVAL_107 <= _EVAL_6;
    end
    if (_EVAL_13) begin
      _EVAL_110 <= 5'h0;
    end else begin
      if (_EVAL_342) begin
        if (_EVAL_164) begin
          if (_EVAL_273) begin
            _EVAL_110 <= _EVAL_348;
          end else begin
            _EVAL_110 <= 5'h0;
          end
        end else begin
          _EVAL_110 <= _EVAL_129;
        end
      end
    end
    if (_EVAL_226) begin
      _EVAL_151 <= _EVAL_12;
    end
    if (_EVAL_226) begin
      _EVAL_176 <= _EVAL_2;
    end
    if (_EVAL_13) begin
      _EVAL_182 <= 5'h0;
    end else begin
      if (_EVAL_392) begin
        if (_EVAL_243) begin
          if (_EVAL_274) begin
            _EVAL_182 <= _EVAL_399;
          end else begin
            _EVAL_182 <= 5'h0;
          end
        end else begin
          _EVAL_182 <= _EVAL_351;
        end
      end
    end
    if (_EVAL_118) begin
      _EVAL_197 <= _EVAL_9;
    end
    if (_EVAL_13) begin
      _EVAL_200 <= 5'h0;
    end else begin
      if (_EVAL_392) begin
        if (_EVAL_146) begin
          if (_EVAL_274) begin
            _EVAL_200 <= _EVAL_399;
          end else begin
            _EVAL_200 <= 5'h0;
          end
        end else begin
          _EVAL_200 <= _EVAL_156;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_223 <= 73'h0;
    end else begin
      _EVAL_223 <= _EVAL_386;
    end
    if (_EVAL_226) begin
      _EVAL_229 <= _EVAL;
    end
    if (_EVAL_118) begin
      _EVAL_292 <= _EVAL_11;
    end
    if (_EVAL_226) begin
      _EVAL_304 <= _EVAL_15;
    end
    if (_EVAL_226) begin
      _EVAL_340 <= _EVAL_17;
    end
    if (_EVAL_226) begin
      _EVAL_379 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef728723)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0d9d9fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5987ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_384) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ecedcc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(916cf201)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b921c045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21f1612f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(184515bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22754c31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a496a0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_346) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5876558d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e0647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(373f159e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_384) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14796d10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21bae347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4ff46a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a637ba43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b824b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(168c2546)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f20acd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_394) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d5d84d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5663f401)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e9e0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c5a9d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b89930b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_329) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d245e171)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5140fcd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_359) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85bfc151)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bad7938b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(992ead0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7adf9d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_356) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b1e5ed4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bb21e26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40142f9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e93781)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e0b4249)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(537460aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_346) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fa059e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3f25940)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ab2ce0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8658ffb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531e9cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(547cd28c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_329) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc426477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c5eb33c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f0b91ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e41482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb6fc2dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(972fbe50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ed85b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25f90f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c143101a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a561846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7997cf4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8cd62c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(396f608c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(443d1e61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d22af7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_356) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fc92477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(def06a6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1487c90c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(753e58d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(223a2ae4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a56f2031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57e41483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1338ba0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d586d83d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a018e4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9332d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70129ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f05d76d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_394) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a28b179f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4626e29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d4ecb57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68082364)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfba56f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(190d195c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeb6793d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbb7b477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2944a1bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b96ce9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d5dcef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65d3ac94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0bdd017)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(864aad3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(321567df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f81b03a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77c301b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3d00270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfa58a05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
