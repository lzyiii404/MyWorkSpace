//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_151(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  output [1:0]  _EVAL_3,
  output        _EVAL_4,
  output [2:0]  _EVAL_5,
  output [2:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [24:0] _EVAL_8,
  input         _EVAL_9,
  output [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  output [24:0] _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  output [2:0]  _EVAL_19,
  output        _EVAL_20,
  output [3:0]  _EVAL_21,
  output        _EVAL_22,
  output [6:0]  _EVAL_23,
  input  [2:0]  _EVAL_24,
  input         _EVAL_25,
  input  [6:0]  _EVAL_26,
  output [6:0]  _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  input  [2:0]  _EVAL_30,
  input         _EVAL_31,
  input  [6:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  output        _EVAL_36,
  output [31:0] _EVAL_37,
  output [31:0] _EVAL_38,
  input  [3:0]  _EVAL_39,
  input         _EVAL_40
);
  assign _EVAL_21 = _EVAL_39;
  assign _EVAL_17 = _EVAL_34;
  assign _EVAL_28 = _EVAL_40;
  assign _EVAL_27 = _EVAL_26;
  assign _EVAL_20 = _EVAL_13;
  assign _EVAL_15 = _EVAL_8;
  assign _EVAL_4 = _EVAL_35;
  assign _EVAL_18 = _EVAL_9;
  assign _EVAL_10 = _EVAL_12;
  assign _EVAL_36 = _EVAL_11;
  assign _EVAL_5 = _EVAL_30;
  assign _EVAL_6 = _EVAL_24;
  assign _EVAL_37 = _EVAL_14;
  assign _EVAL_23 = _EVAL_32;
  assign _EVAL_3 = _EVAL_2;
  assign _EVAL_0 = _EVAL_1;
  assign _EVAL_19 = _EVAL_7;
  assign _EVAL_38 = _EVAL_33;
  assign _EVAL_22 = _EVAL_31;
  assign _EVAL_16 = _EVAL;
endmodule
