//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_307(
  output         _EVAL,
  output         _EVAL_0,
  input          _EVAL_1,
  input  [31:0]  _EVAL_2,
  output         _EVAL_3,
  input          _EVAL_4,
  output [31:0]  _EVAL_5,
  input  [4:0]   _EVAL_6,
  output [1:0]   _EVAL_7,
  output         _EVAL_8,
  output [31:0]  _EVAL_9,
  output [31:0]  _EVAL_10,
  output [1:0]   _EVAL_11,
  output         _EVAL_12,
  output [1:0]   _EVAL_13,
  output [1:0]   _EVAL_14,
  input  [1:0]   _EVAL_15,
  input          _EVAL_16,
  output [1:0]   _EVAL_17,
  output [127:0] _EVAL_18,
  output         _EVAL_19,
  input          _EVAL_20,
  output [31:0]  _EVAL_21,
  input          _EVAL_22,
  input  [127:0] _EVAL_23,
  input          _EVAL_24,
  input  [5:0]   _EVAL_25,
  output         _EVAL_26,
  output         _EVAL_27,
  output         _EVAL_28,
  input          _EVAL_29,
  output         _EVAL_30,
  input          _EVAL_31,
  input          _EVAL_32,
  output         _EVAL_33,
  output         _EVAL_34,
  input          _EVAL_35,
  input          _EVAL_36,
  output [29:0]  _EVAL_37,
  output [1:0]   _EVAL_38,
  input          _EVAL_39,
  input          _EVAL_40,
  output         _EVAL_41,
  output         _EVAL_42,
  output         _EVAL_43,
  output [31:0]  _EVAL_44,
  input          _EVAL_45,
  output [29:0]  _EVAL_46,
  input          _EVAL_47,
  output         _EVAL_48,
  output         _EVAL_49,
  output         _EVAL_50,
  input  [14:0]  _EVAL_51,
  output         _EVAL_52,
  output         _EVAL_53,
  output         _EVAL_54,
  input          _EVAL_55,
  output         _EVAL_56,
  input          _EVAL_57,
  input          _EVAL_58,
  input          _EVAL_59,
  output         _EVAL_60,
  output [29:0]  _EVAL_61,
  output [31:0]  _EVAL_62,
  input          _EVAL_63,
  input  [14:0]  _EVAL_64,
  output         _EVAL_65,
  output [29:0]  _EVAL_66,
  output         _EVAL_67,
  input  [4:0]   _EVAL_68,
  output         _EVAL_69,
  output         _EVAL_70,
  input          _EVAL_71,
  output         _EVAL_72,
  input  [6:0]   _EVAL_73,
  output         _EVAL_74,
  output [2:0]   _EVAL_75,
  input          _EVAL_76,
  output         _EVAL_77,
  input          _EVAL_78,
  output         _EVAL_79,
  input          _EVAL_80,
  input          _EVAL_81,
  output         _EVAL_82,
  output         _EVAL_83,
  input  [2:0]   _EVAL_84,
  output [31:0]  _EVAL_85,
  output         _EVAL_86,
  input          _EVAL_87,
  output [29:0]  _EVAL_88,
  output [29:0]  _EVAL_89,
  input          _EVAL_90,
  input  [4:0]   _EVAL_91,
  input          _EVAL_92,
  output         _EVAL_93,
  output [5:0]   _EVAL_94,
  input          _EVAL_95,
  input  [1:0]   _EVAL_96,
  input  [127:0] _EVAL_97,
  input          _EVAL_98,
  output [2:0]   _EVAL_99,
  output         _EVAL_100,
  output         _EVAL_101,
  input          _EVAL_102,
  output         _EVAL_103,
  input          _EVAL_104,
  input          _EVAL_105,
  input          _EVAL_106,
  input          _EVAL_107,
  input          _EVAL_108,
  output         _EVAL_109,
  input  [31:0]  _EVAL_110,
  input  [5:0]   _EVAL_111,
  output         _EVAL_112,
  output         _EVAL_113,
  output         _EVAL_114,
  input          _EVAL_115,
  output         _EVAL_116,
  output         _EVAL_117,
  output         _EVAL_118,
  input          _EVAL_119,
  output         _EVAL_120,
  input  [6:0]   _EVAL_121,
  input          _EVAL_122,
  output         _EVAL_123,
  output         _EVAL_124,
  output         _EVAL_125,
  output [31:0]  _EVAL_126,
  input          _EVAL_127,
  output         _EVAL_128,
  output         _EVAL_129,
  output         _EVAL_130,
  output         _EVAL_131,
  output [1:0]   _EVAL_132,
  input  [31:0]  _EVAL_133,
  input          _EVAL_134,
  output [1:0]   _EVAL_135,
  output         _EVAL_136,
  input          _EVAL_137,
  input  [31:0]  _EVAL_138,
  output         _EVAL_139,
  output         _EVAL_140,
  input          _EVAL_141,
  input          _EVAL_142,
  output [1:0]   _EVAL_143,
  output         _EVAL_144,
  output         _EVAL_145,
  input          _EVAL_146,
  input          _EVAL_147,
  input          _EVAL_148,
  output         _EVAL_149,
  output         _EVAL_150,
  output [31:0]  _EVAL_151,
  output         _EVAL_152,
  input  [2:0]   _EVAL_153,
  input  [4:0]   _EVAL_154,
  output         _EVAL_155,
  input          _EVAL_156,
  output         _EVAL_157,
  input  [2:0]   _EVAL_158,
  input          _EVAL_159,
  output         _EVAL_160,
  output [1:0]   _EVAL_161,
  output [31:0]  _EVAL_162,
  input          _EVAL_163,
  input          _EVAL_164,
  input          _EVAL_165,
  output [31:0]  _EVAL_166,
  output         _EVAL_167,
  input          _EVAL_168,
  input          _EVAL_169,
  input          _EVAL_170,
  input  [4:0]   _EVAL_171,
  input          _EVAL_172,
  output         _EVAL_173,
  input          _EVAL_174,
  input          _EVAL_175,
  input          _EVAL_176,
  output         _EVAL_177,
  output [1:0]   _EVAL_178,
  input          _EVAL_179,
  input  [4:0]   _EVAL_180,
  output         _EVAL_181,
  output         _EVAL_182,
  input  [2:0]   _EVAL_183,
  input          _EVAL_184,
  output [127:0] _EVAL_185,
  input          _EVAL_186,
  output [31:0]  _EVAL_187,
  input          _EVAL_188,
  output [31:0]  _EVAL_189,
  input          _EVAL_190,
  input  [4:0]   _EVAL_191,
  output         _EVAL_192,
  output         _EVAL_193,
  output [31:0]  _EVAL_194,
  output [31:0]  _EVAL_195,
  input          _EVAL_196,
  output         _EVAL_197,
  input          _EVAL_198,
  output [31:0]  _EVAL_199,
  output [31:0]  _EVAL_200,
  output         _EVAL_201,
  input  [1:0]   _EVAL_202,
  input  [4:0]   _EVAL_203,
  input          _EVAL_204,
  input          _EVAL_205,
  input          _EVAL_206,
  output         _EVAL_207,
  input  [2:0]   _EVAL_208,
  output [31:0]  _EVAL_209,
  output         _EVAL_210,
  output [1:0]   _EVAL_211,
  input          _EVAL_212,
  input          _EVAL_213,
  input          _EVAL_214,
  input          _EVAL_215,
  input          _EVAL_216,
  output [1:0]   _EVAL_217,
  output         _EVAL_218,
  output         _EVAL_219,
  input          _EVAL_220,
  output [1:0]   _EVAL_221,
  input  [2:0]   _EVAL_222,
  output         _EVAL_223,
  input          _EVAL_224,
  output         _EVAL_225,
  input          _EVAL_226,
  output         _EVAL_227,
  output         _EVAL_228,
  output         _EVAL_229,
  output [29:0]  _EVAL_230,
  output         _EVAL_231,
  input          _EVAL_232,
  input          _EVAL_233,
  input  [31:0]  _EVAL_234,
  output         _EVAL_235,
  input          _EVAL_236,
  input          _EVAL_237,
  output [31:0]  _EVAL_238,
  output         _EVAL_239,
  output [31:0]  _EVAL_240,
  output [1:0]   _EVAL_241,
  input          _EVAL_242,
  output         _EVAL_243,
  output         _EVAL_244,
  output         _EVAL_245,
  input          _EVAL_246,
  input          _EVAL_247,
  output [4:0]   _EVAL_248,
  input          _EVAL_249,
  input          _EVAL_250,
  input          _EVAL_251,
  output         _EVAL_252,
  output         _EVAL_253,
  output         _EVAL_254,
  input          _EVAL_255,
  output [1:0]   _EVAL_256,
  output         _EVAL_257,
  output         _EVAL_258,
  input          _EVAL_259,
  input          _EVAL_260,
  input          _EVAL_261,
  output [1:0]   _EVAL_262,
  output [31:0]  _EVAL_263,
  output [29:0]  _EVAL_264,
  input          _EVAL_265,
  output [31:0]  _EVAL_266,
  input          _EVAL_267,
  input          _EVAL_268,
  output [31:0]  _EVAL_269,
  input  [31:0]  _EVAL_270,
  output         _EVAL_271,
  input          _EVAL_272,
  output [31:0]  _EVAL_273,
  input  [4:0]   _EVAL_274,
  output [14:0]  _EVAL_275,
  output         _EVAL_276,
  input          _EVAL_277,
  input          _EVAL_278,
  output         _EVAL_279
);
  wire  fpu__EVAL;
  wire [2:0] fpu__EVAL_0;
  wire  fpu__EVAL_1;
  wire [32:0] fpu__EVAL_2;
  wire [6:0] fpu__EVAL_3;
  wire  fpu__EVAL_4;
  wire [4:0] fpu__EVAL_5;
  wire [32:0] fpu__EVAL_6;
  wire  fpu__EVAL_7;
  wire  fpu__EVAL_8;
  wire [31:0] fpu__EVAL_9;
  wire [2:0] fpu__EVAL_10;
  wire [4:0] fpu__EVAL_11;
  wire  fpu__EVAL_12;
  wire  fpu__EVAL_13;
  wire  fpu__EVAL_14;
  wire  fpu__EVAL_15;
  wire  fpu__EVAL_16;
  wire [6:0] fpu__EVAL_17;
  wire [4:0] fpu__EVAL_18;
  wire [32:0] fpu__EVAL_19;
  wire  fpu__EVAL_20;
  wire [32:0] fpu__EVAL_21;
  wire  fpu__EVAL_22;
  wire [6:0] fpu__EVAL_23;
  wire  fpu__EVAL_24;
  wire [4:0] fpu__EVAL_25;
  wire [4:0] fpu__EVAL_26;
  wire [31:0] fpu__EVAL_27;
  wire [4:0] fpu__EVAL_28;
  wire [4:0] fpu__EVAL_29;
  wire [32:0] fpu__EVAL_30;
  wire [2:0] fpu__EVAL_31;
  wire [32:0] fpu__EVAL_32;
  wire  fpu__EVAL_33;
  wire [2:0] fpu__EVAL_34;
  wire [4:0] fpu__EVAL_35;
  wire  fpu__EVAL_36;
  wire [4:0] fpu__EVAL_37;
  wire  fpu__EVAL_38;
  wire [2:0] fpu__EVAL_39;
  wire  fpu__EVAL_40;
  wire  fpu__EVAL_41;
  wire  fpu__EVAL_42;
  wire [4:0] fpu__EVAL_43;
  wire  fpu__EVAL_44;
  wire [4:0] fpu__EVAL_45;
  wire  fpu__EVAL_46;
  wire [4:0] fpu__EVAL_47;
  wire  fpu__EVAL_48;
  wire  fpu__EVAL_49;
  wire [6:0] fpu__EVAL_50;
  wire [2:0] fpu__EVAL_51;
  wire  fpu__EVAL_52;
  wire  fpu__EVAL_53;
  wire [4:0] fpu__EVAL_54;
  wire  fpu__EVAL_55;
  wire  fpu__EVAL_56;
  wire [4:0] fpu__EVAL_57;
  wire  fpu__EVAL_58;
  wire [6:0] fpu__EVAL_59;
  wire [32:0] fpu__EVAL_60;
  wire  bullet_clock_gate_in;
  wire  bullet_clock_gate_en;
  wire  bullet_clock_gate_out;
  wire  divider__EVAL;
  wire  divider__EVAL_0;
  wire [31:0] divider__EVAL_1;
  wire  divider__EVAL_2;
  wire  divider__EVAL_3;
  wire [3:0] divider__EVAL_4;
  wire [4:0] divider__EVAL_5;
  wire [31:0] divider__EVAL_6;
  wire  divider__EVAL_7;
  wire [31:0] divider__EVAL_8;
  wire  divider__EVAL_9;
  wire  divider__EVAL_10;
  wire [4:0] divider__EVAL_11;
  wire [31:0] csr__EVAL;
  wire [29:0] csr__EVAL_0;
  wire [1:0] csr__EVAL_1;
  wire [31:0] csr__EVAL_2;
  wire  csr__EVAL_3;
  wire [7:0] csr__EVAL_4;
  wire  csr__EVAL_5;
  wire  csr__EVAL_6;
  wire  csr__EVAL_7;
  wire [7:0] csr__EVAL_8;
  wire  csr__EVAL_9;
  wire  csr__EVAL_10;
  wire  csr__EVAL_11;
  wire [1:0] csr__EVAL_12;
  wire  csr__EVAL_13;
  wire [31:0] csr__EVAL_14;
  wire  csr__EVAL_15;
  wire  csr__EVAL_16;
  wire  csr__EVAL_17;
  wire [11:0] csr__EVAL_18;
  wire  csr__EVAL_19;
  wire  csr__EVAL_20;
  wire [1:0] csr__EVAL_21;
  wire [1:0] csr__EVAL_22;
  wire [2:0] csr__EVAL_23;
  wire  csr__EVAL_24;
  wire  csr__EVAL_25;
  wire  csr__EVAL_26;
  wire  csr__EVAL_27;
  wire  csr__EVAL_28;
  wire [1:0] csr__EVAL_29;
  wire [2:0] csr__EVAL_30;
  wire [1:0] csr__EVAL_31;
  wire  csr__EVAL_32;
  wire  csr__EVAL_33;
  wire  csr__EVAL_34;
  wire [1:0] csr__EVAL_35;
  wire  csr__EVAL_36;
  wire [29:0] csr__EVAL_37;
  wire  csr__EVAL_38;
  wire  csr__EVAL_39;
  wire [31:0] csr__EVAL_40;
  wire [1:0] csr__EVAL_41;
  wire  csr__EVAL_42;
  wire [1:0] csr__EVAL_43;
  wire [31:0] csr__EVAL_44;
  wire [1:0] csr__EVAL_45;
  wire  csr__EVAL_46;
  wire  csr__EVAL_47;
  wire  csr__EVAL_48;
  wire [1:0] csr__EVAL_49;
  wire  csr__EVAL_50;
  wire [31:0] csr__EVAL_51;
  wire  csr__EVAL_52;
  wire  csr__EVAL_53;
  wire [29:0] csr__EVAL_54;
  wire [1:0] csr__EVAL_55;
  wire  csr__EVAL_56;
  wire  csr__EVAL_57;
  wire  csr__EVAL_58;
  wire  csr__EVAL_59;
  wire  csr__EVAL_60;
  wire  csr__EVAL_61;
  wire  csr__EVAL_62;
  wire  csr__EVAL_63;
  wire [31:0] csr__EVAL_64;
  wire  csr__EVAL_65;
  wire [29:0] csr__EVAL_66;
  wire  csr__EVAL_67;
  wire [1:0] csr__EVAL_68;
  wire  csr__EVAL_69;
  wire  csr__EVAL_70;
  wire  csr__EVAL_71;
  wire  csr__EVAL_72;
  wire [1:0] csr__EVAL_73;
  wire  csr__EVAL_74;
  wire  csr__EVAL_75;
  wire [1:0] csr__EVAL_76;
  wire  csr__EVAL_77;
  wire [31:0] csr__EVAL_78;
  wire  csr__EVAL_79;
  wire [31:0] csr__EVAL_80;
  wire  csr__EVAL_81;
  wire [1:0] csr__EVAL_82;
  wire [31:0] csr__EVAL_83;
  wire [31:0] csr__EVAL_84;
  wire  csr__EVAL_85;
  wire  csr__EVAL_86;
  wire [31:0] csr__EVAL_87;
  wire [2:0] csr__EVAL_88;
  wire  csr__EVAL_89;
  wire  csr__EVAL_90;
  wire  csr__EVAL_91;
  wire  csr__EVAL_92;
  wire  csr__EVAL_93;
  wire  csr__EVAL_94;
  wire  csr__EVAL_95;
  wire [31:0] csr__EVAL_96;
  wire  csr__EVAL_97;
  wire  csr__EVAL_98;
  wire [2:0] csr__EVAL_99;
  wire [1:0] csr__EVAL_100;
  wire [29:0] csr__EVAL_101;
  wire [11:0] csr__EVAL_102;
  wire  csr__EVAL_103;
  wire  csr__EVAL_104;
  wire  csr__EVAL_105;
  wire  csr__EVAL_106;
  wire  csr__EVAL_107;
  wire  csr__EVAL_108;
  wire  csr__EVAL_109;
  wire  csr__EVAL_110;
  wire  csr__EVAL_111;
  wire  csr__EVAL_112;
  wire [31:0] csr__EVAL_113;
  wire  csr__EVAL_114;
  wire [7:0] csr__EVAL_115;
  wire  csr__EVAL_116;
  wire [31:0] csr__EVAL_117;
  wire [31:0] csr__EVAL_118;
  wire  csr__EVAL_119;
  wire [1:0] csr__EVAL_120;
  wire [1:0] csr__EVAL_121;
  wire  csr__EVAL_122;
  wire [31:0] csr__EVAL_123;
  wire  csr__EVAL_124;
  wire  csr__EVAL_125;
  wire [31:0] csr__EVAL_126;
  wire [26:0] csr__EVAL_127;
  wire  csr__EVAL_128;
  wire  csr__EVAL_129;
  wire  csr__EVAL_130;
  wire  csr__EVAL_131;
  wire [31:0] csr__EVAL_132;
  wire  csr__EVAL_133;
  wire  csr__EVAL_134;
  wire [1:0] csr__EVAL_135;
  wire [31:0] csr__EVAL_136;
  wire  csr__EVAL_137;
  wire [1:0] csr__EVAL_138;
  wire  csr__EVAL_139;
  wire  csr__EVAL_140;
  wire  csr__EVAL_141;
  wire [29:0] csr__EVAL_142;
  wire  csr__EVAL_143;
  wire [4:0] csr__EVAL_144;
  wire [31:0] csr__EVAL_145;
  wire  csr__EVAL_146;
  wire  csr__EVAL_147;
  wire  csr__EVAL_148;
  wire  csr__EVAL_149;
  wire  csr__EVAL_150;
  wire [1:0] csr__EVAL_151;
  wire  csr__EVAL_152;
  wire  csr__EVAL_153;
  wire  csr__EVAL_154;
  wire  csr__EVAL_155;
  wire [29:0] csr__EVAL_156;
  wire  csr__EVAL_157;
  wire [31:0] csr__EVAL_158;
  wire [1:0] csr__EVAL_159;
  wire [31:0] csr__EVAL_160;
  wire  csr__EVAL_161;
  wire [29:0] csr__EVAL_162;
  wire  csr__EVAL_163;
  wire  csr__EVAL_164;
  wire  csr__EVAL_165;
  wire [31:0] csr__EVAL_166;
  wire [31:0] csr__EVAL_167;
  wire  m__EVAL;
  wire [31:0] m__EVAL_0;
  wire  m__EVAL_1;
  wire [31:0] m__EVAL_2;
  wire [3:0] m__EVAL_3;
  wire [31:0] m__EVAL_4;
  wire  m__EVAL_5;
  wire  fpu_clock_gate_in;
  wire  fpu_clock_gate_en;
  wire  fpu_clock_gate_out;
  reg [31:0] _EVAL_708 [0:31];
  reg [31:0] _RAND_0;
  wire [31:0] _EVAL_708__EVAL_709_data;
  wire [4:0] _EVAL_708__EVAL_709_addr;
  wire [31:0] _EVAL_708__EVAL_710_data;
  wire [4:0] _EVAL_708__EVAL_710_addr;
  wire [31:0] _EVAL_708__EVAL_711_data;
  wire [4:0] _EVAL_708__EVAL_711_addr;
  wire [31:0] _EVAL_708__EVAL_712_data;
  wire [4:0] _EVAL_708__EVAL_712_addr;
  wire [31:0] _EVAL_708__EVAL_713_data;
  wire [4:0] _EVAL_708__EVAL_713_addr;
  wire  _EVAL_708__EVAL_713_mask;
  wire  _EVAL_708__EVAL_713_en;
  wire [31:0] _EVAL_708__EVAL_714_data;
  wire [4:0] _EVAL_708__EVAL_714_addr;
  wire  _EVAL_708__EVAL_714_mask;
  wire  _EVAL_708__EVAL_714_en;
  wire [31:0] _EVAL_708__EVAL_715_data;
  wire [4:0] _EVAL_708__EVAL_715_addr;
  wire  _EVAL_708__EVAL_715_mask;
  wire  _EVAL_708__EVAL_715_en;
  reg [32:0] _EVAL_2741 [0:31];
  reg [63:0] _RAND_1;
  wire [32:0] _EVAL_2741__EVAL_2742_data;
  wire [4:0] _EVAL_2741__EVAL_2742_addr;
  wire [32:0] _EVAL_2741__EVAL_2743_data;
  wire [4:0] _EVAL_2741__EVAL_2743_addr;
  wire [32:0] _EVAL_2741__EVAL_2744_data;
  wire [4:0] _EVAL_2741__EVAL_2744_addr;
  wire [32:0] _EVAL_2741__EVAL_2745_data;
  wire [4:0] _EVAL_2741__EVAL_2745_addr;
  wire [32:0] _EVAL_2741__EVAL_2746_data;
  wire [4:0] _EVAL_2741__EVAL_2746_addr;
  wire [32:0] _EVAL_2741__EVAL_2747_data;
  wire [4:0] _EVAL_2741__EVAL_2747_addr;
  wire [32:0] _EVAL_2741__EVAL_2748_data;
  wire [4:0] _EVAL_2741__EVAL_2748_addr;
  wire [32:0] _EVAL_2741__EVAL_2749_data;
  wire [4:0] _EVAL_2741__EVAL_2749_addr;
  wire [32:0] _EVAL_2741__EVAL_2750_data;
  wire [4:0] _EVAL_2741__EVAL_2750_addr;
  wire [32:0] _EVAL_2741__EVAL_2751_data;
  wire [4:0] _EVAL_2741__EVAL_2751_addr;
  wire  _EVAL_2741__EVAL_2751_mask;
  wire  _EVAL_2741__EVAL_2751_en;
  wire [32:0] _EVAL_2741__EVAL_2752_data;
  wire [4:0] _EVAL_2741__EVAL_2752_addr;
  wire  _EVAL_2741__EVAL_2752_mask;
  wire  _EVAL_2741__EVAL_2752_en;
  reg  _EVAL_284;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_313;
  reg [31:0] _RAND_3;
  reg  _EVAL_332;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_350;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_356;
  reg [31:0] _RAND_6;
  reg  _EVAL_366;
  reg [31:0] _RAND_7;
  reg [4:0] _EVAL_375;
  reg [31:0] _RAND_8;
  reg  _EVAL_380;
  reg [31:0] _RAND_9;
  reg  _EVAL_396;
  reg [31:0] _RAND_10;
  reg [4:0] _EVAL_483;
  reg [31:0] _RAND_11;
  reg  _EVAL_490;
  reg [31:0] _RAND_12;
  reg  _EVAL_494;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_498;
  reg [31:0] _RAND_14;
  reg  _EVAL_531;
  reg [31:0] _RAND_15;
  reg  _EVAL_545;
  reg [31:0] _RAND_16;
  reg  _EVAL_601;
  reg [31:0] _RAND_17;
  reg  _EVAL_612;
  reg [31:0] _RAND_18;
  reg [4:0] _EVAL_623;
  reg [31:0] _RAND_19;
  reg  _EVAL_639;
  reg [31:0] _RAND_20;
  reg [4:0] _EVAL_649;
  reg [31:0] _RAND_21;
  reg  _EVAL_653;
  reg [31:0] _RAND_22;
  reg  _EVAL_666;
  reg [31:0] _RAND_23;
  reg  _EVAL_678;
  reg [31:0] _RAND_24;
  reg  _EVAL_690;
  reg [31:0] _RAND_25;
  reg  _EVAL_706;
  reg [31:0] _RAND_26;
  reg [2:0] _EVAL_780;
  reg [31:0] _RAND_27;
  reg  _EVAL_792;
  reg [31:0] _RAND_28;
  reg  _EVAL_811;
  reg [31:0] _RAND_29;
  reg  _EVAL_861;
  reg [31:0] _RAND_30;
  reg  _EVAL_869;
  reg [31:0] _RAND_31;
  reg  _EVAL_896;
  reg [31:0] _RAND_32;
  reg  _EVAL_899;
  reg [31:0] _RAND_33;
  reg  _EVAL_922;
  reg [31:0] _RAND_34;
  reg  _EVAL_925;
  reg [31:0] _RAND_35;
  reg  _EVAL_935;
  reg [31:0] _RAND_36;
  reg  _EVAL_937;
  reg [31:0] _RAND_37;
  reg  _EVAL_946;
  reg [31:0] _RAND_38;
  reg [31:0] _EVAL_949;
  reg [31:0] _RAND_39;
  reg  _EVAL_951;
  reg [31:0] _RAND_40;
  reg [31:0] _EVAL_952;
  reg [31:0] _RAND_41;
  reg  _EVAL_954;
  reg [31:0] _RAND_42;
  reg  _EVAL_971;
  reg [31:0] _RAND_43;
  reg  _EVAL_980;
  reg [31:0] _RAND_44;
  reg [6:0] _EVAL_983;
  reg [31:0] _RAND_45;
  reg  _EVAL_993;
  reg [31:0] _RAND_46;
  reg  _EVAL_1000;
  reg [31:0] _RAND_47;
  reg [2:0] _EVAL_1024;
  reg [31:0] _RAND_48;
  reg  _EVAL_1042;
  reg [31:0] _RAND_49;
  reg [4:0] _EVAL_1059;
  reg [31:0] _RAND_50;
  reg  _EVAL_1097;
  reg [31:0] _RAND_51;
  reg  _EVAL_1103;
  reg [31:0] _RAND_52;
  reg [31:0] _EVAL_1104;
  reg [31:0] _RAND_53;
  reg [31:0] _EVAL_1109;
  reg [31:0] _RAND_54;
  reg  _EVAL_1122;
  reg [31:0] _RAND_55;
  reg  _EVAL_1134;
  reg [31:0] _RAND_56;
  reg [4:0] _EVAL_1146;
  reg [31:0] _RAND_57;
  reg  _EVAL_1149;
  reg [31:0] _RAND_58;
  reg  _EVAL_1187;
  reg [31:0] _RAND_59;
  reg [4:0] _EVAL_1198;
  reg [31:0] _RAND_60;
  reg  _EVAL_1250;
  reg [31:0] _RAND_61;
  reg  _EVAL_1253;
  reg [31:0] _RAND_62;
  reg [31:0] _EVAL_1294;
  reg [31:0] _RAND_63;
  reg  _EVAL_1333;
  reg [31:0] _RAND_64;
  reg [4:0] _EVAL_1347;
  reg [31:0] _RAND_65;
  reg  _EVAL_1352;
  reg [31:0] _RAND_66;
  reg [4:0] _EVAL_1356;
  reg [31:0] _RAND_67;
  reg [2:0] _EVAL_1379;
  reg [31:0] _RAND_68;
  reg [4:0] _EVAL_1415;
  reg [31:0] _RAND_69;
  reg  _EVAL_1446;
  reg [31:0] _RAND_70;
  reg [6:0] _EVAL_1452;
  reg [31:0] _RAND_71;
  reg  _EVAL_1469;
  reg [31:0] _RAND_72;
  reg  _EVAL_1476;
  reg [31:0] _RAND_73;
  reg [4:0] _EVAL_1480;
  reg [31:0] _RAND_74;
  reg  _EVAL_1491;
  reg [31:0] _RAND_75;
  reg  _EVAL_1499;
  reg [31:0] _RAND_76;
  reg  _EVAL_1511;
  reg [31:0] _RAND_77;
  reg  _EVAL_1521;
  reg [31:0] _RAND_78;
  reg  _EVAL_1591;
  reg [31:0] _RAND_79;
  reg  _EVAL_1617;
  reg [31:0] _RAND_80;
  reg [4:0] _EVAL_1641;
  reg [31:0] _RAND_81;
  reg  _EVAL_1647;
  reg [31:0] _RAND_82;
  reg  _EVAL_1654;
  reg [31:0] _RAND_83;
  reg  _EVAL_1671;
  reg [31:0] _RAND_84;
  reg  _EVAL_1699;
  reg [31:0] _RAND_85;
  reg  _EVAL_1702;
  reg [31:0] _RAND_86;
  reg  _EVAL_1724;
  reg [31:0] _RAND_87;
  reg [127:0] _EVAL_1727;
  reg [127:0] _RAND_88;
  reg  _EVAL_1737;
  reg [31:0] _RAND_89;
  reg  _EVAL_1740;
  reg [31:0] _RAND_90;
  reg [4:0] _EVAL_1795;
  reg [31:0] _RAND_91;
  reg  _EVAL_1818;
  reg [31:0] _RAND_92;
  reg [4:0] _EVAL_1827;
  reg [31:0] _RAND_93;
  reg  _EVAL_1828;
  reg [31:0] _RAND_94;
  reg  _EVAL_1854;
  reg [31:0] _RAND_95;
  reg  _EVAL_1895;
  reg [31:0] _RAND_96;
  reg  _EVAL_1896;
  reg [31:0] _RAND_97;
  reg  _EVAL_1908;
  reg [31:0] _RAND_98;
  reg [32:0] _EVAL_1913;
  reg [63:0] _RAND_99;
  reg  _EVAL_1915;
  reg [31:0] _RAND_100;
  reg [31:0] _EVAL_1921;
  reg [31:0] _RAND_101;
  reg  _EVAL_1965;
  reg [31:0] _RAND_102;
  reg  _EVAL_1968;
  reg [31:0] _RAND_103;
  reg [1:0] _EVAL_1972;
  reg [31:0] _RAND_104;
  reg [6:0] _EVAL_2030;
  reg [31:0] _RAND_105;
  reg  _EVAL_2060;
  reg [31:0] _RAND_106;
  reg  _EVAL_2089;
  reg [31:0] _RAND_107;
  reg  _EVAL_2118;
  reg [31:0] _RAND_108;
  reg  _EVAL_2138;
  reg [31:0] _RAND_109;
  reg  _EVAL_2145;
  reg [31:0] _RAND_110;
  reg [1:0] _EVAL_2172;
  reg [31:0] _RAND_111;
  reg  _EVAL_2176;
  reg [31:0] _RAND_112;
  reg [4:0] _EVAL_2193;
  reg [31:0] _RAND_113;
  reg  _EVAL_2219;
  reg [31:0] _RAND_114;
  reg  _EVAL_2244;
  reg [31:0] _RAND_115;
  reg  _EVAL_2258;
  reg [31:0] _RAND_116;
  reg  _EVAL_2268;
  reg [31:0] _RAND_117;
  reg [127:0] _EVAL_2278;
  reg [127:0] _RAND_118;
  reg  _EVAL_2280;
  reg [31:0] _RAND_119;
  reg  _EVAL_2282;
  reg [31:0] _RAND_120;
  reg [4:0] _EVAL_2320;
  reg [31:0] _RAND_121;
  reg  _EVAL_2326;
  reg [31:0] _RAND_122;
  reg  _EVAL_2329;
  reg [31:0] _RAND_123;
  reg [31:0] _EVAL_2331;
  reg [31:0] _RAND_124;
  reg  _EVAL_2369;
  reg [31:0] _RAND_125;
  reg  _EVAL_2371;
  reg [31:0] _RAND_126;
  reg [31:0] _EVAL_2383;
  reg [31:0] _RAND_127;
  reg [31:0] _EVAL_2397;
  reg [31:0] _RAND_128;
  reg  _EVAL_2399;
  reg [31:0] _RAND_129;
  reg  _EVAL_2409;
  reg [31:0] _RAND_130;
  reg [31:0] _EVAL_2423;
  reg [31:0] _RAND_131;
  reg  _EVAL_2424;
  reg [31:0] _RAND_132;
  reg  _EVAL_2443;
  reg [31:0] _RAND_133;
  reg [4:0] _EVAL_2495;
  reg [31:0] _RAND_134;
  reg  _EVAL_2499;
  reg [31:0] _RAND_135;
  reg  _EVAL_2506;
  reg [31:0] _RAND_136;
  reg  _EVAL_2542;
  reg [31:0] _RAND_137;
  reg  _EVAL_2573;
  reg [31:0] _RAND_138;
  reg [4:0] _EVAL_2579;
  reg [31:0] _RAND_139;
  reg  _EVAL_2583;
  reg [31:0] _RAND_140;
  reg [1:0] _EVAL_2587;
  reg [31:0] _RAND_141;
  reg  _EVAL_2596;
  reg [31:0] _RAND_142;
  reg  _EVAL_2603;
  reg [31:0] _RAND_143;
  reg  _EVAL_2624;
  reg [31:0] _RAND_144;
  reg  _EVAL_2644;
  reg [31:0] _RAND_145;
  reg [31:0] _EVAL_2656;
  reg [31:0] _RAND_146;
  reg  _EVAL_2667;
  reg [31:0] _RAND_147;
  reg [4:0] _EVAL_2683;
  reg [31:0] _RAND_148;
  reg  _EVAL_2686;
  reg [31:0] _RAND_149;
  reg  _EVAL_2753;
  reg [31:0] _RAND_150;
  reg [31:0] _EVAL_2758;
  reg [31:0] _RAND_151;
  reg  _EVAL_2765;
  reg [31:0] _RAND_152;
  reg  _EVAL_2794;
  reg [31:0] _RAND_153;
  reg [5:0] _EVAL_2823;
  reg [31:0] _RAND_154;
  reg  _EVAL_2843;
  reg [31:0] _RAND_155;
  reg  _EVAL_2853;
  reg [31:0] _RAND_156;
  reg [31:0] _EVAL_2880;
  reg [31:0] _RAND_157;
  reg  _EVAL_2886;
  reg [31:0] _RAND_158;
  reg  _EVAL_2911;
  reg [31:0] _RAND_159;
  reg [31:0] _EVAL_2912;
  reg [31:0] _RAND_160;
  reg [31:0] _EVAL_2919;
  reg [31:0] _RAND_161;
  reg  _EVAL_2948;
  reg [31:0] _RAND_162;
  reg  _EVAL_2955;
  reg [31:0] _RAND_163;
  reg  _EVAL_2969;
  reg [31:0] _RAND_164;
  reg  _EVAL_2989;
  reg [31:0] _RAND_165;
  reg  _EVAL_3000;
  reg [31:0] _RAND_166;
  reg [127:0] _EVAL_3019;
  reg [127:0] _RAND_167;
  reg [31:0] _EVAL_3025;
  reg [31:0] _RAND_168;
  reg  _EVAL_3029;
  reg [31:0] _RAND_169;
  reg [4:0] _EVAL_3039;
  reg [31:0] _RAND_170;
  reg [4:0] _EVAL_3053;
  reg [31:0] _RAND_171;
  reg [2:0] _EVAL_3064;
  reg [31:0] _RAND_172;
  reg [1:0] _EVAL_3077;
  reg [31:0] _RAND_173;
  reg  _EVAL_3085;
  reg [31:0] _RAND_174;
  reg  _EVAL_3094;
  reg [31:0] _RAND_175;
  reg  _EVAL_3102;
  reg [31:0] _RAND_176;
  reg [4:0] _EVAL_3117;
  reg [31:0] _RAND_177;
  reg [31:0] _EVAL_3132;
  reg [31:0] _RAND_178;
  reg [4:0] _EVAL_3134;
  reg [31:0] _RAND_179;
  reg [31:0] _EVAL_3142;
  reg [31:0] _RAND_180;
  reg  _EVAL_3165;
  reg [31:0] _RAND_181;
  reg  _EVAL_3170;
  reg [31:0] _RAND_182;
  reg  _EVAL_3176;
  reg [31:0] _RAND_183;
  reg [2:0] _EVAL_3178;
  reg [31:0] _RAND_184;
  reg [31:0] _EVAL_3196;
  reg [31:0] _RAND_185;
  reg  _EVAL_3204;
  reg [31:0] _RAND_186;
  reg  _EVAL_3217;
  reg [31:0] _RAND_187;
  reg  _EVAL_3227;
  reg [31:0] _RAND_188;
  reg [6:0] _EVAL_3229;
  reg [31:0] _RAND_189;
  reg  _EVAL_3240;
  reg [31:0] _RAND_190;
  reg [2:0] _EVAL_3270;
  reg [31:0] _RAND_191;
  reg  _EVAL_3276;
  reg [31:0] _RAND_192;
  reg [2:0] _EVAL_3291;
  reg [31:0] _RAND_193;
  reg  _EVAL_3295;
  reg [31:0] _RAND_194;
  reg [2:0] _EVAL_3302;
  reg [31:0] _RAND_195;
  reg [4:0] _EVAL_3309;
  reg [31:0] _RAND_196;
  reg  _EVAL_3355;
  reg [31:0] _RAND_197;
  reg  _EVAL_3362;
  reg [31:0] _RAND_198;
  reg [4:0] _EVAL_3366;
  reg [31:0] _RAND_199;
  reg [4:0] _EVAL_3370;
  reg [31:0] _RAND_200;
  reg [127:0] _EVAL_3384;
  reg [127:0] _RAND_201;
  reg [14:0] _EVAL_3386;
  reg [31:0] _RAND_202;
  reg  _EVAL_3391;
  reg [31:0] _RAND_203;
  reg  _EVAL_3393;
  reg [31:0] _RAND_204;
  reg  _EVAL_3401;
  reg [31:0] _RAND_205;
  reg  _EVAL_3404;
  reg [31:0] _RAND_206;
  reg [31:0] _EVAL_3405;
  reg [31:0] _RAND_207;
  reg  _EVAL_3413;
  reg [31:0] _RAND_208;
  reg  _EVAL_3415;
  reg [31:0] _RAND_209;
  reg  _EVAL_3421;
  reg [31:0] _RAND_210;
  reg [31:0] _EVAL_3432;
  reg [31:0] _RAND_211;
  reg  _EVAL_3448;
  reg [31:0] _RAND_212;
  reg  _EVAL_3476;
  reg [31:0] _RAND_213;
  reg  _EVAL_3481;
  reg [31:0] _RAND_214;
  reg [31:0] _EVAL_3494;
  reg [31:0] _RAND_215;
  reg  _EVAL_3523;
  reg [31:0] _RAND_216;
  reg [4:0] _EVAL_3573;
  reg [31:0] _RAND_217;
  reg  _EVAL_3588;
  reg [31:0] _RAND_218;
  reg  _EVAL_3608;
  reg [31:0] _RAND_219;
  reg  _EVAL_3624;
  reg [31:0] _RAND_220;
  reg  _EVAL_3629;
  reg [31:0] _RAND_221;
  reg  _EVAL_3637;
  reg [31:0] _RAND_222;
  reg [14:0] _EVAL_3645;
  reg [31:0] _RAND_223;
  reg [4:0] _EVAL_3670;
  reg [31:0] _RAND_224;
  reg  _EVAL_3694;
  reg [31:0] _RAND_225;
  reg [4:0] _EVAL_3711;
  reg [31:0] _RAND_226;
  reg  _EVAL_3712;
  reg [31:0] _RAND_227;
  reg [31:0] _EVAL_3727;
  reg [31:0] _RAND_228;
  reg [31:0] _EVAL_3728;
  reg [31:0] _RAND_229;
  reg  _EVAL_3730;
  reg [31:0] _RAND_230;
  reg [4:0] _EVAL_3742;
  reg [31:0] _RAND_231;
  reg  _EVAL_3747;
  reg [31:0] _RAND_232;
  reg  _EVAL_3750;
  reg [31:0] _RAND_233;
  reg [2:0] _EVAL_3752;
  reg [31:0] _RAND_234;
  reg  _EVAL_3771;
  reg [31:0] _RAND_235;
  reg  _EVAL_3798;
  reg [31:0] _RAND_236;
  reg  _EVAL_3814;
  reg [31:0] _RAND_237;
  reg  _EVAL_3840;
  reg [31:0] _RAND_238;
  reg [4:0] _EVAL_3841;
  reg [31:0] _RAND_239;
  reg [31:0] _EVAL_3845;
  reg [31:0] _RAND_240;
  reg [4:0] _EVAL_3851;
  reg [31:0] _RAND_241;
  reg  _EVAL_3858;
  reg [31:0] _RAND_242;
  reg [31:0] _EVAL_3880;
  reg [31:0] _RAND_243;
  reg  _EVAL_3888;
  reg [31:0] _RAND_244;
  reg  _EVAL_3902;
  reg [31:0] _RAND_245;
  reg [2:0] _EVAL_3922;
  reg [31:0] _RAND_246;
  reg  _EVAL_3934;
  reg [31:0] _RAND_247;
  reg  _EVAL_3939;
  reg [31:0] _RAND_248;
  reg [31:0] _EVAL_3940;
  reg [31:0] _RAND_249;
  reg [2:0] _EVAL_3974;
  reg [31:0] _RAND_250;
  reg  _EVAL_3986;
  reg [31:0] _RAND_251;
  reg  _EVAL_3997;
  reg [31:0] _RAND_252;
  reg  _EVAL_4000;
  reg [31:0] _RAND_253;
  reg  _EVAL_4014;
  reg [31:0] _RAND_254;
  reg [6:0] _EVAL_4019;
  reg [31:0] _RAND_255;
  reg  _EVAL_4043;
  reg [31:0] _RAND_256;
  reg [2:0] _EVAL_4064;
  reg [31:0] _RAND_257;
  reg [1:0] _EVAL_4088;
  reg [31:0] _RAND_258;
  reg  _EVAL_4092;
  reg [31:0] _RAND_259;
  reg  _EVAL_4095;
  reg [31:0] _RAND_260;
  reg  _EVAL_4115;
  reg [31:0] _RAND_261;
  reg [4:0] _EVAL_4135;
  reg [31:0] _RAND_262;
  reg [127:0] _EVAL_4154;
  reg [127:0] _RAND_263;
  reg [31:0] _EVAL_4157;
  reg [31:0] _RAND_264;
  reg [63:0] _EVAL_4160;
  reg [63:0] _RAND_265;
  reg [2:0] _EVAL_4162;
  reg [31:0] _RAND_266;
  reg  _EVAL_4167;
  reg [31:0] _RAND_267;
  reg  _EVAL_4168;
  reg [31:0] _RAND_268;
  reg [6:0] _EVAL_4192;
  reg [31:0] _RAND_269;
  reg [31:0] _EVAL_4195;
  reg [31:0] _RAND_270;
  reg [2:0] _EVAL_4201;
  reg [31:0] _RAND_271;
  reg  _EVAL_4203;
  reg [31:0] _RAND_272;
  reg [11:0] _EVAL_4218;
  reg [31:0] _RAND_273;
  reg  _EVAL_4240;
  reg [31:0] _RAND_274;
  reg  _EVAL_4299;
  reg [31:0] _RAND_275;
  reg [31:0] _EVAL_4319;
  reg [31:0] _RAND_276;
  reg [31:0] _EVAL_4322;
  reg [31:0] _RAND_277;
  reg  _EVAL_4360;
  reg [31:0] _RAND_278;
  reg  _EVAL_4362;
  reg [31:0] _RAND_279;
  reg [31:0] _EVAL_4373;
  reg [31:0] _RAND_280;
  reg [4:0] _EVAL_4400;
  reg [31:0] _RAND_281;
  reg  _EVAL_4423;
  reg [31:0] _RAND_282;
  reg  _EVAL_4437;
  reg [31:0] _RAND_283;
  reg [4:0] _EVAL_4460;
  reg [31:0] _RAND_284;
  reg [31:0] _EVAL_4461;
  reg [31:0] _RAND_285;
  reg [31:0] _EVAL_4468;
  reg [31:0] _RAND_286;
  reg [127:0] _EVAL_4481;
  reg [127:0] _RAND_287;
  reg  _EVAL_4512;
  reg [31:0] _RAND_288;
  reg [4:0] _EVAL_4530;
  reg [31:0] _RAND_289;
  reg  _EVAL_4531;
  reg [31:0] _RAND_290;
  reg  _EVAL_4535;
  reg [31:0] _RAND_291;
  reg [2:0] _EVAL_4539;
  reg [31:0] _RAND_292;
  reg [127:0] _EVAL_4550;
  reg [127:0] _RAND_293;
  reg  _EVAL_4562;
  reg [31:0] _RAND_294;
  reg  _EVAL_4596;
  reg [31:0] _RAND_295;
  reg [31:0] _EVAL_4600;
  reg [31:0] _RAND_296;
  reg [2:0] _EVAL_4607;
  reg [31:0] _RAND_297;
  reg [4:0] _EVAL_4614;
  reg [31:0] _RAND_298;
  reg  _EVAL_4620;
  reg [31:0] _RAND_299;
  reg  _EVAL_4632;
  reg [31:0] _RAND_300;
  reg [4:0] _EVAL_4633;
  reg [31:0] _RAND_301;
  reg  _EVAL_4649;
  reg [31:0] _RAND_302;
  reg [31:0] _EVAL_4656;
  reg [31:0] _RAND_303;
  reg [31:0] _EVAL_4679;
  reg [31:0] _RAND_304;
  reg  _EVAL_4684;
  reg [31:0] _RAND_305;
  reg  _EVAL_4692;
  reg [31:0] _RAND_306;
  reg  _EVAL_4698;
  reg [31:0] _RAND_307;
  reg [4:0] _EVAL_4706;
  reg [31:0] _RAND_308;
  reg [4:0] _EVAL_4715;
  reg [31:0] _RAND_309;
  reg  _EVAL_4736;
  reg [31:0] _RAND_310;
  reg [4:0] _EVAL_4745;
  reg [31:0] _RAND_311;
  reg [31:0] _EVAL_4748;
  reg [31:0] _RAND_312;
  reg  _EVAL_4790;
  reg [31:0] _RAND_313;
  reg  _EVAL_4796;
  reg [31:0] _RAND_314;
  reg  _EVAL_4805;
  reg [31:0] _RAND_315;
  reg  _EVAL_4812;
  reg [31:0] _RAND_316;
  reg  _EVAL_4819;
  reg [31:0] _RAND_317;
  reg  _EVAL_4842;
  reg [31:0] _RAND_318;
  reg  _EVAL_4844;
  reg [31:0] _RAND_319;
  reg [31:0] _EVAL_4863;
  reg [31:0] _RAND_320;
  reg [127:0] _EVAL_4915;
  reg [127:0] _RAND_321;
  reg [2:0] _EVAL_4927;
  reg [31:0] _RAND_322;
  reg  _EVAL_4936;
  reg [31:0] _RAND_323;
  reg [4:0] _EVAL_4939;
  reg [31:0] _RAND_324;
  reg  _EVAL_4947;
  reg [31:0] _RAND_325;
  reg  _EVAL_4962;
  reg [31:0] _RAND_326;
  reg [2:0] _EVAL_4968;
  reg [31:0] _RAND_327;
  reg [31:0] _EVAL_5009;
  reg [31:0] _RAND_328;
  reg  _EVAL_5017;
  reg [31:0] _RAND_329;
  reg  _EVAL_5025;
  reg [31:0] _RAND_330;
  reg  _EVAL_5039;
  reg [31:0] _RAND_331;
  reg [31:0] _EVAL_5043;
  reg [31:0] _RAND_332;
  reg  _EVAL_5052;
  reg [31:0] _RAND_333;
  reg  _EVAL_5095;
  reg [31:0] _RAND_334;
  reg [4:0] _EVAL_5099;
  reg [31:0] _RAND_335;
  reg  _EVAL_5178;
  reg [31:0] _RAND_336;
  reg [14:0] _EVAL_5213;
  reg [31:0] _RAND_337;
  reg  _EVAL_5226;
  reg [31:0] _RAND_338;
  reg  _EVAL_5233;
  reg [31:0] _RAND_339;
  reg  _EVAL_5237;
  reg [31:0] _RAND_340;
  reg [2:0] _EVAL_5265;
  reg [31:0] _RAND_341;
  reg  _EVAL_5335;
  reg [31:0] _RAND_342;
  reg  _EVAL_5344;
  reg [31:0] _RAND_343;
  reg [4:0] _EVAL_5363;
  reg [31:0] _RAND_344;
  reg [31:0] _EVAL_5367;
  reg [31:0] _RAND_345;
  reg [31:0] _EVAL_5412;
  reg [31:0] _RAND_346;
  wire  _EVAL_1844;
  wire  _EVAL_5290;
  wire  _EVAL_4710;
  wire  _EVAL_2703;
  wire  _EVAL_1575;
  wire  _EVAL_4848;
  wire  _EVAL_3081;
  wire  _EVAL_315;
  wire [6:0] _EVAL_2400;
  wire  _EVAL_1762;
  wire [1:0] _EVAL_1335;
  wire  _EVAL_4196;
  wire  _EVAL_2393;
  wire [23:0] _EVAL_3538;
  wire  _EVAL_3681;
  wire  _EVAL_1778;
  wire  _EVAL_4721;
  wire  _EVAL_1969;
  wire  _EVAL_3066;
  wire  _EVAL_3904;
  wire  _EVAL_890;
  wire  _EVAL_2868;
  wire  _EVAL_3519;
  wire [1:0] _EVAL_2523;
  wire [1:0] _EVAL_5069;
  wire  _EVAL_1623;
  wire  _EVAL_351;
  wire [4:0] _EVAL_1722;
  wire  _EVAL_1616;
  wire  _EVAL_361;
  wire  _EVAL_1387;
  wire  _EVAL_3820;
  wire  _EVAL_2876;
  wire [4:0] _EVAL_4127;
  wire  _EVAL_2956;
  wire  _EVAL_1608;
  wire  _EVAL_588;
  wire  _EVAL_4623;
  wire  _EVAL_2595;
  wire  _EVAL_3168;
  wire  _EVAL_2133;
  wire  _EVAL_1299;
  wire  _EVAL_1655;
  wire [4:0] _EVAL_3212;
  wire  _EVAL_2594;
  wire  _EVAL_2313;
  wire  _EVAL_1372;
  wire  _EVAL_2025;
  wire  _EVAL_783;
  wire  _EVAL_3808;
  wire  _EVAL_4357;
  wire  _EVAL_3671;
  wire  _EVAL_3116;
  wire  _EVAL_3082;
  wire  _EVAL_631;
  wire  _EVAL_1434;
  wire  _EVAL_3141;
  wire  _EVAL_2321;
  wire  _EVAL_747;
  wire  _EVAL_2394;
  wire  _EVAL_5360;
  wire  _EVAL_4683;
  wire  _EVAL_1255;
  wire  _EVAL_739;
  wire  _EVAL_3346;
  wire  _EVAL_3763;
  wire  _EVAL_2532;
  wire  _EVAL_3962;
  wire  _EVAL_1414;
  wire  _EVAL_1546;
  wire  _EVAL_4528;
  wire  _EVAL_500;
  wire  _EVAL_1570;
  wire  _EVAL_4348;
  wire  _EVAL_2653;
  wire  _EVAL_1158;
  wire  _EVAL_1507;
  wire  _EVAL_2108;
  wire  _EVAL_546;
  wire  _EVAL_408;
  wire  _EVAL_4067;
  wire  _EVAL_584;
  wire  _EVAL_1311;
  wire  _EVAL_1319;
  wire  _EVAL_1952;
  wire  _EVAL_3850;
  wire  _EVAL_4696;
  wire  _EVAL_4197;
  wire  _EVAL_591;
  wire  _EVAL_4963;
  wire  _EVAL_4490;
  wire  _EVAL_821;
  wire  _EVAL_3864;
  wire  _EVAL_4771;
  wire  _EVAL_4260;
  wire  _EVAL_903;
  wire  _EVAL_862;
  wire [11:0] _EVAL_1445;
  wire [1:0] _EVAL_3957;
  wire  _EVAL_1694;
  wire  _EVAL_5111;
  wire  _EVAL_3755;
  wire  _EVAL_1120;
  wire [11:0] _EVAL_5246;
  wire [2:0] _EVAL_2208;
  wire [2:0] _EVAL_4494;
  wire [1:0] _EVAL_4757;
  wire [2:0] _EVAL_5219;
  wire [15:0] _EVAL_818;
  wire  _EVAL_4395;
  wire [1:0] _EVAL_1958;
  wire [2:0] _EVAL_927;
  wire [15:0] _EVAL_1954;
  wire [15:0] _EVAL_1113;
  wire  _EVAL_556;
  wire  _EVAL_3661;
  wire [15:0] _EVAL_2429;
  wire [2:0] _EVAL_2874;
  wire [15:0] _EVAL_3017;
  wire [15:0] _EVAL_2260;
  wire [15:0] _EVAL_5236;
  wire [2:0] _EVAL_3373;
  wire  _EVAL_2034;
  wire [8:0] _EVAL_3232;
  wire [9:0] _EVAL_618;
  wire [7:0] _EVAL_3796;
  wire  _EVAL_3409;
  wire  _EVAL_4001;
  wire  _EVAL_4724;
  wire  _EVAL_1271;
  wire [5:0] _EVAL_1306;
  wire [63:0] _EVAL_2332;
  wire  _EVAL_2488;
  wire  _EVAL_4996;
  wire  _EVAL_813;
  wire  _EVAL_1677;
  wire  _EVAL_3912;
  wire  _EVAL_1477;
  wire  _EVAL_1535;
  wire  _EVAL_2564;
  wire  _EVAL_2509;
  wire  _EVAL_5391;
  wire [5:0] _EVAL_2617;
  wire  _EVAL_1573;
  wire  _EVAL_2120;
  wire  _EVAL_1966;
  wire  _EVAL_296;
  wire  _EVAL_2257;
  wire  _EVAL_423;
  wire  _EVAL_1190;
  wire [5:0] _EVAL_4158;
  wire  _EVAL_2452;
  wire  _EVAL_2942;
  wire  _EVAL_2481;
  wire  _EVAL_1242;
  wire  _EVAL_2524;
  wire [5:0] _EVAL_2316;
  wire [63:0] _EVAL_2301;
  wire  _EVAL_5337;
  wire  _EVAL_3422;
  wire  _EVAL_902;
  wire  _EVAL_1927;
  wire  _EVAL_4388;
  wire  _EVAL_2049;
  wire  _EVAL_3419;
  wire  _EVAL_2549;
  wire  _EVAL_4564;
  wire  _EVAL_3956;
  wire  _EVAL_512;
  wire  _EVAL_2600;
  wire  _EVAL_3679;
  wire [5:0] _EVAL_2954;
  wire [63:0] _EVAL_3509;
  wire  _EVAL_2080;
  wire  _EVAL_1685;
  wire  _EVAL_1167;
  wire  _EVAL_5126;
  wire  _EVAL_4986;
  wire  _EVAL_614;
  wire  _EVAL_2916;
  wire  _EVAL_1670;
  wire  _EVAL_1320;
  wire  _EVAL_4760;
  wire  _EVAL_2638;
  wire  _EVAL_308;
  wire [5:0] _EVAL_2897;
  wire [63:0] _EVAL_1322;
  wire  _EVAL_4769;
  wire  _EVAL_1676;
  wire  _EVAL_1218;
  wire  _EVAL_3492;
  wire  _EVAL_1293;
  wire  _EVAL_1855;
  wire  _EVAL_386;
  wire  _EVAL_2901;
  wire  _EVAL_3027;
  wire  _EVAL_4302;
  wire  _EVAL_3374;
  wire  _EVAL_3256;
  wire  _EVAL_2216;
  wire  _EVAL_2705;
  wire  _EVAL_3231;
  wire  _EVAL_3758;
  wire  _EVAL_4222;
  wire  _EVAL_589;
  wire  _EVAL_2668;
  wire  _EVAL_1241;
  wire [9:0] _EVAL_4033;
  wire  _EVAL_775;
  wire [1:0] _EVAL_524;
  wire  _EVAL_5194;
  wire  _EVAL_4278;
  wire  _EVAL_2243;
  wire  _EVAL_4516;
  wire [2:0] _EVAL_2607;
  wire [20:0] _EVAL_2778;
  wire  _EVAL_2978;
  wire [9:0] _EVAL_1285;
  wire  _EVAL_4259;
  wire [7:0] _EVAL_2173;
  wire [31:0] _EVAL_1628;
  wire  _EVAL_4809;
  wire  _EVAL_3012;
  wire  _EVAL_2359;
  wire  _EVAL_2448;
  wire [11:0] _EVAL_1542;
  wire [2:0] _EVAL_3872;
  wire [2:0] _EVAL_4488;
  wire [1:0] _EVAL_3551;
  wire [2:0] _EVAL_2846;
  wire [15:0] _EVAL_3470;
  wire [2:0] _EVAL_857;
  wire [15:0] _EVAL_4020;
  wire [15:0] _EVAL_3599;
  wire  _EVAL_3126;
  wire  _EVAL_2483;
  wire [15:0] _EVAL_4153;
  wire [3:0] _EVAL_2775;
  wire [15:0] _EVAL_3552;
  wire [15:0] _EVAL_2774;
  wire [15:0] _EVAL_1704;
  wire  _EVAL_850;
  wire  _EVAL_5185;
  wire [15:0] _EVAL_4051;
  wire [15:0] _EVAL_3344;
  wire [15:0] _EVAL_1706;
  wire [15:0] _EVAL_1481;
  wire [15:0] _EVAL_4520;
  wire [15:0] _EVAL_3555;
  wire [15:0] _EVAL_4447;
  wire [15:0] _EVAL_3913;
  wire [15:0] _EVAL_771;
  wire  _EVAL_4093;
  wire  _EVAL_1901;
  wire [19:0] _EVAL_3133;
  wire [19:0] _EVAL_2904;
  wire  _EVAL_2801;
  wire [4:0] _EVAL_1067;
  wire [15:0] _EVAL_2150;
  wire  _EVAL_762;
  wire [11:0] _EVAL_735;
  wire  _EVAL_2512;
  wire [4:0] _EVAL_2998;
  wire [15:0] _EVAL_3862;
  wire [15:0] _EVAL_302;
  wire  _EVAL_3360;
  wire  _EVAL_323;
  wire [15:0] _EVAL_1837;
  wire [15:0] _EVAL_5240;
  wire [15:0] _EVAL_4180;
  wire [15:0] _EVAL_1235;
  wire [15:0] _EVAL_4473;
  wire  _EVAL_3674;
  wire  _EVAL_3347;
  wire  _EVAL_4538;
  wire  _EVAL_4728;
  wire [1:0] _EVAL_5190;
  wire [15:0] _EVAL_3596;
  wire [15:0] _EVAL_507;
  wire [15:0] _EVAL_2898;
  wire  _EVAL_1227;
  wire  _EVAL_4271;
  wire  _EVAL_2673;
  wire [1:0] _EVAL_2128;
  wire [3:0] _EVAL_3490;
  wire  _EVAL_1618;
  wire  _EVAL_4886;
  wire [2:0] _EVAL_809;
  wire [15:0] _EVAL_5250;
  wire [15:0] _EVAL_2609;
  wire [15:0] _EVAL_4122;
  wire [15:0] _EVAL_1473;
  wire [15:0] _EVAL_338;
  wire  _EVAL_3714;
  wire  _EVAL_2090;
  wire  _EVAL_5353;
  wire [2:0] _EVAL_3566;
  wire [1:0] _EVAL_2696;
  wire [15:0] _EVAL_4798;
  wire [1:0] _EVAL_575;
  wire [2:0] _EVAL_2934;
  wire [15:0] _EVAL_3163;
  wire [15:0] _EVAL_4101;
  wire [15:0] _EVAL_1645;
  wire [2:0] _EVAL_4186;
  wire [15:0] _EVAL_909;
  wire [15:0] _EVAL_901;
  wire [15:0] _EVAL_4303;
  wire  _EVAL_2349;
  wire [15:0] _EVAL_1559;
  wire [15:0] _EVAL_452;
  wire [15:0] _EVAL_3530;
  wire [15:0] _EVAL_5225;
  wire [15:0] _EVAL_2910;
  wire [15:0] _EVAL_4374;
  wire [15:0] _EVAL_837;
  wire  _EVAL_2008;
  wire [15:0] _EVAL_4307;
  wire [15:0] _EVAL_421;
  wire [15:0] _EVAL_1540;
  wire [15:0] _EVAL_4257;
  wire [15:0] _EVAL_876;
  wire [15:0] _EVAL_2401;
  wire [15:0] _EVAL_1916;
  wire [15:0] _EVAL_4622;
  wire [15:0] _EVAL_3909;
  wire [15:0] _EVAL_1621;
  wire  _EVAL_4672;
  wire  _EVAL_4818;
  wire  _EVAL_798;
  wire [32:0] _EVAL_1036;
  wire [15:0] _EVAL_1929;
  wire [31:0] _EVAL_2783;
  wire [15:0] _EVAL_3710;
  wire [31:0] _EVAL_5024;
  wire [31:0] _EVAL_4941;
  wire [31:0] _EVAL_3898;
  wire [23:0] _EVAL_3631;
  wire [31:0] _EVAL_3245;
  wire [31:0] _EVAL_4778;
  wire [23:0] _EVAL_336;
  wire [31:0] _EVAL_5332;
  wire [31:0] _EVAL_1625;
  wire [31:0] _EVAL_5106;
  wire [27:0] _EVAL_1132;
  wire [31:0] _EVAL_1133;
  wire [31:0] _EVAL_3317;
  wire [27:0] _EVAL_1658;
  wire [31:0] _EVAL_1912;
  wire [31:0] _EVAL_4335;
  wire [31:0] _EVAL_742;
  wire [29:0] _EVAL_574;
  wire [31:0] _EVAL_533;
  wire [31:0] _EVAL_5218;
  wire [29:0] _EVAL_4318;
  wire [31:0] _EVAL_988;
  wire [31:0] _EVAL_764;
  wire [31:0] _EVAL_3666;
  wire [30:0] _EVAL_704;
  wire [31:0] _EVAL_3881;
  wire [31:0] _EVAL_4973;
  wire [30:0] _EVAL_5305;
  wire [31:0] _EVAL_5284;
  wire [31:0] _EVAL_3980;
  wire [31:0] _EVAL_1478;
  wire [32:0] _EVAL_2935;
  wire [32:0] _EVAL_1307;
  wire  _EVAL_2491;
  wire  _EVAL_3148;
  wire [5:0] _EVAL_4594;
  wire [3:0] _EVAL_3209;
  wire [12:0] _EVAL_4828;
  wire [12:0] _EVAL_3159;
  wire [12:0] _EVAL_1303;
  wire  _EVAL_5370;
  wire [18:0] _EVAL_3852;
  wire [31:0] _EVAL_3471;
  wire [31:0] _EVAL_3463;
  wire [19:0] _EVAL_5389;
  wire [19:0] _EVAL_4334;
  wire  _EVAL_3776;
  wire [7:0] _EVAL_871;
  wire  _EVAL_2127;
  wire [9:0] _EVAL_2295;
  wire [20:0] _EVAL_2044;
  wire [20:0] _EVAL_4431;
  wire [20:0] _EVAL_1194;
  wire  _EVAL_2099;
  wire [10:0] _EVAL_724;
  wire [31:0] _EVAL_4791;
  wire [31:0] _EVAL_2629;
  wire [31:0] _EVAL_1298;
  wire [19:0] _EVAL_2826;
  wire [31:0] _EVAL_3577;
  wire [31:0] _EVAL_547;
  wire [31:0] _EVAL_3676;
  wire [11:0] _EVAL_3086;
  wire [11:0] _EVAL_5083;
  wire [11:0] _EVAL_677;
  wire  _EVAL_2431;
  wire [19:0] _EVAL_1723;
  wire [31:0] _EVAL_3162;
  wire [31:0] _EVAL_5148;
  wire [31:0] _EVAL_2101;
  wire [31:0] _EVAL_2389;
  wire [31:0] _EVAL_3068;
  wire [26:0] _EVAL_611;
  wire [31:0] _EVAL_3166;
  wire [4:0] _EVAL_1728;
  wire [32:0] _EVAL_1064;
  wire [31:0] _EVAL_4879;
  wire [15:0] _EVAL_870;
  wire [31:0] _EVAL_3696;
  wire [15:0] _EVAL_5144;
  wire [31:0] _EVAL_5003;
  wire [31:0] _EVAL_4206;
  wire [31:0] _EVAL_3389;
  wire [23:0] _EVAL_4663;
  wire [31:0] _EVAL_1919;
  wire [31:0] _EVAL_3308;
  wire [23:0] _EVAL_5266;
  wire [31:0] _EVAL_1336;
  wire [31:0] _EVAL_2944;
  wire [31:0] _EVAL_1717;
  wire [27:0] _EVAL_685;
  wire [31:0] _EVAL_560;
  wire [31:0] _EVAL_3591;
  wire [27:0] _EVAL_2626;
  wire [31:0] _EVAL_474;
  wire [31:0] _EVAL_3954;
  wire [31:0] _EVAL_4182;
  wire [29:0] _EVAL_551;
  wire [31:0] _EVAL_5013;
  wire [31:0] _EVAL_3293;
  wire  _EVAL_3243;
  wire  _EVAL_1323;
  wire [2:0] _EVAL_5115;
  wire  _EVAL_2565;
  wire [6:0] _EVAL_1143;
  wire [1:0] _EVAL_1509;
  wire [2:0] _EVAL_4942;
  wire [2:0] _EVAL_3048;
  wire [4:0] _EVAL_4841;
  wire [26:0] _EVAL_1412;
  wire  _EVAL_1631;
  wire [26:0] _EVAL_2447;
  wire [1:0] _EVAL_5401;
  wire [7:0] _EVAL_1367;
  wire [2:0] _EVAL_369;
  wire [4:0] _EVAL_2625;
  wire [27:0] _EVAL_2802;
  wire  _EVAL_2350;
  wire [26:0] _EVAL_2985;
  wire  _EVAL_1023;
  wire [26:0] _EVAL_1474;
  wire  _EVAL_5398;
  wire [26:0] _EVAL_1890;
  wire  _EVAL_2854;
  wire [27:0] _EVAL_4965;
  wire [3:0] _EVAL_5292;
  wire [1:0] _EVAL_738;
  wire [29:0] _EVAL_1528;
  wire [29:0] _EVAL_3228;
  wire [29:0] _EVAL_895;
  wire [29:0] _EVAL_3394;
  wire [29:0] _EVAL_5293;
  wire [29:0] _EVAL_4697;
  wire [29:0] _EVAL_4398;
  wire [29:0] _EVAL_3828;
  wire [31:0] _EVAL_4329;
  wire [31:0] _EVAL_841;
  wire  _EVAL_5130;
  wire  _EVAL_2460;
  wire [1:0] _EVAL_4593;
  wire [1:0] _EVAL_2015;
  wire  _EVAL_3205;
  wire [15:0] _EVAL_2376;
  wire [13:0] _EVAL_2137;
  wire [15:0] _EVAL_4998;
  wire [15:0] _EVAL_1571;
  wire  _EVAL_309;
  wire [15:0] _EVAL_2158;
  wire  _EVAL_2407;
  wire [12:0] _EVAL_1280;
  wire [15:0] _EVAL_1203;
  wire [15:0] _EVAL_2252;
  wire  _EVAL_1604;
  wire  _EVAL_1066;
  wire [15:0] _EVAL_866;
  wire [15:0] _EVAL_3402;
  wire [15:0] _EVAL_3557;
  wire [15:0] _EVAL_1407;
  wire  _EVAL_298;
  wire  _EVAL_2781;
  wire  _EVAL_4245;
  wire  _EVAL_4228;
  wire [19:0] _EVAL_5072;
  wire [19:0] _EVAL_409;
  wire  _EVAL_4086;
  wire  _EVAL_4877;
  wire [1:0] _EVAL_1136;
  wire  _EVAL_2143;
  wire  _EVAL_1761;
  wire  _EVAL_1369;
  wire [2:0] _EVAL_5061;
  wire  _EVAL_3192;
  wire [15:0] _EVAL_4660;
  wire [15:0] _EVAL_4933;
  wire [15:0] _EVAL_828;
  wire [15:0] _EVAL_2721;
  wire [15:0] _EVAL_1703;
  wire  _EVAL_3707;
  wire  _EVAL_1881;
  wire  _EVAL_3233;
  wire  _EVAL_1318;
  wire [4:0] _EVAL_3849;
  wire [15:0] _EVAL_960;
  wire  _EVAL_1825;
  wire  _EVAL_2669;
  wire  _EVAL_4779;
  wire  _EVAL_1290;
  wire  _EVAL_2126;
  wire  _EVAL_4954;
  wire  _EVAL_830;
  wire [2:0] _EVAL_3167;
  wire [15:0] _EVAL_2075;
  wire  _EVAL_2552;
  wire  _EVAL_281;
  wire  _EVAL_3788;
  wire  _EVAL_2602;
  wire  _EVAL_4814;
  wire  _EVAL_3147;
  wire  _EVAL_1188;
  wire [15:0] _EVAL_1842;
  wire [15:0] _EVAL_3656;
  wire [15:0] _EVAL_3684;
  wire [15:0] _EVAL_2732;
  wire [15:0] _EVAL_3507;
  wire  _EVAL_2070;
  wire [2:0] _EVAL_3173;
  wire [15:0] _EVAL_1859;
  wire [2:0] _EVAL_5021;
  wire [15:0] _EVAL_3248;
  wire [15:0] _EVAL_3797;
  wire  _EVAL_522;
  wire  _EVAL_4040;
  wire [15:0] _EVAL_1308;
  wire [3:0] _EVAL_5030;
  wire [15:0] _EVAL_3546;
  wire [15:0] _EVAL_4050;
  wire [15:0] _EVAL_1233;
  wire [15:0] _EVAL_1569;
  wire [15:0] _EVAL_4952;
  wire  _EVAL_3268;
  wire [15:0] _EVAL_2042;
  wire [15:0] _EVAL_2002;
  wire [15:0] _EVAL_776;
  wire [15:0] _EVAL_2716;
  wire [15:0] _EVAL_598;
  wire [15:0] _EVAL_4241;
  wire [15:0] _EVAL_1503;
  wire  _EVAL_424;
  wire  _EVAL_1096;
  wire  _EVAL_1378;
  wire  _EVAL_499;
  wire [4:0] _EVAL_4588;
  wire [15:0] _EVAL_4424;
  wire [15:0] _EVAL_3879;
  wire [15:0] _EVAL_2420;
  wire [15:0] _EVAL_1364;
  wire [15:0] _EVAL_1545;
  wire [15:0] _EVAL_4712;
  wire [15:0] _EVAL_4391;
  wire  _EVAL_388;
  wire  _EVAL_2404;
  wire  _EVAL_3691;
  wire [1:0] _EVAL_4229;
  wire [15:0] _EVAL_2485;
  wire [15:0] _EVAL_2762;
  wire [15:0] _EVAL_5134;
  wire  _EVAL_2958;
  wire  _EVAL_3326;
  wire  _EVAL_4326;
  wire [1:0] _EVAL_864;
  wire [3:0] _EVAL_2550;
  wire  _EVAL_2027;
  wire [15:0] _EVAL_413;
  wire [15:0] _EVAL_3274;
  wire [15:0] _EVAL_1960;
  wire [15:0] _EVAL_5020;
  wire [15:0] _EVAL_3789;
  wire  _EVAL_3759;
  wire  _EVAL_2866;
  wire  _EVAL_613;
  wire [15:0] _EVAL_2720;
  wire [15:0] _EVAL_3897;
  wire [15:0] _EVAL_3638;
  wire [15:0] _EVAL_616;
  wire [15:0] _EVAL_4768;
  wire [15:0] _EVAL_1069;
  wire [15:0] _EVAL_2895;
  wire  _EVAL_2634;
  wire  _EVAL_1208;
  wire [15:0] _EVAL_1090;
  wire [15:0] _EVAL_2872;
  wire [15:0] _EVAL_3964;
  wire [15:0] _EVAL_2347;
  wire [15:0] _EVAL_1534;
  wire [15:0] _EVAL_1615;
  wire [15:0] _EVAL_3804;
  wire [15:0] _EVAL_4522;
  wire [15:0] _EVAL_3990;
  wire [15:0] _EVAL_4396;
  wire [15:0] _EVAL_1039;
  wire [15:0] _EVAL_1630;
  wire [15:0] _EVAL_4295;
  wire [15:0] _EVAL_2903;
  wire [15:0] _EVAL_4418;
  wire [15:0] _EVAL_1949;
  wire [15:0] _EVAL_926;
  wire [15:0] _EVAL_5299;
  wire [15:0] _EVAL_3420;
  wire [15:0] _EVAL_880;
  wire [15:0] _EVAL_4126;
  wire [15:0] _EVAL_4161;
  wire [15:0] _EVAL_1192;
  wire [15:0] _EVAL_5381;
  wire [15:0] _EVAL_2130;
  wire [15:0] _EVAL_5018;
  wire [2:0] _EVAL_1492;
  wire  _EVAL_3226;
  wire [2:0] _EVAL_5197;
  wire  _EVAL_1661;
  wire  _EVAL_327;
  wire  _EVAL_4820;
  wire  _EVAL_3605;
  wire  _EVAL_4811;
  wire  _EVAL_2372;
  wire  _EVAL_3497;
  wire  _EVAL_3528;
  wire  _EVAL_1083;
  wire  _EVAL_4047;
  wire  _EVAL_469;
  wire  _EVAL_1588;
  wire  _EVAL_725;
  wire  _EVAL_405;
  wire  _EVAL_1922;
  wire  _EVAL_1324;
  wire  _EVAL_2977;
  wire [4:0] _EVAL_4832;
  wire  _EVAL_3255;
  wire  _EVAL_5262;
  wire  _EVAL_2162;
  wire  _EVAL_4065;
  wire [31:0] _EVAL_4099;
  wire [31:0] _EVAL_1420;
  wire  _EVAL_5283;
  wire  _EVAL_930;
  wire  _EVAL_4803;
  wire  _EVAL_5082;
  wire [29:0] _EVAL_3160;
  wire [31:0] _EVAL_5181;
  wire [31:0] _EVAL_2215;
  wire [31:0] _EVAL_4983;
  wire [30:0] _EVAL_4752;
  wire  _EVAL_998;
  wire [11:0] _EVAL_4282;
  wire [11:0] _EVAL_1609;
  wire [11:0] _EVAL_3952;
  wire [11:0] _EVAL_3781;
  wire  _EVAL_431;
  wire [19:0] _EVAL_1766;
  wire [31:0] _EVAL_5112;
  wire [31:0] _EVAL_3978;
  wire [31:0] _EVAL_1643;
  wire [31:0] _EVAL_2046;
  wire [26:0] _EVAL_2567;
  wire [31:0] _EVAL_1155;
  wire [31:0] _EVAL_3869;
  wire [31:0] _EVAL_3901;
  wire [32:0] _EVAL_4503;
  wire  _EVAL_3910;
  wire  _EVAL_4705;
  wire  _EVAL_2923;
  wire  _EVAL_1988;
  wire  _EVAL_1400;
  wire  _EVAL_3618;
  wire  _EVAL_345;
  wire  _EVAL_3817;
  wire  _EVAL_873;
  wire  _EVAL_2037;
  wire  _EVAL_1162;
  wire  _EVAL_1291;
  wire  _EVAL_4072;
  wire  _EVAL_4872;
  wire  _EVAL_2237;
  wire  _EVAL_4231;
  wire  _EVAL_286;
  wire  _EVAL_2560;
  wire [14:0] _EVAL_428;
  wire [4:0] _EVAL_1302;
  wire [31:0] _EVAL_4377;
  wire  _EVAL_1125;
  wire  _EVAL_1022;
  wire  _EVAL_4450;
  wire  _EVAL_4483;
  wire  _EVAL_5224;
  wire  _EVAL_4552;
  wire  _EVAL_462;
  wire  _EVAL_3600;
  wire  _EVAL_4719;
  wire  _EVAL_3907;
  wire  _EVAL_2847;
  wire  _EVAL_557;
  wire [11:0] _EVAL_1123;
  wire [11:0] _EVAL_3252;
  wire  _EVAL_2929;
  wire [19:0] _EVAL_938;
  wire [31:0] _EVAL_5254;
  wire [31:0] _EVAL_3324;
  wire [31:0] _EVAL_644;
  wire [31:0] _EVAL_1057;
  wire [26:0] _EVAL_4969;
  wire [31:0] _EVAL_1731;
  wire [31:0] _EVAL_2612;
  wire [31:0] _EVAL_3977;
  wire  _EVAL_4572;
  wire  _EVAL_2471;
  wire [31:0] _EVAL_2951;
  wire [26:0] _EVAL_4659;
  wire [31:0] _EVAL_1483;
  wire  _EVAL_1102;
  wire  _EVAL_354;
  wire  _EVAL_4294;
  wire [15:0] _EVAL_1106;
  wire [15:0] _EVAL_3089;
  wire [15:0] _EVAL_2970;
  wire [15:0] _EVAL_2813;
  wire [15:0] _EVAL_3549;
  wire  _EVAL_3535;
  wire  _EVAL_2106;
  wire  _EVAL_2671;
  wire  _EVAL_3628;
  wire  _EVAL_1220;
  wire [1:0] _EVAL_5186;
  wire  _EVAL_3959;
  wire  _EVAL_2791;
  wire  _EVAL_2430;
  wire [2:0] _EVAL_3499;
  wire  _EVAL_4644;
  wire [15:0] _EVAL_2214;
  wire [15:0] _EVAL_1567;
  wire  _EVAL_1749;
  wire [15:0] _EVAL_4747;
  wire [15:0] _EVAL_4498;
  wire [15:0] _EVAL_2737;
  wire  _EVAL_5195;
  wire  _EVAL_4925;
  wire [1:0] _EVAL_4843;
  wire [1:0] _EVAL_1266;
  wire  _EVAL_1636;
  wire [15:0] _EVAL_3461;
  wire [13:0] _EVAL_2608;
  wire [15:0] _EVAL_4781;
  wire [15:0] _EVAL_2009;
  wire  _EVAL_1551;
  wire [12:0] _EVAL_979;
  wire [15:0] _EVAL_2021;
  wire [15:0] _EVAL_1327;
  wire  _EVAL_1600;
  wire  _EVAL_659;
  wire  _EVAL_4147;
  wire  _EVAL_5065;
  wire  _EVAL_322;
  wire  _EVAL_4615;
  wire  _EVAL_2878;
  wire  _EVAL_4707;
  wire  _EVAL_2475;
  wire  _EVAL_2939;
  wire  _EVAL_3164;
  wire  _EVAL_2599;
  wire  _EVAL_1500;
  wire  _EVAL_1179;
  wire  _EVAL_314;
  wire [15:0] _EVAL_4416;
  wire  _EVAL_603;
  wire  _EVAL_2309;
  wire  _EVAL_1911;
  wire  _EVAL_3561;
  wire  _EVAL_2413;
  wire  _EVAL_3965;
  wire [15:0] _EVAL_2695;
  wire [15:0] _EVAL_4026;
  wire [15:0] _EVAL_3193;
  wire [15:0] _EVAL_4049;
  wire [15:0] _EVAL_3330;
  wire  _EVAL_404;
  wire [15:0] _EVAL_1999;
  wire [15:0] _EVAL_1404;
  wire [15:0] _EVAL_3800;
  wire [15:0] _EVAL_794;
  wire [15:0] _EVAL_2230;
  wire [15:0] _EVAL_1899;
  wire [15:0] _EVAL_461;
  wire [15:0] _EVAL_4591;
  wire [15:0] _EVAL_342;
  wire [15:0] _EVAL_4394;
  wire [15:0] _EVAL_2885;
  wire [15:0] _EVAL_863;
  wire [15:0] _EVAL_3585;
  wire [15:0] _EVAL_4254;
  wire [15:0] _EVAL_4898;
  wire [15:0] _EVAL_5264;
  wire [15:0] _EVAL_4675;
  wire [15:0] _EVAL_577;
  wire [15:0] _EVAL_1914;
  wire [15:0] _EVAL_3992;
  wire [15:0] _EVAL_1032;
  wire [31:0] _EVAL_4961;
  wire  _EVAL_3745;
  wire  _EVAL_1525;
  wire  _EVAL_1527;
  wire  _EVAL_578;
  wire  _EVAL_5093;
  wire  _EVAL_3035;
  wire  _EVAL_1593;
  wire  _EVAL_2785;
  wire  _EVAL_663;
  wire  _EVAL_1868;
  wire  _EVAL_1957;
  wire  _EVAL_1348;
  wire  _EVAL_2077;
  wire  _EVAL_4458;
  wire  _EVAL_2236;
  wire  _EVAL_1010;
  wire  _EVAL_513;
  wire  _EVAL_1690;
  wire  _EVAL_4626;
  wire [2:0] _EVAL_4193;
  wire  _EVAL_1270;
  wire  _EVAL_1970;
  wire  _EVAL_5316;
  wire  _EVAL_4384;
  wire  _EVAL_4448;
  wire  _EVAL_1144;
  wire  _EVAL_2125;
  wire  _EVAL_4339;
  wire  _EVAL_4765;
  wire  _EVAL_1501;
  wire  _EVAL_4726;
  wire [4:0] _EVAL_480;
  wire  _EVAL_5006;
  wire  _EVAL_5163;
  wire  _EVAL_4577;
  wire [4:0] _EVAL_4305;
  wire  _EVAL_1019;
  wire  _EVAL_2718;
  wire  _EVAL_1350;
  wire  _EVAL_2207;
  wire [1:0] _EVAL_727;
  wire  _EVAL_2682;
  wire  _EVAL_2283;
  wire [1:0] _EVAL_941;
  wire  _EVAL_4901;
  wire  _EVAL_4527;
  wire  _EVAL_602;
  wire  _EVAL_2160;
  wire  _EVAL_4451;
  wire  _EVAL_1088;
  wire  _EVAL_5289;
  wire  _EVAL_2256;
  wire  _EVAL_4957;
  wire  _EVAL_2519;
  wire  _EVAL_2908;
  wire  _EVAL_5016;
  wire  _EVAL_3143;
  wire  _EVAL_889;
  wire  _EVAL_5172;
  wire  _EVAL_2582;
  wire  _EVAL_4526;
  wire  _EVAL_2777;
  wire  _EVAL_2659;
  wire  _EVAL_3093;
  wire  _EVAL_3953;
  wire  _EVAL_3859;
  wire  _EVAL_2084;
  wire  _EVAL_1060;
  wire  _EVAL_4382;
  wire  _EVAL_956;
  wire  _EVAL_2221;
  wire  _EVAL_290;
  wire  _EVAL_1920;
  wire  _EVAL_1996;
  wire  _EVAL_2920;
  wire  _EVAL_1442;
  wire  _EVAL_3651;
  wire  _EVAL_2129;
  wire  _EVAL_4311;
  wire  _EVAL_1479;
  wire  _EVAL_3277;
  wire  _EVAL_1178;
  wire  _EVAL_3145;
  wire  _EVAL_1126;
  wire  _EVAL_1714;
  wire  _EVAL_3195;
  wire  _EVAL_5062;
  wire  _EVAL_3155;
  wire  _EVAL_3318;
  wire  _EVAL_3613;
  wire  _EVAL_5281;
  wire  _EVAL_3455;
  wire  _EVAL_4897;
  wire  _EVAL_4525;
  wire  _EVAL_3842;
  wire  _EVAL_4938;
  wire  _EVAL_2640;
  wire  _EVAL_3673;
  wire  _EVAL_3506;
  wire  _EVAL_3033;
  wire  _EVAL_3524;
  wire  _EVAL_5180;
  wire  _EVAL_1349;
  wire [4:0] _EVAL_5129;
  wire  _EVAL_505;
  wire  _EVAL_2902;
  wire  _EVAL_3128;
  wire [4:0] _EVAL_4513;
  wire [11:0] _EVAL_5206;
  wire [11:0] _EVAL_527;
  wire [19:0] _EVAL_2066;
  wire [19:0] _EVAL_4358;
  wire [19:0] _EVAL_5420;
  wire [31:0] _EVAL_1665;
  wire [31:0] _EVAL_4838;
  wire [11:0] _EVAL_1145;
  wire [11:0] _EVAL_2529;
  wire [11:0] _EVAL_2770;
  wire [11:0] _EVAL_1296;
  wire [11:0] _EVAL_1909;
  wire [11:0] _EVAL_3813;
  wire  _EVAL_3737;
  wire [19:0] _EVAL_3069;
  wire [31:0] _EVAL_2417;
  wire [31:0] _EVAL_643;
  wire [31:0] _EVAL_3298;
  wire [31:0] _EVAL_2061;
  wire [31:0] _EVAL_3932;
  wire [26:0] _EVAL_4068;
  wire [31:0] _EVAL_1560;
  wire [31:0] _EVAL_5102;
  wire [31:0] _EVAL_2799;
  wire [29:0] _EVAL_2156;
  wire [6:0] _EVAL_2627;
  wire [127:0] _EVAL_4787;
  wire  _EVAL_2198;
  wire [2:0] _EVAL_2422;
  wire  _EVAL_3639;
  wire [1:0] _EVAL_774;
  wire [3:0] _EVAL_1021;
  wire [7:0] _EVAL_4455;
  wire [2:0] _EVAL_4912;
  wire [4:0] _EVAL_4730;
  wire [27:0] _EVAL_412;
  wire [27:0] _EVAL_1212;
  wire [8:0] _EVAL_3396;
  wire [3:0] _EVAL_3051;
  wire [4:0] _EVAL_1653;
  wire [28:0] _EVAL_390;
  wire  _EVAL_3733;
  wire [4:0] _EVAL_3778;
  wire [24:0] _EVAL_5223;
  wire  _EVAL_4327;
  wire [24:0] _EVAL_3991;
  wire [24:0] _EVAL_3430;
  wire [17:0] _EVAL_3368;
  wire [24:0] _EVAL_911;
  wire [24:0] _EVAL_2474;
  wire [24:0] _EVAL_5282;
  wire [24:0] _EVAL_2149;
  wire [24:0] _EVAL_3091;
  wire [24:0] _EVAL_4446;
  wire [24:0] _EVAL_3650;
  wire [1:0] _EVAL_1577;
  wire [2:0] _EVAL_784;
  wire [27:0] _EVAL_4082;
  wire [27:0] _EVAL_2190;
  wire [28:0] _EVAL_1383;
  wire [25:0] _EVAL_1552;
  wire [28:0] _EVAL_3653;
  wire [28:0] _EVAL_321;
  wire [28:0] _EVAL_3054;
  wire [28:0] _EVAL_1081;
  wire [28:0] _EVAL_3669;
  wire [28:0] _EVAL_294;
  wire [28:0] _EVAL_1711;
  wire [31:0] _EVAL_5114;
  wire  _EVAL_2859;
  wire  _EVAL_2723;
  wire  _EVAL_3485;
  wire  _EVAL_1758;
  wire [26:0] _EVAL_330;
  wire [31:0] _EVAL_1141;
  wire [31:0] _EVAL_3092;
  wire [31:0] _EVAL_3038;
  wire  _EVAL_2578;
  wire [31:0] _EVAL_4578;
  wire [31:0] _EVAL_1142;
  wire [31:0] _EVAL_665;
  wire [2:0] _EVAL_4255;
  wire  _EVAL_854;
  wire  _EVAL_4987;
  wire [1:0] _EVAL_3616;
  wire  _EVAL_1712;
  wire  _EVAL_3105;
  wire  _EVAL_615;
  wire  _EVAL_4328;
  wire  _EVAL_3989;
  wire  _EVAL_2798;
  wire [15:0] _EVAL_1836;
  wire [31:0] _EVAL_3834;
  wire [15:0] _EVAL_2931;
  wire [31:0] _EVAL_759;
  wire [31:0] _EVAL_4492;
  wire [31:0] _EVAL_4066;
  wire [23:0] _EVAL_2790;
  wire [31:0] _EVAL_1117;
  wire [31:0] _EVAL_1154;
  wire [23:0] _EVAL_1449;
  wire [31:0] _EVAL_367;
  wire [31:0] _EVAL_755;
  wire [31:0] _EVAL_4682;
  wire [27:0] _EVAL_3439;
  wire [31:0] _EVAL_5090;
  wire [31:0] _EVAL_3908;
  wire [27:0] _EVAL_640;
  wire [31:0] _EVAL_3357;
  wire [31:0] _EVAL_1936;
  wire [31:0] _EVAL_4873;
  wire  _EVAL_340;
  wire  _EVAL_5318;
  wire  _EVAL_1741;
  wire  _EVAL_3046;
  wire  _EVAL_968;
  wire  _EVAL_1065;
  wire  _EVAL_2719;
  wire  _EVAL_4401;
  wire  _EVAL_4119;
  wire  _EVAL_3743;
  wire  _EVAL_3269;
  wire  _EVAL_5244;
  wire  _EVAL_3299;
  wire [4:0] _EVAL_3598;
  wire  _EVAL_1768;
  wire  _EVAL_4570;
  wire  _EVAL_2094;
  wire  _EVAL_2152;
  wire  _EVAL_4103;
  wire  _EVAL_3119;
  wire  _EVAL_3322;
  wire  _EVAL_2203;
  wire  _EVAL_4630;
  wire [4:0] _EVAL_2059;
  wire  _EVAL_2953;
  wire  _EVAL_4658;
  wire [6:0] _EVAL_416;
  wire [4:0] _EVAL_4859;
  wire [11:0] _EVAL_4045;
  wire [11:0] _EVAL_3911;
  wire  _EVAL_3010;
  wire  _EVAL_3030;
  wire  _EVAL_3703;
  wire  _EVAL_4312;
  wire  _EVAL_2456;
  wire  _EVAL_3377;
  wire  _EVAL_2390;
  wire  _EVAL_4239;
  wire  _EVAL_3175;
  wire  _EVAL_2217;
  wire  _EVAL_1031;
  wire  _EVAL_4907;
  wire  _EVAL_2259;
  wire  _EVAL_5374;
  wire  _EVAL_2660;
  wire  _EVAL_879;
  wire  _EVAL_2817;
  wire  _EVAL_3060;
  wire  _EVAL_4708;
  wire  _EVAL_600;
  wire  _EVAL_4368;
  wire  _EVAL_440;
  wire  _EVAL_3180;
  wire  _EVAL_2685;
  wire  _EVAL_5387;
  wire  _EVAL_2119;
  wire  _EVAL_1985;
  wire  _EVAL_1362;
  wire  _EVAL_4486;
  wire  _EVAL_2995;
  wire  _EVAL_3412;
  wire  _EVAL_5071;
  wire  _EVAL_3787;
  wire  _EVAL_3942;
  wire  _EVAL_449;
  wire  _EVAL_2875;
  wire  _EVAL_4036;
  wire  _EVAL_3111;
  wire  _EVAL_1995;
  wire  _EVAL_2808;
  wire  _EVAL_316;
  wire  _EVAL_4480;
  wire  _EVAL_1275;
  wire  _EVAL_4617;
  wire  _EVAL_5187;
  wire  _EVAL_1408;
  wire  _EVAL_5031;
  wire  _EVAL_1264;
  wire  _EVAL_3971;
  wire  _EVAL_2803;
  wire  _EVAL_4662;
  wire  _EVAL_444;
  wire  _EVAL_4613;
  wire  _EVAL_525;
  wire  _EVAL_2364;
  wire  _EVAL_1127;
  wire  _EVAL_5295;
  wire  _EVAL_2806;
  wire  _EVAL_4244;
  wire  _EVAL_1924;
  wire  _EVAL_5104;
  wire  _EVAL_3565;
  wire  _EVAL_3340;
  wire  _EVAL_4854;
  wire [32:0] _EVAL_3161;
  wire [32:0] _EVAL_3151;
  wire  _EVAL_4098;
  wire  _EVAL_2992;
  wire [32:0] _EVAL_4713;
  wire [32:0] _EVAL_4565;
  wire  _EVAL_1225;
  wire  _EVAL_3208;
  wire  _EVAL_1171;
  wire  _EVAL_3316;
  wire [2:0] _EVAL_2201;
  wire  _EVAL_3188;
  wire  _EVAL_448;
  wire [2:0] _EVAL_2865;
  wire [2:0] _EVAL_3282;
  wire  _EVAL_1812;
  wire  _EVAL_2666;
  wire  _EVAL_4646;
  wire  _EVAL_1973;
  wire  _EVAL_4392;
  wire  _EVAL_2588;
  wire  _EVAL_2937;
  wire  _EVAL_689;
  wire  _EVAL_5023;
  wire  _EVAL_2731;
  wire  _EVAL_4982;
  wire  _EVAL_4583;
  wire  _EVAL_3672;
  wire  _EVAL_4637;
  wire  _EVAL_4643;
  wire  _EVAL_1780;
  wire  _EVAL_2498;
  wire  _EVAL_2810;
  wire  _EVAL_593;
  wire  _EVAL_1523;
  wire  _EVAL_2121;
  wire [2:0] _EVAL_4971;
  wire [1:0] _EVAL_1764;
  wire  _EVAL_750;
  wire  _EVAL_5329;
  wire  _EVAL_799;
  wire [2:0] _EVAL_4091;
  wire  _EVAL_1885;
  wire  _EVAL_1805;
  wire  _EVAL_4786;
  wire [2:0] _EVAL_1274;
  wire [2:0] _EVAL_2679;
  wire  _EVAL_5127;
  wire  _EVAL_1568;
  wire  _EVAL_1775;
  wire  _EVAL_4350;
  wire  _EVAL_3359;
  wire  _EVAL_4183;
  wire  _EVAL_2965;
  wire [4:0] _EVAL_4536;
  wire [2:0] _EVAL_754;
  wire [3:0] _EVAL_1517;
  wire [3:0] _EVAL_3406;
  wire [2:0] _EVAL_945;
  wire [3:0] _EVAL_3515;
  wire [31:0] _EVAL_5091;
  wire [31:0] _EVAL_4238;
  wire  _EVAL_920;
  wire  _EVAL_790;
  wire  _EVAL_3702;
  wire  _EVAL_4284;
  wire  _EVAL_4471;
  wire  _EVAL_5245;
  wire  _EVAL_4048;
  wire  _EVAL_2766;
  wire  _EVAL_4429;
  wire  _EVAL_2848;
  wire  _EVAL_3250;
  wire  _EVAL_3780;
  wire  _EVAL_1263;
  wire  _EVAL_1358;
  wire  _EVAL_4862;
  wire  _EVAL_2406;
  wire  _EVAL_2213;
  wire  _EVAL_5046;
  wire  _EVAL_1396;
  wire  _EVAL_822;
  wire  _EVAL_1018;
  wire  _EVAL_1041;
  wire  _EVAL_671;
  wire  _EVAL_1910;
  wire  _EVAL_4974;
  wire  _EVAL_1659;
  wire  _EVAL_2357;
  wire  _EVAL_1997;
  wire [1:0] _EVAL_3223;
  wire  _EVAL_2164;
  wire [4:0] _EVAL_3943;
  wire  _EVAL_1926;
  wire [4:0] _EVAL_3462;
  wire  _EVAL_5193;
  wire [1:0] _EVAL_2440;
  wire [1:0] _EVAL_2606;
  wire [12:0] _EVAL_558;
  wire  _EVAL_4972;
  wire [5:0] _EVAL_4648;
  wire [3:0] _EVAL_1245;
  wire  _EVAL_3529;
  wire [31:0] _EVAL_4273;
  wire [31:0] _EVAL_2764;
  wire [9:0] _EVAL_3008;
  wire  _EVAL_632;
  wire [1:0] _EVAL_1128;
  wire  _EVAL_3300;
  wire  _EVAL_662;
  wire [2:0] _EVAL_2052;
  wire [20:0] _EVAL_793;
  wire  _EVAL_2026;
  wire [9:0] _EVAL_1951;
  wire  _EVAL_1040;
  wire [7:0] _EVAL_1075;
  wire [31:0] _EVAL_5298;
  wire  _EVAL_5242;
  wire  _EVAL_4995;
  wire  _EVAL_3177;
  wire  _EVAL_3874;
  wire  _EVAL_2265;
  wire  _EVAL_3296;
  wire [2:0] _EVAL_1769;
  wire [2:0] _EVAL_2058;
  wire [2:0] _EVAL_984;
  wire [2:0] _EVAL_1856;
  wire [2:0] _EVAL_1240;
  wire [2:0] _EVAL_1429;
  wire [2:0] _EVAL_3072;
  wire [6:0] _EVAL_1374;
  wire [24:0] _EVAL_310;
  wire [30:0] _EVAL_2038;
  wire  _EVAL_1644;
  wire [30:0] _EVAL_5151;
  wire [30:0] _EVAL_2646;
  wire  _EVAL_1710;
  wire [6:0] _EVAL_2858;
  wire [31:0] _EVAL_2707;
  wire  _EVAL_2601;
  wire [25:0] _EVAL_974;
  wire [30:0] _EVAL_501;
  wire [30:0] _EVAL_1376;
  wire [30:0] _EVAL_1357;
  wire [31:0] _EVAL_1016;
  wire [31:0] _EVAL_1001;
  wire  _EVAL_3716;
  wire [2:0] _EVAL_5339;
  wire [31:0] _EVAL_3810;
  wire [19:0] _EVAL_548;
  wire [31:0] _EVAL_1116;
  wire [31:0] _EVAL_5407;
  wire [31:0] _EVAL_2255;
  wire [31:0] _EVAL_1283;
  wire [31:0] _EVAL_2730;
  wire [31:0] _EVAL_4432;
  wire [31:0] _EVAL_2427;
  wire [31:0] _EVAL_2822;
  wire [31:0] _EVAL_3715;
  wire [31:0] _EVAL_2437;
  wire [31:0] _EVAL_2378;
  wire [31:0] _EVAL_2302;
  wire [4:0] _EVAL_504;
  wire [4:0] _EVAL_5382;
  wire [4:0] _EVAL_1990;
  wire [4:0] _EVAL_1847;
  wire [31:0] _EVAL_3399;
  wire  _EVAL_630;
  wire  _EVAL_4518;
  wire  _EVAL_508;
  wire  _EVAL_3504;
  wire  _EVAL_2915;
  wire  _EVAL_1707;
  wire  _EVAL_4313;
  wire  _EVAL_4992;
  wire  _EVAL_1355;
  wire  _EVAL_3438;
  wire  _EVAL_3246;
  wire  _EVAL_3568;
  wire  _EVAL_3467;
  wire  _EVAL_4150;
  wire [7:0] _EVAL_3894;
  wire  _EVAL_2899;
  wire [22:0] _EVAL_1182;
  wire  _EVAL_299;
  wire  _EVAL_590;
  wire  _EVAL_1450;
  wire [53:0] _EVAL_5334;
  wire [15:0] _EVAL_1870;
  wire [7:0] _EVAL_2006;
  wire [15:0] _EVAL_5309;
  wire [7:0] _EVAL_3960;
  wire [15:0] _EVAL_1917;
  wire [15:0] _EVAL_4935;
  wire [15:0] _EVAL_3495;
  wire [11:0] _EVAL_1810;
  wire [15:0] _EVAL_2670;
  wire [15:0] _EVAL_4496;
  wire [11:0] _EVAL_5267;
  wire [15:0] _EVAL_3056;
  wire [15:0] _EVAL_1160;
  wire [15:0] _EVAL_2628;
  wire [13:0] _EVAL_2815;
  wire [15:0] _EVAL_2459;
  wire [15:0] _EVAL_2819;
  wire [13:0] _EVAL_1642;
  wire [15:0] _EVAL_4121;
  wire [15:0] _EVAL_1224;
  wire [15:0] _EVAL_2739;
  wire [14:0] _EVAL_1017;
  wire [15:0] _EVAL_2642;
  wire [15:0] _EVAL_3741;
  wire [14:0] _EVAL_827;
  wire [15:0] _EVAL_2761;
  wire [15:0] _EVAL_3480;
  wire [15:0] _EVAL_2712;
  wire [6:0] _EVAL_3004;
  wire [3:0] _EVAL_320;
  wire [1:0] _EVAL_1488;
  wire  _EVAL_807;
  wire  _EVAL_3545;
  wire [1:0] _EVAL_4537;
  wire  _EVAL_4910;
  wire  _EVAL_2373;
  wire [2:0] _EVAL_3065;
  wire [1:0] _EVAL_3883;
  wire  _EVAL_2662;
  wire  _EVAL_5200;
  wire  _EVAL_5210;
  wire [22:0] _EVAL_463;
  wire  _EVAL_1377;
  wire  _EVAL_1668;
  wire  _EVAL_840;
  wire  _EVAL_2918;
  wire  _EVAL_5176;
  wire  _EVAL_1382;
  wire  _EVAL_4084;
  wire  _EVAL_2540;
  wire  _EVAL_4407;
  wire  _EVAL_1054;
  wire  _EVAL_1003;
  wire  _EVAL_2202;
  wire  _EVAL_2374;
  wire  _EVAL_2759;
  wire  _EVAL_3786;
  wire  _EVAL_3118;
  wire  _EVAL_4948;
  wire  _EVAL_1375;
  wire  _EVAL_2484;
  wire  _EVAL_4895;
  wire  _EVAL_3040;
  wire  _EVAL_4749;
  wire [4:0] _EVAL_1831;
  wire [4:0] _EVAL_2562;
  wire [4:0] _EVAL_933;
  wire [4:0] _EVAL_4164;
  wire [4:0] _EVAL_3063;
  wire [4:0] _EVAL_3617;
  wire [4:0] _EVAL_741;
  wire [4:0] _EVAL_3484;
  wire [4:0] _EVAL_2674;
  wire [4:0] _EVAL_2314;
  wire [4:0] _EVAL_3941;
  wire [4:0] _EVAL_2633;
  wire [4:0] _EVAL_4321;
  wire [4:0] _EVAL_3871;
  wire [4:0] _EVAL_3993;
  wire [4:0] _EVAL_2183;
  wire [4:0] _EVAL_751;
  wire [4:0] _EVAL_2085;
  wire [4:0] _EVAL_305;
  wire [4:0] _EVAL_1514;
  wire [4:0] _EVAL_2284;
  wire [4:0] _EVAL_596;
  wire [53:0] _EVAL_4625;
  wire [21:0] _EVAL_5257;
  wire [22:0] _EVAL_695;
  wire [22:0] _EVAL_1386;
  wire [24:0] _EVAL_2353;
  wire  _EVAL_4309;
  wire  _EVAL_5252;
  wire  _EVAL_5386;
  wire [4:0] _EVAL_2812;
  wire  _EVAL_743;
  wire  _EVAL_4839;
  wire  _EVAL_3364;
  wire  _EVAL_554;
  wire  _EVAL_3460;
  wire  _EVAL_1228;
  wire  _EVAL_969;
  wire [31:0] _EVAL_4177;
  wire  _EVAL_3271;
  wire  _EVAL_2339;
  wire  _EVAL_523;
  wire [3:0] _EVAL_4191;
  wire [1:0] _EVAL_5168;
  wire [3:0] _EVAL_761;
  wire  _EVAL_451;
  wire [2:0] _EVAL_4892;
  wire  _EVAL_3284;
  wire [1:0] _EVAL_2831;
  wire [3:0] _EVAL_1033;
  wire [7:0] _EVAL_3985;
  wire [2:0] _EVAL_2344;
  wire [4:0] _EVAL_5394;
  wire [4:0] _EVAL_5162;
  wire [27:0] _EVAL_4249;
  wire  _EVAL_4909;
  wire [27:0] _EVAL_1983;
  wire  _EVAL_397;
  wire [2:0] _EVAL_2725;
  wire [2:0] _EVAL_5220;
  wire [8:0] _EVAL_492;
  wire [3:0] _EVAL_4123;
  wire [4:0] _EVAL_550;
  wire [28:0] _EVAL_1675;
  wire  _EVAL_4280;
  wire  _EVAL_2487;
  wire [4:0] _EVAL_475;
  wire [24:0] _EVAL_3144;
  wire  _EVAL_1428;
  wire [24:0] _EVAL_4138;
  wire [24:0] _EVAL_4477;
  wire [17:0] _EVAL_2319;
  wire [24:0] _EVAL_1777;
  wire [24:0] _EVAL_4493;
  wire [24:0] _EVAL_5122;
  wire [24:0] _EVAL_5238;
  wire [24:0] _EVAL_4934;
  wire [24:0] _EVAL_4592;
  wire [24:0] _EVAL_4248;
  wire  _EVAL_5161;
  wire [1:0] _EVAL_3619;
  wire [2:0] _EVAL_978;
  wire [27:0] _EVAL_3777;
  wire  _EVAL_654;
  wire [27:0] _EVAL_2525;
  wire  _EVAL_1897;
  wire [2:0] _EVAL_3643;
  wire [1:0] _EVAL_3935;
  wire [28:0] _EVAL_3738;
  wire [25:0] _EVAL_3327;
  wire [28:0] _EVAL_587;
  wire [28:0] _EVAL_746;
  wire [28:0] _EVAL_982;
  wire [28:0] _EVAL_1756;
  wire [28:0] _EVAL_5191;
  wire [28:0] _EVAL_3878;
  wire [28:0] _EVAL_4470;
  wire [31:0] _EVAL_2522;
  wire [4:0] _EVAL_2637;
  wire  _EVAL_4894;
  wire  _EVAL_2538;
  wire  _EVAL_419;
  wire  _EVAL_2857;
  wire [32:0] _EVAL_1432;
  wire [15:0] _EVAL_1753;
  wire [31:0] _EVAL_4999;
  wire [15:0] _EVAL_962;
  wire [31:0] _EVAL_5156;
  wire [31:0] _EVAL_2124;
  wire [31:0] _EVAL_1578;
  wire [23:0] _EVAL_4320;
  wire [31:0] _EVAL_482;
  wire [31:0] _EVAL_2439;
  wire [23:0] _EVAL_2116;
  wire [31:0] _EVAL_3550;
  wire [31:0] _EVAL_967;
  wire [31:0] _EVAL_3172;
  wire [27:0] _EVAL_343;
  wire [31:0] _EVAL_1581;
  wire [31:0] _EVAL_4061;
  wire [27:0] _EVAL_970;
  wire [31:0] _EVAL_2946;
  wire [31:0] _EVAL_5110;
  wire [31:0] _EVAL_2665;
  wire [29:0] _EVAL_291;
  wire [31:0] _EVAL_2724;
  wire [31:0] _EVAL_852;
  wire [29:0] _EVAL_4850;
  wire [31:0] _EVAL_887;
  wire [31:0] _EVAL_5007;
  wire [31:0] _EVAL_468;
  wire [30:0] _EVAL_4383;
  wire [31:0] _EVAL_620;
  wire [31:0] _EVAL_1599;
  wire [30:0] _EVAL_4403;
  wire [31:0] _EVAL_2032;
  wire [31:0] _EVAL_4604;
  wire [31:0] _EVAL_2571;
  wire [32:0] _EVAL_4116;
  wire [32:0] _EVAL_3593;
  wire [4:0] _EVAL_2192;
  wire [32:0] _EVAL_1005;
  wire [31:0] _EVAL_1735;
  wire [15:0] _EVAL_1774;
  wire [31:0] _EVAL_4144;
  wire [15:0] _EVAL_3150;
  wire [31:0] _EVAL_1012;
  wire [31:0] _EVAL_1467;
  wire [31:0] _EVAL_426;
  wire [23:0] _EVAL_4981;
  wire [31:0] _EVAL_4991;
  wire [31:0] _EVAL_3782;
  wire [23:0] _EVAL_2348;
  wire [31:0] _EVAL_5330;
  wire [31:0] _EVAL_1598;
  wire [31:0] _EVAL_1563;
  wire [27:0] _EVAL_563;
  wire [31:0] _EVAL_496;
  wire [31:0] _EVAL_4234;
  wire [27:0] _EVAL_3665;
  wire [31:0] _EVAL_2526;
  wire [31:0] _EVAL_769;
  wire [31:0] _EVAL_2336;
  wire [29:0] _EVAL_3623;
  wire [31:0] _EVAL_4923;
  wire [31:0] _EVAL_3622;
  wire  _EVAL_3431;
  wire  _EVAL_2197;
  wire  _EVAL_4911;
  wire  _EVAL_4024;
  wire  _EVAL_4034;
  wire  _EVAL_3034;
  wire  _EVAL_3532;
  wire  _EVAL_4474;
  wire  _EVAL_627;
  wire  _EVAL_4774;
  wire  _EVAL_4351;
  wire  _EVAL_3457;
  wire  _EVAL_3876;
  wire  _EVAL_2700;
  wire  _EVAL_1297;
  wire  _EVAL_3273;
  wire [31:0] _EVAL_3279;
  wire [31:0] _EVAL_3187;
  wire [31:0] _EVAL_4993;
  wire [31:0] _EVAL_579;
  wire  _EVAL_3512;
  wire  _EVAL_1789;
  wire  _EVAL_1963;
  wire  _EVAL_4016;
  wire  _EVAL_1030;
  wire  _EVAL_5340;
  wire  _EVAL_1843;
  wire [31:0] _EVAL_4200;
  wire  _EVAL_2144;
  wire  _EVAL_1112;
  wire [6:0] _EVAL_4686;
  wire [1:0] _EVAL_3221;
  wire [4:0] _EVAL_732;
  wire [26:0] _EVAL_636;
  wire [26:0] _EVAL_1893;
  wire [7:0] _EVAL_3983;
  wire [2:0] _EVAL_2807;
  wire [4:0] _EVAL_1806;
  wire [27:0] _EVAL_1006;
  wire [26:0] _EVAL_849;
  wire [26:0] _EVAL_2735;
  wire [26:0] _EVAL_4903;
  wire [27:0] _EVAL_4237;
  wire [3:0] _EVAL_1882;
  wire [1:0] _EVAL_2095;
  wire [29:0] _EVAL_4420;
  wire [29:0] _EVAL_2938;
  wire [29:0] _EVAL_2000;
  wire [29:0] _EVAL_900;
  wire [29:0] _EVAL_4306;
  wire [29:0] _EVAL_1962;
  wire [29:0] _EVAL_529;
  wire [29:0] _EVAL_1708;
  wire [31:0] _EVAL_961;
  wire [31:0] _EVAL_4504;
  wire  _EVAL_2677;
  wire [31:0] _EVAL_2932;
  wire  _EVAL_3328;
  wire  _EVAL_737;
  wire [31:0] _EVAL_2109;
  wire  _EVAL_4549;
  wire  _EVAL_3633;
  wire [31:0] _EVAL_2298;
  wire  _EVAL_2421;
  wire  _EVAL_5184;
  wire [31:0] _EVAL_4454;
  wire  _EVAL_2797;
  wire  _EVAL_1679;
  wire  _EVAL_300;
  wire  _EVAL_1416;
  wire  _EVAL_5408;
  wire  _EVAL_5094;
  wire  _EVAL_700;
  wire  _EVAL_4008;
  wire  _EVAL_3995;
  wire  _EVAL_1292;
  wire  _EVAL_4605;
  wire  _EVAL_3607;
  wire  _EVAL_2242;
  wire  _EVAL_4598;
  wire  _EVAL_3071;
  wire  _EVAL_352;
  wire  _EVAL_387;
  wire  _EVAL_4524;
  wire  _EVAL_4807;
  wire  _EVAL_4476;
  wire  _EVAL_2388;
  wire  _EVAL_2463;
  wire  _EVAL_1281;
  wire  _EVAL_4541;
  wire  _EVAL_4139;
  wire [2:0] _EVAL_3972;
  wire  _EVAL_717;
  wire  _EVAL_3580;
  wire [2:0] _EVAL_4847;
  wire [2:0] _EVAL_791;
  wire [31:0] _EVAL_2442;
  wire [31:0] _EVAL_1746;
  wire [31:0] _EVAL_1063;
  wire [26:0] _EVAL_929;
  wire [31:0] _EVAL_2983;
  wire  _EVAL_2271;
  wire [1:0] _EVAL_459;
  wire [7:0] _EVAL_3646;
  wire [7:0] _EVAL_3966;
  wire [8:0] _EVAL_4547;
  wire  _EVAL_280;
  wire  _EVAL_2818;
  wire  _EVAL_3534;
  wire [2:0] _EVAL_3511;
  wire [29:0] _EVAL_1557;
  wire [31:0] _EVAL_2643;
  wire [29:0] _EVAL_1156;
  wire [31:0] _EVAL_1047;
  wire [31:0] _EVAL_1981;
  wire [29:0] _EVAL_5413;
  wire [31:0] _EVAL_1824;
  wire [31:0] _EVAL_2472;
  wire [31:0] _EVAL_1193;
  wire [30:0] _EVAL_748;
  wire [31:0] _EVAL_540;
  wire [31:0] _EVAL_5054;
  wire  _EVAL_2990;
  wire  _EVAL_2717;
  wire  _EVAL_2263;
  wire [31:0] _EVAL_458;
  wire [31:0] _EVAL_2072;
  wire [31:0] _EVAL_1992;
  wire [26:0] _EVAL_1105;
  wire [32:0] _EVAL_4109;
  wire [31:0] _EVAL_2333;
  wire [31:0] _EVAL_3734;
  wire [32:0] _EVAL_4813;
  wire [32:0] _EVAL_4514;
  wire [31:0] _EVAL_1230;
  wire [31:0] _EVAL_4210;
  wire [1:0] _EVAL_5217;
  wire  _EVAL_4230;
  wire [31:0] _EVAL_5138;
  wire  _EVAL_4031;
  wire  _EVAL_806;
  wire  _EVAL_3709;
  wire  _EVAL_3230;
  wire  _EVAL_3724;
  wire  _EVAL_4574;
  wire  _EVAL_5086;
  wire  _EVAL_3886;
  wire  _EVAL_3575;
  wire [31:0] _EVAL_923;
  wire [31:0] _EVAL_5380;
  wire  _EVAL_1048;
  wire  _EVAL_3927;
  wire [31:0] _EVAL_4888;
  wire [31:0] _EVAL_1140;
  wire  _EVAL_3823;
  wire [31:0] _EVAL_3238;
  wire [31:0] _EVAL_2454;
  wire [31:0] _EVAL_3443;
  wire [31:0] _EVAL_2306;
  wire [31:0] _EVAL_3713;
  wire  _EVAL_2102;
  wire [30:0] _EVAL_1231;
  wire [31:0] _EVAL_2926;
  wire [31:0] _EVAL_2558;
  wire [31:0] _EVAL_1830;
  wire [31:0] _EVAL_2694;
  wire [31:0] _EVAL_3265;
  wire [31:0] _EVAL_3526;
  wire [31:0] _EVAL_4737;
  wire [31:0] _EVAL_1932;
  wire  _EVAL_5288;
  wire  _EVAL_1180;
  wire  _EVAL_719;
  wire  _EVAL_2327;
  wire [31:0] _EVAL_3331;
  wire  _EVAL_373;
  wire  _EVAL_5271;
  wire  _EVAL_1815;
  wire  _EVAL_1558;
  wire [2:0] _EVAL_5056;
  wire  _EVAL_4544;
  wire  _EVAL_3258;
  wire  _EVAL_1098;
  wire  _EVAL_3522;
  wire  _EVAL_5055;
  wire  _EVAL_358;
  wire  _EVAL_5010;
  wire [32:0] _EVAL_2289;
  wire [31:0] _EVAL_2266;
  wire [30:0] _EVAL_1373;
  wire [31:0] _EVAL_2726;
  wire [31:0] _EVAL_3635;
  wire [31:0] _EVAL_1880;
  wire [32:0] _EVAL_1801;
  wire [32:0] _EVAL_1427;
  wire [4:0] _EVAL_3283;
  wire [32:0] _EVAL_803;
  wire [31:0] _EVAL_1505;
  wire [15:0] _EVAL_3885;
  wire  _EVAL_2892;
  wire  _EVAL_2973;
  wire  _EVAL_2041;
  wire [2:0] _EVAL_4089;
  wire [3:0] _EVAL_2636;
  wire [3:0] _EVAL_5321;
  wire [2:0] _EVAL_3379;
  wire [3:0] _EVAL_2303;
  wire  _EVAL_4755;
  wire  _EVAL_5232;
  wire  _EVAL_4880;
  wire  _EVAL_4361;
  wire [2:0] _EVAL_3578;
  wire [3:0] _EVAL_3961;
  wire [3:0] _EVAL_364;
  wire [2:0] _EVAL_991;
  wire [3:0] _EVAL_311;
  wire  _EVAL_4517;
  wire  _EVAL_5411;
  wire  _EVAL_585;
  wire [4:0] _EVAL_3924;
  wire  _EVAL_4298;
  wire [5:0] _EVAL_5377;
  wire [3:0] _EVAL_470;
  wire [12:0] _EVAL_2249;
  wire [12:0] _EVAL_4890;
  wire [12:0] _EVAL_884;
  wire  _EVAL_2317;
  wire  _EVAL_772;
  wire  _EVAL_3057;
  wire  _EVAL_5157;
  wire  _EVAL_607;
  wire  _EVAL_2387;
  wire  _EVAL_4264;
  wire  _EVAL_2768;
  wire  _EVAL_1304;
  wire  _EVAL_5142;
  wire  _EVAL_3947;
  wire  _EVAL_826;
  wire  _EVAL_3356;
  wire  _EVAL_4172;
  wire  _EVAL_3107;
  wire  _EVAL_2693;
  wire [7:0] _EVAL_2577;
  wire  _EVAL_5338;
  wire  _EVAL_5241;
  wire [15:0] _EVAL_4545;
  wire [15:0] _EVAL_3474;
  wire  _EVAL_2436;
  wire  _EVAL_3948;
  wire  _EVAL_2620;
  wire  _EVAL_3783;
  wire  _EVAL_5097;
  wire  _EVAL_4580;
  wire [5:0] _EVAL_1950;
  wire [63:0] _EVAL_4951;
  wire  _EVAL_4865;
  wire  _EVAL_5274;
  wire  _EVAL_4421;
  wire  _EVAL_2246;
  wire  _EVAL_3124;
  wire  _EVAL_1093;
  wire  _EVAL_1345;
  wire  _EVAL_2569;
  wire  _EVAL_667;
  wire  _EVAL_4039;
  wire  _EVAL_532;
  wire  _EVAL_4634;
  wire  _EVAL_5120;
  wire  _EVAL_3856;
  wire  _EVAL_3456;
  wire  _EVAL_2477;
  wire  _EVAL_3854;
  wire  _EVAL_2733;
  wire  _EVAL_2467;
  wire  _EVAL_4227;
  wire  _EVAL_740;
  wire  _EVAL_4714;
  wire  _EVAL_4729;
  wire  _EVAL_4920;
  wire [32:0] _EVAL_4208;
  wire  _EVAL_2914;
  wire  _EVAL_2884;
  wire  _EVAL_1607;
  wire  _EVAL_2727;
  wire  _EVAL_3700;
  wire  _EVAL_4266;
  wire  _EVAL_4353;
  wire  _EVAL_2054;
  wire  _EVAL_3525;
  wire  _EVAL_1484;
  wire  _EVAL_4018;
  wire  _EVAL_5326;
  wire  _EVAL_1934;
  wire  _EVAL_3353;
  wire  _EVAL_4970;
  wire  _EVAL_4433;
  wire  _EVAL_4406;
  wire  _EVAL_4060;
  wire  _EVAL_3157;
  wire  _EVAL_5315;
  wire  _EVAL_1068;
  wire  _EVAL_4587;
  wire  _EVAL_5198;
  wire  _EVAL_4780;
  wire  _EVAL_3304;
  wire  _EVAL_2141;
  wire  _EVAL_650;
  wire [2:0] _EVAL_2157;
  wire [2:0] _EVAL_4439;
  wire [2:0] _EVAL_4104;
  wire [1:0] _EVAL_2111;
  wire [2:0] _EVAL_4794;
  wire [3:0] _EVAL_4595;
  wire  _EVAL_4214;
  wire  _EVAL_5373;
  wire  _EVAL_5248;
  wire  _EVAL_1905;
  wire  _EVAL_1002;
  wire  _EVAL_3746;
  wire  _EVAL_2159;
  wire  _EVAL_1857;
  wire  _EVAL_1713;
  wire  _EVAL_1729;
  wire  _EVAL_3884;
  wire  _EVAL_2365;
  wire  _EVAL_3440;
  wire  _EVAL_779;
  wire  _EVAL_4007;
  wire  _EVAL_1849;
  wire  _EVAL_4376;
  wire  _EVAL_1215;
  wire  _EVAL_918;
  wire  _EVAL_1529;
  wire  _EVAL_5203;
  wire  _EVAL_377;
  wire  _EVAL_3123;
  wire  _EVAL_1397;
  wire  _EVAL_1458;
  wire  _EVAL_4608;
  wire  _EVAL_5324;
  wire  _EVAL_3387;
  wire  _EVAL_5222;
  wire  _EVAL_2925;
  wire  _EVAL_2593;
  wire  _EVAL_2358;
  wire  _EVAL_2828;
  wire  _EVAL_1587;
  wire  _EVAL_3917;
  wire  _EVAL_981;
  wire  _EVAL_2416;
  wire  _EVAL_5261;
  wire  _EVAL_4152;
  wire  _EVAL_1823;
  wire  _EVAL_5034;
  wire  _EVAL_977;
  wire  _EVAL_781;
  wire  _EVAL_1697;
  wire  _EVAL_2287;
  wire  _EVAL_1497;
  wire  _EVAL_4937;
  wire  _EVAL_3423;
  wire  _EVAL_3915;
  wire  _EVAL_796;
  wire  _EVAL_2654;
  wire  _EVAL_2551;
  wire  _EVAL_1405;
  wire  _EVAL_1742;
  wire  _EVAL_478;
  wire  _EVAL_3825;
  wire  _EVAL_3896;
  wire  _EVAL_2231;
  wire  _EVAL_1776;
  wire  _EVAL_1721;
  wire  _EVAL_520;
  wire  _EVAL_1444;
  wire  _EVAL_2318;
  wire  _EVAL_2943;
  wire  _EVAL_3202;
  wire  _EVAL_2023;
  wire  _EVAL_4816;
  wire  _EVAL_4341;
  wire  _EVAL_4521;
  wire  _EVAL_2779;
  wire  _EVAL_384;
  wire  _EVAL_1524;
  wire  _EVAL_1366;
  wire  _EVAL_5026;
  wire  _EVAL_4801;
  wire  _EVAL_4741;
  wire  _EVAL_347;
  wire  _EVAL_415;
  wire  _EVAL_3100;
  wire  _EVAL_1759;
  wire  _EVAL_400;
  wire  _EVAL_1279;
  wire  _EVAL_4171;
  wire  _EVAL_2053;
  wire  _EVAL_2547;
  wire  _EVAL_519;
  wire  _EVAL_3843;
  wire  _EVAL_5423;
  wire  _EVAL_4124;
  wire  _EVAL_2274;
  wire  _EVAL_897;
  wire  _EVAL_1564;
  wire  _EVAL_836;
  wire  _EVAL_5158;
  wire  _EVAL_5143;
  wire  _EVAL_4506;
  wire [3:0] _EVAL_2528;
  wire  _EVAL_1576;
  wire  _EVAL_3220;
  wire  _EVAL_647;
  wire  _EVAL_1086;
  wire  _EVAL_5395;
  wire  _EVAL_1813;
  wire  _EVAL_4641;
  wire  _EVAL_4921;
  wire  _EVAL_4456;
  wire  _EVAL_3458;
  wire  _EVAL_1635;
  wire  _EVAL_3286;
  wire  _EVAL_5192;
  wire  _EVAL_1441;
  wire  _EVAL_2166;
  wire  _EVAL_2167;
  wire  _EVAL_5164;
  wire  _EVAL_4687;
  wire  _EVAL_1413;
  wire  _EVAL_1651;
  wire  _EVAL_2196;
  wire  _EVAL_3215;
  wire  _EVAL_4112;
  wire  _EVAL_4795;
  wire  _EVAL_1510;
  wire  _EVAL_2976;
  wire  _EVAL_5302;
  wire  _EVAL_2691;
  wire  _EVAL_1310;
  wire  _EVAL_464;
  wire  _EVAL_3103;
  wire  _EVAL_5047;
  wire  _EVAL_5002;
  wire  _EVAL_3594;
  wire  _EVAL_552;
  wire  _EVAL_4510;
  wire  _EVAL_2337;
  wire  _EVAL_1869;
  wire  _EVAL_1424;
  wire  _EVAL_2330;
  wire  _EVAL_4100;
  wire  _EVAL_4864;
  wire  _EVAL_1698;
  wire  _EVAL_1808;
  wire  _EVAL_2461;
  wire  _EVAL_5066;
  wire [3:0] _EVAL_567;
  wire  _EVAL_3174;
  wire  _EVAL_1632;
  wire  _EVAL_5355;
  wire  _EVAL_1640;
  wire  _EVAL_3632;
  wire  _EVAL_4247;
  wire  _EVAL_1646;
  wire  _EVAL_1547;
  wire  _EVAL_518;
  wire  _EVAL_3015;
  wire  _EVAL_324;
  wire  _EVAL_3951;
  wire  _EVAL_1672;
  wire  _EVAL_1979;
  wire  _EVAL_1894;
  wire  _EVAL_5383;
  wire  _EVAL_4849;
  wire  _EVAL_1451;
  wire  _EVAL_1046;
  wire  _EVAL_5319;
  wire  _EVAL_538;
  wire  _EVAL_4386;
  wire  _EVAL_2345;
  wire  _EVAL_3498;
  wire  _EVAL_2734;
  wire [1:0] _EVAL_2064;
  wire  _EVAL_2003;
  wire [1:0] _EVAL_4751;
  wire [2:0] _EVAL_4776;
  wire  _EVAL_2927;
  wire  _EVAL_766;
  wire  _EVAL_626;
  wire [4:0] _EVAL_3184;
  wire [1:0] _EVAL_2655;
  wire [1:0] _EVAL_3253;
  wire [12:0] _EVAL_1159;
  wire  _EVAL_4702;
  wire [5:0] _EVAL_453;
  wire [3:0] _EVAL_2381;
  wire  _EVAL_2949;
  wire [31:0] _EVAL_814;
  wire [31:0] _EVAL_3351;
  wire [31:0] _EVAL_2071;
  wire  _EVAL_3131;
  wire  _EVAL_3655;
  wire  _EVAL_555;
  wire  _EVAL_4857;
  wire  _EVAL_4198;
  wire  _EVAL_3657;
  wire [2:0] _EVAL_975;
  wire [2:0] _EVAL_2684;
  wire [2:0] _EVAL_4037;
  wire [2:0] _EVAL_1498;
  wire [2:0] _EVAL_1254;
  wire [6:0] _EVAL_1391;
  wire [24:0] _EVAL_4487;
  wire [30:0] _EVAL_5304;
  wire  _EVAL_5125;
  wire [30:0] _EVAL_733;
  wire [30:0] _EVAL_2623;
  wire  _EVAL_1797;
  wire [6:0] _EVAL_1410;
  wire [31:0] _EVAL_2462;
  wire  _EVAL_5359;
  wire [25:0] _EVAL_628;
  wire [30:0] _EVAL_4619;
  wire [30:0] _EVAL_5308;
  wire [30:0] _EVAL_679;
  wire [31:0] _EVAL_1317;
  wire [31:0] _EVAL_795;
  wire  _EVAL_2324;
  wire [31:0] _EVAL_4563;
  wire [14:0] _EVAL_5365;
  wire [31:0] _EVAL_1313;
  wire [19:0] _EVAL_2521;
  wire [31:0] _EVAL_5078;
  wire [31:0] _EVAL_1353;
  wire [31:0] _EVAL_2247;
  wire [31:0] _EVAL_2253;
  wire [31:0] _EVAL_2204;
  wire [31:0] _EVAL_705;
  wire [31:0] _EVAL_3257;
  wire [31:0] _EVAL_3261;
  wire [31:0] _EVAL_4584;
  wire [31:0] _EVAL_4856;
  wire [31:0] _EVAL_1475;
  wire [31:0] _EVAL_4855;
  wire  _EVAL_1262;
  wire  _EVAL_2224;
  wire [15:0] _EVAL_5291;
  wire  _EVAL_2964;
  wire [31:0] _EVAL_2619;
  wire  _EVAL_1244;
  wire [31:0] _EVAL_1049;
  wire [31:0] _EVAL_517;
  wire  _EVAL_4226;
  wire  _EVAL_2146;
  wire [4:0] _EVAL_1555;
  wire  _EVAL_5414;
  wire  _EVAL_346;
  wire  _EVAL_5393;
  wire  _EVAL_3372;
  wire  _EVAL_1426;
  wire  _EVAL_3416;
  wire  _EVAL_5042;
  wire  _EVAL_2185;
  wire  _EVAL_4568;
  wire  _EVAL_4793;
  wire  _EVAL_3680;
  wire  _EVAL_2515;
  wire  _EVAL_848;
  wire  _EVAL_1015;
  wire  _EVAL_1246;
  wire [22:0] _EVAL_2110;
  wire  _EVAL_3088;
  wire  _EVAL_768;
  wire [1:0] _EVAL_2449;
  wire  _EVAL_757;
  wire [31:0] _EVAL_3705;
  wire [4:0] _EVAL_4869;
  wire  _EVAL_544;
  wire [4:0] _EVAL_3171;
  wire  _EVAL_2180;
  wire [4:0] _EVAL_2991;
  wire [4:0] _EVAL_2074;
  wire [4:0] _EVAL_3806;
  wire [4:0] _EVAL_675;
  wire [4:0] _EVAL_4252;
  wire  _EVAL_1206;
  wire  _EVAL_2763;
  wire  _EVAL_3149;
  wire  _EVAL_4688;
  wire  _EVAL_5378;
  wire [3:0] _EVAL_2012;
  wire [3:0] _EVAL_5087;
  wire  _EVAL_1940;
  wire  _EVAL_4215;
  wire  _EVAL_2135;
  wire  _EVAL_4823;
  wire [1:0] _EVAL_1139;
  wire  _EVAL_2134;
  wire [31:0] _EVAL_3641;
  wire [31:0] _EVAL_4885;
  wire  _EVAL_597;
  wire  _EVAL_4221;
  wire  _EVAL_3210;
  wire [31:0] _EVAL_2867;
  wire  _EVAL_3930;
  wire  _EVAL_1603;
  wire  _EVAL_2940;
  wire  _EVAL_5385;
  wire  _EVAL_3075;
  wire  _EVAL_641;
  wire [3:0] _EVAL_331;
  wire [31:0] _EVAL_1079;
  wire [31:0] _EVAL_5297;
  wire [31:0] _EVAL_2346;
  wire [31:0] _EVAL_1138;
  wire  _EVAL_4085;
  wire  _EVAL_2229;
  wire  _EVAL_2435;
  wire [2:0] _EVAL_4624;
  wire  _EVAL_2922;
  wire [1:0] _EVAL_3831;
  wire  _EVAL_4163;
  wire  _EVAL_4044;
  wire  _EVAL_5167;
  wire [2:0] _EVAL_5170;
  wire [2:0] _EVAL_4699;
  wire [2:0] _EVAL_1300;
  wire  _EVAL_707;
  wire  _EVAL_1100;
  wire  _EVAL_1487;
  wire  _EVAL_1533;
  wire  _EVAL_3540;
  wire  _EVAL_629;
  wire  _EVAL_5183;
  wire  _EVAL_2869;
  wire  _EVAL_702;
  wire [32:0] _EVAL_3037;
  wire [32:0] _EVAL_2782;
  wire [31:0] _EVAL_3892;
  wire [31:0] _EVAL_5117;
  wire [1:0] _EVAL_1101;
  wire  _EVAL_1941;
  wire  _EVAL_782;
  wire  _EVAL_3938;
  wire  _EVAL_2647;
  wire  _EVAL_1494;
  wire  _EVAL_4413;
  wire  _EVAL_3031;
  wire  _EVAL_5015;
  wire  _EVAL_696;
  wire [31:0] _EVAL_2151;
  wire [31:0] _EVAL_1119;
  wire [31:0] _EVAL_4585;
  wire  _EVAL_718;
  wire  _EVAL_676;
  wire  _EVAL_681;
  wire [32:0] _EVAL_4668;
  wire [15:0] _EVAL_3186;
  wire [31:0] _EVAL_4612;
  wire [15:0] _EVAL_4211;
  wire [31:0] _EVAL_2796;
  wire [31:0] _EVAL_744;
  wire [31:0] _EVAL_4586;
  wire [23:0] _EVAL_562;
  wire [31:0] _EVAL_4017;
  wire [31:0] _EVAL_4763;
  wire [23:0] _EVAL_4861;
  wire [31:0] _EVAL_1078;
  wire [31:0] _EVAL_2142;
  wire [31:0] _EVAL_1633;
  wire [27:0] _EVAL_3905;
  wire [31:0] _EVAL_1745;
  wire [31:0] _EVAL_656;
  wire [27:0] _EVAL_1657;
  wire [31:0] _EVAL_5333;
  wire [31:0] _EVAL_1898;
  wire [31:0] _EVAL_3521;
  wire [29:0] _EVAL_1550;
  wire [31:0] _EVAL_5038;
  wire [31:0] _EVAL_1365;
  wire [29:0] _EVAL_3967;
  wire [31:0] _EVAL_688;
  wire [31:0] _EVAL_4853;
  wire [31:0] _EVAL_3446;
  wire [30:0] _EVAL_1848;
  wire [31:0] _EVAL_1197;
  wire [31:0] _EVAL_2896;
  wire [30:0] _EVAL_3998;
  wire [31:0] _EVAL_3251;
  wire [31:0] _EVAL_4408;
  wire [31:0] _EVAL_3547;
  wire [32:0] _EVAL_3866;
  wire [32:0] _EVAL_303;
  wire [4:0] _EVAL_3683;
  wire [32:0] _EVAL_2894;
  wire [31:0] _EVAL_1866;
  wire [31:0] _EVAL_5215;
  wire  _EVAL_1944;
  wire [15:0] _EVAL_5328;
  wire [31:0] _EVAL_2264;
  wire [15:0] _EVAL_3615;
  wire [31:0] _EVAL_5124;
  wire [31:0] _EVAL_3601;
  wire [31:0] _EVAL_4371;
  wire [23:0] _EVAL_2516;
  wire [31:0] _EVAL_4412;
  wire [31:0] _EVAL_1331;
  wire [23:0] _EVAL_2520;
  wire [31:0] _EVAL_5336;
  wire [31:0] _EVAL_668;
  wire [31:0] _EVAL_3182;
  wire [27:0] _EVAL_5231;
  wire [31:0] _EVAL_4958;
  wire [31:0] _EVAL_3572;
  wire [27:0] _EVAL_642;
  wire [31:0] _EVAL_1312;
  wire [31:0] _EVAL_5033;
  wire [31:0] _EVAL_3337;
  wire [29:0] _EVAL_3564;
  wire [31:0] _EVAL_4616;
  wire [31:0] _EVAL_3833;
  wire [29:0] _EVAL_3189;
  wire [31:0] _EVAL_658;
  wire [31:0] _EVAL_2663;
  wire [31:0] _EVAL_4342;
  wire [30:0] _EVAL_2984;
  wire [31:0] _EVAL_3397;
  wire [31:0] _EVAL_553;
  wire [30:0] _EVAL_2392;
  wire [31:0] _EVAL_1265;
  wire [31:0] _EVAL_3891;
  wire [31:0] _EVAL_3749;
  wire [31:0] _EVAL_572;
  wire [31:0] _EVAL_3726;
  wire [31:0] _EVAL_1495;
  wire [31:0] _EVAL_2845;
  wire [31:0] _EVAL_4399;
  wire  _EVAL_924;
  wire  _EVAL_1891;
  wire  _EVAL_3378;
  wire [32:0] _EVAL_4870;
  wire [32:0] _EVAL_1715;
  wire [32:0] _EVAL_943;
  wire [31:0] _EVAL_4330;
  wire [31:0] _EVAL_363;
  wire [1:0] _EVAL_1784;
  wire  _EVAL_986;
  wire  _EVAL_4946;
  wire  _EVAL_3729;
  wire  _EVAL_3756;
  wire  _EVAL_1841;
  wire [31:0] _EVAL_2947;
  wire [31:0] _EVAL_1489;
  wire  _EVAL_4717;
  wire  _EVAL_4651;
  wire [31:0] _EVAL_2950;
  wire [31:0] _EVAL_3447;
  wire  _EVAL_1662;
  wire [31:0] _EVAL_1791;
  wire [31:0] _EVAL_2179;
  wire [31:0] _EVAL_1833;
  wire [31:0] _EVAL_2769;
  wire  _EVAL_4694;
  wire [31:0] _EVAL_3487;
  wire  _EVAL_698;
  wire [31:0] _EVAL_1720;
  wire [15:0] _EVAL_571;
  wire [31:0] _EVAL_3136;
  wire [31:0] _EVAL_1295;
  wire [31:0] _EVAL_484;
  wire [23:0] _EVAL_2418;
  wire [31:0] _EVAL_5119;
  wire [31:0] _EVAL_2713;
  wire [23:0] _EVAL_1663;
  wire [31:0] _EVAL_4777;
  wire [31:0] _EVAL_4784;
  wire [31:0] _EVAL_385;
  wire [27:0] _EVAL_638;
  wire [31:0] _EVAL_4331;
  wire [31:0] _EVAL_3206;
  wire [27:0] _EVAL_1554;
  wire [31:0] _EVAL_4315;
  wire [31:0] _EVAL_4529;
  wire [31:0] _EVAL_2837;
  wire [29:0] _EVAL_4868;
  wire [31:0] _EVAL_2433;
  wire [31:0] _EVAL_3773;
  wire [29:0] _EVAL_1058;
  wire [31:0] _EVAL_825;
  wire [31:0] _EVAL_5005;
  wire [31:0] _EVAL_3179;
  wire [30:0] _EVAL_4922;
  wire [31:0] _EVAL_4434;
  wire [31:0] _EVAL_5028;
  wire [30:0] _EVAL_2755;
  wire [31:0] _EVAL_4076;
  wire [31:0] _EVAL_3437;
  wire [31:0] _EVAL_2240;
  wire [31:0] _EVAL_4258;
  wire [31:0] _EVAL_3595;
  wire [31:0] _EVAL_3125;
  wire [31:0] _EVAL_942;
  wire [31:0] _EVAL_3923;
  wire  _EVAL_2039;
  wire  _EVAL_932;
  wire  _EVAL_1961;
  wire  _EVAL_5350;
  wire  _EVAL_5092;
  wire  _EVAL_4599;
  wire [31:0] _EVAL_3185;
  wire [31:0] _EVAL_1044;
  wire [31:0] _EVAL_2877;
  wire [31:0] _EVAL_3262;
  wire [31:0] _EVAL_2199;
  wire  _EVAL_2004;
  wire [23:0] _EVAL_5323;
  wire  _EVAL_1803;
  wire  _EVAL_450;
  wire [1:0] _EVAL_3790;
  wire  _EVAL_4114;
  wire  _EVAL_660;
  wire  _EVAL_4426;
  wire  _EVAL_2871;
  wire  _EVAL_5263;
  wire  _EVAL_4235;
  wire  _EVAL_1549;
  wire  _EVAL_2689;
  wire  _EVAL_3811;
  wire  _EVAL_2829;
  wire  _EVAL_4988;
  wire  _EVAL_4661;
  wire  _EVAL_5409;
  wire  _EVAL_4117;
  wire  _EVAL_4325;
  wire  _EVAL_3207;
  wire  _EVAL_357;
  wire  _EVAL_2115;
  wire  _EVAL_576;
  wire  _EVAL_3349;
  wire  _EVAL_3807;
  wire  _EVAL_2616;
  wire  _EVAL_2438;
  wire  _EVAL_905;
  wire  _EVAL_1821;
  wire  _EVAL_5419;
  wire  _EVAL_2850;
  wire  _EVAL_703;
  wire  _EVAL_5417;
  wire  _EVAL_4023;
  wire  _EVAL_4078;
  wire  _EVAL_4209;
  wire  _EVAL_1061;
  wire  _EVAL_3190;
  wire  _EVAL_3644;
  wire  _EVAL_2233;
  wire  _EVAL_2403;
  wire  _EVAL_2013;
  wire  _EVAL_5208;
  wire  _EVAL_4141;
  wire  _EVAL_5201;
  wire  _EVAL_1196;
  wire  _EVAL_4449;
  wire [2:0] _EVAL_5022;
  wire  _EVAL_5107;
  wire  _EVAL_2545;
  wire  _EVAL_4826;
  wire  _EVAL_1243;
  wire  _EVAL_3533;
  wire  _EVAL_1267;
  wire  _EVAL_2079;
  wire  _EVAL_1273;
  wire  _EVAL_3113;
  wire [32:0] _EVAL_1490;
  wire [32:0] _EVAL_2200;
  wire  _EVAL_1165;
  wire  _EVAL_2226;
  wire [32:0] _EVAL_2174;
  wire [32:0] _EVAL_5327;
  wire  _EVAL_3979;
  wire [1:0] _EVAL_3682;
  wire  _EVAL_1330;
  wire  _EVAL_910;
  wire  _EVAL_4056;
  wire  _EVAL_838;
  wire  _EVAL_3452;
  wire  _EVAL_3658;
  wire [2:0] _EVAL_2270;
  wire  _EVAL_664;
  wire  _EVAL_2457;
  wire  _EVAL_4680;
  wire  _EVAL_2434;
  wire  _EVAL_1864;
  wire  _EVAL_2076;
  wire  _EVAL_4170;
  wire  _EVAL_2480;
  wire  _EVAL_1448;
  wire  _EVAL_5113;
  wire  _EVAL_430;
  wire  _EVAL_4129;
  wire  _EVAL_815;
  wire  _EVAL_4069;
  wire  _EVAL_3753;
  wire  _EVAL_4789;
  wire  _EVAL_1887;
  wire  _EVAL_3853;
  wire  _EVAL_1430;
  wire  _EVAL_2649;
  wire  _EVAL_581;
  wire  _EVAL_1221;
  wire  _EVAL_4410;
  wire  _EVAL_5354;
  wire  _EVAL_3689;
  wire  _EVAL_1543;
  wire  _EVAL_3847;
  wire  _EVAL_2635;
  wire  _EVAL_4279;
  wire  _EVAL_2335;
  wire  _EVAL_917;
  wire  _EVAL_1726;
  wire  _EVAL_4840;
  wire  _EVAL_2148;
  wire  _EVAL_4874;
  wire  _EVAL_4846;
  wire  _EVAL_4159;
  wire  _EVAL_2228;
  wire  _EVAL_1530;
  wire  _EVAL_2844;
  wire  _EVAL_1177;
  wire  _EVAL_2773;
  wire  _EVAL_1515;
  wire  _EVAL_853;
  wire  _EVAL_5101;
  wire  _EVAL_4766;
  wire  _EVAL_1388;
  wire  _EVAL_1718;
  wire  _EVAL_2341;
  wire  _EVAL_1620;
  wire  _EVAL_3626;
  wire  _EVAL_964;
  wire  _EVAL_801;
  wire  _EVAL_5141;
  wire  _EVAL_4499;
  wire  _EVAL_1767;
  wire  _EVAL_2827;
  wire  _EVAL_1183;
  wire  _EVAL_992;
  wire  _EVAL_4654;
  wire  _EVAL_442;
  wire  _EVAL_875;
  wire  _EVAL_1858;
  wire  _EVAL_3408;
  wire  _EVAL_4485;
  wire  _EVAL_1315;
  wire  _EVAL_1877;
  wire  _EVAL_5063;
  wire  _EVAL_1888;
  wire  _EVAL_3527;
  wire  _EVAL_467;
  wire  _EVAL_5204;
  wire  _EVAL_2007;
  wire  _EVAL_2279;
  wire  _EVAL_370;
  wire  _EVAL_5347;
  wire  _EVAL_1594;
  wire  _EVAL_2986;
  wire  _EVAL_4184;
  wire  _EVAL_3464;
  wire  _EVAL_2468;
  wire  _EVAL_4276;
  wire  _EVAL_2639;
  wire  _EVAL_1693;
  wire  _EVAL_1073;
  wire  _EVAL_4557;
  wire  _EVAL_1440;
  wire  _EVAL_503;
  wire  _EVAL_438;
  wire  _EVAL_1229;
  wire  _EVAL_2889;
  wire  _EVAL_4317;
  wire  _EVAL_1301;
  wire  _EVAL_1993;
  wire  _EVAL_1682;
  wire  _EVAL_2618;
  wire  _EVAL_5103;
  wire  _EVAL_699;
  wire  _EVAL_1980;
  wire  _EVAL_2482;
  wire  _EVAL_3139;
  wire  _EVAL_3799;
  wire  _EVAL_3514;
  wire  _EVAL_770;
  wire [32:0] _EVAL_1839;
  wire [31:0] _EVAL_3792;
  wire [32:0] _EVAL_1987;
  wire [32:0] _EVAL_5199;
  wire [31:0] _EVAL_3860;
  wire [31:0] _EVAL_2830;
  wire [1:0] _EVAL_2211;
  wire  _EVAL_2432;
  wire  _EVAL_4366;
  wire  _EVAL_3478;
  wire  _EVAL_592;
  wire  _EVAL_1986;
  wire  _EVAL_491;
  wire  _EVAL_2010;
  wire  _EVAL_1092;
  wire  _EVAL_3640;
  wire  _EVAL_3058;
  wire [31:0] _EVAL_3929;
  wire [31:0] _EVAL_5137;
  wire  _EVAL_3664;
  wire  _EVAL_2610;
  wire [31:0] _EVAL_4268;
  wire [31:0] _EVAL_2988;
  wire  _EVAL_1673;
  wire [31:0] _EVAL_2248;
  wire [31:0] _EVAL_4739;
  wire [31:0] _EVAL_1343;
  wire [31:0] _EVAL_1739;
  wire  _EVAL_1666;
  wire [31:0] _EVAL_3468;
  wire  _EVAL_4134;
  wire [29:0] _EVAL_3916;
  wire [31:0] _EVAL_2473;
  wire [31:0] _EVAL_1217;
  wire [31:0] _EVAL_720;
  wire [30:0] _EVAL_5080;
  wire [31:0] _EVAL_4323;
  wire [31:0] _EVAL_3410;
  wire [30:0] _EVAL_2792;
  wire [31:0] _EVAL_2702;
  wire [31:0] _EVAL_381;
  wire [31:0] _EVAL_3411;
  wire [31:0] _EVAL_1512;
  wire [31:0] _EVAL_5361;
  wire [31:0] _EVAL_1572;
  wire  _EVAL_2073;
  wire  _EVAL_4207;
  wire  _EVAL_436;
  wire  _EVAL_1205;
  wire  _EVAL_4824;
  wire  _EVAL_820;
  wire  _EVAL_5189;
  wire  _EVAL_2478;
  wire  _EVAL_391;
  wire  _EVAL_1129;
  wire  _EVAL_4097;
  wire  _EVAL_2971;
  wire  _EVAL_1485;
  wire  _EVAL_4810;
  wire  _EVAL_3801;
  wire  _EVAL_4977;
  wire  _EVAL_4046;
  wire  _EVAL_2464;
  wire [31:0] _EVAL_1853;
  wire [31:0] _EVAL_5376;
  wire [31:0] _EVAL_5310;
  wire [31:0] _EVAL_568;
  wire [31:0] _EVAL_4878;
  wire [31:0] _EVAL_1457;
  wire [31:0] _EVAL_1974;
  wire [31:0] _EVAL_1288;
  wire [31:0] _EVAL_1257;
  wire [31:0] _EVAL_886;
  wire [31:0] _EVAL_1431;
  wire  _EVAL_3135;
  wire  _EVAL_4405;
  wire  _EVAL_4292;
  wire  _EVAL_3083;
  wire  _EVAL_3426;
  wire  _EVAL_5075;
  wire  _EVAL_3723;
  wire  _EVAL_2652;
  wire  _EVAL_3581;
  wire  _EVAL_4571;
  wire  _EVAL_3870;
  wire  _EVAL_4978;
  wire  _EVAL_2963;
  wire  _EVAL_3028;
  wire  _EVAL_1020;
  wire [4:0] _EVAL_2784;
  wire  _EVAL_1114;
  wire  _EVAL_2414;
  wire  _EVAL_445;
  wire  _EVAL_3336;
  wire  _EVAL_4554;
  wire  _EVAL_1937;
  wire  _EVAL_2598;
  wire  _EVAL_5317;
  wire  _EVAL_765;
  wire  _EVAL_3837;
  wire  _EVAL_1975;
  wire  _EVAL_5177;
  wire  _EVAL_2824;
  wire  _EVAL_1094;
  wire  _EVAL_3442;
  wire  _EVAL_1029;
  wire  _EVAL_5053;
  wire  _EVAL_1089;
  wire  _EVAL_2367;
  wire  _EVAL_3199;
  wire  _EVAL_1406;
  wire  _EVAL_2273;
  wire [4:0] _EVAL_4009;
  wire  _EVAL_2276;
  wire  _EVAL_1873;
  wire  _EVAL_4438;
  wire  _EVAL_4502;
  wire  _EVAL_3612;
  wire  _EVAL_3945;
  wire  _EVAL_2993;
  wire  _EVAL_786;
  wire  _EVAL_4293;
  wire  _EVAL_812;
  wire  _EVAL_2078;
  wire  _EVAL_4012;
  wire  _EVAL_2334;
  wire  _EVAL_4990;
  wire  _EVAL_3084;
  wire  _EVAL_4511;
  wire  _EVAL_4681;
  wire  _EVAL_4058;
  wire  _EVAL_4263;
  wire  _EVAL_4579;
  wire  _EVAL_479;
  wire  _EVAL_2672;
  wire  _EVAL_1892;
  wire  _EVAL_4835;
  wire  _EVAL_3698;
  wire  _EVAL_2411;
  wire  _EVAL_1686;
  wire [4:0] _EVAL_521;
  wire  _EVAL_4006;
  wire  _EVAL_1872;
  wire  _EVAL_4775;
  wire  _EVAL_745;
  wire  _EVAL_2385;
  wire  _EVAL_1945;
  wire  _EVAL_987;
  wire  _EVAL_5421;
  wire  _EVAL_1314;
  wire  _EVAL_2293;
  wire  _EVAL_1211;
  wire  _EVAL_3562;
  wire  _EVAL_682;
  wire  _EVAL_1586;
  wire  _EVAL_4029;
  wire  _EVAL_4013;
  wire  _EVAL_2212;
  wire  _EVAL_2288;
  wire  _EVAL_4509;
  wire  _EVAL_3654;
  wire  _EVAL_5118;
  wire  _EVAL_5322;
  wire  _EVAL_5402;
  wire  _EVAL_5415;
  wire  _EVAL_4369;
  wire  _EVAL_4265;
  wire  _EVAL_427;
  wire  _EVAL_2580;
  wire  _EVAL_3970;
  wire  _EVAL_1371;
  wire  _EVAL_3129;
  wire  _EVAL_1669;
  wire  _EVAL_805;
  wire  _EVAL_3699;
  wire  _EVAL_2492;
  wire  _EVAL_3835;
  wire  _EVAL_2728;
  wire  _EVAL_1743;
  wire  _EVAL_4916;
  wire  _EVAL_4111;
  wire  _EVAL_3303;
  wire  _EVAL_773;
  wire  _EVAL_4187;
  wire  _EVAL_1900;
  wire  _EVAL_3348;
  wire  _EVAL_1252;
  wire  _EVAL_1906;
  wire  _EVAL_293;
  wire  _EVAL_2531;
  wire  _EVAL_2170;
  wire  _EVAL_5346;
  wire  _EVAL_435;
  wire  _EVAL_3343;
  wire  _EVAL_4042;
  wire  _EVAL_4071;
  wire  _EVAL_5040;
  wire  _EVAL_4821;
  wire  _EVAL_3779;
  wire  _EVAL_2891;
  wire  _EVAL_5116;
  wire  _EVAL_4381;
  wire  _EVAL_4137;
  wire  _EVAL_5098;
  wire  _EVAL_1131;
  wire  _EVAL_3761;
  wire  _EVAL_5147;
  wire  _EVAL_2789;
  wire  _EVAL_3589;
  wire  _EVAL_4057;
  wire  _EVAL_3895;
  wire  _EVAL_4582;
  wire  _EVAL_4286;
  wire  _EVAL_868;
  wire  _EVAL_2182;
  wire  _EVAL_1584;
  wire  _EVAL_4250;
  wire  _EVAL_1422;
  wire  _EVAL_3213;
  wire  _EVAL_3264;
  wire  _EVAL_2574;
  wire  _EVAL_4243;
  wire  _EVAL_4852;
  wire  _EVAL_2585;
  wire  _EVAL_5287;
  wire  _EVAL_1258;
  wire  _EVAL_3647;
  wire  _EVAL_4742;
  wire  _EVAL_3486;
  wire  _EVAL_1008;
  wire  _EVAL_1667;
  wire  _EVAL_4156;
  wire  _EVAL_3234;
  wire  _EVAL_344;
  wire  _EVAL_2917;
  wire  _EVAL_4792;
  wire  _EVAL_5345;
  wire  _EVAL_1799;
  wire  _EVAL_4500;
  wire  _EVAL_2597;
  wire  _EVAL_4650;
  wire  _EVAL_594;
  wire  _EVAL_3809;
  wire  _EVAL_966;
  wire  _EVAL_3501;
  wire  _EVAL_3739;
  wire  _EVAL_2028;
  wire  _EVAL_3290;
  wire  _EVAL_4136;
  wire  _EVAL_3541;
  wire  _EVAL_4441;
  wire  _EVAL_1234;
  wire  _EVAL_2987;
  wire  _EVAL_3812;
  wire  _EVAL_4055;
  wire  _EVAL_1011;
  wire [4:0] _EVAL_2839;
  wire [4:0] _EVAL_3158;
  wire [19:0] _EVAL_4169;
  wire [19:0] _EVAL_997;
  wire  _EVAL_4665;
  wire  _EVAL_3928;
  wire  _EVAL_1334;
  wire  _EVAL_4467;
  wire  _EVAL_4175;
  wire  _EVAL_1519;
  wire  _EVAL_1804;
  wire  _EVAL_1278;
  wire  _EVAL_2710;
  wire  _EVAL_856;
  wire  _EVAL_3659;
  wire  _EVAL_417;
  wire [31:0] _EVAL_1556;
  wire [32:0] _EVAL_2936;
  wire [32:0] _EVAL_2262;
  wire [32:0] _EVAL_1385;
  wire  _EVAL_476;
  wire  _EVAL_3043;
  wire  _EVAL_5032;
  wire  _EVAL_1071;
  wire  _EVAL_4716;
  wire  _EVAL_3444;
  wire  _EVAL_1998;
  wire  _EVAL_2019;
  wire  _EVAL_3191;
  wire  _EVAL_3857;
  wire  _EVAL_2163;
  wire  _EVAL_5303;
  wire  _EVAL_5255;
  wire  _EVAL_4032;
  wire  _EVAL_1566;
  wire  _EVAL_2340;
  wire  _EVAL_4930;
  wire  _EVAL_599;
  wire  _EVAL_4867;
  wire  _EVAL_4677;
  wire  _EVAL_2882;
  wire  _EVAL_395;
  wire  _EVAL_4753;
  wire  _EVAL_2069;
  wire  _EVAL_940;
  wire  _EVAL_2235;
  wire  _EVAL_3154;
  wire  _EVAL_4199;
  wire  _EVAL_2097;
  wire  _EVAL_1565;
  wire  _EVAL_3061;
  wire  _EVAL_3390;
  wire  _EVAL_5035;
  wire  _EVAL_804;
  wire  _EVAL_3768;
  wire  _EVAL_691;
  wire  _EVAL_5174;
  wire  _EVAL_2972;
  wire  _EVAL_1700;
  wire  _EVAL_958;
  wire  _EVAL_4767;
  wire  _EVAL_2979;
  wire  _EVAL_842;
  wire  _EVAL_4893;
  wire  _EVAL_2704;
  wire  _EVAL_1170;
  wire  _EVAL_2771;
  wire  _EVAL_4555;
  wire  _EVAL_4691;
  wire  _EVAL_2210;
  wire  _EVAL_4428;
  wire  _EVAL_1437;
  wire  _EVAL_570;
  wire  _EVAL_3263;
  wire  _EVAL_4627;
  wire  _EVAL_1946;
  wire  _EVAL_3949;
  wire  _EVAL_3059;
  wire  _EVAL_3717;
  wire  _EVAL_5273;
  wire  _EVAL_2177;
  wire  _EVAL_2408;
  wire  _EVAL_1935;
  wire  _EVAL_606;
  wire  _EVAL_1851;
  wire  _EVAL_1800;
  wire  _EVAL_4479;
  wire  _EVAL_2045;
  wire  _EVAL_2855;
  wire  _EVAL_3224;
  wire  _EVAL_334;
  wire  _EVAL_891;
  wire  _EVAL_5375;
  wire  _EVAL_1108;
  wire  _EVAL_823;
  wire  _EVAL_5234;
  wire  _EVAL_1977;
  wire  _EVAL_4349;
  wire  _EVAL_2530;
  wire  _EVAL_465;
  wire  _EVAL_3996;
  wire  _EVAL_1346;
  wire  _EVAL_1595;
  wire  _EVAL_1861;
  wire  _EVAL_3466;
  wire  _EVAL_1925;
  wire  _EVAL_4281;
  wire  _EVAL_3244;
  wire  _EVAL_1725;
  wire  _EVAL_1496;
  wire  _EVAL_989;
  wire  _EVAL_1989;
  wire  _EVAL_2738;
  wire [11:0] _EVAL_1363;
  wire [11:0] _EVAL_4559;
  wire [11:0] _EVAL_285;
  wire [11:0] _EVAL_4338;
  wire [11:0] _EVAL_4202;
  wire [11:0] _EVAL_3570;
  wire  _EVAL_2576;
  wire [31:0] _EVAL_5041;
  wire  _EVAL_5243;
  wire  _EVAL_4359;
  wire  _EVAL_1329;
  wire  _EVAL_3450;
  wire  _EVAL_878;
  wire  _EVAL_3890;
  wire [31:0] _EVAL_2020;
  wire [5:0] _EVAL_1701;
  wire [63:0] _EVAL_1161;
  wire  _EVAL_4772;
  wire  _EVAL_4324;
  wire  _EVAL_5216;
  wire  _EVAL_2893;
  wire  _EVAL_3237;
  wire  _EVAL_3493;
  wire  _EVAL_4628;
  wire  _EVAL_4542;
  wire  _EVAL_972;
  wire  _EVAL_4507;
  wire  _EVAL_1173;
  wire  _EVAL_3183;
  wire  _EVAL_2809;
  wire  _EVAL_4151;
  wire  _EVAL_1650;
  wire  _EVAL_4666;
  wire  _EVAL_1135;
  wire  _EVAL_282;
  wire  _EVAL_3936;
  wire  _EVAL_1592;
  wire  _EVAL_2136;
  wire  _EVAL_5279;
  wire  _EVAL_2861;
  wire  _EVAL_3722;
  wire  _EVAL_2622;
  wire  _EVAL_3055;
  wire  _EVAL_1683;
  wire  _EVAL_5369;
  wire  _EVAL_1582;
  wire  _EVAL_2614;
  wire  _EVAL_3130;
  wire  _EVAL_3751;
  wire  _EVAL_3275;
  wire  _EVAL_1239;
  wire  _EVAL_2756;
  wire  _EVAL_319;
  wire  _EVAL_1287;
  wire  _EVAL_2535;
  wire  _EVAL_5320;
  wire  _EVAL_2057;
  wire  _EVAL_2687;
  wire  _EVAL_434;
  wire  _EVAL_4597;
  wire  _EVAL_1695;
  wire  _EVAL_3341;
  wire  _EVAL_1247;
  wire  _EVAL_1209;
  wire  _EVAL_5352;
  wire  _EVAL_657;
  wire  _EVAL_3350;
  wire  _EVAL_2795;
  wire  _EVAL_2188;
  wire  _EVAL_1809;
  wire  _EVAL_3339;
  wire  _EVAL_3832;
  wire [2:0] _EVAL_2047;
  wire  _EVAL_2277;
  wire  _EVAL_3312;
  wire  _EVAL_5076;
  wire  _EVAL_4900;
  wire [4:0] _EVAL_3688;
  wire [1:0] _EVAL_2338;
  wire [1:0] _EVAL_4808;
  wire [1:0] _EVAL_1150;
  wire  _EVAL_4718;
  wire  _EVAL_4205;
  wire  _EVAL_3889;
  wire  _EVAL_3510;
  wire [1:0] _EVAL_2842;
  wire [1:0] _EVAL_5081;
  wire [1:0] _EVAL_5286;
  wire  _EVAL_2234;
  wire  _EVAL_3428;
  wire  _EVAL_5019;
  wire  _EVAL_1624;
  wire  _EVAL_3663;
  wire  _EVAL_1562;
  wire  _EVAL_5088;
  wire  _EVAL_976;
  wire  _EVAL_1014;
  wire  _EVAL_729;
  wire  _EVAL_2994;
  wire  _EVAL_3920;
  wire  _EVAL_3918;
  wire  _EVAL_4953;
  wire  _EVAL_2930;
  wire  _EVAL_5368;
  wire  _EVAL_2206;
  wire  _EVAL_3417;
  wire  _EVAL_4140;
  wire  _EVAL_817;
  wire  _EVAL_2561;
  wire  _EVAL_4166;
  wire  _EVAL_3944;
  wire  _EVAL_816;
  wire  _EVAL_4347;
  wire  _EVAL_881;
  wire  _EVAL_4216;
  wire  _EVAL_1085;
  wire  _EVAL_4845;
  wire  _EVAL_317;
  wire  _EVAL_1520;
  wire  _EVAL_1091;
  wire  _EVAL_1455;
  wire  _EVAL_2888;
  wire  _EVAL_5366;
  wire  _EVAL_2022;
  wire  _EVAL_3222;
  wire  _EVAL_4015;
  wire  _EVAL_389;
  wire  _EVAL_2821;
  wire  _EVAL_4422;
  wire  _EVAL_4463;
  wire  _EVAL_2544;
  wire  _EVAL_1518;
  wire  _EVAL_730;
  wire  _EVAL_5146;
  wire  _EVAL_736;
  wire  _EVAL_3001;
  wire  _EVAL_847;
  wire  _EVAL_2139;
  wire  _EVAL_4073;
  wire  _EVAL_1865;
  wire  _EVAL_4546;
  wire  _EVAL_2825;
  wire  _EVAL_3329;
  wire  _EVAL_3531;
  wire [31:0] _EVAL_1214;
  wire [31:0] _EVAL_4515;
  wire [31:0] _EVAL_4770;
  wire [31:0] _EVAL_872;
  wire [31:0] _EVAL_4561;
  wire [31:0] _EVAL_2412;
  wire [31:0] _EVAL_1471;
  wire [31:0] _EVAL_422;
  wire  _EVAL_2363;
  wire  _EVAL_4316;
  wire  _EVAL_2096;
  wire  _EVAL_3867;
  wire  _EVAL_4489;
  wire [1:0] _EVAL_4287;
  wire  _EVAL_906;
  wire  _EVAL_429;
  wire  _EVAL_5300;
  wire  _EVAL_4453;
  wire  _EVAL_1486;
  wire  _EVAL_3614;
  wire  _EVAL_2952;
  wire  _EVAL_2453;
  wire  _EVAL_3602;
  wire [1:0] _EVAL_307;
  wire [2:0] _EVAL_3579;
  wire  _EVAL_2981;
  wire [2:0] _EVAL_3677;
  wire  _EVAL_1627;
  wire [31:0] _EVAL_634;
  wire  _EVAL_2227;
  wire [31:0] _EVAL_2104;
  wire  _EVAL_2419;
  wire  _EVAL_3946;
  wire [31:0] _EVAL_3836;
  wire  _EVAL_2458;
  wire  _EVAL_4754;
  wire [31:0] _EVAL_1684;
  wire  _EVAL_2553;
  wire  _EVAL_3323;
  wire  _EVAL_5150;
  wire  _EVAL_5214;
  wire [31:0] _EVAL_3049;
  wire  _EVAL_502;
  wire  _EVAL_4352;
  wire [4:0] _EVAL_2980;
  wire  _EVAL_4105;
  wire  _EVAL_1802;
  wire [8:0] _EVAL_1502;
  wire [8:0] _EVAL_5372;
  wire [8:0] _EVAL_335;
  wire [8:0] _EVAL_3963;
  wire [9:0] _EVAL_1687;
  wire [2:0] _EVAL_2959;
  wire [2:0] _EVAL_3926;
  wire  _EVAL_959;
  wire  _EVAL_965;
  wire  _EVAL_721;
  wire  _EVAL_3937;
  wire [3:0] _EVAL_1553;
  wire [3:0] _EVAL_5132;
  wire  _EVAL_2155;
  wire  _EVAL_1648;
  wire  _EVAL_393;
  wire  _EVAL_3026;
  wire [1:0] _EVAL_2715;
  wire  _EVAL_471;
  wire [31:0] _EVAL_3919;
  wire  _EVAL_3882;
  wire  _EVAL_3697;
  wire  _EVAL_4233;
  wire  _EVAL_1792;
  wire  _EVAL_4964;
  wire  _EVAL_3875;
  wire  _EVAL_5169;
  wire  _EVAL_2356;
  wire  _EVAL_2272;
  wire [3:0] _EVAL_2883;
  wire [31:0] _EVAL_1798;
  wire [31:0] _EVAL_3846;
  wire [31:0] _EVAL_5027;
  wire [31:0] _EVAL_1418;
  wire  _EVAL_4569;
  wire  _EVAL_2105;
  wire  _EVAL_1269;
  wire  _EVAL_5229;
  wire  _EVAL_4782;
  wire  _EVAL_1009;
  wire  _EVAL_4261;
  wire  _EVAL_3218;
  wire  _EVAL_1817;
  wire  _EVAL_834;
  wire  _EVAL_2100;
  wire  _EVAL_4459;
  wire  _EVAL_1967;
  wire [31:0] _EVAL_561;
  wire  _EVAL_3278;
  wire  _EVAL_472;
  wire  _EVAL_1832;
  wire  _EVAL_2114;
  wire  _EVAL_418;
  wire  _EVAL_3604;
  wire  _EVAL_3007;
  wire  _EVAL_948;
  wire [31:0] _EVAL_1425;
  wire [31:0] _EVAL_5313;
  wire [31:0] _EVAL_3044;
  wire  _EVAL_4645;
  wire  _EVAL_2611;
  wire  _EVAL_3414;
  wire  _EVAL_4190;
  wire  _EVAL_995;
  wire  _EVAL_3736;
  wire  _EVAL_1597;
  wire  _EVAL_3047;
  wire  _EVAL_4176;
  wire  _EVAL_3496;
  wire [1:0] _EVAL_3649;
  wire  _EVAL_4896;
  wire  _EVAL_2996;
  wire  _EVAL_4943;
  wire  _EVAL_4389;
  wire  _EVAL_3050;
  wire  _EVAL_2676;
  wire  _EVAL_1691;
  wire  _EVAL_686;
  wire  _EVAL_646;
  wire  _EVAL_2557;
  wire  _EVAL_1982;
  wire  _EVAL_4223;
  wire [8:0] _EVAL_1889;
  wire [17:0] _EVAL_2065;
  wire [23:0] _EVAL_2864;
  wire [23:0] _EVAL_362;
  wire [5:0] _EVAL_2605;
  wire [63:0] _EVAL_3584;
  wire  _EVAL_1754;
  wire  _EVAL_3542;
  wire  _EVAL_2697;
  wire  _EVAL_2186;
  wire  _EVAL_4397;
  wire [31:0] _EVAL_1793;
  wire [31:0] _EVAL_2140;
  wire [31:0] _EVAL_2091;
  wire [31:0] _EVAL_3830;
  wire [31:0] _EVAL_3704;
  wire [1:0] _EVAL_907;
  wire [31:0] _EVAL_4430;
  wire [31:0] _EVAL_1928;
  wire  _EVAL_348;
  wire [31:0] _EVAL_5067;
  wire  _EVAL_1755;
  wire  _EVAL_1807;
  wire [31:0] _EVAL_3435;
  wire  _EVAL_4344;
  wire  _EVAL_1933;
  wire [31:0] _EVAL_2005;
  wire  _EVAL_2714;
  wire  _EVAL_3254;
  wire [31:0] _EVAL_4685;
  wire  _EVAL_3214;
  wire  _EVAL_2928;
  wire [31:0] _EVAL_1226;
  wire  _EVAL_5396;
  wire  _EVAL_2736;
  wire  _EVAL_2251;
  wire  _EVAL_1923;
  wire [31:0] _EVAL_3014;
  wire  _EVAL_4340;
  wire [31:0] _EVAL_3096;
  wire  _EVAL_2323;
  wire  _EVAL_2083;
  wire  _EVAL_1421;
  wire  _EVAL_5342;
  wire [31:0] _EVAL_3762;
  wire  _EVAL_2294;
  wire  _EVAL_3554;
  wire [31:0] _EVAL_4267;
  wire  _EVAL_2907;
  wire  _EVAL_536;
  wire [31:0] _EVAL_835;
  wire  _EVAL_2267;
  wire  _EVAL_785;
  wire  _EVAL_1332;
  wire [31:0] _EVAL_5331;
  wire  _EVAL_4304;
  wire [31:0] _EVAL_4275;
  wire  _EVAL_604;
  wire  _EVAL_410;
  wire  _EVAL_4128;
  wire [31:0] _EVAL_2957;
  wire  _EVAL_5294;
  wire  _EVAL_2444;
  wire  _EVAL_3465;
  wire  _EVAL_3868;
  wire [31:0] _EVAL_1419;
  wire  _EVAL_4081;
  wire  _EVAL_4647;
  wire [4:0] _EVAL_3765;
  wire  _EVAL_2754;
  wire  _EVAL_3744;
  wire [31:0] _EVAL_1964;
  wire  _EVAL_4610;
  wire  _EVAL_3721;
  wire [4:0] _EVAL_5405;
  wire  _EVAL_3289;
  wire  _EVAL_2123;
  wire  _EVAL_800;
  wire  _EVAL_1185;
  wire  _EVAL_692;
  wire [4:0] _EVAL_3558;
  wire [4:0] _EVAL_5153;
  wire [4:0] _EVAL_4611;
  wire [4:0] _EVAL_4179;
  wire [4:0] _EVAL_1443;
  wire  _EVAL_2366;
  wire  _EVAL_4673;
  wire [18:0] _EVAL_1730;
  wire [31:0] _EVAL_5128;
  wire [31:0] _EVAL_2701;
  wire  _EVAL_1736;
  wire  _EVAL_3969;
  wire [7:0] _EVAL_2489;
  wire [9:0] _EVAL_4425;
  wire [20:0] _EVAL_2641;
  wire [20:0] _EVAL_1991;
  wire [20:0] _EVAL_1674;
  wire  _EVAL_1688;
  wire [10:0] _EVAL_1390;
  wire [31:0] _EVAL_3981;
  wire [31:0] _EVAL_672;
  wire [31:0] _EVAL_407;
  wire  _EVAL_455;
  wire  _EVAL_2500;
  wire [19:0] _EVAL_3288;
  wire [31:0] _EVAL_326;
  wire [31:0] _EVAL_3021;
  wire [31:0] _EVAL_3095;
  wire  _EVAL_4602;
  wire  _EVAL_3080;
  wire  _EVAL_3583;
  wire  _EVAL_583;
  wire [11:0] _EVAL_2048;
  wire  _EVAL_4800;
  wire [19:0] _EVAL_1978;
  wire [31:0] _EVAL_1765;
  wire [31:0] _EVAL_4232;
  wire [31:0] _EVAL_1886;
  wire  _EVAL_1344;
  wire  _EVAL_683;
  wire  _EVAL_5179;
  wire  _EVAL_3042;
  wire  _EVAL_2081;
  wire [31:0] _EVAL_1464;
  wire [31:0] _EVAL_514;
  wire [31:0] _EVAL_4929;
  wire [31:0] _EVAL_4744;
  wire [31:0] _EVAL_2029;
  wire [31:0] _EVAL_2194;
  wire  _EVAL_4174;
  wire  _EVAL_3609;
  wire  _EVAL_1656;
  wire  _EVAL_4417;
  wire [31:0] _EVAL_3197;
  wire [31:0] _EVAL_3695;
  wire [31:0] _EVAL_425;
  wire [31:0] _EVAL_481;
  wire [31:0] _EVAL_2933;
  wire  _EVAL_2425;
  wire  _EVAL_4734;
  wire  _EVAL_3662;
  wire  _EVAL_3074;
  wire  _EVAL_2632;
  wire  _EVAL_749;
  wire [31:0] _EVAL_4709;
  wire  _EVAL_3078;
  wire  _EVAL_3630;
  wire  _EVAL_1025;
  wire  _EVAL_3345;
  wire  _EVAL_2377;
  wire  _EVAL_2184;
  wire [5:0] _EVAL_5045;
  wire [63:0] _EVAL_5403;
  wire  _EVAL_3921;
  wire  _EVAL_4337;
  wire  _EVAL_4310;
  wire  _EVAL_2292;
  wire  _EVAL_337;
  wire  _EVAL_1459;
  wire  _EVAL_1199;
  wire  _EVAL_1056;
  wire  _EVAL_4657;
  wire  _EVAL_1395;
  wire  _EVAL_3576;
  wire  _EVAL_2165;
  wire  _EVAL_3287;
  wire  _EVAL_2311;
  wire  _EVAL_2410;
  wire  _EVAL_3152;
  wire  _EVAL_4478;
  wire  _EVAL_3097;
  wire  _EVAL_4346;
  wire  _EVAL_3267;
  wire  _EVAL_2398;
  wire  _EVAL_2539;
  wire  _EVAL_3235;
  wire  _EVAL_5160;
  wire  _EVAL_1204;
  wire  _EVAL_1176;
  wire  _EVAL_2402;
  wire  _EVAL_950;
  wire  _EVAL_2017;
  wire  _EVAL_2168;
  wire  _EVAL_1360;
  wire  _EVAL_824;
  wire  _EVAL_1846;
  wire  _EVAL_2479;
  wire  _EVAL_4285;
  wire  _EVAL_5251;
  wire  _EVAL_2905;
  wire  _EVAL_3380;
  wire  _EVAL_2708;
  wire  _EVAL_3013;
  wire  _EVAL_4815;
  wire  _EVAL_855;
  wire  _EVAL_2881;
  wire  _EVAL_1118;
  wire  _EVAL_1115;
  wire [4:0] _EVAL_2117;
  wire  _EVAL_4074;
  wire  _EVAL_5008;
  wire  _EVAL_1055;
  wire  _EVAL_1664;
  wire [1:0] _EVAL_2154;
  wire [2:0] _EVAL_4913;
  wire [3:0] _EVAL_1045;
  wire [3:0] _EVAL_3826;
  wire [2:0] _EVAL_4603;
  wire [3:0] _EVAL_1202;
  wire [3:0] _EVAL_3543;
  wire [31:0] _EVAL_4642;
  wire [31:0] _EVAL_1834;
  wire  _EVAL_5306;
  wire  _EVAL_2681;
  wire  _EVAL_2342;
  wire  _EVAL_506;
  wire  _EVAL_2040;
  wire  _EVAL_5154;
  wire  _EVAL_2709;
  wire  _EVAL_5239;
  wire  _EVAL_5133;
  wire  _EVAL_2122;
  wire  _EVAL_716;
  wire  _EVAL_4435;
  wire  _EVAL_3052;
  wire  _EVAL_3520;
  wire [11:0] _EVAL_5341;
  wire [11:0] _EVAL_1462;
  wire [11:0] _EVAL_2450;
  wire  _EVAL_5050;
  wire [19:0] _EVAL_833;
  wire [31:0] _EVAL_4472;
  wire [31:0] _EVAL_4333;
  wire  _EVAL_4960;
  wire  _EVAL_3434;
  wire  _EVAL_4882;
  wire [31:0] _EVAL_2153;
  wire [31:0] _EVAL_1152;
  wire [31:0] _EVAL_4041;
  wire [31:0] _EVAL_2351;
  wire [31:0] _EVAL_944;
  wire [31:0] _EVAL_4967;
  wire [6:0] _EVAL_2546;
  wire [127:0] _EVAL_297;
  wire [127:0] _EVAL_5349;
  wire  _EVAL_1943;
  wire  _EVAL_1248;
  wire  _EVAL_3319;
  wire  _EVAL_3073;
  wire  _EVAL_4079;
  wire  _EVAL_4106;
  wire  _EVAL_3259;
  wire [3:0] _EVAL_985;
  wire [3:0] _EVAL_1466;
  wire  _EVAL_655;
  wire  _EVAL_3571;
  wire  _EVAL_1411;
  wire  _EVAL_4217;
  wire  _EVAL_497;
  wire  _EVAL_3844;
  wire  _EVAL_4689;
  wire [3:0] _EVAL_2852;
  wire [31:0] _EVAL_420;
  wire [31:0] _EVAL_368;
  wire [31:0] _EVAL_4533;
  wire [31:0] _EVAL_1368;
  wire  _EVAL_2082;
  wire  _EVAL_2036;
  wire  _EVAL_2575;
  wire  _EVAL_1222;
  wire [1:0] _EVAL_2879;
  wire  _EVAL_5259;
  wire  _EVAL_394;
  wire  _EVAL_947;
  wire [2:0] _EVAL_1038;
  wire [2:0] _EVAL_4291;
  wire [5:0] _EVAL_4075;
  wire [22:0] _EVAL_3606;
  wire [32:0] _EVAL_1004;
  wire  _EVAL_3732;
  wire [2:0] _EVAL_625;
  wire [2:0] _EVAL_2035;
  wire  _EVAL_2661;
  wire  _EVAL_2787;
  wire  _EVAL_5173;
  wire  _EVAL_2286;
  wire  _EVAL_5384;
  wire  _EVAL_4932;
  wire  _EVAL_1153;
  wire  _EVAL_1238;
  wire [12:0] _EVAL_2841;
  wire [1:0] _EVAL_1883;
  wire  _EVAL_1602;
  wire  _EVAL_3795;
  wire  _EVAL_4133;
  wire  _EVAL_2445;
  wire  _EVAL_4356;
  wire  _EVAL_4132;
  wire  _EVAL_1579;
  wire [3:0] _EVAL_4700;
  wire  _EVAL_5136;
  wire [31:0] _EVAL_3693;
  wire [31:0] _EVAL_4601;
  wire  _EVAL_5388;
  wire  _EVAL_5171;
  wire  _EVAL_4236;
  wire  _EVAL_3032;
  wire [31:0] _EVAL_1454;
  wire  _EVAL_292;
  wire  _EVAL_414;
  wire  _EVAL_4165;
  wire [31:0] _EVAL_1316;
  wire  _EVAL_1907;
  wire  _EVAL_2232;
  wire [31:0] _EVAL_1738;
  wire  _EVAL_4314;
  wire  _EVAL_5109;
  wire [31:0] _EVAL_2043;
  wire  _EVAL_1622;
  wire  _EVAL_3553;
  wire  _EVAL_3433;
  wire  _EVAL_582;
  wire [31:0] _EVAL_4884;
  wire  _EVAL_2760;
  wire [31:0] _EVAL_3332;
  wire  _EVAL_4253;
  wire  _EVAL_4332;
  wire [31:0] _EVAL_3479;
  wire  _EVAL_3388;
  wire  _EVAL_2312;
  wire [31:0] _EVAL_1456;
  wire  _EVAL_3563;
  wire  _EVAL_1814;
  wire [31:0] _EVAL_371;
  wire  _EVAL_1689;
  wire  _EVAL_3371;
  wire [31:0] _EVAL_2024;
  wire  _EVAL_4096;
  wire  _EVAL_5014;
  wire  _EVAL_1538;
  wire  _EVAL_1867;
  wire [31:0] _EVAL_4797;
  wire  _EVAL_4107;
  wire [31:0] _EVAL_4631;
  wire  _EVAL_4738;
  wire  _EVAL_4618;
  wire [31:0] _EVAL_860;
  wire  _EVAL_1195;
  wire  _EVAL_549;
  wire  _EVAL_892;
  wire  _EVAL_4652;
  wire [31:0] _EVAL_4090;
  wire  _EVAL_5149;
  wire  _EVAL_2220;
  wire  _EVAL_1359;
  wire  _EVAL_916;
  wire  _EVAL_2465;
  wire  _EVAL_5371;
  wire  _EVAL_3611;
  wire  _EVAL_1207;
  wire  _EVAL_1942;
  wire  _EVAL_4002;
  wire  _EVAL_5404;
  wire  _EVAL_1051;
  wire  _EVAL_2370;
  wire  _EVAL_2496;
  wire  _EVAL_1871;
  wire  _EVAL_2291;
  wire [31:0] _EVAL_4956;
  wire [31:0] _EVAL_1087;
  wire [31:0] _EVAL_3449;
  wire [31:0] _EVAL_5001;
  wire  _EVAL_1829;
  wire  _EVAL_2269;
  wire  _EVAL_1277;
  wire  _EVAL_2112;
  wire [2:0] _EVAL_2352;
  wire [3:0] _EVAL_3219;
  wire  _EVAL_3819;
  wire  _EVAL_1463;
  wire [2:0] _EVAL_4436;
  wire  _EVAL_3958;
  wire [31:0] _EVAL_2711;
  wire  _EVAL_534;
  wire  _EVAL_3592;
  wire  _EVAL_2767;
  wire [1:0] _EVAL_728;
  wire  _EVAL_3445;
  wire  _EVAL_3398;
  wire  _EVAL_2067;
  wire [3:0] _EVAL_372;
  wire  _EVAL_1904;
  wire  _EVAL_4955;
  wire [2:0] _EVAL_2974;
  wire [3:0] _EVAL_3002;
  wire [3:0] _EVAL_5406;
  wire [2:0] _EVAL_1453;
  wire [3:0] _EVAL_3794;
  wire [3:0] _EVAL_2690;
  wire [12:0] _EVAL_2862;
  wire  _EVAL_3022;
  wire  _EVAL_4130;
  wire  _EVAL_1216;
  wire  _EVAL_3260;
  wire  _EVAL_1157;
  wire  _EVAL_3459;
  wire  _EVAL_1398;
  wire  _EVAL_3009;
  wire [28:0] _EVAL_5230;
  wire  _EVAL_1601;
  wire  _EVAL_996;
  wire  _EVAL_3818;
  wire  _EVAL_3597;
  wire  _EVAL_3361;
  wire  _EVAL_2740;
  wire  _EVAL_1380;
  wire  _EVAL_486;
  wire  _EVAL_2945;
  wire  _EVAL_4944;
  wire  _EVAL_1504;
  wire  _EVAL_1181;
  wire  _EVAL_325;
  wire  _EVAL_2921;
  wire  _EVAL_839;
  wire  _EVAL_5068;
  wire [1:0] _EVAL_359;
  wire  _EVAL_5260;
  wire  _EVAL_3517;
  wire  _EVAL_4475;
  wire  _EVAL_4365;
  wire  _EVAL_5275;
  wire  _EVAL_283;
  wire  _EVAL_4270;
  wire  _EVAL_4025;
  wire  _EVAL_4534;
  wire  _EVAL_5175;
  wire  _EVAL_1705;
  wire  _EVAL_565;
  wire  _EVAL_569;
  wire  _EVAL_5123;
  wire  _EVAL_1589;
  wire [15:0] _EVAL_1526;
  wire [15:0] _EVAL_477;
  wire [31:0] _EVAL_4256;
  wire  _EVAL_1860;
  wire  _EVAL_3301;
  wire  _EVAL_1082;
  wire  _EVAL_4301;
  wire  _EVAL_1326;
  wire  _EVAL_1536;
  wire  _EVAL_934;
  wire  _EVAL_2250;
  wire  _EVAL_4118;
  wire  _EVAL_5152;
  wire  _EVAL_3297;
  wire  _EVAL_2466;
  wire  _EVAL_3513;
  wire  _EVAL_1561;
  wire  _EVAL_2664;
  wire  _EVAL_4560;
  wire  _EVAL_3285;
  wire  _EVAL_4409;
  wire  _EVAL_2566;
  wire  _EVAL_1788;
  wire  _EVAL_3011;
  wire  _EVAL_4393;
  wire [31:0] _EVAL_2092;
  wire  _EVAL_5358;
  wire  _EVAL_2999;
  wire  _EVAL_2451;
  wire  _EVAL_3153;
  wire  _EVAL_3675;
  wire  _EVAL_2534;
  wire  _EVAL_1389;
  wire  _EVAL_2147;
  wire  _EVAL_5155;
  wire  _EVAL_670;
  wire  _EVAL_3582;
  wire  _EVAL_3903;
  wire  _EVAL_4928;
  wire  _EVAL_734;
  wire  _EVAL_2011;
  wire  _EVAL_1137;
  wire  _EVAL_3491;
  wire  _EVAL_1585;
  wire  _EVAL_4875;
  wire  _EVAL_399;
  wire  _EVAL_756;
  wire  _EVAL_1461;
  wire  _EVAL_3757;
  wire  _EVAL_3121;
  wire  _EVAL_4980;
  wire  _EVAL_697;
  wire  _EVAL_1750;
  wire  _EVAL_2205;
  wire  _EVAL_3539;
  wire  _EVAL_1612;
  wire  _EVAL_3292;
  wire  _EVAL_3863;
  wire  _EVAL_1381;
  wire  _EVAL_1249;
  wire  _EVAL_329;
  wire  _EVAL_3815;
  wire  _EVAL_1309;
  wire  _EVAL_1539;
  wire  _EVAL_4194;
  wire  _EVAL_2299;
  wire  _EVAL_2379;
  wire  _EVAL_4225;
  wire  _EVAL_2510;
  wire  _EVAL_4573;
  wire  _EVAL_4788;
  wire  _EVAL_539;
  wire  _EVAL_2001;
  wire  _EVAL_2508;
  wire  _EVAL_1013;
  wire  _EVAL_4827;
  wire  _EVAL_3587;
  wire  _EVAL_2239;
  wire  _EVAL_1124;
  wire  _EVAL_4701;
  wire  _EVAL_1770;
  wire  _EVAL_3725;
  wire [4:0] _EVAL_3201;
  wire [4:0] _EVAL_5277;
  wire [4:0] _EVAL_3321;
  wire [5:0] _EVAL_3070;
  wire [23:0] _EVAL_701;
  wire  _EVAL_2354;
  wire [4:0] _EVAL_3112;
  wire  _EVAL_3873;
  wire  _EVAL_4671;
  wire  _EVAL_4005;
  wire  _EVAL_1840;
  wire [8:0] _EVAL_3973;
  wire  _EVAL_1734;
  wire  _EVAL_4300;
  wire  _EVAL_1862;
  wire  _EVAL_4491;
  wire  _EVAL_4908;
  wire  _EVAL_3216;
  wire  _EVAL_3731;
  wire  _EVAL_5311;
  wire  _EVAL_4639;
  wire  _EVAL_810;
  wire  _EVAL_4902;
  wire  _EVAL_635;
  wire  _EVAL_2967;
  wire  _EVAL_4297;
  wire  _EVAL_2913;
  wire  _EVAL_609;
  wire  _EVAL_402;
  wire  _EVAL_4831;
  wire  _EVAL_1392;
  wire  _EVAL_2507;
  wire  _EVAL_1460;
  wire  _EVAL_1747;
  wire  _EVAL_5399;
  wire  _EVAL_4372;
  wire  _EVAL_4914;
  wire  _EVAL_559;
  wire  _EVAL_4272;
  wire  _EVAL_1402;
  wire [4:0] _EVAL_2343;
  wire [4:0] _EVAL_3333;
  wire [1:0] _EVAL_5278;
  wire  _EVAL_2840;
  wire  _EVAL_4802;
  wire [4:0] _EVAL_1610;
  wire  _EVAL_4783;
  wire  _EVAL_1052;
  wire [31:0] _EVAL_4690;
  wire [31:0] _EVAL_1223;
  wire  _EVAL_2275;
  wire  _EVAL_1874;
  wire [2:0] _EVAL_5418;
  wire [3:0] _EVAL_953;
  wire [3:0] _EVAL_4743;
  wire [3:0] _EVAL_2189;
  wire [3:0] _EVAL_2493;
  wire  _EVAL_3313;
  wire  _EVAL_4011;
  wire [4:0] _EVAL_5084;
  wire  _EVAL_3955;
  wire  _EVAL_3900;
  wire  _EVAL_4959;
  wire  _EVAL_5059;
  wire  _EVAL_893;
  wire  _EVAL_1763;
  wire  _EVAL_617;
  wire  _EVAL_3784;
  wire  _EVAL_3020;
  wire  _EVAL_1522;
  wire  _EVAL_2428;
  wire  _EVAL_1200;
  wire  _EVAL_1191;
  wire  _EVAL_2591;
  wire  _EVAL_526;
  wire  _EVAL_2975;
  wire  _EVAL_3367;
  wire  _EVAL_4387;
  wire  _EVAL_1976;
  wire  _EVAL_2706;
  wire  _EVAL_3620;
  wire  _EVAL_4540;
  wire  _EVAL_1947;
  wire  _EVAL_4414;
  wire  _EVAL_3392;
  wire  _EVAL_3933;
  wire  _EVAL_398;
  wire  _EVAL_885;
  wire  _EVAL_2469;
  wire  _EVAL_1629;
  wire  _EVAL_1341;
  wire  _EVAL_3764;
  wire  _EVAL_3242;
  wire  _EVAL_2511;
  wire  _EVAL_3376;
  wire  _EVAL_726;
  wire  _EVAL_406;
  wire  _EVAL_973;
  wire  _EVAL_4242;
  wire  _EVAL_1261;
  wire  _EVAL_2308;
  wire  _EVAL_1259;
  wire  _EVAL_1189;
  wire  _EVAL_4189;
  wire  _EVAL_4415;
  wire  _EVAL_4125;
  wire  _EVAL_2541;
  wire [17:0] _EVAL_5070;
  wire  _EVAL_5422;
  wire [2:0] _EVAL_318;
  wire  _EVAL_1340;
  wire  _EVAL_2851;
  wire  _EVAL_454;
  wire [1:0] _EVAL_1305;
  wire  _EVAL_401;
  wire  _EVAL_4653;
  wire  _EVAL_4851;
  wire  _EVAL_1236;
  wire  _EVAL_4931;
  wire  _EVAL_753;
  wire  _EVAL_1660;
  wire  _EVAL_4465;
  wire  _EVAL_2604;
  wire  _EVAL_2415;
  wire [11:0] _EVAL_3610;
  wire  _EVAL_1948;
  wire [11:0] _EVAL_1370;
  wire  _EVAL_2087;
  wire  _EVAL_2543;
  wire  _EVAL_4926;
  wire [4:0] _EVAL_3023;
  wire  _EVAL_1531;
  wire  _EVAL_2581;
  wire  _EVAL_2554;
  wire  _EVAL_487;
  wire [2:0] _EVAL_3325;
  wire [2:0] _EVAL_3931;
  wire  _EVAL_1794;
  wire  _EVAL_595;
  wire  _EVAL_2805;
  wire  _EVAL_687;
  wire  _EVAL_843;
  wire  _EVAL_3502;
  wire  _EVAL_4825;
  wire  _EVAL_543;
  wire  _EVAL_788;
  wire  _EVAL_1508;
  wire  _EVAL_1548;
  wire  _EVAL_5221;
  wire  _EVAL_888;
  wire  _EVAL_5060;
  wire  _EVAL_4905;
  wire  _EVAL_2088;
  wire  _EVAL_3305;
  wire  _EVAL_1074;
  wire  _EVAL_3076;
  wire [2:0] _EVAL_4146;
  wire  _EVAL_3334;
  wire [2:0] _EVAL_1953;
  wire [2:0] _EVAL_2536;
  wire  _EVAL_4532;
  wire  _EVAL_2555;
  wire  _EVAL_4670;
  wire  _EVAL_5188;
  wire  _EVAL_1282;
  wire  _EVAL_4575;
  wire  _EVAL_2722;
  wire  _EVAL_2062;
  wire  _EVAL_3975;
  wire  _EVAL_3984;
  wire  _EVAL_5270;
  wire  _EVAL_1470;
  wire  _EVAL_541;
  wire  _EVAL_4345;
  wire  _EVAL_3382;
  wire  _EVAL_912;
  wire  _EVAL_4363;
  wire  _EVAL_883;
  wire  _EVAL_3358;
  wire  _EVAL_2187;
  wire  _EVAL_2941;
  wire  _EVAL_360;
  wire  _EVAL_1210;
  wire  _EVAL_2171;
  wire  _EVAL_4143;
  wire  _EVAL_3369;
  wire  _EVAL_3488;
  wire  _EVAL_2589;
  wire  _EVAL_846;
  wire [3:0] _EVAL_4077;
  wire [3:0] _EVAL_2375;
  wire [1:0] _EVAL_4246;
  wire  _EVAL_4860;
  wire  _EVAL_1757;
  wire  _EVAL_4979;
  wire  _EVAL_2559;
  wire  _EVAL_2961;
  wire  _EVAL_4378;
  wire  _EVAL_3194;
  wire [63:0] _EVAL_4379;
  wire [63:0] _EVAL_3127;
  wire  _EVAL_4149;
  wire  _EVAL_5121;
  wire [11:0] _EVAL_3400;
  wire [2:0] _EVAL_2849;
  wire  _EVAL_3829;
  wire  _EVAL_2698;
  wire  _EVAL_5416;
  wire  _EVAL_2870;
  wire  _EVAL_4523;
  wire  _EVAL_1493;
  wire [31:0] _EVAL_1076;
  wire [31:0] _EVAL_4482;
  wire [31:0] _EVAL_4444;
  wire [31:0] _EVAL_955;
  wire  _EVAL_4906;
  wire [2:0] _EVAL_1037;
  wire [1:0] _EVAL_3692;
  wire [2:0] _EVAL_509;
  wire  _EVAL_566;
  wire  _EVAL_333;
  wire  _EVAL_4188;
  wire  _EVAL_2909;
  wire [2:0] _EVAL_5400;
  wire [2:0] _EVAL_4837;
  wire  _EVAL_4145;
  wire  _EVAL_3685;
  wire  _EVAL_4213;
  wire  _EVAL_5296;
  wire  _EVAL_1438;
  wire  _EVAL_2396;
  wire  _EVAL_1771;
  wire  _EVAL_1637;
  wire  _EVAL_3427;
  wire [7:0] _EVAL_2470;
  wire [7:0] _EVAL_4785;
  wire [7:0] _EVAL_5139;
  wire [24:0] _EVAL_1043;
  wire [23:0] _EVAL_466;
  wire [4:0] _EVAL_3770;
  wire [4:0] _EVAL_5343;
  wire [23:0] _EVAL_4501;
  wire [22:0] _EVAL_2675;
  wire [22:0] _EVAL_1796;
  wire [22:0] _EVAL_1751;
  wire [22:0] _EVAL_3899;
  wire [31:0] _EVAL_4035;
  wire  _EVAL_3791;
  wire  _EVAL_1072;
  wire  _EVAL_5357;
  wire  _EVAL_4094;
  wire [1:0] _EVAL_1394;
  wire  _EVAL_306;
  wire  _EVAL_2834;
  wire  _EVAL_4830;
  wire  _EVAL_1151;
  wire  _EVAL_3861;
  wire  _EVAL_3018;
  wire  _EVAL_4704;
  wire  _EVAL_1289;
  wire [1:0] _EVAL_2304;
  wire  _EVAL_1361;
  wire  _EVAL_4556;
  wire  _EVAL_2169;
  wire  _EVAL_3816;
  wire  _EVAL_4108;
  wire  _EVAL_1284;
  wire  _EVAL_939;
  wire  _EVAL_4102;
  wire  _EVAL_3469;
  wire  _EVAL_3006;
  wire  _EVAL_3690;
  wire  _EVAL_2887;
  wire  _EVAL_4997;
  wire  _EVAL_5096;
  wire  _EVAL_2191;
  wire  _EVAL_999;
  wire  _EVAL_3280;
  wire  _EVAL_493;
  wire  _EVAL_3824;
  wire  _EVAL_3306;
  wire  _EVAL_4940;
  wire  _EVAL_5012;
  wire  _EVAL_4296;
  wire  _EVAL_328;
  wire  _EVAL_5280;
  wire  _EVAL_802;
  wire  _EVAL_3098;
  wire [4:0] _EVAL_2093;
  wire [4:0] _EVAL_3320;
  wire [4:0] _EVAL_2729;
  wire [4:0] _EVAL_3067;
  wire [4:0] _EVAL_1339;
  wire [4:0] _EVAL_4635;
  wire [4:0] _EVAL_5228;
  wire [4:0] _EVAL_3110;
  wire  _EVAL_3489;
  wire  _EVAL_684;
  wire [63:0] _EVAL_4629;
  wire [11:0] _EVAL_2223;
  wire [11:0] _EVAL_1435;
  wire  _EVAL_4762;
  wire  _EVAL_2300;
  wire  _EVAL_3537;
  wire  _EVAL_1050;
  wire  _EVAL_3483;
  wire  _EVAL_1506;
  wire  _EVAL_4950;
  wire  _EVAL_5410;
  wire  _EVAL_5037;
  wire  _EVAL_288;
  wire  _EVAL_3735;
  wire  _EVAL_4508;
  wire  _EVAL_4740;
  wire  _EVAL_2218;
  wire  _EVAL_3429;
  wire  _EVAL_1820;
  wire  _EVAL_3407;
  wire [32:0] _EVAL_3560;
  wire [32:0] _EVAL_1148;
  wire [32:0] _EVAL_2570;
  wire  _EVAL_2590;
  wire [31:0] _EVAL_4083;
  wire  _EVAL_1955;
  wire  _EVAL_4484;
  wire  _EVAL_3914;
  wire  _EVAL_353;
  wire  _EVAL_921;
  wire  _EVAL_4010;
  wire  _EVAL_2086;
  wire  _EVAL_4667;
  wire  _EVAL_2181;
  wire [4:0] _EVAL_4606;
  wire [2:0] _EVAL_4703;
  wire  _EVAL_4080;
  wire  _EVAL_5235;
  wire  _EVAL_3793;
  wire  _EVAL_2426;
  wire [31:0] _EVAL_4589;
  wire [31:0] _EVAL_3848;
  wire  _EVAL_2982;
  wire  _EVAL_915;
  wire  _EVAL_1760;
  wire  _EVAL_433;
  wire  _EVAL_3307;
  wire  _EVAL_4519;
  wire [2:0] _EVAL_4219;
  wire [3:0] _EVAL_3569;
  wire [3:0] _EVAL_3418;
  wire  _EVAL_1080;
  wire [3:0] _EVAL_5029;
  wire [3:0] _EVAL_378;
  wire [3:0] _EVAL_4385;
  wire [31:0] _EVAL_4053;
  wire [31:0] _EVAL_341;
  wire [31:0] _EVAL_1026;
  wire [31:0] _EVAL_4761;
  wire [32:0] _EVAL_4548;
  wire [32:0] _EVAL_3024;
  wire [32:0] _EVAL_3625;
  wire [31:0] _EVAL_5397;
  wire  _EVAL_3342;
  wire  _EVAL_4829;
  wire [31:0] _EVAL_1175;
  wire [31:0] _EVAL_5000;
  wire [31:0] _EVAL_489;
  wire [31:0] _EVAL_4733;
  wire [31:0] _EVAL_5364;
  wire  _EVAL_379;
  wire  _EVAL_2503;
  wire  _EVAL_2307;
  wire  _EVAL_5105;
  wire  _EVAL_832;
  wire  _EVAL_3236;
  wire  _EVAL_2860;
  wire  _EVAL_1384;
  wire  _EVAL_4308;
  wire  _EVAL_680;
  wire  _EVAL_4725;
  wire  _EVAL_2107;
  wire  _EVAL_1482;
  wire [19:0] _EVAL_4462;
  wire [19:0] _EVAL_1787;
  wire  _EVAL_5312;
  wire  _EVAL_1779;
  wire  _EVAL_4858;
  wire [11:0] _EVAL_1107;
  wire  _EVAL_3877;
  wire [19:0] _EVAL_3472;
  wire [31:0] _EVAL_1121;
  wire [31:0] _EVAL_2533;
  wire  _EVAL_1852;
  wire  _EVAL_5108;
  wire  _EVAL_2820;
  wire  _EVAL_573;
  wire  _EVAL_4773;
  wire  _EVAL_845;
  wire  _EVAL_2800;
  wire  _EVAL_5272;
  wire  _EVAL_957;
  wire  _EVAL_460;
  wire  _EVAL_4543;
  wire  _EVAL_2486;
  wire  _EVAL_819;
  wire  _EVAL_4693;
  wire  _EVAL_5249;
  wire  _EVAL_1034;
  wire  _EVAL_4638;
  wire [4:0] _EVAL_4070;
  wire [10:0] _EVAL_2613;
  wire [23:0] _EVAL_2645;
  wire  _EVAL_437;
  wire  _EVAL_1744;
  wire [32:0] _EVAL_3536;
  wire  _EVAL_2835;
  wire  _EVAL_1321;
  wire  _EVAL_3375;
  wire  _EVAL_4062;
  wire  _EVAL_4375;
  wire  _EVAL_1613;
  wire  _EVAL_2103;
  wire  _EVAL_510;
  wire [31:0] _EVAL_3805;
  wire [31:0] _EVAL_4290;
  wire [31:0] _EVAL_1931;
  wire [4:0] _EVAL_535;
  wire  _EVAL_2776;
  wire [31:0] _EVAL_3249;
  wire  _EVAL_3748;
  wire  _EVAL_1403;
  wire  _EVAL_4022;
  wire  _EVAL_4919;
  wire  _EVAL_4440;
  wire  _EVAL_1786;
  wire [3:0] _EVAL_5011;
  wire  _EVAL_1163;
  wire [1:0] _EVAL_1845;
  wire [3:0] _EVAL_4975;
  wire [3:0] _EVAL_5211;
  wire [3:0] _EVAL_1903;
  wire  _EVAL_651;
  wire  _EVAL_4027;
  wire  _EVAL_5100;
  wire [19:0] _EVAL_3090;
  wire [31:0] _EVAL_4224;
  wire [31:0] _EVAL_5073;
  wire [31:0] _EVAL_831;
  wire  _EVAL_2175;
  wire [31:0] _EVAL_829;
  wire [31:0] _EVAL_1938;
  wire [31:0] _EVAL_4442;
  wire  _EVAL_528;
  wire [4:0] _EVAL_3708;
  wire [4:0] _EVAL_2178;
  wire [4:0] _EVAL_3574;
  wire [4:0] _EVAL_4370;
  wire  _EVAL_990;
  wire [4:0] _EVAL_1095;
  wire  _EVAL_4354;
  wire  _EVAL_3821;
  wire [1:0] _EVAL_5253;
  wire  _EVAL_4367;
  wire  _EVAL_5276;
  wire  _EVAL_4994;
  wire  _EVAL_392;
  wire  _EVAL_1716;
  wire  _EVAL_4553;
  wire  _EVAL_5074;
  wire [1:0] _EVAL_674;
  wire  _EVAL_1826;
  wire  _EVAL_1678;
  wire  _EVAL_2962;
  wire  _EVAL_1433;
  wire  _EVAL_1733;
  wire  _EVAL_1169;
  wire  _EVAL_4003;
  wire  _EVAL_3548;
  wire [31:0] _EVAL_4251;
  wire  _EVAL_516;
  wire  _EVAL_2098;
  wire  _EVAL_3425;
  wire [1:0] _EVAL_3395;
  wire [1:0] _EVAL_2572;
  wire  _EVAL_2832;
  wire [23:0] _EVAL_530;
  wire  _EVAL_511;
  wire  _EVAL_4269;
  wire  _EVAL_5207;
  wire  _EVAL_4735;
  wire [31:0] _EVAL_3775;
  wire [31:0] _EVAL_3169;
  wire  _EVAL_4581;
  wire  _EVAL_3865;
  wire  _EVAL_669;
  wire  _EVAL_2563;
  wire  _EVAL_1268;
  wire  _EVAL_3987;
  wire  _EVAL_1875;
  wire  _EVAL_2405;
  wire [2:0] _EVAL_447;
  wire [3:0] _EVAL_1918;
  wire [3:0] _EVAL_4277;
  wire [2:0] _EVAL_867;
  wire [3:0] _EVAL_1959;
  wire  _EVAL_4142;
  wire  _EVAL_928;
  wire  _EVAL_619;
  wire  _EVAL_2050;
  wire  _EVAL_5209;
  wire  _EVAL_1423;
  wire [4:0] _EVAL_4836;
  wire [4:0] _EVAL_894;
  wire [4:0] _EVAL_919;
  wire [4:0] _EVAL_2836;
  wire [4:0] _EVAL_3225;
  wire  _EVAL_908;
  wire  _EVAL_456;
  wire [31:0] _EVAL_3477;
  wire  _EVAL_383;
  wire  _EVAL_4343;
  wire  _EVAL_931;
  wire  _EVAL_2384;
  wire [1:0] _EVAL_4063;
  wire [4:0] _EVAL_1201;
  wire  _EVAL_301;
  wire  _EVAL_4148;
  wire  _EVAL_365;
  wire  _EVAL_2658;
  wire  _EVAL_4759;
  wire  _EVAL_3518;
  wire  _EVAL_3925;
  wire  _EVAL_2297;
  wire  _EVAL_859;
  wire  _EVAL_1939;
  wire  _EVAL_1174;
  wire  _EVAL_1186;
  wire [23:0] _EVAL_339;
  wire  _EVAL_1130;
  wire [32:0] _EVAL_1574;
  wire [31:0] _EVAL_2772;
  wire  _EVAL_5285;
  wire  _EVAL_673;
  wire  _EVAL_439;
  wire  _EVAL_1835;
  wire [32:0] _EVAL_1773;
  wire [32:0] _EVAL_3122;
  wire [32:0] _EVAL_4758;
  wire  _EVAL_1876;
  wire  _EVAL_5051;
  wire  _EVAL_633;
  wire  _EVAL_767;
  wire  _EVAL_3706;
  wire  _EVAL_4883;
  wire  _EVAL_4636;
  wire  _EVAL_1652;
  wire  _EVAL_1732;
  wire  _EVAL_3621;
  wire  _EVAL_4567;
  wire  _EVAL_2548;
  wire  _EVAL_3994;
  wire  _EVAL_4732;
  wire  _EVAL_3045;
  wire  _EVAL_5057;
  wire  _EVAL_4402;
  wire  _EVAL_2494;
  wire  _EVAL_4355;
  wire [31:0] _EVAL_1028;
  wire [63:0] _EVAL_2296;
  wire [63:0] _EVAL_5089;
  wire [63:0] _EVAL_3272;
  wire  _EVAL_2556;
  wire  _EVAL_789;
  wire  _EVAL_515;
  wire  _EVAL_2537;
  wire  _EVAL_1070;
  wire  _EVAL_874;
  wire  _EVAL_3365;
  wire [32:0] _EVAL_2325;
  wire  _EVAL_4731;
  wire  _EVAL_5268;
  wire  _EVAL_3453;
  wire  _EVAL_4173;
  wire  _EVAL_3041;
  wire  _EVAL_4452;
  wire [31:0] _EVAL_722;
  wire  _EVAL_4059;
  wire  _EVAL_1099;
  wire  _EVAL_3906;
  wire  _EVAL_2699;
  wire [4:0] _EVAL_3769;
  wire  _EVAL_2631;
  wire [4:0] _EVAL_4640;
  wire [31:0] _EVAL_4457;
  wire [19:0] _EVAL_3785;
  wire [31:0] _EVAL_3354;
  wire [31:0] _EVAL_1680;
  wire [31:0] _EVAL_3822;
  wire [31:0] _EVAL_1468;
  wire [31:0] _EVAL_693;
  wire  _EVAL_3338;
  wire  _EVAL_4336;
  wire  _EVAL_3241;
  wire  _EVAL_1838;
  wire [63:0] _EVAL_1709;
  wire [63:0] _EVAL_4750;
  wire [63:0] _EVAL_2630;
  wire [63:0] _EVAL_3104;
  wire [63:0] _EVAL_2504;
  wire [23:0] _EVAL_3003;
  wire  _EVAL_3559;
  wire  _EVAL_4204;
  wire  _EVAL_2497;
  wire [2:0] _EVAL_5077;
  wire  _EVAL_4274;
  wire  _EVAL_3988;
  wire  _EVAL_4443;
  wire  _EVAL_1062;
  wire  _EVAL_4945;
  wire [1:0] _EVAL_2161;
  wire [5:0] _EVAL_4804;
  wire [3:0] _EVAL_5202;
  wire  _EVAL_4030;
  wire [31:0] _EVAL_797;
  wire [15:0] _EVAL_4404;
  wire [31:0] _EVAL_382;
  wire [31:0] _EVAL_2322;
  wire [31:0] _EVAL_3211;
  wire [31:0] _EVAL_1748;
  wire [31:0] _EVAL_2621;
  wire  _EVAL_2056;
  wire  _EVAL_5135;
  wire  _EVAL_851;
  wire  _EVAL_4676;
  wire  _EVAL_4917;
  wire  _EVAL_3310;
  wire  _EVAL_4871;
  wire  _EVAL_1399;
  wire  _EVAL_1465;
  wire [1:0] _EVAL_904;
  wire  _EVAL_882;
  wire  _EVAL_5131;
  wire [3:0] _EVAL_1614;
  wire [31:0] _EVAL_2997;
  wire  _EVAL_1782;
  wire  _EVAL_4834;
  wire  _EVAL_3181;
  wire  _EVAL_4052;
  wire  _EVAL_2195;
  wire  _EVAL_2132;
  wire  _EVAL_2514;
  wire  _EVAL_624;
  wire  _EVAL_2238;
  wire  _EVAL_2063;
  wire  _EVAL_605;
  wire  _EVAL_5049;
  wire  _EVAL_637;
  wire  _EVAL_4756;
  wire [7:0] _EVAL_586;
  wire [31:0] _EVAL_1338;
  wire [31:0] _EVAL_1971;
  wire [32:0] _EVAL_2584;
  wire  _EVAL_1790;
  wire [31:0] _EVAL_2873;
  wire [28:0] _EVAL_2386;
  wire  _EVAL_2924;
  wire [31:0] _EVAL_5145;
  wire [31:0] _EVAL_3403;
  wire  _EVAL_994;
  wire  _EVAL_1328;
  wire  _EVAL_3603;
  wire  _EVAL_4390;
  wire  _EVAL_403;
  wire  _EVAL_2863;
  wire [31:0] _EVAL_5348;
  wire [31:0] _EVAL_2838;
  wire  _EVAL_936;
  wire  _EVAL_2355;
  wire  _EVAL_4212;
  wire  _EVAL_4590;
  wire [31:0] _EVAL_3106;
  wire [10:0] _EVAL_4178;
  wire [23:0] _EVAL_2031;
  wire [23:0] _EVAL_2446;
  wire [31:0] _EVAL_723;
  wire [31:0] _EVAL_3016;
  wire [31:0] _EVAL_1822;
  wire [4:0] _EVAL_1260;
  wire  _EVAL_2592;
  wire  _EVAL_5227;
  wire [31:0] _EVAL_2455;
  wire [127:0] _EVAL_4669;
  wire  _EVAL_1605;
  wire [31:0] _EVAL_3108;
  wire [31:0] _EVAL_1166;
  wire [31:0] _EVAL_2517;
  wire  _EVAL_3754;
  wire [23:0] _EVAL_4985;
  wire  _EVAL_4021;
  wire [31:0] _EVAL_4220;
  wire  _EVAL_2051;
  wire  _EVAL_2890;
  wire  _EVAL_1994;
  wire [31:0] _EVAL_1619;
  wire [31:0] _EVAL_777;
  wire [31:0] _EVAL_4576;
  wire  _EVAL_4427;
  wire  _EVAL_1902;
  wire  _EVAL_2068;
  wire [1:0] _EVAL_3311;
  wire  _EVAL_443;
  wire  _EVAL_2906;
  wire  _EVAL_2281;
  wire  _EVAL_3198;
  wire  _EVAL_4038;
  wire  _EVAL_3385;
  wire [31:0] _EVAL_3381;
  wire  _EVAL_2305;
  wire [5:0] _EVAL_3109;
  wire  _EVAL_4764;
  wire [32:0] _EVAL_758;
  wire [32:0] _EVAL_4918;
  wire [32:0] _EVAL_3855;
  wire [31:0] _EVAL_4723;
  wire  _EVAL_1583;
  wire [3:0] _EVAL_5356;
  wire  _EVAL_3383;
  wire [31:0] _EVAL_3200;
  wire [31:0] _EVAL_1007;
  wire [6:0] _EVAL_4889;
  wire  _EVAL_4806;
  wire [3:0] _EVAL_3115;
  wire  _EVAL_1634;
  wire [23:0] _EVAL_4131;
  wire  _EVAL_2245;
  wire [23:0] _EVAL_3803;
  wire [23:0] _EVAL_661;
  wire [31:0] _EVAL_3473;
  wire [31:0] _EVAL_3247;
  wire [31:0] _EVAL_4887;
  wire  _EVAL_5004;
  wire [31:0] _EVAL_5362;
  wire [31:0] _EVAL_537;
  wire [23:0] _EVAL_4004;
  wire  _EVAL_1027;
  wire [23:0] _EVAL_4924;
  wire [31:0] _EVAL_1325;
  wire [4:0] _EVAL_2804;
  wire  _EVAL_3138;
  wire [31:0] _EVAL_5269;
  SiFive__EVAL_303 fpu (
    ._EVAL(fpu__EVAL),
    ._EVAL_0(fpu__EVAL_0),
    ._EVAL_1(fpu__EVAL_1),
    ._EVAL_2(fpu__EVAL_2),
    ._EVAL_3(fpu__EVAL_3),
    ._EVAL_4(fpu__EVAL_4),
    ._EVAL_5(fpu__EVAL_5),
    ._EVAL_6(fpu__EVAL_6),
    ._EVAL_7(fpu__EVAL_7),
    ._EVAL_8(fpu__EVAL_8),
    ._EVAL_9(fpu__EVAL_9),
    ._EVAL_10(fpu__EVAL_10),
    ._EVAL_11(fpu__EVAL_11),
    ._EVAL_12(fpu__EVAL_12),
    ._EVAL_13(fpu__EVAL_13),
    ._EVAL_14(fpu__EVAL_14),
    ._EVAL_15(fpu__EVAL_15),
    ._EVAL_16(fpu__EVAL_16),
    ._EVAL_17(fpu__EVAL_17),
    ._EVAL_18(fpu__EVAL_18),
    ._EVAL_19(fpu__EVAL_19),
    ._EVAL_20(fpu__EVAL_20),
    ._EVAL_21(fpu__EVAL_21),
    ._EVAL_22(fpu__EVAL_22),
    ._EVAL_23(fpu__EVAL_23),
    ._EVAL_24(fpu__EVAL_24),
    ._EVAL_25(fpu__EVAL_25),
    ._EVAL_26(fpu__EVAL_26),
    ._EVAL_27(fpu__EVAL_27),
    ._EVAL_28(fpu__EVAL_28),
    ._EVAL_29(fpu__EVAL_29),
    ._EVAL_30(fpu__EVAL_30),
    ._EVAL_31(fpu__EVAL_31),
    ._EVAL_32(fpu__EVAL_32),
    ._EVAL_33(fpu__EVAL_33),
    ._EVAL_34(fpu__EVAL_34),
    ._EVAL_35(fpu__EVAL_35),
    ._EVAL_36(fpu__EVAL_36),
    ._EVAL_37(fpu__EVAL_37),
    ._EVAL_38(fpu__EVAL_38),
    ._EVAL_39(fpu__EVAL_39),
    ._EVAL_40(fpu__EVAL_40),
    ._EVAL_41(fpu__EVAL_41),
    ._EVAL_42(fpu__EVAL_42),
    ._EVAL_43(fpu__EVAL_43),
    ._EVAL_44(fpu__EVAL_44),
    ._EVAL_45(fpu__EVAL_45),
    ._EVAL_46(fpu__EVAL_46),
    ._EVAL_47(fpu__EVAL_47),
    ._EVAL_48(fpu__EVAL_48),
    ._EVAL_49(fpu__EVAL_49),
    ._EVAL_50(fpu__EVAL_50),
    ._EVAL_51(fpu__EVAL_51),
    ._EVAL_52(fpu__EVAL_52),
    ._EVAL_53(fpu__EVAL_53),
    ._EVAL_54(fpu__EVAL_54),
    ._EVAL_55(fpu__EVAL_55),
    ._EVAL_56(fpu__EVAL_56),
    ._EVAL_57(fpu__EVAL_57),
    ._EVAL_58(fpu__EVAL_58),
    ._EVAL_59(fpu__EVAL_59),
    ._EVAL_60(fpu__EVAL_60)
  );
  EICG_wrapper bullet_clock_gate (
    .in(bullet_clock_gate_in),
    .en(bullet_clock_gate_en),
    .out(bullet_clock_gate_out)
  );
  SiFive__EVAL_305 divider (
    ._EVAL(divider__EVAL),
    ._EVAL_0(divider__EVAL_0),
    ._EVAL_1(divider__EVAL_1),
    ._EVAL_2(divider__EVAL_2),
    ._EVAL_3(divider__EVAL_3),
    ._EVAL_4(divider__EVAL_4),
    ._EVAL_5(divider__EVAL_5),
    ._EVAL_6(divider__EVAL_6),
    ._EVAL_7(divider__EVAL_7),
    ._EVAL_8(divider__EVAL_8),
    ._EVAL_9(divider__EVAL_9),
    ._EVAL_10(divider__EVAL_10),
    ._EVAL_11(divider__EVAL_11)
  );
  SiFive__EVAL_304 csr (
    ._EVAL(csr__EVAL),
    ._EVAL_0(csr__EVAL_0),
    ._EVAL_1(csr__EVAL_1),
    ._EVAL_2(csr__EVAL_2),
    ._EVAL_3(csr__EVAL_3),
    ._EVAL_4(csr__EVAL_4),
    ._EVAL_5(csr__EVAL_5),
    ._EVAL_6(csr__EVAL_6),
    ._EVAL_7(csr__EVAL_7),
    ._EVAL_8(csr__EVAL_8),
    ._EVAL_9(csr__EVAL_9),
    ._EVAL_10(csr__EVAL_10),
    ._EVAL_11(csr__EVAL_11),
    ._EVAL_12(csr__EVAL_12),
    ._EVAL_13(csr__EVAL_13),
    ._EVAL_14(csr__EVAL_14),
    ._EVAL_15(csr__EVAL_15),
    ._EVAL_16(csr__EVAL_16),
    ._EVAL_17(csr__EVAL_17),
    ._EVAL_18(csr__EVAL_18),
    ._EVAL_19(csr__EVAL_19),
    ._EVAL_20(csr__EVAL_20),
    ._EVAL_21(csr__EVAL_21),
    ._EVAL_22(csr__EVAL_22),
    ._EVAL_23(csr__EVAL_23),
    ._EVAL_24(csr__EVAL_24),
    ._EVAL_25(csr__EVAL_25),
    ._EVAL_26(csr__EVAL_26),
    ._EVAL_27(csr__EVAL_27),
    ._EVAL_28(csr__EVAL_28),
    ._EVAL_29(csr__EVAL_29),
    ._EVAL_30(csr__EVAL_30),
    ._EVAL_31(csr__EVAL_31),
    ._EVAL_32(csr__EVAL_32),
    ._EVAL_33(csr__EVAL_33),
    ._EVAL_34(csr__EVAL_34),
    ._EVAL_35(csr__EVAL_35),
    ._EVAL_36(csr__EVAL_36),
    ._EVAL_37(csr__EVAL_37),
    ._EVAL_38(csr__EVAL_38),
    ._EVAL_39(csr__EVAL_39),
    ._EVAL_40(csr__EVAL_40),
    ._EVAL_41(csr__EVAL_41),
    ._EVAL_42(csr__EVAL_42),
    ._EVAL_43(csr__EVAL_43),
    ._EVAL_44(csr__EVAL_44),
    ._EVAL_45(csr__EVAL_45),
    ._EVAL_46(csr__EVAL_46),
    ._EVAL_47(csr__EVAL_47),
    ._EVAL_48(csr__EVAL_48),
    ._EVAL_49(csr__EVAL_49),
    ._EVAL_50(csr__EVAL_50),
    ._EVAL_51(csr__EVAL_51),
    ._EVAL_52(csr__EVAL_52),
    ._EVAL_53(csr__EVAL_53),
    ._EVAL_54(csr__EVAL_54),
    ._EVAL_55(csr__EVAL_55),
    ._EVAL_56(csr__EVAL_56),
    ._EVAL_57(csr__EVAL_57),
    ._EVAL_58(csr__EVAL_58),
    ._EVAL_59(csr__EVAL_59),
    ._EVAL_60(csr__EVAL_60),
    ._EVAL_61(csr__EVAL_61),
    ._EVAL_62(csr__EVAL_62),
    ._EVAL_63(csr__EVAL_63),
    ._EVAL_64(csr__EVAL_64),
    ._EVAL_65(csr__EVAL_65),
    ._EVAL_66(csr__EVAL_66),
    ._EVAL_67(csr__EVAL_67),
    ._EVAL_68(csr__EVAL_68),
    ._EVAL_69(csr__EVAL_69),
    ._EVAL_70(csr__EVAL_70),
    ._EVAL_71(csr__EVAL_71),
    ._EVAL_72(csr__EVAL_72),
    ._EVAL_73(csr__EVAL_73),
    ._EVAL_74(csr__EVAL_74),
    ._EVAL_75(csr__EVAL_75),
    ._EVAL_76(csr__EVAL_76),
    ._EVAL_77(csr__EVAL_77),
    ._EVAL_78(csr__EVAL_78),
    ._EVAL_79(csr__EVAL_79),
    ._EVAL_80(csr__EVAL_80),
    ._EVAL_81(csr__EVAL_81),
    ._EVAL_82(csr__EVAL_82),
    ._EVAL_83(csr__EVAL_83),
    ._EVAL_84(csr__EVAL_84),
    ._EVAL_85(csr__EVAL_85),
    ._EVAL_86(csr__EVAL_86),
    ._EVAL_87(csr__EVAL_87),
    ._EVAL_88(csr__EVAL_88),
    ._EVAL_89(csr__EVAL_89),
    ._EVAL_90(csr__EVAL_90),
    ._EVAL_91(csr__EVAL_91),
    ._EVAL_92(csr__EVAL_92),
    ._EVAL_93(csr__EVAL_93),
    ._EVAL_94(csr__EVAL_94),
    ._EVAL_95(csr__EVAL_95),
    ._EVAL_96(csr__EVAL_96),
    ._EVAL_97(csr__EVAL_97),
    ._EVAL_98(csr__EVAL_98),
    ._EVAL_99(csr__EVAL_99),
    ._EVAL_100(csr__EVAL_100),
    ._EVAL_101(csr__EVAL_101),
    ._EVAL_102(csr__EVAL_102),
    ._EVAL_103(csr__EVAL_103),
    ._EVAL_104(csr__EVAL_104),
    ._EVAL_105(csr__EVAL_105),
    ._EVAL_106(csr__EVAL_106),
    ._EVAL_107(csr__EVAL_107),
    ._EVAL_108(csr__EVAL_108),
    ._EVAL_109(csr__EVAL_109),
    ._EVAL_110(csr__EVAL_110),
    ._EVAL_111(csr__EVAL_111),
    ._EVAL_112(csr__EVAL_112),
    ._EVAL_113(csr__EVAL_113),
    ._EVAL_114(csr__EVAL_114),
    ._EVAL_115(csr__EVAL_115),
    ._EVAL_116(csr__EVAL_116),
    ._EVAL_117(csr__EVAL_117),
    ._EVAL_118(csr__EVAL_118),
    ._EVAL_119(csr__EVAL_119),
    ._EVAL_120(csr__EVAL_120),
    ._EVAL_121(csr__EVAL_121),
    ._EVAL_122(csr__EVAL_122),
    ._EVAL_123(csr__EVAL_123),
    ._EVAL_124(csr__EVAL_124),
    ._EVAL_125(csr__EVAL_125),
    ._EVAL_126(csr__EVAL_126),
    ._EVAL_127(csr__EVAL_127),
    ._EVAL_128(csr__EVAL_128),
    ._EVAL_129(csr__EVAL_129),
    ._EVAL_130(csr__EVAL_130),
    ._EVAL_131(csr__EVAL_131),
    ._EVAL_132(csr__EVAL_132),
    ._EVAL_133(csr__EVAL_133),
    ._EVAL_134(csr__EVAL_134),
    ._EVAL_135(csr__EVAL_135),
    ._EVAL_136(csr__EVAL_136),
    ._EVAL_137(csr__EVAL_137),
    ._EVAL_138(csr__EVAL_138),
    ._EVAL_139(csr__EVAL_139),
    ._EVAL_140(csr__EVAL_140),
    ._EVAL_141(csr__EVAL_141),
    ._EVAL_142(csr__EVAL_142),
    ._EVAL_143(csr__EVAL_143),
    ._EVAL_144(csr__EVAL_144),
    ._EVAL_145(csr__EVAL_145),
    ._EVAL_146(csr__EVAL_146),
    ._EVAL_147(csr__EVAL_147),
    ._EVAL_148(csr__EVAL_148),
    ._EVAL_149(csr__EVAL_149),
    ._EVAL_150(csr__EVAL_150),
    ._EVAL_151(csr__EVAL_151),
    ._EVAL_152(csr__EVAL_152),
    ._EVAL_153(csr__EVAL_153),
    ._EVAL_154(csr__EVAL_154),
    ._EVAL_155(csr__EVAL_155),
    ._EVAL_156(csr__EVAL_156),
    ._EVAL_157(csr__EVAL_157),
    ._EVAL_158(csr__EVAL_158),
    ._EVAL_159(csr__EVAL_159),
    ._EVAL_160(csr__EVAL_160),
    ._EVAL_161(csr__EVAL_161),
    ._EVAL_162(csr__EVAL_162),
    ._EVAL_163(csr__EVAL_163),
    ._EVAL_164(csr__EVAL_164),
    ._EVAL_165(csr__EVAL_165),
    ._EVAL_166(csr__EVAL_166),
    ._EVAL_167(csr__EVAL_167)
  );
  SiFive__EVAL_306 m (
    ._EVAL(m__EVAL),
    ._EVAL_0(m__EVAL_0),
    ._EVAL_1(m__EVAL_1),
    ._EVAL_2(m__EVAL_2),
    ._EVAL_3(m__EVAL_3),
    ._EVAL_4(m__EVAL_4),
    ._EVAL_5(m__EVAL_5)
  );
  EICG_wrapper fpu_clock_gate (
    .in(fpu_clock_gate_in),
    .en(fpu_clock_gate_en),
    .out(fpu_clock_gate_out)
  );
  assign _EVAL_708__EVAL_709_addr = _EVAL_274;
  assign _EVAL_708__EVAL_709_data = _EVAL_708[_EVAL_708__EVAL_709_addr];
  assign _EVAL_708__EVAL_710_addr = _EVAL_180;
  assign _EVAL_708__EVAL_710_data = _EVAL_708[_EVAL_708__EVAL_710_addr];
  assign _EVAL_708__EVAL_711_addr = _EVAL_154;
  assign _EVAL_708__EVAL_711_data = _EVAL_708[_EVAL_708__EVAL_711_addr];
  assign _EVAL_708__EVAL_712_addr = _EVAL_68;
  assign _EVAL_708__EVAL_712_data = _EVAL_708[_EVAL_708__EVAL_712_addr];
  assign _EVAL_708__EVAL_713_data = _EVAL_4863;
  assign _EVAL_708__EVAL_713_addr = _EVAL_5099;
  assign _EVAL_708__EVAL_713_mask = 1'h1;
  assign _EVAL_708__EVAL_713_en = _EVAL_4774 & _EVAL_332;
  assign _EVAL_708__EVAL_714_data = _EVAL_2257 ? divider__EVAL_8 : _EVAL_3279;
  assign _EVAL_708__EVAL_714_addr = _EVAL_2257 ? divider__EVAL_11 : _EVAL_4939;
  assign _EVAL_708__EVAL_714_mask = 1'h1;
  assign _EVAL_708__EVAL_714_en = _EVAL_5252 & _EVAL_5386;
  assign _EVAL_708__EVAL_715_data = 32'h0;
  assign _EVAL_708__EVAL_715_addr = 5'h0;
  assign _EVAL_708__EVAL_715_mask = 1'h1;
  assign _EVAL_708__EVAL_715_en = 1'h1;
  assign _EVAL_2741__EVAL_2742_addr = _EVAL_4400;
  assign _EVAL_2741__EVAL_2742_data = _EVAL_2741[_EVAL_2741__EVAL_2742_addr];
  assign _EVAL_2741__EVAL_2743_addr = _EVAL_1795;
  assign _EVAL_2741__EVAL_2743_data = _EVAL_2741[_EVAL_2741__EVAL_2743_addr];
  assign _EVAL_2741__EVAL_2744_addr = _EVAL_3851;
  assign _EVAL_2741__EVAL_2744_data = _EVAL_2741[_EVAL_2741__EVAL_2744_addr];
  assign _EVAL_2741__EVAL_2745_addr = _EVAL_2320;
  assign _EVAL_2741__EVAL_2745_data = _EVAL_2741[_EVAL_2741__EVAL_2745_addr];
  assign _EVAL_2741__EVAL_2746_addr = _EVAL_375;
  assign _EVAL_2741__EVAL_2746_data = _EVAL_2741[_EVAL_2741__EVAL_2746_addr];
  assign _EVAL_2741__EVAL_2747_addr = _EVAL_1356;
  assign _EVAL_2741__EVAL_2747_data = _EVAL_2741[_EVAL_2741__EVAL_2747_addr];
  assign _EVAL_2741__EVAL_2748_addr = _EVAL_1480;
  assign _EVAL_2741__EVAL_2748_data = _EVAL_2741[_EVAL_2741__EVAL_2748_addr];
  assign _EVAL_2741__EVAL_2749_addr = _EVAL_4745;
  assign _EVAL_2741__EVAL_2749_data = _EVAL_2741[_EVAL_2741__EVAL_2749_addr];
  assign _EVAL_2741__EVAL_2750_addr = _EVAL_3711;
  assign _EVAL_2741__EVAL_2750_data = _EVAL_2741[_EVAL_2741__EVAL_2750_addr];
  assign _EVAL_2741__EVAL_2751_data = {_EVAL_3115,_EVAL_5230};
  assign _EVAL_2741__EVAL_2751_addr = _EVAL_5099;
  assign _EVAL_2741__EVAL_2751_mask = 1'h1;
  assign _EVAL_2741__EVAL_2751_en = _EVAL_4774 & _EVAL_4362;
  assign _EVAL_2741__EVAL_2752_data = fpu__EVAL_21;
  assign _EVAL_2741__EVAL_2752_addr = fpu__EVAL_29;
  assign _EVAL_2741__EVAL_2752_mask = 1'h1;
  assign _EVAL_2741__EVAL_2752_en = fpu__EVAL_12 & fpu__EVAL_55;
  assign _EVAL_1844 = _EVAL_98 == 1'h0;
  assign _EVAL_5290 = _EVAL_176 == 1'h0;
  assign _EVAL_4710 = _EVAL_1844 & _EVAL_5290;
  assign _EVAL_2703 = _EVAL_247 == 1'h0;
  assign _EVAL_1575 = _EVAL_98 & _EVAL_2703;
  assign _EVAL_4848 = _EVAL_4710 | _EVAL_1575;
  assign _EVAL_3081 = _EVAL_90 & _EVAL_236;
  assign _EVAL_315 = _EVAL_4848 | _EVAL_3081;
  assign _EVAL_2400 = _EVAL_315 ? _EVAL_73 : _EVAL_121;
  assign _EVAL_1762 = _EVAL_2400[0];
  assign _EVAL_1335 = csr__EVAL_14[1:0];
  assign _EVAL_4196 = _EVAL_1335 == 2'h1;
  assign _EVAL_2393 = _EVAL_4167 | _EVAL_4168;
  assign _EVAL_3538 = csr__EVAL_14[31:8];
  assign _EVAL_3681 = _EVAL_3538[0];
  assign _EVAL_1778 = _EVAL_490 == 1'h0;
  assign _EVAL_4721 = _EVAL_4000 & _EVAL_1778;
  assign _EVAL_1969 = _EVAL_4721 & _EVAL_1134;
  assign _EVAL_3066 = _EVAL_3681 ? _EVAL_1647 : _EVAL_1969;
  assign _EVAL_3904 = _EVAL_2443 == 1'h0;
  assign _EVAL_890 = _EVAL_612 & _EVAL_3904;
  assign _EVAL_2868 = _EVAL_890 & _EVAL_3523;
  assign _EVAL_3519 = _EVAL_3681 ? 1'h0 : _EVAL_2868;
  assign _EVAL_2523 = _EVAL_3066 + _EVAL_3519;
  assign _EVAL_5069 = _EVAL_4196 ? {{1'd0}, _EVAL_2393} : _EVAL_2523;
  assign _EVAL_1623 = fpu__EVAL_34 > 3'h1;
  assign _EVAL_351 = fpu__EVAL_8 & fpu__EVAL_24;
  assign _EVAL_1722 = fpu__EVAL_57;
  assign _EVAL_1616 = _EVAL_154 == _EVAL_1722;
  assign _EVAL_361 = _EVAL_148 & _EVAL_1616;
  assign _EVAL_1387 = _EVAL_68 == _EVAL_1722;
  assign _EVAL_3820 = _EVAL_179 & _EVAL_1387;
  assign _EVAL_2876 = _EVAL_361 | _EVAL_3820;
  assign _EVAL_4127 = _EVAL_121[6:2];
  assign _EVAL_2956 = _EVAL_4127 == _EVAL_1722;
  assign _EVAL_1608 = _EVAL_119 & _EVAL_2956;
  assign _EVAL_588 = _EVAL_2876 | _EVAL_1608;
  assign _EVAL_4623 = _EVAL_351 & _EVAL_588;
  assign _EVAL_2595 = _EVAL_274 == _EVAL_1722;
  assign _EVAL_3168 = _EVAL_39 & _EVAL_2595;
  assign _EVAL_2133 = _EVAL_180 == _EVAL_1722;
  assign _EVAL_1299 = _EVAL_188 & _EVAL_2133;
  assign _EVAL_1655 = _EVAL_3168 | _EVAL_1299;
  assign _EVAL_3212 = _EVAL_73[6:2];
  assign _EVAL_2594 = _EVAL_3212 == _EVAL_1722;
  assign _EVAL_2313 = _EVAL_260 & _EVAL_2594;
  assign _EVAL_1372 = _EVAL_1655 | _EVAL_2313;
  assign _EVAL_2025 = _EVAL_351 & _EVAL_1372;
  assign _EVAL_783 = _EVAL_315 ? _EVAL_4623 : _EVAL_2025;
  assign _EVAL_3808 = _EVAL_1623 & _EVAL_783;
  assign _EVAL_4357 = _EVAL_315 ? _EVAL_16 : _EVAL_58;
  assign _EVAL_3671 = _EVAL_315 ? _EVAL_39 : _EVAL_148;
  assign _EVAL_3116 = _EVAL_4357 | _EVAL_3671;
  assign _EVAL_3082 = fpu__EVAL_54 == 5'h7;
  assign _EVAL_631 = fpu__EVAL_13 & _EVAL_3082;
  assign _EVAL_1434 = _EVAL_3116 & _EVAL_631;
  assign _EVAL_3141 = _EVAL_16 & _EVAL_4299;
  assign _EVAL_2321 = _EVAL_214 & _EVAL_4692;
  assign _EVAL_747 = _EVAL_3141 | _EVAL_2321;
  assign _EVAL_2394 = _EVAL_171 == _EVAL_4135;
  assign _EVAL_5360 = _EVAL_747 & _EVAL_2394;
  assign _EVAL_4683 = _EVAL_58 & _EVAL_4299;
  assign _EVAL_1255 = _EVAL_268 & _EVAL_4692;
  assign _EVAL_739 = _EVAL_4683 | _EVAL_1255;
  assign _EVAL_3346 = _EVAL_91 == _EVAL_4135;
  assign _EVAL_3763 = _EVAL_739 & _EVAL_3346;
  assign _EVAL_2532 = _EVAL_315 ? _EVAL_5360 : _EVAL_3763;
  assign _EVAL_3962 = _EVAL_4240 & _EVAL_2532;
  assign _EVAL_1414 = _EVAL_315 ? _EVAL_3962 : _EVAL_3962;
  assign _EVAL_1546 = _EVAL_1414 & _EVAL_4299;
  assign _EVAL_4528 = _EVAL_1434 | _EVAL_1546;
  assign _EVAL_500 = _EVAL_16 & _EVAL_2573;
  assign _EVAL_1570 = _EVAL_214 & _EVAL_1724;
  assign _EVAL_4348 = _EVAL_500 | _EVAL_1570;
  assign _EVAL_2653 = _EVAL_171 == _EVAL_3670;
  assign _EVAL_1158 = _EVAL_4348 & _EVAL_2653;
  assign _EVAL_1507 = _EVAL_58 & _EVAL_2573;
  assign _EVAL_2108 = _EVAL_268 & _EVAL_1724;
  assign _EVAL_546 = _EVAL_1507 | _EVAL_2108;
  assign _EVAL_408 = _EVAL_91 == _EVAL_3670;
  assign _EVAL_4067 = _EVAL_546 & _EVAL_408;
  assign _EVAL_584 = _EVAL_315 ? _EVAL_1158 : _EVAL_4067;
  assign _EVAL_1311 = _EVAL_3624 & _EVAL_584;
  assign _EVAL_1319 = _EVAL_315 ? _EVAL_1311 : _EVAL_1311;
  assign _EVAL_1952 = _EVAL_1319 & _EVAL_2573;
  assign _EVAL_3850 = fpu__EVAL_4;
  assign _EVAL_4696 = _EVAL_1952 & _EVAL_3850;
  assign _EVAL_4197 = _EVAL_4528 | _EVAL_4696;
  assign _EVAL_591 = fpu__EVAL_13;
  assign _EVAL_4963 = _EVAL_591 & _EVAL_16;
  assign _EVAL_4490 = _EVAL_171 == fpu__EVAL_37;
  assign _EVAL_821 = _EVAL_4963 & _EVAL_4490;
  assign _EVAL_3864 = _EVAL_591 & _EVAL_58;
  assign _EVAL_4771 = _EVAL_91 == fpu__EVAL_37;
  assign _EVAL_4260 = _EVAL_3864 & _EVAL_4771;
  assign _EVAL_903 = _EVAL_315 ? _EVAL_821 : _EVAL_4260;
  assign _EVAL_862 = _EVAL_4197 | _EVAL_903;
  assign _EVAL_1445 = {_EVAL_4019,_EVAL_4706};
  assign _EVAL_3957 = _EVAL_1445[4:3];
  assign _EVAL_1694 = _EVAL_5344 == 1'h0;
  assign _EVAL_5111 = _EVAL_1694 | _EVAL_2145;
  assign _EVAL_3755 = _EVAL_4201[0];
  assign _EVAL_1120 = _EVAL_4715[3];
  assign _EVAL_5246 = {_EVAL_4019,_EVAL_1198};
  assign _EVAL_2208 = _EVAL_5246[5:3];
  assign _EVAL_4494 = _EVAL_4715[2:0];
  assign _EVAL_4757 = _EVAL_5246[7:6];
  assign _EVAL_5219 = _EVAL_4706[2:0];
  assign _EVAL_818 = {3'h3,_EVAL_2208,_EVAL_4494,_EVAL_4757,_EVAL_5219,2'h0};
  assign _EVAL_4395 = _EVAL_5246[5];
  assign _EVAL_1958 = _EVAL_5246[4:3];
  assign _EVAL_927 = _EVAL_5246[8:6];
  assign _EVAL_1954 = {3'h3,_EVAL_4395,_EVAL_4706,_EVAL_1958,_EVAL_927,2'h2};
  assign _EVAL_1113 = _EVAL_1120 ? _EVAL_818 : _EVAL_1954;
  assign _EVAL_556 = _EVAL_5246[2];
  assign _EVAL_3661 = _EVAL_5246[6];
  assign _EVAL_2429 = {3'h2,_EVAL_2208,_EVAL_4494,_EVAL_556,_EVAL_3661,_EVAL_5219,2'h0};
  assign _EVAL_2874 = _EVAL_5246[4:2];
  assign _EVAL_3017 = {3'h2,_EVAL_4395,_EVAL_4706,_EVAL_2874,_EVAL_4757,2'h2};
  assign _EVAL_2260 = _EVAL_1120 ? _EVAL_2429 : _EVAL_3017;
  assign _EVAL_5236 = _EVAL_3755 ? _EVAL_1113 : _EVAL_2260;
  assign _EVAL_3373 = _EVAL_21[15:13];
  assign _EVAL_2034 = _EVAL_3373 == 3'h5;
  assign _EVAL_3232 = _EVAL_1913[31:23];
  assign _EVAL_618 = {1'b0,$signed(_EVAL_3232)};
  assign _EVAL_3796 = _EVAL_618[7:0];
  assign _EVAL_3409 = _EVAL_4962 & _EVAL_188;
  assign _EVAL_4001 = _EVAL_1333 & _EVAL_250;
  assign _EVAL_4724 = _EVAL_3409 | _EVAL_4001;
  assign _EVAL_1271 = _EVAL_268 | _EVAL_58;
  assign _EVAL_1306 = {_EVAL_58,_EVAL_91};
  assign _EVAL_2332 = _EVAL_4160 >> _EVAL_1306;
  assign _EVAL_2488 = _EVAL_2332[0];
  assign _EVAL_4996 = _EVAL_1103 == 1'h0;
  assign _EVAL_813 = _EVAL_3814 & _EVAL_4996;
  assign _EVAL_1677 = _EVAL_3771 == 1'h0;
  assign _EVAL_3912 = _EVAL_813 & _EVAL_1677;
  assign _EVAL_1477 = _EVAL_4805 == 1'h0;
  assign _EVAL_1535 = _EVAL_3912 & _EVAL_1477;
  assign _EVAL_2564 = _EVAL_2823 == _EVAL_1306;
  assign _EVAL_2509 = _EVAL_1535 & _EVAL_2564;
  assign _EVAL_5391 = _EVAL_2488 | _EVAL_2509;
  assign _EVAL_2617 = {{1'd0}, divider__EVAL_5};
  assign _EVAL_1573 = _EVAL_2617 == _EVAL_1306;
  assign _EVAL_2120 = divider__EVAL_2 & _EVAL_1573;
  assign _EVAL_1966 = _EVAL_5391 | _EVAL_2120;
  assign _EVAL_296 = divider__EVAL == 1'h0;
  assign _EVAL_2257 = divider__EVAL_0 & divider__EVAL_3;
  assign _EVAL_423 = _EVAL_2257 == 1'h0;
  assign _EVAL_1190 = _EVAL_296 & _EVAL_423;
  assign _EVAL_4158 = {{1'd0}, divider__EVAL_11};
  assign _EVAL_2452 = _EVAL_4158 == _EVAL_1306;
  assign _EVAL_2942 = _EVAL_1190 & _EVAL_2452;
  assign _EVAL_2481 = _EVAL_1966 | _EVAL_2942;
  assign _EVAL_1242 = _EVAL_1271 & _EVAL_2481;
  assign _EVAL_2524 = _EVAL_1 | _EVAL_148;
  assign _EVAL_2316 = {_EVAL_148,_EVAL_154};
  assign _EVAL_2301 = _EVAL_4160 >> _EVAL_2316;
  assign _EVAL_5337 = _EVAL_2301[0];
  assign _EVAL_3422 = _EVAL_2823 == _EVAL_2316;
  assign _EVAL_902 = _EVAL_1535 & _EVAL_3422;
  assign _EVAL_1927 = _EVAL_5337 | _EVAL_902;
  assign _EVAL_4388 = _EVAL_2617 == _EVAL_2316;
  assign _EVAL_2049 = divider__EVAL_2 & _EVAL_4388;
  assign _EVAL_3419 = _EVAL_1927 | _EVAL_2049;
  assign _EVAL_2549 = _EVAL_4158 == _EVAL_2316;
  assign _EVAL_4564 = _EVAL_1190 & _EVAL_2549;
  assign _EVAL_3956 = _EVAL_3419 | _EVAL_4564;
  assign _EVAL_512 = _EVAL_2524 & _EVAL_3956;
  assign _EVAL_2600 = _EVAL_1242 | _EVAL_512;
  assign _EVAL_3679 = _EVAL_141 | _EVAL_179;
  assign _EVAL_2954 = {_EVAL_179,_EVAL_68};
  assign _EVAL_3509 = _EVAL_4160 >> _EVAL_2954;
  assign _EVAL_2080 = _EVAL_3509[0];
  assign _EVAL_1685 = _EVAL_2823 == _EVAL_2954;
  assign _EVAL_1167 = _EVAL_1535 & _EVAL_1685;
  assign _EVAL_5126 = _EVAL_2080 | _EVAL_1167;
  assign _EVAL_4986 = _EVAL_2617 == _EVAL_2954;
  assign _EVAL_614 = divider__EVAL_2 & _EVAL_4986;
  assign _EVAL_2916 = _EVAL_5126 | _EVAL_614;
  assign _EVAL_1670 = _EVAL_4158 == _EVAL_2954;
  assign _EVAL_1320 = _EVAL_1190 & _EVAL_1670;
  assign _EVAL_4760 = _EVAL_2916 | _EVAL_1320;
  assign _EVAL_2638 = _EVAL_3679 & _EVAL_4760;
  assign _EVAL_308 = _EVAL_2600 | _EVAL_2638;
  assign _EVAL_2897 = {_EVAL_119,_EVAL_4127};
  assign _EVAL_1322 = _EVAL_4160 >> _EVAL_2897;
  assign _EVAL_4769 = _EVAL_1322[0];
  assign _EVAL_1676 = _EVAL_2823 == _EVAL_2897;
  assign _EVAL_1218 = _EVAL_1535 & _EVAL_1676;
  assign _EVAL_3492 = _EVAL_4769 | _EVAL_1218;
  assign _EVAL_1293 = _EVAL_2617 == _EVAL_2897;
  assign _EVAL_1855 = divider__EVAL_2 & _EVAL_1293;
  assign _EVAL_386 = _EVAL_3492 | _EVAL_1855;
  assign _EVAL_2901 = _EVAL_4158 == _EVAL_2897;
  assign _EVAL_3027 = _EVAL_1190 & _EVAL_2901;
  assign _EVAL_4302 = _EVAL_386 | _EVAL_3027;
  assign _EVAL_3374 = _EVAL_119 & _EVAL_4302;
  assign _EVAL_3256 = _EVAL_308 | _EVAL_3374;
  assign _EVAL_2216 = _EVAL_4135 == _EVAL_274;
  assign _EVAL_2705 = _EVAL_4692 & _EVAL_2216;
  assign _EVAL_3231 = _EVAL_4240 & _EVAL_2705;
  assign _EVAL_3758 = _EVAL_4135 == _EVAL_154;
  assign _EVAL_4222 = _EVAL_4692 & _EVAL_3758;
  assign _EVAL_589 = _EVAL_4240 & _EVAL_4222;
  assign _EVAL_2668 = _EVAL_315 ? _EVAL_3231 : _EVAL_589;
  assign _EVAL_1241 = _EVAL_269[12];
  assign _EVAL_4033 = _EVAL_1241 ? 10'h3ff : 10'h0;
  assign _EVAL_775 = _EVAL_269[8];
  assign _EVAL_524 = _EVAL_269[10:9];
  assign _EVAL_5194 = _EVAL_269[6];
  assign _EVAL_4278 = _EVAL_269[7];
  assign _EVAL_2243 = _EVAL_269[2];
  assign _EVAL_4516 = _EVAL_269[11];
  assign _EVAL_2607 = _EVAL_269[5:3];
  assign _EVAL_2778 = {_EVAL_4033,_EVAL_775,_EVAL_524,_EVAL_5194,_EVAL_4278,_EVAL_2243,_EVAL_4516,_EVAL_2607,1'h0};
  assign _EVAL_2978 = _EVAL_2778[20];
  assign _EVAL_1285 = _EVAL_2778[10:1];
  assign _EVAL_4259 = _EVAL_2778[11];
  assign _EVAL_2173 = _EVAL_2778[19:12];
  assign _EVAL_1628 = {_EVAL_2978,_EVAL_1285,_EVAL_4259,_EVAL_2173,5'h1,7'h6f};
  assign _EVAL_4809 = _EVAL_5099 == _EVAL_1480;
  assign _EVAL_3012 = _EVAL_4614 == 5'ha;
  assign _EVAL_2359 = _EVAL_1024[0];
  assign _EVAL_2448 = _EVAL_5363[3];
  assign _EVAL_1542 = {_EVAL_3229,_EVAL_3742};
  assign _EVAL_3872 = _EVAL_1542[5:3];
  assign _EVAL_4488 = _EVAL_5363[2:0];
  assign _EVAL_3551 = _EVAL_1542[7:6];
  assign _EVAL_2846 = _EVAL_1641[2:0];
  assign _EVAL_3470 = {3'h7,_EVAL_3872,_EVAL_4488,_EVAL_3551,_EVAL_2846,2'h0};
  assign _EVAL_857 = _EVAL_1542[8:6];
  assign _EVAL_4020 = {3'h7,_EVAL_3872,_EVAL_857,_EVAL_1641,2'h2};
  assign _EVAL_3599 = _EVAL_2448 ? _EVAL_3470 : _EVAL_4020;
  assign _EVAL_3126 = _EVAL_1542[2];
  assign _EVAL_2483 = _EVAL_1542[6];
  assign _EVAL_4153 = {3'h6,_EVAL_3872,_EVAL_4488,_EVAL_3126,_EVAL_2483,_EVAL_2846,2'h0};
  assign _EVAL_2775 = _EVAL_1542[5:2];
  assign _EVAL_3552 = {3'h6,_EVAL_2775,_EVAL_3551,_EVAL_1641,2'h2};
  assign _EVAL_2774 = _EVAL_2448 ? _EVAL_4153 : _EVAL_3552;
  assign _EVAL_1704 = _EVAL_2359 ? _EVAL_3599 : _EVAL_2774;
  assign _EVAL_850 = _EVAL_4614 == 5'h9;
  assign _EVAL_5185 = _EVAL_1024[1];
  assign _EVAL_4051 = {3'h5,_EVAL_3872,_EVAL_4488,_EVAL_3551,_EVAL_2846,2'h0};
  assign _EVAL_3344 = {3'h5,_EVAL_3872,_EVAL_857,_EVAL_1641,2'h2};
  assign _EVAL_1706 = _EVAL_2448 ? _EVAL_4051 : _EVAL_3344;
  assign _EVAL_1481 = {3'h7,_EVAL_3872,_EVAL_4488,_EVAL_3126,_EVAL_2483,_EVAL_2846,2'h0};
  assign _EVAL_4520 = {3'h7,_EVAL_2775,_EVAL_3551,_EVAL_1641,2'h2};
  assign _EVAL_3555 = _EVAL_2448 ? _EVAL_1481 : _EVAL_4520;
  assign _EVAL_4447 = _EVAL_2359 ? _EVAL_1706 : _EVAL_3555;
  assign _EVAL_3913 = {3'h4,_EVAL_3872,_EVAL_4488,_EVAL_3126,_EVAL_2483,_EVAL_2846,2'h0};
  assign _EVAL_771 = _EVAL_5185 ? _EVAL_4447 : _EVAL_3913;
  assign _EVAL_4093 = _EVAL_4614 == 5'h8;
  assign _EVAL_1901 = _EVAL_4614 == 5'h7;
  assign _EVAL_3133 = {_EVAL_3229,_EVAL_1641,_EVAL_5363,_EVAL_1024};
  assign _EVAL_2904 = $signed(_EVAL_3133);
  assign _EVAL_2801 = _EVAL_2904[19];
  assign _EVAL_1067 = _EVAL_2904[4:0];
  assign _EVAL_2150 = {3'h3,_EVAL_2801,_EVAL_3742,_EVAL_1067,2'h1};
  assign _EVAL_762 = _EVAL_4614 == 5'h6;
  assign _EVAL_735 = {_EVAL_3229,_EVAL_1641};
  assign _EVAL_2512 = _EVAL_735[5];
  assign _EVAL_2998 = _EVAL_735[4:0];
  assign _EVAL_3862 = {3'h4,_EVAL_2512,2'h0,_EVAL_4488,_EVAL_2998,2'h1};
  assign _EVAL_302 = _EVAL_3862 | 16'h800;
  assign _EVAL_3360 = _EVAL_1024[2];
  assign _EVAL_323 = _EVAL_3229[5];
  assign _EVAL_1837 = _EVAL_3862 | 16'h400;
  assign _EVAL_5240 = _EVAL_323 ? _EVAL_1837 : _EVAL_3862;
  assign _EVAL_4180 = {3'h0,_EVAL_2512,_EVAL_3742,_EVAL_2998,2'h2};
  assign _EVAL_1235 = _EVAL_3360 ? _EVAL_5240 : _EVAL_4180;
  assign _EVAL_4473 = _EVAL_5185 ? _EVAL_302 : _EVAL_1235;
  assign _EVAL_3674 = _EVAL_5363[1];
  assign _EVAL_3347 = _EVAL_735[9];
  assign _EVAL_4538 = _EVAL_735[4];
  assign _EVAL_4728 = _EVAL_735[6];
  assign _EVAL_5190 = _EVAL_735[8:7];
  assign _EVAL_3596 = {3'h3,_EVAL_3347,_EVAL_3742,_EVAL_4538,_EVAL_4728,_EVAL_5190,_EVAL_2512,2'h1};
  assign _EVAL_507 = {3'h2,_EVAL_2512,_EVAL_3742,_EVAL_2998,2'h1};
  assign _EVAL_2898 = _EVAL_3674 ? _EVAL_3596 : _EVAL_507;
  assign _EVAL_1227 = _EVAL_3742[3];
  assign _EVAL_4271 = _EVAL_2448 == 1'h0;
  assign _EVAL_2673 = _EVAL_1227 & _EVAL_4271;
  assign _EVAL_2128 = _EVAL_735[5:4];
  assign _EVAL_3490 = _EVAL_735[9:6];
  assign _EVAL_1618 = _EVAL_735[2];
  assign _EVAL_4886 = _EVAL_735[3];
  assign _EVAL_809 = _EVAL_3742[2:0];
  assign _EVAL_5250 = {3'h0,_EVAL_2128,_EVAL_3490,_EVAL_1618,_EVAL_4886,_EVAL_809,2'h0};
  assign _EVAL_2609 = {3'h0,_EVAL_2512,_EVAL_3742,_EVAL_2998,2'h1};
  assign _EVAL_4122 = _EVAL_2673 ? _EVAL_5250 : _EVAL_2609;
  assign _EVAL_1473 = _EVAL_2060 ? _EVAL_2898 : _EVAL_4122;
  assign _EVAL_338 = _EVAL_2359 ? _EVAL_4473 : _EVAL_1473;
  assign _EVAL_3714 = _EVAL_4614 == 5'h5;
  assign _EVAL_2090 = _EVAL_4614 == 5'h4;
  assign _EVAL_5353 = _EVAL_4614 == 5'h3;
  assign _EVAL_3566 = _EVAL_735[5:3];
  assign _EVAL_2696 = _EVAL_735[7:6];
  assign _EVAL_4798 = {3'h1,_EVAL_3566,_EVAL_4488,_EVAL_2696,_EVAL_809,2'h0};
  assign _EVAL_575 = _EVAL_735[4:3];
  assign _EVAL_2934 = _EVAL_735[8:6];
  assign _EVAL_3163 = {3'h1,_EVAL_2512,_EVAL_3742,_EVAL_575,_EVAL_2934,2'h2};
  assign _EVAL_4101 = _EVAL_2448 ? _EVAL_4798 : _EVAL_3163;
  assign _EVAL_1645 = {3'h3,_EVAL_3566,_EVAL_4488,_EVAL_1618,_EVAL_4728,_EVAL_809,2'h0};
  assign _EVAL_4186 = _EVAL_735[4:2];
  assign _EVAL_909 = {3'h3,_EVAL_2512,_EVAL_3742,_EVAL_4186,_EVAL_2696,2'h2};
  assign _EVAL_901 = _EVAL_2448 ? _EVAL_1645 : _EVAL_909;
  assign _EVAL_4303 = _EVAL_2359 ? _EVAL_4101 : _EVAL_901;
  assign _EVAL_2349 = _EVAL_4614 == 5'h2;
  assign _EVAL_1559 = {3'h3,_EVAL_3566,_EVAL_4488,_EVAL_2696,_EVAL_809,2'h0};
  assign _EVAL_452 = {3'h3,_EVAL_2512,_EVAL_3742,_EVAL_575,_EVAL_2934,2'h2};
  assign _EVAL_3530 = _EVAL_2448 ? _EVAL_1559 : _EVAL_452;
  assign _EVAL_5225 = {3'h2,_EVAL_3566,_EVAL_4488,_EVAL_1618,_EVAL_4728,_EVAL_809,2'h0};
  assign _EVAL_2910 = {3'h2,_EVAL_2512,_EVAL_3742,_EVAL_4186,_EVAL_2696,2'h2};
  assign _EVAL_4374 = _EVAL_2448 ? _EVAL_5225 : _EVAL_2910;
  assign _EVAL_837 = _EVAL_2359 ? _EVAL_3530 : _EVAL_4374;
  assign _EVAL_2008 = _EVAL_4614 == 5'h1;
  assign _EVAL_4307 = _EVAL_2008 ? _EVAL_4303 : _EVAL_837;
  assign _EVAL_421 = _EVAL_2349 ? _EVAL_837 : _EVAL_4307;
  assign _EVAL_1540 = _EVAL_5353 ? _EVAL_4303 : _EVAL_421;
  assign _EVAL_4257 = _EVAL_2090 ? _EVAL_338 : _EVAL_1540;
  assign _EVAL_876 = _EVAL_3714 ? _EVAL_2150 : _EVAL_4257;
  assign _EVAL_2401 = _EVAL_762 ? _EVAL_338 : _EVAL_876;
  assign _EVAL_1916 = _EVAL_1901 ? _EVAL_2150 : _EVAL_2401;
  assign _EVAL_4622 = _EVAL_4093 ? _EVAL_1704 : _EVAL_1916;
  assign _EVAL_3909 = _EVAL_850 ? _EVAL_771 : _EVAL_4622;
  assign _EVAL_1621 = _EVAL_3012 ? _EVAL_1704 : _EVAL_3909;
  assign _EVAL_4672 = _EVAL_780[2];
  assign _EVAL_4818 = _EVAL_4322[31];
  assign _EVAL_798 = _EVAL_4632 & _EVAL_4818;
  assign _EVAL_1036 = {_EVAL_798,_EVAL_4322};
  assign _EVAL_1929 = _EVAL_4322[31:16];
  assign _EVAL_2783 = {{16'd0}, _EVAL_1929};
  assign _EVAL_3710 = _EVAL_4322[15:0];
  assign _EVAL_5024 = {_EVAL_3710, 16'h0};
  assign _EVAL_4941 = _EVAL_5024 & 32'hffff0000;
  assign _EVAL_3898 = _EVAL_2783 | _EVAL_4941;
  assign _EVAL_3631 = _EVAL_3898[31:8];
  assign _EVAL_3245 = {{8'd0}, _EVAL_3631};
  assign _EVAL_4778 = _EVAL_3245 & 32'hff00ff;
  assign _EVAL_336 = _EVAL_3898[23:0];
  assign _EVAL_5332 = {_EVAL_336, 8'h0};
  assign _EVAL_1625 = _EVAL_5332 & 32'hff00ff00;
  assign _EVAL_5106 = _EVAL_4778 | _EVAL_1625;
  assign _EVAL_1132 = _EVAL_5106[31:4];
  assign _EVAL_1133 = {{4'd0}, _EVAL_1132};
  assign _EVAL_3317 = _EVAL_1133 & 32'hf0f0f0f;
  assign _EVAL_1658 = _EVAL_5106[27:0];
  assign _EVAL_1912 = {_EVAL_1658, 4'h0};
  assign _EVAL_4335 = _EVAL_1912 & 32'hf0f0f0f0;
  assign _EVAL_742 = _EVAL_3317 | _EVAL_4335;
  assign _EVAL_574 = _EVAL_742[31:2];
  assign _EVAL_533 = {{2'd0}, _EVAL_574};
  assign _EVAL_5218 = _EVAL_533 & 32'h33333333;
  assign _EVAL_4318 = _EVAL_742[29:0];
  assign _EVAL_988 = {_EVAL_4318, 2'h0};
  assign _EVAL_764 = _EVAL_988 & 32'hcccccccc;
  assign _EVAL_3666 = _EVAL_5218 | _EVAL_764;
  assign _EVAL_704 = _EVAL_3666[31:1];
  assign _EVAL_3881 = {{1'd0}, _EVAL_704};
  assign _EVAL_4973 = _EVAL_3881 & 32'h55555555;
  assign _EVAL_5305 = _EVAL_3666[30:0];
  assign _EVAL_5284 = {_EVAL_5305, 1'h0};
  assign _EVAL_3980 = _EVAL_5284 & 32'haaaaaaaa;
  assign _EVAL_1478 = _EVAL_4973 | _EVAL_3980;
  assign _EVAL_2935 = _EVAL_4672 ? _EVAL_1036 : {{1'd0}, _EVAL_1478};
  assign _EVAL_1307 = $signed(_EVAL_2935);
  assign _EVAL_2491 = _EVAL_4192[6];
  assign _EVAL_3148 = _EVAL_4135[0];
  assign _EVAL_4594 = _EVAL_4192[5:0];
  assign _EVAL_3209 = _EVAL_4135[4:1];
  assign _EVAL_4828 = {_EVAL_2491,_EVAL_3148,_EVAL_4594,_EVAL_3209,1'h0};
  assign _EVAL_3159 = $signed(_EVAL_4828);
  assign _EVAL_1303 = $unsigned(_EVAL_3159);
  assign _EVAL_5370 = _EVAL_1303[12];
  assign _EVAL_3852 = _EVAL_5370 ? 19'h7ffff : 19'h0;
  assign _EVAL_3471 = {_EVAL_3852,_EVAL_1303};
  assign _EVAL_3463 = _EVAL_4092 ? _EVAL_3471 : 32'h0;
  assign _EVAL_5389 = {_EVAL_4192,_EVAL_623,_EVAL_3053,_EVAL_1379};
  assign _EVAL_4334 = $signed(_EVAL_5389);
  assign _EVAL_3776 = _EVAL_4334[19];
  assign _EVAL_871 = _EVAL_4334[7:0];
  assign _EVAL_2127 = _EVAL_4334[8];
  assign _EVAL_2295 = _EVAL_4334[18:9];
  assign _EVAL_2044 = {_EVAL_3776,_EVAL_871,_EVAL_2127,_EVAL_2295,1'h0};
  assign _EVAL_4431 = $signed(_EVAL_2044);
  assign _EVAL_1194 = $unsigned(_EVAL_4431);
  assign _EVAL_2099 = _EVAL_1194[20];
  assign _EVAL_724 = _EVAL_2099 ? 11'h7ff : 11'h0;
  assign _EVAL_4791 = {_EVAL_724,_EVAL_1194};
  assign _EVAL_2629 = _EVAL_1915 ? _EVAL_4791 : 32'h0;
  assign _EVAL_1298 = _EVAL_3463 | _EVAL_2629;
  assign _EVAL_2826 = $unsigned(_EVAL_4334);
  assign _EVAL_3577 = {_EVAL_2826, 12'h0};
  assign _EVAL_547 = _EVAL_4684 ? _EVAL_3577 : 32'h0;
  assign _EVAL_3676 = _EVAL_1298 | _EVAL_547;
  assign _EVAL_3086 = {_EVAL_4192,_EVAL_623};
  assign _EVAL_5083 = $signed(_EVAL_3086);
  assign _EVAL_677 = $unsigned(_EVAL_5083);
  assign _EVAL_2431 = _EVAL_677[11];
  assign _EVAL_1723 = _EVAL_2431 ? 20'hfffff : 20'h0;
  assign _EVAL_3162 = {_EVAL_1723,_EVAL_677};
  assign _EVAL_5148 = _EVAL_2794 ? _EVAL_3162 : 32'h0;
  assign _EVAL_2101 = _EVAL_3676 | _EVAL_5148;
  assign _EVAL_2389 = _EVAL_494 ? _EVAL_3880 : 32'h0;
  assign _EVAL_3068 = _EVAL_2101 | _EVAL_2389;
  assign _EVAL_611 = _EVAL_3068[31:5];
  assign _EVAL_3166 = {_EVAL_611,_EVAL_498};
  assign _EVAL_1728 = _EVAL_3166[4:0];
  assign _EVAL_1064 = $signed(_EVAL_1307) >>> _EVAL_1728;
  assign _EVAL_4879 = _EVAL_1064[31:0];
  assign _EVAL_870 = _EVAL_4879[31:16];
  assign _EVAL_3696 = {{16'd0}, _EVAL_870};
  assign _EVAL_5144 = _EVAL_4879[15:0];
  assign _EVAL_5003 = {_EVAL_5144, 16'h0};
  assign _EVAL_4206 = _EVAL_5003 & 32'hffff0000;
  assign _EVAL_3389 = _EVAL_3696 | _EVAL_4206;
  assign _EVAL_4663 = _EVAL_3389[31:8];
  assign _EVAL_1919 = {{8'd0}, _EVAL_4663};
  assign _EVAL_3308 = _EVAL_1919 & 32'hff00ff;
  assign _EVAL_5266 = _EVAL_3389[23:0];
  assign _EVAL_1336 = {_EVAL_5266, 8'h0};
  assign _EVAL_2944 = _EVAL_1336 & 32'hff00ff00;
  assign _EVAL_1717 = _EVAL_3308 | _EVAL_2944;
  assign _EVAL_685 = _EVAL_1717[31:4];
  assign _EVAL_560 = {{4'd0}, _EVAL_685};
  assign _EVAL_3591 = _EVAL_560 & 32'hf0f0f0f;
  assign _EVAL_2626 = _EVAL_1717[27:0];
  assign _EVAL_474 = {_EVAL_2626, 4'h0};
  assign _EVAL_3954 = _EVAL_474 & 32'hf0f0f0f0;
  assign _EVAL_4182 = _EVAL_3591 | _EVAL_3954;
  assign _EVAL_551 = _EVAL_4182[29:0];
  assign _EVAL_5013 = {_EVAL_551, 2'h0};
  assign _EVAL_3293 = _EVAL_5013 & 32'hcccccccc;
  assign _EVAL_3243 = _EVAL_3373 == 3'h7;
  assign _EVAL_1323 = _EVAL_21[5];
  assign _EVAL_5115 = _EVAL_21[12:10];
  assign _EVAL_2565 = _EVAL_21[6];
  assign _EVAL_1143 = {_EVAL_1323,_EVAL_5115,_EVAL_2565,2'h0};
  assign _EVAL_1509 = _EVAL_1143[6:5];
  assign _EVAL_4942 = _EVAL_21[4:2];
  assign _EVAL_3048 = _EVAL_21[9:7];
  assign _EVAL_4841 = _EVAL_1143[4:0];
  assign _EVAL_1412 = {_EVAL_1509,2'h1,_EVAL_4942,2'h1,_EVAL_3048,3'h2,_EVAL_4841,7'h27};
  assign _EVAL_1631 = _EVAL_3373 == 3'h6;
  assign _EVAL_2447 = {_EVAL_1509,2'h1,_EVAL_4942,2'h1,_EVAL_3048,3'h2,_EVAL_4841,7'h23};
  assign _EVAL_5401 = _EVAL_21[6:5];
  assign _EVAL_1367 = {_EVAL_5401,_EVAL_5115,3'h0};
  assign _EVAL_369 = _EVAL_1367[7:5];
  assign _EVAL_2625 = _EVAL_1367[4:0];
  assign _EVAL_2802 = {_EVAL_369,2'h1,_EVAL_4942,2'h1,_EVAL_3048,3'h3,_EVAL_2625,7'h27};
  assign _EVAL_2350 = _EVAL_3373 == 3'h4;
  assign _EVAL_2985 = {_EVAL_1509,2'h1,_EVAL_4942,2'h1,_EVAL_3048,3'h0,_EVAL_4841,7'h27};
  assign _EVAL_1023 = _EVAL_3373 == 3'h3;
  assign _EVAL_1474 = {_EVAL_1323,_EVAL_5115,_EVAL_2565,2'h0,2'h1,_EVAL_3048,3'h2,2'h1,_EVAL_4942,7'h7};
  assign _EVAL_5398 = _EVAL_3373 == 3'h2;
  assign _EVAL_1890 = {_EVAL_1323,_EVAL_5115,_EVAL_2565,2'h0,2'h1,_EVAL_3048,3'h2,2'h1,_EVAL_4942,7'h3};
  assign _EVAL_2854 = _EVAL_3373 == 3'h1;
  assign _EVAL_4965 = {_EVAL_5401,_EVAL_5115,3'h0,2'h1,_EVAL_3048,3'h3,2'h1,_EVAL_4942,7'h7};
  assign _EVAL_5292 = _EVAL_21[10:7];
  assign _EVAL_738 = _EVAL_21[12:11];
  assign _EVAL_1528 = {_EVAL_5292,_EVAL_738,_EVAL_1323,_EVAL_2565,2'h0,5'h2,3'h0,2'h1,_EVAL_4942,7'h13};
  assign _EVAL_3228 = _EVAL_2854 ? {{2'd0}, _EVAL_4965} : _EVAL_1528;
  assign _EVAL_895 = _EVAL_5398 ? {{3'd0}, _EVAL_1890} : _EVAL_3228;
  assign _EVAL_3394 = _EVAL_1023 ? {{3'd0}, _EVAL_1474} : _EVAL_895;
  assign _EVAL_5293 = _EVAL_2350 ? {{3'd0}, _EVAL_2985} : _EVAL_3394;
  assign _EVAL_4697 = _EVAL_2034 ? {{2'd0}, _EVAL_2802} : _EVAL_5293;
  assign _EVAL_4398 = _EVAL_1631 ? {{3'd0}, _EVAL_2447} : _EVAL_4697;
  assign _EVAL_3828 = _EVAL_3243 ? {{3'd0}, _EVAL_1412} : _EVAL_4398;
  assign _EVAL_4329 = {2'h0,_EVAL_3828};
  assign _EVAL_841 = _EVAL_4329 & 32'h28;
  assign _EVAL_5130 = _EVAL_3309 == 5'h1a;
  assign _EVAL_2460 = _EVAL_1445[8];
  assign _EVAL_4593 = _EVAL_1445[7:6];
  assign _EVAL_2015 = _EVAL_1445[2:1];
  assign _EVAL_3205 = _EVAL_1445[5];
  assign _EVAL_2376 = {3'h6,_EVAL_2460,_EVAL_3957,_EVAL_4494,_EVAL_4593,_EVAL_2015,_EVAL_3205,2'h1};
  assign _EVAL_2137 = {_EVAL_3755, 13'h0};
  assign _EVAL_4998 = {{2'd0}, _EVAL_2137};
  assign _EVAL_1571 = _EVAL_2376 | _EVAL_4998;
  assign _EVAL_309 = _EVAL_3309 == 5'h19;
  assign _EVAL_2158 = {4'h8,_EVAL_4715,_EVAL_1198,2'h2};
  assign _EVAL_2407 = _EVAL_4706[0];
  assign _EVAL_1280 = {_EVAL_2407, 12'h0};
  assign _EVAL_1203 = {{3'd0}, _EVAL_1280};
  assign _EVAL_2252 = _EVAL_2158 | _EVAL_1203;
  assign _EVAL_1604 = _EVAL_3309 == 5'h18;
  assign _EVAL_1066 = _EVAL_3309 == 5'h17;
  assign _EVAL_866 = ~ _EVAL_2158;
  assign _EVAL_3402 = _EVAL_866 | 16'h4;
  assign _EVAL_3557 = ~ _EVAL_3402;
  assign _EVAL_1407 = _EVAL_3557 | 16'h1000;
  assign _EVAL_298 = _EVAL_3309 == 5'h16;
  assign _EVAL_2781 = _EVAL_3309 == 5'h15;
  assign _EVAL_4245 = _EVAL_3309 == 5'h14;
  assign _EVAL_4228 = _EVAL_3309 == 5'h13;
  assign _EVAL_5072 = {_EVAL_4019,_EVAL_1198,_EVAL_4715,_EVAL_4201};
  assign _EVAL_409 = $signed(_EVAL_5072);
  assign _EVAL_4086 = _EVAL_409[19];
  assign _EVAL_4877 = _EVAL_409[12];
  assign _EVAL_1136 = _EVAL_409[17:16];
  assign _EVAL_2143 = _EVAL_409[18];
  assign _EVAL_1761 = _EVAL_409[14];
  assign _EVAL_1369 = _EVAL_409[15];
  assign _EVAL_5061 = _EVAL_409[11:9];
  assign _EVAL_3192 = _EVAL_409[13];
  assign _EVAL_4660 = {3'h5,_EVAL_4086,_EVAL_4877,_EVAL_1136,_EVAL_2143,_EVAL_1761,_EVAL_1369,_EVAL_5061,_EVAL_3192,2'h1};
  assign _EVAL_4933 = ~ _EVAL_4660;
  assign _EVAL_828 = {_EVAL_2407, 15'h0};
  assign _EVAL_2721 = _EVAL_4933 | _EVAL_828;
  assign _EVAL_1703 = ~ _EVAL_2721;
  assign _EVAL_3707 = _EVAL_3309 == 5'h12;
  assign _EVAL_1881 = _EVAL_3309 == 5'h11;
  assign _EVAL_3233 = _EVAL_3309 == 5'h10;
  assign _EVAL_1318 = _EVAL_3309 == 5'hf;
  assign _EVAL_3849 = _EVAL_409[4:0];
  assign _EVAL_960 = {3'h3,_EVAL_4086,_EVAL_4706,_EVAL_3849,2'h1};
  assign _EVAL_1825 = _EVAL_3309 == 5'he;
  assign _EVAL_2669 = _EVAL_4201[1];
  assign _EVAL_4779 = _EVAL_2669 == 1'h0;
  assign _EVAL_1290 = _EVAL_4019[5];
  assign _EVAL_2126 = _EVAL_1290 == 1'h0;
  assign _EVAL_4954 = _EVAL_4779 & _EVAL_2126;
  assign _EVAL_830 = _EVAL_3755 | _EVAL_4954;
  assign _EVAL_3167 = _EVAL_1198[2:0];
  assign _EVAL_2075 = {6'h27,_EVAL_4494,_EVAL_2669,_EVAL_830,_EVAL_3167,2'h1};
  assign _EVAL_2552 = _EVAL_3309 == 5'hd;
  assign _EVAL_281 = _EVAL_3309 == 5'hc;
  assign _EVAL_3788 = _EVAL_4201[2];
  assign _EVAL_2602 = _EVAL_3788 & _EVAL_1120;
  assign _EVAL_4814 = _EVAL_2602 | _EVAL_1290;
  assign _EVAL_3147 = _EVAL_4779 & _EVAL_3788;
  assign _EVAL_1188 = _EVAL_3755 | _EVAL_3147;
  assign _EVAL_1842 = {6'h23,_EVAL_4494,_EVAL_2669,_EVAL_1188,_EVAL_3167,2'h1};
  assign _EVAL_3656 = {4'h8,_EVAL_4706,_EVAL_1198,2'h2};
  assign _EVAL_3684 = _EVAL_3656 | 16'h1000;
  assign _EVAL_2732 = _EVAL_3788 ? _EVAL_3656 : _EVAL_3684;
  assign _EVAL_3507 = _EVAL_4814 ? _EVAL_1842 : _EVAL_2732;
  assign _EVAL_2070 = _EVAL_3309 == 5'hb;
  assign _EVAL_3173 = _EVAL_1445[5:3];
  assign _EVAL_1859 = {3'h5,_EVAL_3173,_EVAL_4494,_EVAL_4593,_EVAL_3167,2'h0};
  assign _EVAL_5021 = _EVAL_1445[8:6];
  assign _EVAL_3248 = {3'h5,_EVAL_3173,_EVAL_5021,_EVAL_1198,2'h2};
  assign _EVAL_3797 = _EVAL_1120 ? _EVAL_1859 : _EVAL_3248;
  assign _EVAL_522 = _EVAL_1445[2];
  assign _EVAL_4040 = _EVAL_1445[6];
  assign _EVAL_1308 = {3'h7,_EVAL_3173,_EVAL_4494,_EVAL_522,_EVAL_4040,_EVAL_3167,2'h0};
  assign _EVAL_5030 = _EVAL_1445[5:2];
  assign _EVAL_3546 = {3'h7,_EVAL_5030,_EVAL_4593,_EVAL_1198,2'h2};
  assign _EVAL_4050 = _EVAL_1120 ? _EVAL_1308 : _EVAL_3546;
  assign _EVAL_1233 = _EVAL_3755 ? _EVAL_3797 : _EVAL_4050;
  assign _EVAL_1569 = {3'h4,_EVAL_3173,_EVAL_4494,_EVAL_522,_EVAL_4040,_EVAL_3167,2'h0};
  assign _EVAL_4952 = _EVAL_2669 ? _EVAL_1233 : _EVAL_1569;
  assign _EVAL_3268 = _EVAL_3309 == 5'ha;
  assign _EVAL_2042 = {3'h7,_EVAL_3173,_EVAL_4494,_EVAL_4593,_EVAL_3167,2'h0};
  assign _EVAL_2002 = {3'h7,_EVAL_3173,_EVAL_5021,_EVAL_1198,2'h2};
  assign _EVAL_776 = _EVAL_1120 ? _EVAL_2042 : _EVAL_2002;
  assign _EVAL_2716 = {3'h6,_EVAL_3173,_EVAL_4494,_EVAL_522,_EVAL_4040,_EVAL_3167,2'h0};
  assign _EVAL_598 = {3'h6,_EVAL_5030,_EVAL_4593,_EVAL_1198,2'h2};
  assign _EVAL_4241 = _EVAL_1120 ? _EVAL_2716 : _EVAL_598;
  assign _EVAL_1503 = _EVAL_3755 ? _EVAL_776 : _EVAL_4241;
  assign _EVAL_424 = _EVAL_3309 == 5'h9;
  assign _EVAL_1096 = _EVAL_3309 == 5'h8;
  assign _EVAL_1378 = _EVAL_3309 == 5'h7;
  assign _EVAL_499 = _EVAL_3309 == 5'h6;
  assign _EVAL_4588 = _EVAL_5246[4:0];
  assign _EVAL_4424 = {3'h4,_EVAL_4395,2'h0,_EVAL_4494,_EVAL_4588,2'h1};
  assign _EVAL_3879 = _EVAL_4424 | 16'h800;
  assign _EVAL_2420 = _EVAL_4424 | 16'h400;
  assign _EVAL_1364 = _EVAL_1290 ? _EVAL_2420 : _EVAL_4424;
  assign _EVAL_1545 = {3'h0,_EVAL_4395,_EVAL_4706,_EVAL_4588,2'h2};
  assign _EVAL_4712 = _EVAL_3788 ? _EVAL_1364 : _EVAL_1545;
  assign _EVAL_4391 = _EVAL_2669 ? _EVAL_3879 : _EVAL_4712;
  assign _EVAL_388 = _EVAL_4715[1];
  assign _EVAL_2404 = _EVAL_5246[9];
  assign _EVAL_3691 = _EVAL_5246[4];
  assign _EVAL_4229 = _EVAL_5246[8:7];
  assign _EVAL_2485 = {3'h3,_EVAL_2404,_EVAL_4706,_EVAL_3691,_EVAL_3661,_EVAL_4229,_EVAL_4395,2'h1};
  assign _EVAL_2762 = {3'h2,_EVAL_4395,_EVAL_4706,_EVAL_4588,2'h1};
  assign _EVAL_5134 = _EVAL_388 ? _EVAL_2485 : _EVAL_2762;
  assign _EVAL_2958 = _EVAL_4706[3];
  assign _EVAL_3326 = _EVAL_1120 == 1'h0;
  assign _EVAL_4326 = _EVAL_2958 & _EVAL_3326;
  assign _EVAL_864 = _EVAL_5246[5:4];
  assign _EVAL_2550 = _EVAL_5246[9:6];
  assign _EVAL_2027 = _EVAL_5246[3];
  assign _EVAL_413 = {3'h0,_EVAL_864,_EVAL_2550,_EVAL_556,_EVAL_2027,_EVAL_5219,2'h0};
  assign _EVAL_3274 = {3'h0,_EVAL_4395,_EVAL_4706,_EVAL_4588,2'h1};
  assign _EVAL_1960 = _EVAL_4326 ? _EVAL_413 : _EVAL_3274;
  assign _EVAL_5020 = _EVAL_4796 ? _EVAL_5134 : _EVAL_1960;
  assign _EVAL_3789 = _EVAL_3755 ? _EVAL_4391 : _EVAL_5020;
  assign _EVAL_3759 = _EVAL_3309 == 5'h5;
  assign _EVAL_2866 = _EVAL_3309 == 5'h4;
  assign _EVAL_613 = _EVAL_3309 == 5'h3;
  assign _EVAL_2720 = {3'h1,_EVAL_2208,_EVAL_4494,_EVAL_4757,_EVAL_5219,2'h0};
  assign _EVAL_3897 = {3'h1,_EVAL_4395,_EVAL_4706,_EVAL_1958,_EVAL_927,2'h2};
  assign _EVAL_3638 = _EVAL_1120 ? _EVAL_2720 : _EVAL_3897;
  assign _EVAL_616 = {3'h3,_EVAL_2208,_EVAL_4494,_EVAL_556,_EVAL_3661,_EVAL_5219,2'h0};
  assign _EVAL_4768 = {3'h3,_EVAL_4395,_EVAL_4706,_EVAL_2874,_EVAL_4757,2'h2};
  assign _EVAL_1069 = _EVAL_1120 ? _EVAL_616 : _EVAL_4768;
  assign _EVAL_2895 = _EVAL_3755 ? _EVAL_3638 : _EVAL_1069;
  assign _EVAL_2634 = _EVAL_3309 == 5'h2;
  assign _EVAL_1208 = _EVAL_3309 == 5'h1;
  assign _EVAL_1090 = _EVAL_1208 ? _EVAL_2895 : _EVAL_5236;
  assign _EVAL_2872 = _EVAL_2634 ? _EVAL_5236 : _EVAL_1090;
  assign _EVAL_3964 = _EVAL_613 ? _EVAL_2895 : _EVAL_2872;
  assign _EVAL_2347 = _EVAL_2866 ? _EVAL_3789 : _EVAL_3964;
  assign _EVAL_1534 = _EVAL_3759 ? _EVAL_960 : _EVAL_2347;
  assign _EVAL_1615 = _EVAL_499 ? _EVAL_3789 : _EVAL_1534;
  assign _EVAL_3804 = _EVAL_1378 ? _EVAL_960 : _EVAL_1615;
  assign _EVAL_4522 = _EVAL_1096 ? _EVAL_1503 : _EVAL_3804;
  assign _EVAL_3990 = _EVAL_424 ? _EVAL_4952 : _EVAL_4522;
  assign _EVAL_4396 = _EVAL_3268 ? _EVAL_1503 : _EVAL_3990;
  assign _EVAL_1039 = _EVAL_2070 ? _EVAL_4952 : _EVAL_4396;
  assign _EVAL_1630 = _EVAL_281 ? _EVAL_3507 : _EVAL_1039;
  assign _EVAL_4295 = _EVAL_2552 ? _EVAL_960 : _EVAL_1630;
  assign _EVAL_2903 = _EVAL_1825 ? _EVAL_2075 : _EVAL_4295;
  assign _EVAL_4418 = _EVAL_1318 ? _EVAL_960 : _EVAL_2903;
  assign _EVAL_1949 = _EVAL_3233 ? _EVAL_1571 : _EVAL_4418;
  assign _EVAL_926 = _EVAL_1881 ? _EVAL_2252 : _EVAL_1949;
  assign _EVAL_5299 = _EVAL_3707 ? _EVAL_1571 : _EVAL_926;
  assign _EVAL_3420 = _EVAL_4228 ? _EVAL_1703 : _EVAL_5299;
  assign _EVAL_880 = _EVAL_4245 ? _EVAL_1407 : _EVAL_3420;
  assign _EVAL_4126 = _EVAL_2781 ? _EVAL_1407 : _EVAL_880;
  assign _EVAL_4161 = _EVAL_298 ? _EVAL_1407 : _EVAL_4126;
  assign _EVAL_1192 = _EVAL_1066 ? _EVAL_1407 : _EVAL_4161;
  assign _EVAL_5381 = _EVAL_1604 ? _EVAL_1571 : _EVAL_1192;
  assign _EVAL_2130 = _EVAL_309 ? _EVAL_2252 : _EVAL_5381;
  assign _EVAL_5018 = _EVAL_5130 ? _EVAL_1571 : _EVAL_2130;
  assign _EVAL_1492 = _EVAL_191[4:2];
  assign _EVAL_3226 = _EVAL_1492 == 3'h7;
  assign _EVAL_5197 = _EVAL_6[4:2];
  assign _EVAL_1661 = _EVAL_5197 == 3'h7;
  assign _EVAL_327 = _EVAL_315 ? _EVAL_3226 : _EVAL_1661;
  assign _EVAL_4820 = _EVAL_2118 | _EVAL_4240;
  assign _EVAL_3605 = _EVAL_4820 | _EVAL_2326;
  assign _EVAL_4811 = _EVAL_3605 | _EVAL_3624;
  assign _EVAL_2372 = _EVAL_4811 | _EVAL_2506;
  assign _EVAL_3497 = _EVAL_2372 | _EVAL_3227;
  assign _EVAL_3528 = _EVAL_327 & _EVAL_3497;
  assign _EVAL_1083 = _EVAL_3608 | _EVAL_2853;
  assign _EVAL_4047 = _EVAL_5197 == 3'h6;
  assign _EVAL_469 = _EVAL_1492 == 3'h6;
  assign _EVAL_1588 = _EVAL_315 ? _EVAL_4047 : _EVAL_469;
  assign _EVAL_725 = _EVAL_315 ? _EVAL_205 : _EVAL_1;
  assign _EVAL_405 = _EVAL_725 == 1'h0;
  assign _EVAL_1922 = _EVAL_315 ? _EVAL_250 : _EVAL_141;
  assign _EVAL_1324 = _EVAL_405 | _EVAL_1922;
  assign _EVAL_2977 = _EVAL_1588 & _EVAL_1324;
  assign _EVAL_4832 = _EVAL_315 ? _EVAL_6 : _EVAL_191;
  assign _EVAL_3255 = _EVAL_4832[3];
  assign _EVAL_5262 = _EVAL_3255 == 1'h0;
  assign _EVAL_2162 = _EVAL_405 & _EVAL_5262;
  assign _EVAL_4065 = _EVAL_2977 | _EVAL_2162;
  assign _EVAL_4099 = _EVAL_315 ? _EVAL_2 : _EVAL_138;
  assign _EVAL_1420 = _EVAL_4065 ? _EVAL_4099 : 32'h0;
  assign _EVAL_5283 = _EVAL_6[4];
  assign _EVAL_930 = _EVAL_653 | _EVAL_3747;
  assign _EVAL_4803 = _EVAL_2118 & _EVAL_930;
  assign _EVAL_5082 = fpu__EVAL_26 == _EVAL_4745;
  assign _EVAL_3160 = _EVAL_4182[31:2];
  assign _EVAL_5181 = {{2'd0}, _EVAL_3160};
  assign _EVAL_2215 = _EVAL_5181 & 32'h33333333;
  assign _EVAL_4983 = _EVAL_2215 | _EVAL_3293;
  assign _EVAL_4752 = _EVAL_4983[30:0];
  assign _EVAL_998 = fpu__EVAL_29 == _EVAL_4745;
  assign _EVAL_4282 = $signed(_EVAL_1445);
  assign _EVAL_1609 = $signed(_EVAL_5246);
  assign _EVAL_3952 = _EVAL_3858 ? $signed(_EVAL_4282) : $signed(_EVAL_1609);
  assign _EVAL_3781 = $unsigned(_EVAL_3952);
  assign _EVAL_431 = _EVAL_3781[11];
  assign _EVAL_1766 = _EVAL_431 ? 20'hfffff : 20'h0;
  assign _EVAL_5112 = {_EVAL_1766,_EVAL_3781};
  assign _EVAL_3978 = _EVAL_5017 ? _EVAL_5112 : 32'h0;
  assign _EVAL_1643 = _EVAL_3415 ? _EVAL_4748 : 32'h0;
  assign _EVAL_2046 = _EVAL_3978 | _EVAL_1643;
  assign _EVAL_2567 = _EVAL_2046[31:5];
  assign _EVAL_1155 = {_EVAL_2567,_EVAL_1415};
  assign _EVAL_3869 = ~ _EVAL_1155;
  assign _EVAL_3901 = _EVAL_2282 ? _EVAL_3869 : _EVAL_1155;
  assign _EVAL_4503 = {_EVAL_3901,_EVAL_2282};
  assign _EVAL_3910 = _EVAL_3309[4];
  assign _EVAL_4705 = _EVAL_3910 == 1'h0;
  assign _EVAL_2923 = _EVAL_3309[3];
  assign _EVAL_1988 = _EVAL_4705 & _EVAL_2923;
  assign _EVAL_1400 = _EVAL_3309[1];
  assign _EVAL_3618 = _EVAL_1400 == 1'h0;
  assign _EVAL_345 = _EVAL_1988 & _EVAL_3618;
  assign _EVAL_3817 = _EVAL_1446 & _EVAL_345;
  assign _EVAL_873 = _EVAL_3309[0];
  assign _EVAL_2037 = _EVAL_345 & _EVAL_873;
  assign _EVAL_1162 = _EVAL_1446 & _EVAL_2037;
  assign _EVAL_1291 = _EVAL_1162 == 1'h0;
  assign _EVAL_4072 = _EVAL_3817 & _EVAL_1291;
  assign _EVAL_4872 = _EVAL_1452[0];
  assign _EVAL_2237 = _EVAL_4299 & _EVAL_119;
  assign _EVAL_4231 = _EVAL_4127 == _EVAL_4135;
  assign _EVAL_286 = _EVAL_2237 & _EVAL_4231;
  assign _EVAL_2560 = _EVAL_21[12];
  assign _EVAL_428 = _EVAL_2560 ? 15'h7fff : 15'h0;
  assign _EVAL_1302 = _EVAL_21[6:2];
  assign _EVAL_4377 = {_EVAL_428,_EVAL_1302,12'h0};
  assign _EVAL_1125 = _EVAL_58 & _EVAL_3747;
  assign _EVAL_1022 = _EVAL_268 & _EVAL_653;
  assign _EVAL_4450 = _EVAL_1125 | _EVAL_1022;
  assign _EVAL_4483 = _EVAL_91 == _EVAL_2579;
  assign _EVAL_5224 = _EVAL_4450 & _EVAL_4483;
  assign _EVAL_4552 = _EVAL_16 & _EVAL_3747;
  assign _EVAL_462 = _EVAL_214 & _EVAL_653;
  assign _EVAL_3600 = _EVAL_4552 | _EVAL_462;
  assign _EVAL_4719 = _EVAL_171 == _EVAL_2579;
  assign _EVAL_3907 = _EVAL_3600 & _EVAL_4719;
  assign _EVAL_2847 = _EVAL_315 ? _EVAL_5224 : _EVAL_3907;
  assign _EVAL_557 = _EVAL_4064[0];
  assign _EVAL_1123 = $signed(_EVAL_735);
  assign _EVAL_3252 = $unsigned(_EVAL_1123);
  assign _EVAL_2929 = _EVAL_3252[11];
  assign _EVAL_938 = _EVAL_2929 ? 20'hfffff : 20'h0;
  assign _EVAL_5254 = {_EVAL_938,_EVAL_3252};
  assign _EVAL_3324 = _EVAL_380 ? _EVAL_5254 : 32'h0;
  assign _EVAL_644 = _EVAL_4790 ? _EVAL_4373 : 32'h0;
  assign _EVAL_1057 = _EVAL_3324 | _EVAL_644;
  assign _EVAL_4969 = _EVAL_1057[31:5];
  assign _EVAL_1731 = {_EVAL_4969,_EVAL_3370};
  assign _EVAL_2612 = ~ _EVAL_1731;
  assign _EVAL_3977 = _EVAL_1818 ? _EVAL_2612 : _EVAL_1731;
  assign _EVAL_4572 = _EVAL_3977[31];
  assign _EVAL_2471 = _EVAL_4572 == 1'h0;
  assign _EVAL_2951 = _EVAL_1699 ? _EVAL_5043 : _EVAL_2758;
  assign _EVAL_4659 = _EVAL_2951[31:5];
  assign _EVAL_1483 = {_EVAL_4659,_EVAL_2683};
  assign _EVAL_1102 = _EVAL_1483[31];
  assign _EVAL_354 = _EVAL_557 ? _EVAL_2471 : _EVAL_1102;
  assign _EVAL_4294 = _EVAL_4614 == 5'h1f;
  assign _EVAL_1106 = {4'h8,_EVAL_5363,_EVAL_1641,2'h2};
  assign _EVAL_3089 = ~ _EVAL_1106;
  assign _EVAL_2970 = _EVAL_3089 | 16'h4;
  assign _EVAL_2813 = ~ _EVAL_2970;
  assign _EVAL_3549 = _EVAL_2813 | 16'h1000;
  assign _EVAL_3535 = _EVAL_4614 == 5'h1e;
  assign _EVAL_2106 = _EVAL_4614 == 5'h1d;
  assign _EVAL_2671 = _EVAL_4614 == 5'h1c;
  assign _EVAL_3628 = _EVAL_4614 == 5'h1b;
  assign _EVAL_1220 = _EVAL_2904[12];
  assign _EVAL_5186 = _EVAL_2904[17:16];
  assign _EVAL_3959 = _EVAL_2904[18];
  assign _EVAL_2791 = _EVAL_2904[14];
  assign _EVAL_2430 = _EVAL_2904[15];
  assign _EVAL_3499 = _EVAL_2904[11:9];
  assign _EVAL_4644 = _EVAL_2904[13];
  assign _EVAL_2214 = {3'h5,_EVAL_2801,_EVAL_1220,_EVAL_5186,_EVAL_3959,_EVAL_2791,_EVAL_2430,_EVAL_3499,_EVAL_4644,2'h1};
  assign _EVAL_1567 = ~ _EVAL_2214;
  assign _EVAL_1749 = _EVAL_3742[0];
  assign _EVAL_4747 = {_EVAL_1749, 15'h0};
  assign _EVAL_4498 = _EVAL_1567 | _EVAL_4747;
  assign _EVAL_2737 = ~ _EVAL_4498;
  assign _EVAL_5195 = _EVAL_4614 == 5'h1a;
  assign _EVAL_4925 = _EVAL_1542[8];
  assign _EVAL_4843 = _EVAL_1542[4:3];
  assign _EVAL_1266 = _EVAL_1542[2:1];
  assign _EVAL_1636 = _EVAL_1542[5];
  assign _EVAL_3461 = {3'h6,_EVAL_4925,_EVAL_4843,_EVAL_4488,_EVAL_3551,_EVAL_1266,_EVAL_1636,2'h1};
  assign _EVAL_2608 = {_EVAL_2359, 13'h0};
  assign _EVAL_4781 = {{2'd0}, _EVAL_2608};
  assign _EVAL_2009 = _EVAL_3461 | _EVAL_4781;
  assign _EVAL_1551 = _EVAL_4614 == 5'h19;
  assign _EVAL_979 = {_EVAL_1749, 12'h0};
  assign _EVAL_2021 = {{3'd0}, _EVAL_979};
  assign _EVAL_1327 = _EVAL_1106 | _EVAL_2021;
  assign _EVAL_1600 = _EVAL_4614 == 5'h18;
  assign _EVAL_659 = _EVAL_4614 == 5'h17;
  assign _EVAL_4147 = _EVAL_4614 == 5'h16;
  assign _EVAL_5065 = _EVAL_4614 == 5'h15;
  assign _EVAL_322 = _EVAL_4614 == 5'h14;
  assign _EVAL_4615 = _EVAL_4614 == 5'h13;
  assign _EVAL_2878 = _EVAL_4614 == 5'h12;
  assign _EVAL_4707 = _EVAL_4614 == 5'h11;
  assign _EVAL_2475 = _EVAL_4614 == 5'h10;
  assign _EVAL_2939 = _EVAL_4614 == 5'hf;
  assign _EVAL_3164 = _EVAL_4614 == 5'he;
  assign _EVAL_2599 = _EVAL_5185 == 1'h0;
  assign _EVAL_1500 = _EVAL_323 == 1'h0;
  assign _EVAL_1179 = _EVAL_2599 & _EVAL_1500;
  assign _EVAL_314 = _EVAL_2359 | _EVAL_1179;
  assign _EVAL_4416 = {6'h27,_EVAL_4488,_EVAL_5185,_EVAL_314,_EVAL_2846,2'h1};
  assign _EVAL_603 = _EVAL_4614 == 5'hd;
  assign _EVAL_2309 = _EVAL_4614 == 5'hc;
  assign _EVAL_1911 = _EVAL_3360 & _EVAL_2448;
  assign _EVAL_3561 = _EVAL_1911 | _EVAL_323;
  assign _EVAL_2413 = _EVAL_2599 & _EVAL_3360;
  assign _EVAL_3965 = _EVAL_2359 | _EVAL_2413;
  assign _EVAL_2695 = {6'h23,_EVAL_4488,_EVAL_5185,_EVAL_3965,_EVAL_2846,2'h1};
  assign _EVAL_4026 = {4'h8,_EVAL_3742,_EVAL_1641,2'h2};
  assign _EVAL_3193 = _EVAL_4026 | 16'h1000;
  assign _EVAL_4049 = _EVAL_3360 ? _EVAL_4026 : _EVAL_3193;
  assign _EVAL_3330 = _EVAL_3561 ? _EVAL_2695 : _EVAL_4049;
  assign _EVAL_404 = _EVAL_4614 == 5'hb;
  assign _EVAL_1999 = _EVAL_404 ? _EVAL_771 : _EVAL_1621;
  assign _EVAL_1404 = _EVAL_2309 ? _EVAL_3330 : _EVAL_1999;
  assign _EVAL_3800 = _EVAL_603 ? _EVAL_2150 : _EVAL_1404;
  assign _EVAL_794 = _EVAL_3164 ? _EVAL_4416 : _EVAL_3800;
  assign _EVAL_2230 = _EVAL_2939 ? _EVAL_2150 : _EVAL_794;
  assign _EVAL_1899 = _EVAL_2475 ? _EVAL_2009 : _EVAL_2230;
  assign _EVAL_461 = _EVAL_4707 ? _EVAL_1327 : _EVAL_1899;
  assign _EVAL_4591 = _EVAL_2878 ? _EVAL_2009 : _EVAL_461;
  assign _EVAL_342 = _EVAL_4615 ? _EVAL_2737 : _EVAL_4591;
  assign _EVAL_4394 = _EVAL_322 ? _EVAL_3549 : _EVAL_342;
  assign _EVAL_2885 = _EVAL_5065 ? _EVAL_3549 : _EVAL_4394;
  assign _EVAL_863 = _EVAL_4147 ? _EVAL_3549 : _EVAL_2885;
  assign _EVAL_3585 = _EVAL_659 ? _EVAL_3549 : _EVAL_863;
  assign _EVAL_4254 = _EVAL_1600 ? _EVAL_2009 : _EVAL_3585;
  assign _EVAL_4898 = _EVAL_1551 ? _EVAL_1327 : _EVAL_4254;
  assign _EVAL_5264 = _EVAL_5195 ? _EVAL_2009 : _EVAL_4898;
  assign _EVAL_4675 = _EVAL_3628 ? _EVAL_2737 : _EVAL_5264;
  assign _EVAL_577 = _EVAL_2671 ? _EVAL_3549 : _EVAL_4675;
  assign _EVAL_1914 = _EVAL_2106 ? _EVAL_3549 : _EVAL_577;
  assign _EVAL_3992 = _EVAL_3535 ? _EVAL_3549 : _EVAL_1914;
  assign _EVAL_1032 = _EVAL_4294 ? _EVAL_3549 : _EVAL_3992;
  assign _EVAL_4961 = {_EVAL_3229,_EVAL_1641,_EVAL_5363,_EVAL_1024,_EVAL_3742,_EVAL_4614,2'h3};
  assign _EVAL_3745 = _EVAL_2573 & _EVAL_148;
  assign _EVAL_1525 = _EVAL_1724 & _EVAL_1;
  assign _EVAL_1527 = _EVAL_3745 | _EVAL_1525;
  assign _EVAL_578 = _EVAL_3742 == _EVAL_2193;
  assign _EVAL_5093 = _EVAL_2219 & _EVAL_578;
  assign _EVAL_3035 = _EVAL_98 ? _EVAL_165 : _EVAL_204;
  assign _EVAL_1593 = _EVAL_98 ? _EVAL_212 : _EVAL_92;
  assign _EVAL_2785 = _EVAL_3035 | _EVAL_1593;
  assign _EVAL_663 = _EVAL_98 ? _EVAL_32 : _EVAL_80;
  assign _EVAL_1868 = _EVAL_2785 | _EVAL_663;
  assign _EVAL_1957 = _EVAL_98 ? _EVAL_172 : _EVAL_213;
  assign _EVAL_1348 = _EVAL_1868 | _EVAL_1957;
  assign _EVAL_2077 = _EVAL_98 ? _EVAL_40 : _EVAL_59;
  assign _EVAL_4458 = _EVAL_2077 == 1'h0;
  assign _EVAL_2236 = _EVAL_98 ? _EVAL_58 : _EVAL_16;
  assign _EVAL_1010 = _EVAL_98 ? _EVAL_148 : _EVAL_39;
  assign _EVAL_513 = _EVAL_2236 | _EVAL_1010;
  assign _EVAL_1690 = _EVAL_98 ? _EVAL_179 : _EVAL_188;
  assign _EVAL_4626 = _EVAL_513 | _EVAL_1690;
  assign _EVAL_4193 = _EVAL_98 ? _EVAL_153 : _EVAL_84;
  assign _EVAL_1270 = _EVAL_4193 == 3'h5;
  assign _EVAL_1970 = _EVAL_4193 == 3'h6;
  assign _EVAL_5316 = _EVAL_1270 | _EVAL_1970;
  assign _EVAL_4384 = csr__EVAL_134 | _EVAL_5316;
  assign _EVAL_4448 = _EVAL_4193 == 3'h7;
  assign _EVAL_1144 = csr__EVAL_99 >= 3'h5;
  assign _EVAL_2125 = _EVAL_4448 & _EVAL_1144;
  assign _EVAL_4339 = _EVAL_4384 | _EVAL_2125;
  assign _EVAL_4765 = _EVAL_4626 & _EVAL_4339;
  assign _EVAL_1501 = _EVAL_4458 | _EVAL_4765;
  assign _EVAL_4726 = _EVAL_98 ? _EVAL_1 : _EVAL_205;
  assign _EVAL_480 = _EVAL_98 ? _EVAL_154 : _EVAL_274;
  assign _EVAL_5006 = _EVAL_480 != _EVAL_480;
  assign _EVAL_5163 = _EVAL_4726 & _EVAL_5006;
  assign _EVAL_4577 = _EVAL_98 ? _EVAL_141 : _EVAL_250;
  assign _EVAL_4305 = _EVAL_98 ? _EVAL_68 : _EVAL_180;
  assign _EVAL_1019 = _EVAL_4305 != _EVAL_4305;
  assign _EVAL_2718 = _EVAL_4577 & _EVAL_1019;
  assign _EVAL_1350 = _EVAL_5163 | _EVAL_2718;
  assign _EVAL_2207 = _EVAL_1501 | _EVAL_1350;
  assign _EVAL_727 = _EVAL_153[1:0];
  assign _EVAL_2682 = _EVAL_727 != 2'h0;
  assign _EVAL_2283 = _EVAL_3226 & _EVAL_2682;
  assign _EVAL_941 = _EVAL_84[1:0];
  assign _EVAL_4901 = _EVAL_941 != 2'h0;
  assign _EVAL_4527 = _EVAL_1661 & _EVAL_4901;
  assign _EVAL_602 = _EVAL_98 ? _EVAL_2283 : _EVAL_4527;
  assign _EVAL_2160 = _EVAL_153[1];
  assign _EVAL_4451 = _EVAL_3226 & _EVAL_2160;
  assign _EVAL_1088 = _EVAL_154 == 5'h0;
  assign _EVAL_5289 = _EVAL_4451 & _EVAL_1088;
  assign _EVAL_2256 = _EVAL_84[1];
  assign _EVAL_4957 = _EVAL_1661 & _EVAL_2256;
  assign _EVAL_2519 = _EVAL_274 == 5'h0;
  assign _EVAL_2908 = _EVAL_4957 & _EVAL_2519;
  assign _EVAL_5016 = _EVAL_98 ? _EVAL_5289 : _EVAL_2908;
  assign _EVAL_3143 = _EVAL_5016 == 1'h0;
  assign _EVAL_889 = _EVAL_3143 & csr__EVAL_42;
  assign _EVAL_5172 = csr__EVAL_90 | _EVAL_889;
  assign _EVAL_2582 = _EVAL_602 & _EVAL_5172;
  assign _EVAL_4526 = _EVAL_2207 | _EVAL_2582;
  assign _EVAL_2777 = _EVAL_98 ? _EVAL_3226 : _EVAL_1661;
  assign _EVAL_2659 = _EVAL_602 == 1'h0;
  assign _EVAL_3093 = _EVAL_2777 & _EVAL_2659;
  assign _EVAL_3953 = _EVAL_3093 & csr__EVAL_85;
  assign _EVAL_3859 = _EVAL_4526 | _EVAL_3953;
  assign _EVAL_2084 = _EVAL_1348 | _EVAL_3859;
  assign _EVAL_1060 = _EVAL_55 & _EVAL_2084;
  assign _EVAL_4382 = _EVAL_601 == 1'h0;
  assign _EVAL_956 = _EVAL_1060 & _EVAL_4382;
  assign _EVAL_2221 = _EVAL_3608 & _EVAL_148;
  assign _EVAL_290 = _EVAL_4043 & _EVAL_1;
  assign _EVAL_1920 = _EVAL_2221 | _EVAL_290;
  assign _EVAL_1996 = _EVAL_154 == _EVAL_3117;
  assign _EVAL_2920 = _EVAL_1920 & _EVAL_1996;
  assign _EVAL_1442 = _EVAL_3608 & _EVAL_179;
  assign _EVAL_3651 = _EVAL_4043 & _EVAL_141;
  assign _EVAL_2129 = _EVAL_1442 | _EVAL_3651;
  assign _EVAL_4311 = _EVAL_68 == _EVAL_3117;
  assign _EVAL_1479 = _EVAL_2129 & _EVAL_4311;
  assign _EVAL_3277 = _EVAL_2920 | _EVAL_1479;
  assign _EVAL_1178 = _EVAL_3608 & _EVAL_119;
  assign _EVAL_3145 = _EVAL_4127 == _EVAL_3117;
  assign _EVAL_1126 = _EVAL_1178 & _EVAL_3145;
  assign _EVAL_1714 = _EVAL_3277 | _EVAL_1126;
  assign _EVAL_3195 = _EVAL_3608 & _EVAL_39;
  assign _EVAL_5062 = _EVAL_4043 & _EVAL_205;
  assign _EVAL_3155 = _EVAL_3195 | _EVAL_5062;
  assign _EVAL_3318 = _EVAL_274 == _EVAL_3117;
  assign _EVAL_3613 = _EVAL_3155 & _EVAL_3318;
  assign _EVAL_5281 = _EVAL_3608 & _EVAL_188;
  assign _EVAL_3455 = _EVAL_4043 & _EVAL_250;
  assign _EVAL_4897 = _EVAL_5281 | _EVAL_3455;
  assign _EVAL_4525 = _EVAL_180 == _EVAL_3117;
  assign _EVAL_3842 = _EVAL_4897 & _EVAL_4525;
  assign _EVAL_4938 = _EVAL_3613 | _EVAL_3842;
  assign _EVAL_2640 = _EVAL_3608 & _EVAL_260;
  assign _EVAL_3673 = _EVAL_3212 == _EVAL_3117;
  assign _EVAL_3506 = _EVAL_2640 & _EVAL_3673;
  assign _EVAL_3033 = _EVAL_4938 | _EVAL_3506;
  assign _EVAL_3524 = _EVAL_315 ? _EVAL_1714 : _EVAL_3033;
  assign _EVAL_5180 = _EVAL_2326 & _EVAL_3524;
  assign _EVAL_1349 = _EVAL_315 ? _EVAL_5180 : _EVAL_5180;
  assign _EVAL_5129 = fpu__EVAL_37;
  assign _EVAL_505 = _EVAL_3212 == _EVAL_5129;
  assign _EVAL_2902 = _EVAL_260 & _EVAL_505;
  assign _EVAL_3128 = _EVAL_116 == 1'h0;
  assign _EVAL_4513 = _EVAL_315 ? _EVAL_180 : _EVAL_68;
  assign _EVAL_5206 = {_EVAL_2400,_EVAL_4513};
  assign _EVAL_527 = $signed(_EVAL_5206);
  assign _EVAL_2066 = {_EVAL_983,_EVAL_1347,_EVAL_3134,_EVAL_4539};
  assign _EVAL_4358 = $signed(_EVAL_2066);
  assign _EVAL_5420 = $unsigned(_EVAL_4358);
  assign _EVAL_1665 = {_EVAL_5420, 12'h0};
  assign _EVAL_4838 = _EVAL_3840 ? _EVAL_1665 : 32'h0;
  assign _EVAL_1145 = {_EVAL_983,_EVAL_2579};
  assign _EVAL_2529 = $signed(_EVAL_1145);
  assign _EVAL_2770 = {_EVAL_983,_EVAL_1347};
  assign _EVAL_1296 = $signed(_EVAL_2770);
  assign _EVAL_1909 = _EVAL_2686 ? $signed(_EVAL_2529) : $signed(_EVAL_1296);
  assign _EVAL_3813 = $unsigned(_EVAL_1909);
  assign _EVAL_3737 = _EVAL_3813[11];
  assign _EVAL_3069 = _EVAL_3737 ? 20'hfffff : 20'h0;
  assign _EVAL_2417 = {_EVAL_3069,_EVAL_3813};
  assign _EVAL_643 = _EVAL_792 ? _EVAL_2417 : 32'h0;
  assign _EVAL_3298 = _EVAL_4838 | _EVAL_643;
  assign _EVAL_2061 = _EVAL_3481 ? _EVAL_949 : 32'h0;
  assign _EVAL_3932 = _EVAL_3298 | _EVAL_2061;
  assign _EVAL_4068 = _EVAL_3932[31:5];
  assign _EVAL_1560 = {_EVAL_4068,_EVAL_350};
  assign _EVAL_5102 = ~ _EVAL_1560;
  assign _EVAL_2799 = _EVAL_315 ? _EVAL_138 : _EVAL_2;
  assign _EVAL_2156 = _EVAL_2799[31:2];
  assign _EVAL_2627 = _EVAL_2156[6:0];
  assign _EVAL_4787 = _EVAL_3019 >> _EVAL_2627;
  assign _EVAL_2198 = _EVAL_4787[0];
  assign _EVAL_2422 = {_EVAL_2560,_EVAL_5401};
  assign _EVAL_3639 = _EVAL_2422 == 3'h4;
  assign _EVAL_774 = _EVAL_21[8:7];
  assign _EVAL_1021 = _EVAL_21[12:9];
  assign _EVAL_4455 = {_EVAL_774,_EVAL_1021,2'h0};
  assign _EVAL_4912 = _EVAL_4455[7:5];
  assign _EVAL_4730 = _EVAL_4455[4:0];
  assign _EVAL_412 = {_EVAL_4912,_EVAL_1302,5'h2,3'h2,_EVAL_4730,7'h27};
  assign _EVAL_1212 = {_EVAL_4912,_EVAL_1302,5'h2,3'h2,_EVAL_4730,7'h23};
  assign _EVAL_3396 = {_EVAL_3048,_EVAL_5115,3'h0};
  assign _EVAL_3051 = _EVAL_3396[8:5];
  assign _EVAL_1653 = _EVAL_3396[4:0];
  assign _EVAL_390 = {_EVAL_3051,_EVAL_1302,5'h2,3'h3,_EVAL_1653,7'h27};
  assign _EVAL_3733 = _EVAL_1302 != 5'h0;
  assign _EVAL_3778 = _EVAL_21[11:7];
  assign _EVAL_5223 = {_EVAL_1302,_EVAL_3778,3'h0,_EVAL_3778,7'h33};
  assign _EVAL_4327 = _EVAL_3778 != 5'h0;
  assign _EVAL_3991 = {_EVAL_1302,_EVAL_3778,3'h0,12'he7};
  assign _EVAL_3430 = {_EVAL_1302,_EVAL_3778,3'h0,12'h67};
  assign _EVAL_3368 = _EVAL_3430[24:7];
  assign _EVAL_911 = {_EVAL_3368,7'h73};
  assign _EVAL_2474 = _EVAL_911 | 25'h100000;
  assign _EVAL_5282 = _EVAL_4327 ? _EVAL_3991 : _EVAL_2474;
  assign _EVAL_2149 = _EVAL_3733 ? _EVAL_5223 : _EVAL_5282;
  assign _EVAL_3091 = {_EVAL_1302,5'h0,3'h4,_EVAL_3778,7'h33};
  assign _EVAL_4446 = _EVAL_3733 ? _EVAL_3091 : _EVAL_3430;
  assign _EVAL_3650 = _EVAL_2560 ? _EVAL_2149 : _EVAL_4446;
  assign _EVAL_1577 = _EVAL_21[3:2];
  assign _EVAL_784 = _EVAL_21[6:4];
  assign _EVAL_4082 = {_EVAL_1577,_EVAL_2560,_EVAL_784,2'h0,5'h2,3'h2,_EVAL_3778,7'h7};
  assign _EVAL_2190 = {_EVAL_1577,_EVAL_2560,_EVAL_784,2'h0,5'h2,3'h2,_EVAL_3778,7'h3};
  assign _EVAL_1383 = {_EVAL_4942,_EVAL_2560,_EVAL_5401,3'h0,5'h2,3'h3,_EVAL_3778,7'h7};
  assign _EVAL_1552 = {_EVAL_2560,_EVAL_1302,_EVAL_3778,3'h1,_EVAL_3778,7'h13};
  assign _EVAL_3653 = _EVAL_2854 ? _EVAL_1383 : {{3'd0}, _EVAL_1552};
  assign _EVAL_321 = _EVAL_5398 ? {{1'd0}, _EVAL_2190} : _EVAL_3653;
  assign _EVAL_3054 = _EVAL_1023 ? {{1'd0}, _EVAL_4082} : _EVAL_321;
  assign _EVAL_1081 = _EVAL_2350 ? {{4'd0}, _EVAL_3650} : _EVAL_3054;
  assign _EVAL_3669 = _EVAL_2034 ? _EVAL_390 : _EVAL_1081;
  assign _EVAL_294 = _EVAL_1631 ? {{1'd0}, _EVAL_1212} : _EVAL_3669;
  assign _EVAL_1711 = _EVAL_3243 ? {{1'd0}, _EVAL_412} : _EVAL_294;
  assign _EVAL_5114 = {3'h0,_EVAL_1711};
  assign _EVAL_2859 = _EVAL_4162[2];
  assign _EVAL_2723 = _EVAL_4162[0];
  assign _EVAL_3485 = _EVAL_2723 == 1'h0;
  assign _EVAL_1758 = _EVAL_2859 & _EVAL_3485;
  assign _EVAL_330 = _EVAL_5412[31:5];
  assign _EVAL_1141 = {_EVAL_330,_EVAL_1827};
  assign _EVAL_3092 = _EVAL_1141 ^ _EVAL_3901;
  assign _EVAL_3038 = _EVAL_1758 ? _EVAL_3092 : 32'h0;
  assign _EVAL_2578 = _EVAL_4162 >= 3'h6;
  assign _EVAL_4578 = _EVAL_1141 & _EVAL_3901;
  assign _EVAL_1142 = _EVAL_2578 ? _EVAL_4578 : 32'h0;
  assign _EVAL_665 = _EVAL_3038 | _EVAL_1142;
  assign _EVAL_4255 = _EVAL_4614[4:2];
  assign _EVAL_854 = _EVAL_4255 == 3'h7;
  assign _EVAL_4987 = _EVAL_3227 & _EVAL_854;
  assign _EVAL_3616 = _EVAL_4832[1:0];
  assign _EVAL_1712 = _EVAL_3616 == 2'h0;
  assign _EVAL_3105 = _EVAL_1588 & _EVAL_1712;
  assign _EVAL_615 = _EVAL_315 ? _EVAL_57 : _EVAL_20;
  assign _EVAL_4328 = _EVAL_615 == 1'h0;
  assign _EVAL_3989 = _EVAL_3105 & _EVAL_4328;
  assign _EVAL_2798 = _EVAL_315 ? _EVAL_236 : _EVAL_176;
  assign _EVAL_1836 = _EVAL_2758[31:16];
  assign _EVAL_3834 = {{16'd0}, _EVAL_1836};
  assign _EVAL_2931 = _EVAL_2758[15:0];
  assign _EVAL_759 = {_EVAL_2931, 16'h0};
  assign _EVAL_4492 = _EVAL_759 & 32'hffff0000;
  assign _EVAL_4066 = _EVAL_3834 | _EVAL_4492;
  assign _EVAL_2790 = _EVAL_4066[31:8];
  assign _EVAL_1117 = {{8'd0}, _EVAL_2790};
  assign _EVAL_1154 = _EVAL_1117 & 32'hff00ff;
  assign _EVAL_1449 = _EVAL_4066[23:0];
  assign _EVAL_367 = {_EVAL_1449, 8'h0};
  assign _EVAL_755 = _EVAL_367 & 32'hff00ff00;
  assign _EVAL_4682 = _EVAL_1154 | _EVAL_755;
  assign _EVAL_3439 = _EVAL_4682[31:4];
  assign _EVAL_5090 = {{4'd0}, _EVAL_3439};
  assign _EVAL_3908 = _EVAL_5090 & 32'hf0f0f0f;
  assign _EVAL_640 = _EVAL_4682[27:0];
  assign _EVAL_3357 = {_EVAL_640, 4'h0};
  assign _EVAL_1936 = _EVAL_3357 & 32'hf0f0f0f0;
  assign _EVAL_4873 = _EVAL_3908 | _EVAL_1936;
  assign _EVAL_340 = _EVAL_4596 == 1'h0;
  assign _EVAL_5318 = _EVAL_274 == _EVAL_3670;
  assign _EVAL_1741 = _EVAL_205 & _EVAL_5318;
  assign _EVAL_3046 = _EVAL_4633[4];
  assign _EVAL_968 = _EVAL_3046 == 1'h0;
  assign _EVAL_1065 = _EVAL_4633[3];
  assign _EVAL_2719 = _EVAL_968 & _EVAL_1065;
  assign _EVAL_4401 = _EVAL_4633[1];
  assign _EVAL_4119 = _EVAL_4401 == 1'h0;
  assign _EVAL_3743 = _EVAL_2719 & _EVAL_4119;
  assign _EVAL_3269 = _EVAL_545 & _EVAL_3743;
  assign _EVAL_5244 = _EVAL_2118 & _EVAL_3269;
  assign _EVAL_3299 = _EVAL_315 ? _EVAL_170 : _EVAL_242;
  assign _EVAL_3598 = _EVAL_315 ? _EVAL_191 : _EVAL_6;
  assign _EVAL_1768 = _EVAL_3598[4];
  assign _EVAL_4570 = _EVAL_1768 == 1'h0;
  assign _EVAL_2094 = _EVAL_3598[3];
  assign _EVAL_2152 = _EVAL_4570 & _EVAL_2094;
  assign _EVAL_4103 = _EVAL_3598[1];
  assign _EVAL_3119 = _EVAL_4103 == 1'h0;
  assign _EVAL_3322 = _EVAL_2152 & _EVAL_3119;
  assign _EVAL_2203 = _EVAL_3299 & _EVAL_3322;
  assign _EVAL_4630 = _EVAL_5244 & _EVAL_2203;
  assign _EVAL_2059 = _EVAL_315 ? _EVAL_154 : _EVAL_274;
  assign _EVAL_2953 = _EVAL_3134 == _EVAL_2059;
  assign _EVAL_4658 = _EVAL_4630 & _EVAL_2953;
  assign _EVAL_416 = _EVAL_315 ? _EVAL_121 : _EVAL_73;
  assign _EVAL_4859 = _EVAL_315 ? _EVAL_91 : _EVAL_171;
  assign _EVAL_4045 = {_EVAL_416,_EVAL_4859};
  assign _EVAL_3911 = $signed(_EVAL_4045);
  assign _EVAL_3010 = $signed(_EVAL_2529) == $signed(_EVAL_3911);
  assign _EVAL_3030 = _EVAL_4658 & _EVAL_3010;
  assign _EVAL_3703 = _EVAL_3747 & _EVAL_39;
  assign _EVAL_4312 = _EVAL_653 & _EVAL_205;
  assign _EVAL_2456 = _EVAL_3703 | _EVAL_4312;
  assign _EVAL_3377 = _EVAL_274 == _EVAL_2579;
  assign _EVAL_2390 = _EVAL_2456 & _EVAL_3377;
  assign _EVAL_4239 = _EVAL_3747 & _EVAL_188;
  assign _EVAL_3175 = _EVAL_653 & _EVAL_250;
  assign _EVAL_2217 = _EVAL_4239 | _EVAL_3175;
  assign _EVAL_1031 = _EVAL_180 == _EVAL_2579;
  assign _EVAL_4907 = _EVAL_2217 & _EVAL_1031;
  assign _EVAL_2259 = _EVAL_2390 | _EVAL_4907;
  assign _EVAL_5374 = _EVAL_3747 & _EVAL_260;
  assign _EVAL_2660 = _EVAL_3212 == _EVAL_2579;
  assign _EVAL_879 = _EVAL_5374 & _EVAL_2660;
  assign _EVAL_2817 = _EVAL_2259 | _EVAL_879;
  assign _EVAL_3060 = _EVAL_3747 & _EVAL_148;
  assign _EVAL_4708 = _EVAL_653 & _EVAL_1;
  assign _EVAL_600 = _EVAL_3060 | _EVAL_4708;
  assign _EVAL_4368 = _EVAL_154 == _EVAL_2579;
  assign _EVAL_440 = _EVAL_600 & _EVAL_4368;
  assign _EVAL_3180 = _EVAL_3747 & _EVAL_179;
  assign _EVAL_2685 = _EVAL_653 & _EVAL_141;
  assign _EVAL_5387 = _EVAL_3180 | _EVAL_2685;
  assign _EVAL_2119 = _EVAL_68 == _EVAL_2579;
  assign _EVAL_1985 = _EVAL_5387 & _EVAL_2119;
  assign _EVAL_1362 = _EVAL_440 | _EVAL_1985;
  assign _EVAL_4486 = _EVAL_3747 & _EVAL_119;
  assign _EVAL_2995 = _EVAL_4127 == _EVAL_2579;
  assign _EVAL_3412 = _EVAL_4486 & _EVAL_2995;
  assign _EVAL_5071 = _EVAL_1362 | _EVAL_3412;
  assign _EVAL_3787 = _EVAL_315 ? _EVAL_2817 : _EVAL_5071;
  assign _EVAL_3942 = _EVAL_2118 & _EVAL_3787;
  assign _EVAL_449 = _EVAL_315 ? _EVAL_3942 : _EVAL_3942;
  assign _EVAL_2875 = _EVAL_449 & _EVAL_3747;
  assign _EVAL_4036 = _EVAL_58 | _EVAL_148;
  assign _EVAL_3111 = _EVAL_4036 | _EVAL_179;
  assign _EVAL_1995 = _EVAL_2923 == 1'h0;
  assign _EVAL_2808 = _EVAL_4705 & _EVAL_1995;
  assign _EVAL_316 = _EVAL_2808 & _EVAL_3618;
  assign _EVAL_4480 = _EVAL_1446 & _EVAL_316;
  assign _EVAL_1275 = _EVAL_4299 & _EVAL_188;
  assign _EVAL_4617 = _EVAL_4692 & _EVAL_250;
  assign _EVAL_5187 = _EVAL_1275 | _EVAL_4617;
  assign _EVAL_1408 = _EVAL_2422 == 3'h3;
  assign _EVAL_5031 = _EVAL_2268 == 1'h0;
  assign _EVAL_1264 = _EVAL_2506 & _EVAL_5031;
  assign _EVAL_3971 = _EVAL_2506 & _EVAL_1446;
  assign _EVAL_2803 = _EVAL_3971 & _EVAL_196;
  assign _EVAL_4662 = _EVAL_3421 | _EVAL_2803;
  assign _EVAL_444 = _EVAL_3971 & _EVAL_122;
  assign _EVAL_4613 = _EVAL_4662 | _EVAL_444;
  assign _EVAL_525 = _EVAL_3971 & _EVAL_175;
  assign _EVAL_2364 = _EVAL_4613 | _EVAL_525;
  assign _EVAL_1127 = _EVAL_3971 & _EVAL_146;
  assign _EVAL_5295 = _EVAL_2364 | _EVAL_1127;
  assign _EVAL_2806 = _EVAL_3971 & _EVAL_249;
  assign _EVAL_4244 = _EVAL_5295 | _EVAL_2806;
  assign _EVAL_1924 = _EVAL_3971 & _EVAL_255;
  assign _EVAL_5104 = _EVAL_4244 | _EVAL_1924;
  assign _EVAL_3565 = _EVAL_1264 & _EVAL_5104;
  assign _EVAL_3340 = _EVAL_2758[31];
  assign _EVAL_4854 = _EVAL_5185 | _EVAL_3340;
  assign _EVAL_3161 = {_EVAL_4854,_EVAL_2758};
  assign _EVAL_3151 = $signed(_EVAL_3161);
  assign _EVAL_4098 = _EVAL_4373[31];
  assign _EVAL_2992 = _EVAL_5185 | _EVAL_4098;
  assign _EVAL_4713 = {_EVAL_2992,_EVAL_4373};
  assign _EVAL_4565 = $signed(_EVAL_4713);
  assign _EVAL_1225 = $signed(_EVAL_3151) < $signed(_EVAL_4565);
  assign _EVAL_3208 = _EVAL_3227 & _EVAL_5052;
  assign _EVAL_1171 = _EVAL_2644 == 1'h0;
  assign _EVAL_3316 = _EVAL_3208 & _EVAL_1171;
  assign _EVAL_2201 = _EVAL_3316 ? _EVAL_1024 : 3'h2;
  assign _EVAL_3188 = _EVAL_3208 & _EVAL_1250;
  assign _EVAL_448 = _EVAL_3188 & _EVAL_1171;
  assign _EVAL_2865 = {{2'd0}, _EVAL_448};
  assign _EVAL_3282 = _EVAL_2201 ^ _EVAL_2865;
  assign _EVAL_1812 = _EVAL_3282[0];
  assign _EVAL_2666 = _EVAL_3282[2];
  assign _EVAL_4646 = _EVAL_1812 ^ _EVAL_2666;
  assign _EVAL_1973 = _EVAL_2758 == _EVAL_4373;
  assign _EVAL_4392 = _EVAL_2666 == 1'h0;
  assign _EVAL_2588 = _EVAL_3282[1];
  assign _EVAL_2937 = _EVAL_2588 == 1'h0;
  assign _EVAL_689 = _EVAL_4392 & _EVAL_2937;
  assign _EVAL_5023 = _EVAL_1812 ^ _EVAL_689;
  assign _EVAL_2731 = _EVAL_1973 ? _EVAL_5023 : _EVAL_1812;
  assign _EVAL_4982 = _EVAL_1225 ? _EVAL_4646 : _EVAL_2731;
  assign _EVAL_4583 = _EVAL_4982 == 1'h0;
  assign _EVAL_3672 = _EVAL_3565 & _EVAL_4583;
  assign _EVAL_4637 = _EVAL_3672 | csr__EVAL_89;
  assign _EVAL_4643 = _EVAL_1333 | _EVAL_4962;
  assign _EVAL_1780 = _EVAL_3971 & _EVAL_4643;
  assign _EVAL_2498 = _EVAL_163 == 1'h0;
  assign _EVAL_2810 = _EVAL_1780 & _EVAL_2498;
  assign _EVAL_593 = _EVAL_3404 == 1'h0;
  assign _EVAL_1523 = _EVAL_2810 & _EVAL_593;
  assign _EVAL_2121 = _EVAL_4637 | _EVAL_1523;
  assign _EVAL_4971 = _EVAL_5043[2:0];
  assign _EVAL_1764 = _EVAL_4614[1:0];
  assign _EVAL_750 = _EVAL_1764 == 2'h0;
  assign _EVAL_5329 = _EVAL_1699 & _EVAL_750;
  assign _EVAL_799 = _EVAL_3227 & _EVAL_5329;
  assign _EVAL_4091 = _EVAL_799 ? _EVAL_1024 : 3'h2;
  assign _EVAL_1885 = _EVAL_3227 & _EVAL_1699;
  assign _EVAL_1805 = _EVAL_750 == 1'h0;
  assign _EVAL_4786 = _EVAL_1885 & _EVAL_1805;
  assign _EVAL_1274 = {{2'd0}, _EVAL_4786};
  assign _EVAL_2679 = _EVAL_4091 ^ _EVAL_1274;
  assign _EVAL_5127 = _EVAL_2679[2];
  assign _EVAL_1568 = _EVAL_5127 == 1'h0;
  assign _EVAL_1775 = _EVAL_68 != _EVAL_68;
  assign _EVAL_4350 = _EVAL_3039[4];
  assign _EVAL_3359 = _EVAL_4350 == 1'h0;
  assign _EVAL_4183 = _EVAL_3039[2];
  assign _EVAL_2965 = _EVAL_3359 & _EVAL_4183;
  assign _EVAL_4536 = _EVAL_5114[24:20];
  assign _EVAL_754 = _EVAL_4562 ? 3'h4 : 3'h6;
  assign _EVAL_1517 = _EVAL_4562 ? 4'h6 : 4'h8;
  assign _EVAL_3406 = _EVAL_5233 ? {{1'd0}, _EVAL_754} : _EVAL_1517;
  assign _EVAL_945 = _EVAL_4562 ? 3'h2 : 3'h4;
  assign _EVAL_3515 = _EVAL_4423 ? _EVAL_3406 : {{1'd0}, _EVAL_945};
  assign _EVAL_5091 = {{28'd0}, _EVAL_3515};
  assign _EVAL_4238 = _EVAL_4157 + _EVAL_5091;
  assign _EVAL_920 = _EVAL_16 & _EVAL_4962;
  assign _EVAL_790 = _EVAL_214 & _EVAL_1333;
  assign _EVAL_3702 = _EVAL_920 | _EVAL_790;
  assign _EVAL_4284 = _EVAL_4362 & _EVAL_148;
  assign _EVAL_4471 = _EVAL_332 & _EVAL_1;
  assign _EVAL_5245 = _EVAL_4284 | _EVAL_4471;
  assign _EVAL_4048 = _EVAL_154 == _EVAL_5099;
  assign _EVAL_2766 = _EVAL_5245 & _EVAL_4048;
  assign _EVAL_4429 = _EVAL_4362 & _EVAL_179;
  assign _EVAL_2848 = _EVAL_332 & _EVAL_141;
  assign _EVAL_3250 = _EVAL_4429 | _EVAL_2848;
  assign _EVAL_3780 = _EVAL_68 == _EVAL_5099;
  assign _EVAL_1263 = _EVAL_3250 & _EVAL_3780;
  assign _EVAL_1358 = _EVAL_2766 | _EVAL_1263;
  assign _EVAL_4862 = _EVAL_4362 & _EVAL_119;
  assign _EVAL_2406 = _EVAL_4127 == _EVAL_5099;
  assign _EVAL_2213 = _EVAL_4862 & _EVAL_2406;
  assign _EVAL_5046 = _EVAL_1358 | _EVAL_2213;
  assign _EVAL_1396 = _EVAL_1065 == 1'h0;
  assign _EVAL_822 = _EVAL_968 & _EVAL_1396;
  assign _EVAL_1018 = _EVAL_822 & _EVAL_4119;
  assign _EVAL_1041 = _EVAL_545 & _EVAL_1018;
  assign _EVAL_671 = _EVAL_2719 & _EVAL_4401;
  assign _EVAL_1910 = _EVAL_545 & _EVAL_671;
  assign _EVAL_4974 = _EVAL_1041 | _EVAL_1910;
  assign _EVAL_1659 = _EVAL_2118 & _EVAL_4974;
  assign _EVAL_2357 = _EVAL_259 == 1'h0;
  assign _EVAL_1997 = _EVAL_1659 & _EVAL_2357;
  assign _EVAL_3223 = _EVAL_21[1:0];
  assign _EVAL_2164 = _EVAL_3223 == 2'h2;
  assign _EVAL_3943 = _EVAL_5114[11:7];
  assign _EVAL_1926 = _EVAL_3223 == 2'h1;
  assign _EVAL_3462 = _EVAL_2560 ? 5'h1f : 5'h0;
  assign _EVAL_5193 = _EVAL_21[2];
  assign _EVAL_2440 = _EVAL_21[11:10];
  assign _EVAL_2606 = _EVAL_21[4:3];
  assign _EVAL_558 = {_EVAL_3462,_EVAL_5401,_EVAL_5193,_EVAL_2440,_EVAL_2606,1'h0};
  assign _EVAL_4972 = _EVAL_558[12];
  assign _EVAL_4648 = _EVAL_558[10:5];
  assign _EVAL_1245 = _EVAL_558[4:1];
  assign _EVAL_3529 = _EVAL_558[11];
  assign _EVAL_4273 = {_EVAL_4972,_EVAL_4648,5'h0,2'h1,_EVAL_3048,3'h1,_EVAL_1245,_EVAL_3529,7'h63};
  assign _EVAL_2764 = {_EVAL_4972,_EVAL_4648,5'h0,2'h1,_EVAL_3048,3'h0,_EVAL_1245,_EVAL_3529,7'h63};
  assign _EVAL_3008 = _EVAL_2560 ? 10'h3ff : 10'h0;
  assign _EVAL_632 = _EVAL_21[8];
  assign _EVAL_1128 = _EVAL_21[10:9];
  assign _EVAL_3300 = _EVAL_21[7];
  assign _EVAL_662 = _EVAL_21[11];
  assign _EVAL_2052 = _EVAL_21[5:3];
  assign _EVAL_793 = {_EVAL_3008,_EVAL_632,_EVAL_1128,_EVAL_2565,_EVAL_3300,_EVAL_5193,_EVAL_662,_EVAL_2052,1'h0};
  assign _EVAL_2026 = _EVAL_793[20];
  assign _EVAL_1951 = _EVAL_793[10:1];
  assign _EVAL_1040 = _EVAL_793[11];
  assign _EVAL_1075 = _EVAL_793[19:12];
  assign _EVAL_5298 = {_EVAL_2026,_EVAL_1951,_EVAL_1040,_EVAL_1075,5'h0,7'h6f};
  assign _EVAL_5242 = _EVAL_2440 == 2'h3;
  assign _EVAL_4995 = _EVAL_2422 == 3'h7;
  assign _EVAL_3177 = _EVAL_2422 == 3'h6;
  assign _EVAL_3874 = _EVAL_2422 == 3'h5;
  assign _EVAL_2265 = _EVAL_2422 == 3'h2;
  assign _EVAL_3296 = _EVAL_2422 == 3'h1;
  assign _EVAL_1769 = _EVAL_3296 ? 3'h4 : 3'h0;
  assign _EVAL_2058 = _EVAL_2265 ? 3'h6 : _EVAL_1769;
  assign _EVAL_984 = _EVAL_1408 ? 3'h7 : _EVAL_2058;
  assign _EVAL_1856 = _EVAL_3639 ? 3'h0 : _EVAL_984;
  assign _EVAL_1240 = _EVAL_3874 ? 3'h0 : _EVAL_1856;
  assign _EVAL_1429 = _EVAL_3177 ? 3'h2 : _EVAL_1240;
  assign _EVAL_3072 = _EVAL_4995 ? 3'h3 : _EVAL_1429;
  assign _EVAL_1374 = _EVAL_2560 ? 7'h3b : 7'h33;
  assign _EVAL_310 = {2'h1,_EVAL_4942,2'h1,_EVAL_3048,_EVAL_3072,2'h1,_EVAL_3048,_EVAL_1374};
  assign _EVAL_2038 = {{6'd0}, _EVAL_310};
  assign _EVAL_1644 = _EVAL_5401 == 2'h0;
  assign _EVAL_5151 = {_EVAL_1644, 30'h0};
  assign _EVAL_2646 = _EVAL_2038 | _EVAL_5151;
  assign _EVAL_1710 = _EVAL_2440 == 2'h2;
  assign _EVAL_2858 = _EVAL_2560 ? 7'h7f : 7'h0;
  assign _EVAL_2707 = {_EVAL_2858,_EVAL_1302,2'h1,_EVAL_3048,3'h7,2'h1,_EVAL_3048,7'h13};
  assign _EVAL_2601 = _EVAL_2440 == 2'h1;
  assign _EVAL_974 = {_EVAL_2560,_EVAL_1302,2'h1,_EVAL_3048,3'h5,2'h1,_EVAL_3048,7'h13};
  assign _EVAL_501 = {{5'd0}, _EVAL_974};
  assign _EVAL_1376 = _EVAL_501 | 31'h40000000;
  assign _EVAL_1357 = _EVAL_2601 ? _EVAL_1376 : {{5'd0}, _EVAL_974};
  assign _EVAL_1016 = _EVAL_1710 ? _EVAL_2707 : {{1'd0}, _EVAL_1357};
  assign _EVAL_1001 = _EVAL_5242 ? {{1'd0}, _EVAL_2646} : _EVAL_1016;
  assign _EVAL_3716 = _EVAL_3778 == 5'h2;
  assign _EVAL_5339 = _EVAL_2560 ? 3'h7 : 3'h0;
  assign _EVAL_3810 = {_EVAL_5339,_EVAL_2606,_EVAL_1323,_EVAL_5193,_EVAL_2565,4'h0,_EVAL_3778,3'h0,_EVAL_3778,7'h13};
  assign _EVAL_548 = _EVAL_4377[31:12];
  assign _EVAL_1116 = {_EVAL_548,_EVAL_3778,7'h37};
  assign _EVAL_5407 = _EVAL_3716 ? _EVAL_3810 : _EVAL_1116;
  assign _EVAL_2255 = {_EVAL_2858,_EVAL_1302,5'h0,3'h0,_EVAL_3778,7'h13};
  assign _EVAL_1283 = {_EVAL_2026,_EVAL_1951,_EVAL_1040,_EVAL_1075,5'h1,7'h6f};
  assign _EVAL_2730 = {_EVAL_2858,_EVAL_1302,_EVAL_3778,3'h0,_EVAL_3778,7'h13};
  assign _EVAL_4432 = _EVAL_2854 ? _EVAL_1283 : _EVAL_2730;
  assign _EVAL_2427 = _EVAL_5398 ? _EVAL_2255 : _EVAL_4432;
  assign _EVAL_2822 = _EVAL_1023 ? _EVAL_5407 : _EVAL_2427;
  assign _EVAL_3715 = _EVAL_2350 ? _EVAL_1001 : _EVAL_2822;
  assign _EVAL_2437 = _EVAL_2034 ? _EVAL_5298 : _EVAL_3715;
  assign _EVAL_2378 = _EVAL_1631 ? _EVAL_2764 : _EVAL_2437;
  assign _EVAL_2302 = _EVAL_3243 ? _EVAL_4273 : _EVAL_2378;
  assign _EVAL_504 = _EVAL_2302[11:7];
  assign _EVAL_5382 = _EVAL_4329[11:7];
  assign _EVAL_1990 = _EVAL_1926 ? _EVAL_504 : _EVAL_5382;
  assign _EVAL_1847 = _EVAL_2164 ? _EVAL_3943 : _EVAL_1990;
  assign _EVAL_3399 = csr__EVAL_160;
  assign _EVAL_630 = _EVAL_1333 & _EVAL_205;
  assign _EVAL_4518 = _EVAL_4614[4];
  assign _EVAL_508 = _EVAL_4518 == 1'h0;
  assign _EVAL_3504 = _EVAL_4614[2];
  assign _EVAL_2915 = _EVAL_508 & _EVAL_3504;
  assign _EVAL_1707 = _EVAL_4614[3];
  assign _EVAL_4313 = _EVAL_2915 & _EVAL_1707;
  assign _EVAL_4992 = _EVAL_4614[0];
  assign _EVAL_1355 = _EVAL_4992 == 1'h0;
  assign _EVAL_3438 = _EVAL_4313 & _EVAL_1355;
  assign _EVAL_3246 = _EVAL_3229[0];
  assign _EVAL_3568 = _EVAL_3438 & _EVAL_3246;
  assign _EVAL_3467 = _EVAL_3360 == 1'h0;
  assign _EVAL_4150 = _EVAL_3568 & _EVAL_3467;
  assign _EVAL_3894 = _EVAL_2912[30:23];
  assign _EVAL_2899 = _EVAL_3894 == 8'h0;
  assign _EVAL_1182 = _EVAL_2912[22:0];
  assign _EVAL_299 = _EVAL_1182 == 23'h0;
  assign _EVAL_590 = _EVAL_2899 & _EVAL_299;
  assign _EVAL_1450 = _EVAL_590 == 1'h0;
  assign _EVAL_5334 = {{31'd0}, _EVAL_1182};
  assign _EVAL_1870 = _EVAL_1182[15:0];
  assign _EVAL_2006 = _EVAL_1870[15:8];
  assign _EVAL_5309 = {{8'd0}, _EVAL_2006};
  assign _EVAL_3960 = _EVAL_1870[7:0];
  assign _EVAL_1917 = {_EVAL_3960, 8'h0};
  assign _EVAL_4935 = _EVAL_1917 & 16'hff00;
  assign _EVAL_3495 = _EVAL_5309 | _EVAL_4935;
  assign _EVAL_1810 = _EVAL_3495[15:4];
  assign _EVAL_2670 = {{4'd0}, _EVAL_1810};
  assign _EVAL_4496 = _EVAL_2670 & 16'hf0f;
  assign _EVAL_5267 = _EVAL_3495[11:0];
  assign _EVAL_3056 = {_EVAL_5267, 4'h0};
  assign _EVAL_1160 = _EVAL_3056 & 16'hf0f0;
  assign _EVAL_2628 = _EVAL_4496 | _EVAL_1160;
  assign _EVAL_2815 = _EVAL_2628[15:2];
  assign _EVAL_2459 = {{2'd0}, _EVAL_2815};
  assign _EVAL_2819 = _EVAL_2459 & 16'h3333;
  assign _EVAL_1642 = _EVAL_2628[13:0];
  assign _EVAL_4121 = {_EVAL_1642, 2'h0};
  assign _EVAL_1224 = _EVAL_4121 & 16'hcccc;
  assign _EVAL_2739 = _EVAL_2819 | _EVAL_1224;
  assign _EVAL_1017 = _EVAL_2739[15:1];
  assign _EVAL_2642 = {{1'd0}, _EVAL_1017};
  assign _EVAL_3741 = _EVAL_2642 & 16'h5555;
  assign _EVAL_827 = _EVAL_2739[14:0];
  assign _EVAL_2761 = {_EVAL_827, 1'h0};
  assign _EVAL_3480 = _EVAL_2761 & 16'haaaa;
  assign _EVAL_2712 = _EVAL_3741 | _EVAL_3480;
  assign _EVAL_3004 = _EVAL_1182[22:16];
  assign _EVAL_320 = _EVAL_3004[3:0];
  assign _EVAL_1488 = _EVAL_320[1:0];
  assign _EVAL_807 = _EVAL_1488[0];
  assign _EVAL_3545 = _EVAL_1488[1];
  assign _EVAL_4537 = _EVAL_320[3:2];
  assign _EVAL_4910 = _EVAL_4537[0];
  assign _EVAL_2373 = _EVAL_4537[1];
  assign _EVAL_3065 = _EVAL_3004[6:4];
  assign _EVAL_3883 = _EVAL_3065[1:0];
  assign _EVAL_2662 = _EVAL_3883[0];
  assign _EVAL_5200 = _EVAL_3883[1];
  assign _EVAL_5210 = _EVAL_3065[2];
  assign _EVAL_463 = {_EVAL_2712,_EVAL_807,_EVAL_3545,_EVAL_4910,_EVAL_2373,_EVAL_2662,_EVAL_5200,_EVAL_5210};
  assign _EVAL_1377 = _EVAL_463[0];
  assign _EVAL_1668 = _EVAL_463[1];
  assign _EVAL_840 = _EVAL_463[2];
  assign _EVAL_2918 = _EVAL_463[3];
  assign _EVAL_5176 = _EVAL_463[4];
  assign _EVAL_1382 = _EVAL_463[5];
  assign _EVAL_4084 = _EVAL_463[6];
  assign _EVAL_2540 = _EVAL_463[7];
  assign _EVAL_4407 = _EVAL_463[8];
  assign _EVAL_1054 = _EVAL_463[9];
  assign _EVAL_1003 = _EVAL_463[10];
  assign _EVAL_2202 = _EVAL_463[11];
  assign _EVAL_2374 = _EVAL_463[12];
  assign _EVAL_2759 = _EVAL_463[13];
  assign _EVAL_3786 = _EVAL_463[14];
  assign _EVAL_3118 = _EVAL_463[15];
  assign _EVAL_4948 = _EVAL_463[16];
  assign _EVAL_1375 = _EVAL_463[17];
  assign _EVAL_2484 = _EVAL_463[18];
  assign _EVAL_4895 = _EVAL_463[19];
  assign _EVAL_3040 = _EVAL_463[20];
  assign _EVAL_4749 = _EVAL_463[21];
  assign _EVAL_1831 = _EVAL_4749 ? 5'h15 : 5'h16;
  assign _EVAL_2562 = _EVAL_3040 ? 5'h14 : _EVAL_1831;
  assign _EVAL_933 = _EVAL_4895 ? 5'h13 : _EVAL_2562;
  assign _EVAL_4164 = _EVAL_2484 ? 5'h12 : _EVAL_933;
  assign _EVAL_3063 = _EVAL_1375 ? 5'h11 : _EVAL_4164;
  assign _EVAL_3617 = _EVAL_4948 ? 5'h10 : _EVAL_3063;
  assign _EVAL_741 = _EVAL_3118 ? 5'hf : _EVAL_3617;
  assign _EVAL_3484 = _EVAL_3786 ? 5'he : _EVAL_741;
  assign _EVAL_2674 = _EVAL_2759 ? 5'hd : _EVAL_3484;
  assign _EVAL_2314 = _EVAL_2374 ? 5'hc : _EVAL_2674;
  assign _EVAL_3941 = _EVAL_2202 ? 5'hb : _EVAL_2314;
  assign _EVAL_2633 = _EVAL_1003 ? 5'ha : _EVAL_3941;
  assign _EVAL_4321 = _EVAL_1054 ? 5'h9 : _EVAL_2633;
  assign _EVAL_3871 = _EVAL_4407 ? 5'h8 : _EVAL_4321;
  assign _EVAL_3993 = _EVAL_2540 ? 5'h7 : _EVAL_3871;
  assign _EVAL_2183 = _EVAL_4084 ? 5'h6 : _EVAL_3993;
  assign _EVAL_751 = _EVAL_1382 ? 5'h5 : _EVAL_2183;
  assign _EVAL_2085 = _EVAL_5176 ? 5'h4 : _EVAL_751;
  assign _EVAL_305 = _EVAL_2918 ? 5'h3 : _EVAL_2085;
  assign _EVAL_1514 = _EVAL_840 ? 5'h2 : _EVAL_305;
  assign _EVAL_2284 = _EVAL_1668 ? 5'h1 : _EVAL_1514;
  assign _EVAL_596 = _EVAL_1377 ? 5'h0 : _EVAL_2284;
  assign _EVAL_4625 = _EVAL_5334 << _EVAL_596;
  assign _EVAL_5257 = _EVAL_4625[21:0];
  assign _EVAL_695 = {_EVAL_5257, 1'h0};
  assign _EVAL_1386 = _EVAL_2899 ? _EVAL_695 : _EVAL_1182;
  assign _EVAL_2353 = {1'h0,_EVAL_1450,_EVAL_1386};
  assign _EVAL_4309 = _EVAL_3405 == 32'hc;
  assign _EVAL_5252 = _EVAL_2257 ? 1'h1 : _EVAL_612;
  assign _EVAL_5386 = _EVAL_2257 ? 1'h1 : _EVAL_4844;
  assign _EVAL_2812 = _EVAL_2257 ? divider__EVAL_11 : _EVAL_4939;
  assign _EVAL_743 = _EVAL_2812 == _EVAL_154;
  assign _EVAL_4839 = _EVAL_5386 & _EVAL_743;
  assign _EVAL_3364 = _EVAL_5252 & _EVAL_4839;
  assign _EVAL_554 = _EVAL_2812 == _EVAL_274;
  assign _EVAL_3460 = _EVAL_5386 & _EVAL_554;
  assign _EVAL_1228 = _EVAL_5252 & _EVAL_3460;
  assign _EVAL_969 = _EVAL_315 ? _EVAL_3364 : _EVAL_1228;
  assign _EVAL_4177 = _EVAL_5114 & 32'h50;
  assign _EVAL_3271 = _EVAL_4177 == 32'h10;
  assign _EVAL_2339 = csr__EVAL_15;
  assign _EVAL_523 = csr__EVAL_131;
  assign _EVAL_4191 = {_EVAL_2339,1'h0,1'h0,_EVAL_523};
  assign _EVAL_5168 = csr__EVAL_76;
  assign _EVAL_761 = _EVAL_4191 >> _EVAL_5168;
  assign _EVAL_451 = _EVAL_761[0];
  assign _EVAL_4892 = _EVAL_269[15:13];
  assign _EVAL_3284 = _EVAL_4892 == 3'h7;
  assign _EVAL_2831 = _EVAL_269[8:7];
  assign _EVAL_1033 = _EVAL_269[12:9];
  assign _EVAL_3985 = {_EVAL_2831,_EVAL_1033,2'h0};
  assign _EVAL_2344 = _EVAL_3985[7:5];
  assign _EVAL_5394 = _EVAL_269[6:2];
  assign _EVAL_5162 = _EVAL_3985[4:0];
  assign _EVAL_4249 = {_EVAL_2344,_EVAL_5394,5'h2,3'h2,_EVAL_5162,7'h27};
  assign _EVAL_4909 = _EVAL_4892 == 3'h6;
  assign _EVAL_1983 = {_EVAL_2344,_EVAL_5394,5'h2,3'h2,_EVAL_5162,7'h23};
  assign _EVAL_397 = _EVAL_4892 == 3'h5;
  assign _EVAL_2725 = _EVAL_269[9:7];
  assign _EVAL_5220 = _EVAL_269[12:10];
  assign _EVAL_492 = {_EVAL_2725,_EVAL_5220,3'h0};
  assign _EVAL_4123 = _EVAL_492[8:5];
  assign _EVAL_550 = _EVAL_492[4:0];
  assign _EVAL_1675 = {_EVAL_4123,_EVAL_5394,5'h2,3'h3,_EVAL_550,7'h27};
  assign _EVAL_4280 = _EVAL_4892 == 3'h4;
  assign _EVAL_2487 = _EVAL_5394 != 5'h0;
  assign _EVAL_475 = _EVAL_269[11:7];
  assign _EVAL_3144 = {_EVAL_5394,_EVAL_475,3'h0,_EVAL_475,7'h33};
  assign _EVAL_1428 = _EVAL_475 != 5'h0;
  assign _EVAL_4138 = {_EVAL_5394,_EVAL_475,3'h0,12'he7};
  assign _EVAL_4477 = {_EVAL_5394,_EVAL_475,3'h0,12'h67};
  assign _EVAL_2319 = _EVAL_4477[24:7];
  assign _EVAL_1777 = {_EVAL_2319,7'h73};
  assign _EVAL_4493 = _EVAL_1777 | 25'h100000;
  assign _EVAL_5122 = _EVAL_1428 ? _EVAL_4138 : _EVAL_4493;
  assign _EVAL_5238 = _EVAL_2487 ? _EVAL_3144 : _EVAL_5122;
  assign _EVAL_4934 = {_EVAL_5394,5'h0,3'h4,_EVAL_475,7'h33};
  assign _EVAL_4592 = _EVAL_2487 ? _EVAL_4934 : _EVAL_4477;
  assign _EVAL_4248 = _EVAL_1241 ? _EVAL_5238 : _EVAL_4592;
  assign _EVAL_5161 = _EVAL_4892 == 3'h3;
  assign _EVAL_3619 = _EVAL_269[3:2];
  assign _EVAL_978 = _EVAL_269[6:4];
  assign _EVAL_3777 = {_EVAL_3619,_EVAL_1241,_EVAL_978,2'h0,5'h2,3'h2,_EVAL_475,7'h7};
  assign _EVAL_654 = _EVAL_4892 == 3'h2;
  assign _EVAL_2525 = {_EVAL_3619,_EVAL_1241,_EVAL_978,2'h0,5'h2,3'h2,_EVAL_475,7'h3};
  assign _EVAL_1897 = _EVAL_4892 == 3'h1;
  assign _EVAL_3643 = _EVAL_269[4:2];
  assign _EVAL_3935 = _EVAL_269[6:5];
  assign _EVAL_3738 = {_EVAL_3643,_EVAL_1241,_EVAL_3935,3'h0,5'h2,3'h3,_EVAL_475,7'h7};
  assign _EVAL_3327 = {_EVAL_1241,_EVAL_5394,_EVAL_475,3'h1,_EVAL_475,7'h13};
  assign _EVAL_587 = _EVAL_1897 ? _EVAL_3738 : {{3'd0}, _EVAL_3327};
  assign _EVAL_746 = _EVAL_654 ? {{1'd0}, _EVAL_2525} : _EVAL_587;
  assign _EVAL_982 = _EVAL_5161 ? {{1'd0}, _EVAL_3777} : _EVAL_746;
  assign _EVAL_1756 = _EVAL_4280 ? {{4'd0}, _EVAL_4248} : _EVAL_982;
  assign _EVAL_5191 = _EVAL_397 ? _EVAL_1675 : _EVAL_1756;
  assign _EVAL_3878 = _EVAL_4909 ? {{1'd0}, _EVAL_1983} : _EVAL_5191;
  assign _EVAL_4470 = _EVAL_3284 ? {{1'd0}, _EVAL_4249} : _EVAL_3878;
  assign _EVAL_2522 = {3'h0,_EVAL_4470};
  assign _EVAL_2637 = _EVAL_2522[11:7];
  assign _EVAL_4894 = _EVAL_2637 != 5'h0;
  assign _EVAL_2538 = _EVAL_313[2];
  assign _EVAL_419 = _EVAL_4468[31];
  assign _EVAL_2857 = _EVAL_5237 & _EVAL_419;
  assign _EVAL_1432 = {_EVAL_2857,_EVAL_4468};
  assign _EVAL_1753 = _EVAL_4468[31:16];
  assign _EVAL_4999 = {{16'd0}, _EVAL_1753};
  assign _EVAL_962 = _EVAL_4468[15:0];
  assign _EVAL_5156 = {_EVAL_962, 16'h0};
  assign _EVAL_2124 = _EVAL_5156 & 32'hffff0000;
  assign _EVAL_1578 = _EVAL_4999 | _EVAL_2124;
  assign _EVAL_4320 = _EVAL_1578[31:8];
  assign _EVAL_482 = {{8'd0}, _EVAL_4320};
  assign _EVAL_2439 = _EVAL_482 & 32'hff00ff;
  assign _EVAL_2116 = _EVAL_1578[23:0];
  assign _EVAL_3550 = {_EVAL_2116, 8'h0};
  assign _EVAL_967 = _EVAL_3550 & 32'hff00ff00;
  assign _EVAL_3172 = _EVAL_2439 | _EVAL_967;
  assign _EVAL_343 = _EVAL_3172[31:4];
  assign _EVAL_1581 = {{4'd0}, _EVAL_343};
  assign _EVAL_4061 = _EVAL_1581 & 32'hf0f0f0f;
  assign _EVAL_970 = _EVAL_3172[27:0];
  assign _EVAL_2946 = {_EVAL_970, 4'h0};
  assign _EVAL_5110 = _EVAL_2946 & 32'hf0f0f0f0;
  assign _EVAL_2665 = _EVAL_4061 | _EVAL_5110;
  assign _EVAL_291 = _EVAL_2665[31:2];
  assign _EVAL_2724 = {{2'd0}, _EVAL_291};
  assign _EVAL_852 = _EVAL_2724 & 32'h33333333;
  assign _EVAL_4850 = _EVAL_2665[29:0];
  assign _EVAL_887 = {_EVAL_4850, 2'h0};
  assign _EVAL_5007 = _EVAL_887 & 32'hcccccccc;
  assign _EVAL_468 = _EVAL_852 | _EVAL_5007;
  assign _EVAL_4383 = _EVAL_468[31:1];
  assign _EVAL_620 = {{1'd0}, _EVAL_4383};
  assign _EVAL_1599 = _EVAL_620 & 32'h55555555;
  assign _EVAL_4403 = _EVAL_468[30:0];
  assign _EVAL_2032 = {_EVAL_4403, 1'h0};
  assign _EVAL_4604 = _EVAL_2032 & 32'haaaaaaaa;
  assign _EVAL_2571 = _EVAL_1599 | _EVAL_4604;
  assign _EVAL_4116 = _EVAL_2538 ? _EVAL_1432 : {{1'd0}, _EVAL_2571};
  assign _EVAL_3593 = $signed(_EVAL_4116);
  assign _EVAL_2192 = _EVAL_1560[4:0];
  assign _EVAL_1005 = $signed(_EVAL_3593) >>> _EVAL_2192;
  assign _EVAL_1735 = _EVAL_1005[31:0];
  assign _EVAL_1774 = _EVAL_1735[31:16];
  assign _EVAL_4144 = {{16'd0}, _EVAL_1774};
  assign _EVAL_3150 = _EVAL_1735[15:0];
  assign _EVAL_1012 = {_EVAL_3150, 16'h0};
  assign _EVAL_1467 = _EVAL_1012 & 32'hffff0000;
  assign _EVAL_426 = _EVAL_4144 | _EVAL_1467;
  assign _EVAL_4981 = _EVAL_426[31:8];
  assign _EVAL_4991 = {{8'd0}, _EVAL_4981};
  assign _EVAL_3782 = _EVAL_4991 & 32'hff00ff;
  assign _EVAL_2348 = _EVAL_426[23:0];
  assign _EVAL_5330 = {_EVAL_2348, 8'h0};
  assign _EVAL_1598 = _EVAL_5330 & 32'hff00ff00;
  assign _EVAL_1563 = _EVAL_3782 | _EVAL_1598;
  assign _EVAL_563 = _EVAL_1563[31:4];
  assign _EVAL_496 = {{4'd0}, _EVAL_563};
  assign _EVAL_4234 = _EVAL_496 & 32'hf0f0f0f;
  assign _EVAL_3665 = _EVAL_1563[27:0];
  assign _EVAL_2526 = {_EVAL_3665, 4'h0};
  assign _EVAL_769 = _EVAL_2526 & 32'hf0f0f0f0;
  assign _EVAL_2336 = _EVAL_4234 | _EVAL_769;
  assign _EVAL_3623 = _EVAL_2336[29:0];
  assign _EVAL_4923 = {_EVAL_3623, 2'h0};
  assign _EVAL_3622 = _EVAL_4923 & 32'hcccccccc;
  assign _EVAL_3431 = _EVAL_4043 | _EVAL_3608;
  assign _EVAL_2197 = _EVAL_2121 | _EVAL_147;
  assign _EVAL_4911 = _EVAL_3888 | _EVAL_2268;
  assign _EVAL_4024 = _EVAL_2506 & _EVAL_4911;
  assign _EVAL_4034 = _EVAL_1352 | _EVAL_951;
  assign _EVAL_3034 = _EVAL_3227 & _EVAL_4034;
  assign _EVAL_3532 = _EVAL_4024 | _EVAL_3034;
  assign _EVAL_4474 = _EVAL_2197 | _EVAL_3532;
  assign _EVAL_627 = _EVAL_58 & _EVAL_2369;
  assign _EVAL_4774 = _EVAL_3094 ? 1'h1 : _EVAL_4000;
  assign _EVAL_4351 = _EVAL_5099 == _EVAL_4460;
  assign _EVAL_3457 = _EVAL_332 & _EVAL_4351;
  assign _EVAL_3876 = _EVAL_4774 & _EVAL_3457;
  assign _EVAL_2700 = _EVAL_2812 == _EVAL_4460;
  assign _EVAL_1297 = _EVAL_5386 & _EVAL_2700;
  assign _EVAL_3273 = _EVAL_5252 & _EVAL_1297;
  assign _EVAL_3279 = _EVAL_3629 ? fpu__EVAL_9 : _EVAL_3727;
  assign _EVAL_3187 = _EVAL_2257 ? divider__EVAL_8 : _EVAL_3279;
  assign _EVAL_4993 = _EVAL_3273 ? _EVAL_3187 : _EVAL_2919;
  assign _EVAL_579 = _EVAL_3876 ? _EVAL_4863 : _EVAL_4993;
  assign _EVAL_3512 = _EVAL_5099 == _EVAL_2495;
  assign _EVAL_1789 = _EVAL_3742 == _EVAL_274;
  assign _EVAL_1963 = _EVAL_2219 & _EVAL_1789;
  assign _EVAL_4016 = _EVAL_780 == 3'h5;
  assign _EVAL_1030 = _EVAL_315 ? _EVAL_119 : _EVAL_260;
  assign _EVAL_5340 = _EVAL_315 ? _EVAL_179 : _EVAL_188;
  assign _EVAL_1843 = _EVAL_1030 ? 1'h1 : _EVAL_5340;
  assign _EVAL_4200 = {{31'd0}, _EVAL_127};
  assign _EVAL_2144 = _EVAL_180 == _EVAL_91;
  assign _EVAL_1112 = _EVAL_269[5];
  assign _EVAL_4686 = {_EVAL_1112,_EVAL_5220,_EVAL_5194,2'h0};
  assign _EVAL_3221 = _EVAL_4686[6:5];
  assign _EVAL_732 = _EVAL_4686[4:0];
  assign _EVAL_636 = {_EVAL_3221,2'h1,_EVAL_3643,2'h1,_EVAL_2725,3'h2,_EVAL_732,7'h27};
  assign _EVAL_1893 = {_EVAL_3221,2'h1,_EVAL_3643,2'h1,_EVAL_2725,3'h2,_EVAL_732,7'h23};
  assign _EVAL_3983 = {_EVAL_3935,_EVAL_5220,3'h0};
  assign _EVAL_2807 = _EVAL_3983[7:5];
  assign _EVAL_1806 = _EVAL_3983[4:0];
  assign _EVAL_1006 = {_EVAL_2807,2'h1,_EVAL_3643,2'h1,_EVAL_2725,3'h3,_EVAL_1806,7'h27};
  assign _EVAL_849 = {_EVAL_3221,2'h1,_EVAL_3643,2'h1,_EVAL_2725,3'h0,_EVAL_732,7'h27};
  assign _EVAL_2735 = {_EVAL_1112,_EVAL_5220,_EVAL_5194,2'h0,2'h1,_EVAL_2725,3'h2,2'h1,_EVAL_3643,7'h7};
  assign _EVAL_4903 = {_EVAL_1112,_EVAL_5220,_EVAL_5194,2'h0,2'h1,_EVAL_2725,3'h2,2'h1,_EVAL_3643,7'h3};
  assign _EVAL_4237 = {_EVAL_3935,_EVAL_5220,3'h0,2'h1,_EVAL_2725,3'h3,2'h1,_EVAL_3643,7'h7};
  assign _EVAL_1882 = _EVAL_269[10:7];
  assign _EVAL_2095 = _EVAL_269[12:11];
  assign _EVAL_4420 = {_EVAL_1882,_EVAL_2095,_EVAL_1112,_EVAL_5194,2'h0,5'h2,3'h0,2'h1,_EVAL_3643,7'h13};
  assign _EVAL_2938 = _EVAL_1897 ? {{2'd0}, _EVAL_4237} : _EVAL_4420;
  assign _EVAL_2000 = _EVAL_654 ? {{3'd0}, _EVAL_4903} : _EVAL_2938;
  assign _EVAL_900 = _EVAL_5161 ? {{3'd0}, _EVAL_2735} : _EVAL_2000;
  assign _EVAL_4306 = _EVAL_4280 ? {{3'd0}, _EVAL_849} : _EVAL_900;
  assign _EVAL_1962 = _EVAL_397 ? {{2'd0}, _EVAL_1006} : _EVAL_4306;
  assign _EVAL_529 = _EVAL_4909 ? {{3'd0}, _EVAL_1893} : _EVAL_1962;
  assign _EVAL_1708 = _EVAL_3284 ? {{3'd0}, _EVAL_636} : _EVAL_529;
  assign _EVAL_961 = {2'h0,_EVAL_1708};
  assign _EVAL_4504 = _EVAL_961 & 32'h64;
  assign _EVAL_2677 = _EVAL_4504 == 32'h0;
  assign _EVAL_2932 = _EVAL_961 & 32'h50;
  assign _EVAL_3328 = _EVAL_2932 == 32'h10;
  assign _EVAL_737 = _EVAL_2677 | _EVAL_3328;
  assign _EVAL_2109 = _EVAL_961 & 32'h2024;
  assign _EVAL_4549 = _EVAL_2109 == 32'h24;
  assign _EVAL_3633 = _EVAL_737 | _EVAL_4549;
  assign _EVAL_2298 = _EVAL_961 & 32'h28;
  assign _EVAL_2421 = _EVAL_2298 == 32'h28;
  assign _EVAL_5184 = _EVAL_3633 | _EVAL_2421;
  assign _EVAL_4454 = _EVAL_961 & 32'h30;
  assign _EVAL_2797 = _EVAL_4454 == 32'h30;
  assign _EVAL_1679 = _EVAL_5184 | _EVAL_2797;
  assign _EVAL_300 = _EVAL_4982 ? 1'h0 : _EVAL_2506;
  assign _EVAL_1416 = _EVAL_3672 ? 1'h0 : _EVAL_300;
  assign _EVAL_5408 = _EVAL_1523 ? 1'h1 : _EVAL_3888;
  assign _EVAL_5094 = _EVAL_2506 == 1'h0;
  assign _EVAL_700 = _EVAL_5094 | _EVAL_3421;
  assign _EVAL_4008 = _EVAL_700 | _EVAL_2268;
  assign _EVAL_3995 = _EVAL_4008 == 1'h0;
  assign _EVAL_1292 = _EVAL_3995 ? 1'h1 : _EVAL_2268;
  assign _EVAL_4605 = _EVAL_147 ? _EVAL_1292 : _EVAL_2268;
  assign _EVAL_3607 = _EVAL_5408 | _EVAL_4605;
  assign _EVAL_2242 = _EVAL_1416 & _EVAL_3607;
  assign _EVAL_4598 = csr__EVAL_102[1];
  assign _EVAL_3071 = _EVAL_4598 == 1'h0;
  assign _EVAL_352 = csr__EVAL_89 & _EVAL_3071;
  assign _EVAL_387 = _EVAL_2644 ? 1'h0 : _EVAL_3227;
  assign _EVAL_4524 = _EVAL_147 ? _EVAL_387 : _EVAL_3227;
  assign _EVAL_4807 = _EVAL_2644 ? 1'h0 : _EVAL_4524;
  assign _EVAL_4476 = _EVAL_1523 ? _EVAL_4807 : _EVAL_4524;
  assign _EVAL_2388 = _EVAL_2644 ? 1'h0 : _EVAL_4476;
  assign _EVAL_2463 = _EVAL_3672 ? _EVAL_2388 : _EVAL_4476;
  assign _EVAL_1281 = _EVAL_352 ? 1'h0 : _EVAL_2463;
  assign _EVAL_4541 = _EVAL_1281 & _EVAL_4034;
  assign _EVAL_4139 = _EVAL_2242 | _EVAL_4541;
  assign _EVAL_3972 = {_EVAL_1241,_EVAL_3935};
  assign _EVAL_717 = _EVAL_3972 == 3'h2;
  assign _EVAL_3580 = _EVAL_3972 == 3'h1;
  assign _EVAL_4847 = _EVAL_3580 ? 3'h4 : 3'h0;
  assign _EVAL_791 = _EVAL_717 ? 3'h6 : _EVAL_4847;
  assign _EVAL_2442 = _EVAL_1617 ? _EVAL_3940 : 32'h0;
  assign _EVAL_1746 = _EVAL_4095 ? _EVAL_4468 : 32'h0;
  assign _EVAL_1063 = _EVAL_2442 | _EVAL_1746;
  assign _EVAL_929 = _EVAL_1063[31:5];
  assign _EVAL_2983 = {_EVAL_929,_EVAL_3366};
  assign _EVAL_2271 = _EVAL_3039[3];
  assign _EVAL_459 = _EVAL_2899 ? 2'h2 : 2'h1;
  assign _EVAL_3646 = {{6'd0}, _EVAL_459};
  assign _EVAL_3966 = 8'h80 | _EVAL_3646;
  assign _EVAL_4547 = {{1'd0}, _EVAL_3966};
  assign _EVAL_280 = _EVAL_49 == 1'h0;
  assign _EVAL_2818 = _EVAL_123 & _EVAL_280;
  assign _EVAL_3534 = _EVAL_2818;
  assign _EVAL_3511 = _EVAL_1241 ? 3'h7 : 3'h0;
  assign _EVAL_1557 = _EVAL_2880[31:2];
  assign _EVAL_2643 = _EVAL_2522 & 32'h2024;
  assign _EVAL_1156 = _EVAL_4873[31:2];
  assign _EVAL_1047 = {{2'd0}, _EVAL_1156};
  assign _EVAL_1981 = _EVAL_1047 & 32'h33333333;
  assign _EVAL_5413 = _EVAL_4873[29:0];
  assign _EVAL_1824 = {_EVAL_5413, 2'h0};
  assign _EVAL_2472 = _EVAL_1824 & 32'hcccccccc;
  assign _EVAL_1193 = _EVAL_1981 | _EVAL_2472;
  assign _EVAL_748 = _EVAL_1193[31:1];
  assign _EVAL_540 = {{1'd0}, _EVAL_748};
  assign _EVAL_5054 = _EVAL_5114 & 32'h2024;
  assign _EVAL_2990 = _EVAL_5054 == 32'h24;
  assign _EVAL_2717 = _EVAL_4014 | _EVAL_3588;
  assign _EVAL_2263 = _EVAL_780 == 3'h0;
  assign _EVAL_458 = _EVAL_1968 ? _EVAL_3432 : 32'h0;
  assign _EVAL_2072 = _EVAL_1737 ? _EVAL_4322 : 32'h0;
  assign _EVAL_1992 = _EVAL_458 | _EVAL_2072;
  assign _EVAL_1105 = _EVAL_1992[31:5];
  assign _EVAL_4109 = {_EVAL_1105,_EVAL_483,1'h1};
  assign _EVAL_2333 = ~ _EVAL_3166;
  assign _EVAL_3734 = _EVAL_4632 ? _EVAL_2333 : _EVAL_3166;
  assign _EVAL_4813 = {_EVAL_3734,_EVAL_4632};
  assign _EVAL_4514 = _EVAL_4109 + _EVAL_4813;
  assign _EVAL_1230 = _EVAL_4514[32:1];
  assign _EVAL_4210 = _EVAL_2263 ? _EVAL_1230 : 32'h0;
  assign _EVAL_5217 = _EVAL_780[2:1];
  assign _EVAL_4230 = _EVAL_5217 == 2'h1;
  assign _EVAL_5138 = {_EVAL_1105,_EVAL_483};
  assign _EVAL_4031 = _EVAL_5138[31];
  assign _EVAL_806 = _EVAL_3734[31];
  assign _EVAL_3709 = _EVAL_4031 ^ _EVAL_806;
  assign _EVAL_3230 = _EVAL_1230[31];
  assign _EVAL_3724 = _EVAL_780[0];
  assign _EVAL_4574 = _EVAL_806 == 1'h0;
  assign _EVAL_5086 = _EVAL_3724 ? _EVAL_4574 : _EVAL_4031;
  assign _EVAL_3886 = _EVAL_3709 ? _EVAL_3230 : _EVAL_5086;
  assign _EVAL_3575 = _EVAL_4230 & _EVAL_3886;
  assign _EVAL_923 = {{31'd0}, _EVAL_3575};
  assign _EVAL_5380 = _EVAL_4210 | _EVAL_923;
  assign _EVAL_1048 = _EVAL_3724 == 1'h0;
  assign _EVAL_3927 = _EVAL_4672 & _EVAL_1048;
  assign _EVAL_4888 = _EVAL_5138 ^ _EVAL_3734;
  assign _EVAL_1140 = _EVAL_3927 ? _EVAL_4888 : 32'h0;
  assign _EVAL_3823 = _EVAL_780 >= 3'h6;
  assign _EVAL_3238 = _EVAL_5138 & _EVAL_3734;
  assign _EVAL_2454 = _EVAL_3823 ? _EVAL_3238 : 32'h0;
  assign _EVAL_3443 = _EVAL_1140 | _EVAL_2454;
  assign _EVAL_2306 = _EVAL_5380 | _EVAL_3443;
  assign _EVAL_3713 = _EVAL_4016 ? _EVAL_4879 : 32'h0;
  assign _EVAL_2102 = _EVAL_780 == 3'h1;
  assign _EVAL_1231 = _EVAL_4983[31:1];
  assign _EVAL_2926 = {{1'd0}, _EVAL_1231};
  assign _EVAL_2558 = _EVAL_2926 & 32'h55555555;
  assign _EVAL_1830 = {_EVAL_4752, 1'h0};
  assign _EVAL_2694 = _EVAL_1830 & 32'haaaaaaaa;
  assign _EVAL_3265 = _EVAL_2558 | _EVAL_2694;
  assign _EVAL_3526 = _EVAL_2102 ? _EVAL_3265 : 32'h0;
  assign _EVAL_4737 = _EVAL_3713 | _EVAL_3526;
  assign _EVAL_1932 = _EVAL_2306 | _EVAL_4737;
  assign _EVAL_5288 = _EVAL_2573 & _EVAL_179;
  assign _EVAL_1180 = _EVAL_171 == _EVAL_3742;
  assign _EVAL_719 = csr__EVAL_70 & _EVAL_869;
  assign _EVAL_2327 = _EVAL_2326 | _EVAL_3624;
  assign _EVAL_3331 = _EVAL_2583 ? _EVAL_3132 : _EVAL_4157;
  assign _EVAL_373 = _EVAL_2423 != _EVAL_3331;
  assign _EVAL_5271 = _EVAL_2327 & _EVAL_373;
  assign _EVAL_1815 = _EVAL_719 | _EVAL_5271;
  assign _EVAL_1558 = _EVAL_2326 | _EVAL_1815;
  assign _EVAL_5056 = _EVAL_3232[8:6];
  assign _EVAL_4544 = _EVAL_5056 == 3'h0;
  assign _EVAL_3258 = _EVAL_4544 == 1'h0;
  assign _EVAL_1098 = _EVAL_3742 == _EVAL_180;
  assign _EVAL_3522 = _EVAL_2219 & _EVAL_1098;
  assign _EVAL_5055 = _EVAL_3227 & _EVAL_3522;
  assign _EVAL_358 = _EVAL_4064[2];
  assign _EVAL_5010 = _EVAL_1818 & _EVAL_3340;
  assign _EVAL_2289 = {_EVAL_5010,_EVAL_2758};
  assign _EVAL_2266 = _EVAL_540 & 32'h55555555;
  assign _EVAL_1373 = _EVAL_1193[30:0];
  assign _EVAL_2726 = {_EVAL_1373, 1'h0};
  assign _EVAL_3635 = _EVAL_2726 & 32'haaaaaaaa;
  assign _EVAL_1880 = _EVAL_2266 | _EVAL_3635;
  assign _EVAL_1801 = _EVAL_358 ? _EVAL_2289 : {{1'd0}, _EVAL_1880};
  assign _EVAL_1427 = $signed(_EVAL_1801);
  assign _EVAL_3283 = _EVAL_1731[4:0];
  assign _EVAL_803 = $signed(_EVAL_1427) >>> _EVAL_3283;
  assign _EVAL_1505 = _EVAL_803[31:0];
  assign _EVAL_3885 = _EVAL_1505[31:16];
  assign _EVAL_2892 = _EVAL_315 ? _EVAL_251 : _EVAL_115;
  assign _EVAL_2973 = _EVAL_315 ? _EVAL_71 : _EVAL_106;
  assign _EVAL_2041 = _EVAL_315 ? _EVAL_78 : _EVAL_186;
  assign _EVAL_4089 = _EVAL_2041 ? 3'h4 : 3'h6;
  assign _EVAL_2636 = _EVAL_2041 ? 4'h6 : 4'h8;
  assign _EVAL_5321 = _EVAL_2973 ? {{1'd0}, _EVAL_4089} : _EVAL_2636;
  assign _EVAL_3379 = _EVAL_2041 ? 3'h2 : 3'h4;
  assign _EVAL_2303 = _EVAL_2892 ? _EVAL_5321 : {{1'd0}, _EVAL_3379};
  assign _EVAL_4755 = _EVAL_2303 == 4'h2;
  assign _EVAL_5232 = _EVAL_315 ? _EVAL_115 : _EVAL_251;
  assign _EVAL_4880 = _EVAL_315 ? _EVAL_106 : _EVAL_71;
  assign _EVAL_4361 = _EVAL_315 ? _EVAL_186 : _EVAL_78;
  assign _EVAL_3578 = _EVAL_4361 ? 3'h4 : 3'h6;
  assign _EVAL_3961 = _EVAL_4361 ? 4'h6 : 4'h8;
  assign _EVAL_364 = _EVAL_4880 ? {{1'd0}, _EVAL_3578} : _EVAL_3961;
  assign _EVAL_991 = _EVAL_4361 ? 3'h2 : 3'h4;
  assign _EVAL_311 = _EVAL_5232 ? _EVAL_364 : {{1'd0}, _EVAL_991};
  assign _EVAL_4517 = _EVAL_311 == 4'h2;
  assign _EVAL_5411 = _EVAL_4755 & _EVAL_4517;
  assign _EVAL_585 = _EVAL_2400[6];
  assign _EVAL_3924 = _EVAL_315 ? _EVAL_171 : _EVAL_91;
  assign _EVAL_4298 = _EVAL_3924[0];
  assign _EVAL_5377 = _EVAL_2400[5:0];
  assign _EVAL_470 = _EVAL_3924[4:1];
  assign _EVAL_2249 = {_EVAL_585,_EVAL_4298,_EVAL_5377,_EVAL_470,1'h0};
  assign _EVAL_4890 = $signed(_EVAL_2249);
  assign _EVAL_884 = $unsigned(_EVAL_4890);
  assign _EVAL_2317 = _EVAL_884 == 13'h4;
  assign _EVAL_772 = _EVAL_5411 & _EVAL_2317;
  assign _EVAL_3057 = _EVAL_311 == 4'h4;
  assign _EVAL_5157 = _EVAL_4755 & _EVAL_3057;
  assign _EVAL_607 = _EVAL_884 == 13'h6;
  assign _EVAL_2387 = _EVAL_5157 & _EVAL_607;
  assign _EVAL_4264 = _EVAL_772 | _EVAL_2387;
  assign _EVAL_2768 = _EVAL_2303 == 4'h4;
  assign _EVAL_1304 = _EVAL_2768 & _EVAL_4517;
  assign _EVAL_5142 = _EVAL_1304 & _EVAL_607;
  assign _EVAL_3947 = _EVAL_4264 | _EVAL_5142;
  assign _EVAL_826 = _EVAL_2768 & _EVAL_3057;
  assign _EVAL_3356 = _EVAL_884 == 13'h8;
  assign _EVAL_4172 = _EVAL_826 & _EVAL_3356;
  assign _EVAL_3107 = _EVAL_3947 | _EVAL_4172;
  assign _EVAL_2693 = _EVAL_3107 == 1'h0;
  assign _EVAL_2577 = _EVAL_3796 - 8'h81;
  assign _EVAL_5338 = _EVAL_3309 == 5'h1c;
  assign _EVAL_5241 = _EVAL_3309 == 5'h1b;
  assign _EVAL_4545 = _EVAL_5241 ? _EVAL_1703 : _EVAL_5018;
  assign _EVAL_3474 = _EVAL_5338 ? _EVAL_1407 : _EVAL_4545;
  assign _EVAL_2436 = _EVAL_1 & _EVAL_1996;
  assign _EVAL_3948 = _EVAL_4043 & _EVAL_2436;
  assign _EVAL_2620 = _EVAL_205 & _EVAL_3318;
  assign _EVAL_3783 = _EVAL_4043 & _EVAL_2620;
  assign _EVAL_5097 = _EVAL_315 ? _EVAL_3948 : _EVAL_3783;
  assign _EVAL_4580 = _EVAL_4240 & _EVAL_946;
  assign _EVAL_1950 = {_EVAL_260,_EVAL_3212};
  assign _EVAL_4951 = _EVAL_4160 >> _EVAL_1950;
  assign _EVAL_4865 = _EVAL_4951[0];
  assign _EVAL_5274 = _EVAL_2823 == _EVAL_1950;
  assign _EVAL_4421 = _EVAL_1535 & _EVAL_5274;
  assign _EVAL_2246 = _EVAL_4865 | _EVAL_4421;
  assign _EVAL_3124 = _EVAL_2617 == _EVAL_1950;
  assign _EVAL_1093 = divider__EVAL_2 & _EVAL_3124;
  assign _EVAL_1345 = _EVAL_2246 | _EVAL_1093;
  assign _EVAL_2569 = _EVAL_4158 == _EVAL_1950;
  assign _EVAL_667 = _EVAL_1190 & _EVAL_2569;
  assign _EVAL_4039 = _EVAL_1345 | _EVAL_667;
  assign _EVAL_532 = _EVAL_260 & _EVAL_4039;
  assign _EVAL_4634 = _EVAL_4614[1];
  assign _EVAL_5120 = _EVAL_1699 & _EVAL_4634;
  assign _EVAL_3856 = _EVAL_58 & _EVAL_4962;
  assign _EVAL_3456 = _EVAL_268 & _EVAL_1333;
  assign _EVAL_2477 = _EVAL_3856 | _EVAL_3456;
  assign _EVAL_3854 = _EVAL_91 == _EVAL_4706;
  assign _EVAL_2733 = _EVAL_2477 & _EVAL_3854;
  assign _EVAL_2467 = _EVAL_171 == _EVAL_4706;
  assign _EVAL_4227 = _EVAL_3702 & _EVAL_2467;
  assign _EVAL_740 = _EVAL_315 ? _EVAL_2733 : _EVAL_4227;
  assign _EVAL_4714 = _EVAL_2506 & _EVAL_740;
  assign _EVAL_4729 = fpu__EVAL_12 & fpu__EVAL_55;
  assign _EVAL_4920 = _EVAL_4729 & _EVAL_998;
  assign _EVAL_4208 = _EVAL_4920 ? fpu__EVAL_21 : _EVAL_2741__EVAL_2749_data;
  assign _EVAL_2914 = _EVAL_2573 & _EVAL_39;
  assign _EVAL_2884 = _EVAL_1724 & _EVAL_205;
  assign _EVAL_1607 = _EVAL_2914 | _EVAL_2884;
  assign _EVAL_2727 = _EVAL_1607 & _EVAL_5318;
  assign _EVAL_3700 = _EVAL_2573 & _EVAL_188;
  assign _EVAL_4266 = _EVAL_1724 & _EVAL_250;
  assign _EVAL_4353 = _EVAL_3700 | _EVAL_4266;
  assign _EVAL_2054 = _EVAL_180 == _EVAL_3670;
  assign _EVAL_3525 = _EVAL_4353 & _EVAL_2054;
  assign _EVAL_1484 = _EVAL_2727 | _EVAL_3525;
  assign _EVAL_4018 = _EVAL_2573 & _EVAL_260;
  assign _EVAL_5326 = _EVAL_3212 == _EVAL_3670;
  assign _EVAL_1934 = _EVAL_4018 & _EVAL_5326;
  assign _EVAL_3353 = _EVAL_1484 | _EVAL_1934;
  assign _EVAL_4970 = _EVAL_154 == _EVAL_3670;
  assign _EVAL_4433 = _EVAL_1527 & _EVAL_4970;
  assign _EVAL_4406 = _EVAL_1724 & _EVAL_141;
  assign _EVAL_4060 = _EVAL_5288 | _EVAL_4406;
  assign _EVAL_3157 = _EVAL_68 == _EVAL_3670;
  assign _EVAL_5315 = _EVAL_4060 & _EVAL_3157;
  assign _EVAL_1068 = _EVAL_4433 | _EVAL_5315;
  assign _EVAL_4587 = _EVAL_2573 & _EVAL_119;
  assign _EVAL_5198 = _EVAL_4127 == _EVAL_3670;
  assign _EVAL_4780 = _EVAL_4587 & _EVAL_5198;
  assign _EVAL_3304 = _EVAL_1068 | _EVAL_4780;
  assign _EVAL_2141 = _EVAL_315 ? _EVAL_3353 : _EVAL_3304;
  assign _EVAL_650 = _EVAL_3624 & _EVAL_2141;
  assign _EVAL_2157 = _EVAL_4203 ? 3'h2 : 3'h4;
  assign _EVAL_4439 = _EVAL_4203 ? 3'h4 : 3'h6;
  assign _EVAL_4104 = _EVAL_2060 ? _EVAL_2157 : _EVAL_4439;
  assign _EVAL_2111 = _EVAL_4203 ? 2'h0 : 2'h2;
  assign _EVAL_4794 = _EVAL_2603 ? _EVAL_4104 : {{1'd0}, _EVAL_2111};
  assign _EVAL_4595 = _EVAL_4971 + _EVAL_4794;
  assign _EVAL_4214 = _EVAL_154 == _EVAL_5129;
  assign _EVAL_5373 = _EVAL_148 & _EVAL_4214;
  assign _EVAL_5248 = _EVAL_261 == 1'h0;
  assign _EVAL_1905 = _EVAL_5248 | _EVAL_118;
  assign _EVAL_1002 = _EVAL_1905 == 1'h0;
  assign _EVAL_3746 = _EVAL_3421 == 1'h0;
  assign _EVAL_2159 = _EVAL_3405 == 32'h3;
  assign _EVAL_1857 = _EVAL_3405 == 32'h1;
  assign _EVAL_1713 = _EVAL_2159 | _EVAL_1857;
  assign _EVAL_1729 = _EVAL_1713 | _EVAL_4309;
  assign _EVAL_3884 = _EVAL_3746 | _EVAL_1729;
  assign _EVAL_2365 = _EVAL_649[4];
  assign _EVAL_3440 = _EVAL_2365 == 1'h0;
  assign _EVAL_779 = _EVAL_649[3];
  assign _EVAL_4007 = _EVAL_3440 & _EVAL_779;
  assign _EVAL_1849 = _EVAL_649[1];
  assign _EVAL_4376 = _EVAL_1849 == 1'h0;
  assign _EVAL_1215 = _EVAL_4007 & _EVAL_4376;
  assign _EVAL_918 = _EVAL_2965 & _EVAL_2271;
  assign _EVAL_1529 = _EVAL_3039[0];
  assign _EVAL_5203 = _EVAL_1529 == 1'h0;
  assign _EVAL_377 = _EVAL_918 & _EVAL_5203;
  assign _EVAL_3123 = _EVAL_4192[0];
  assign _EVAL_1397 = _EVAL_377 & _EVAL_3123;
  assign _EVAL_1458 = _EVAL_1379[2];
  assign _EVAL_4608 = _EVAL_1397 & _EVAL_1458;
  assign _EVAL_5324 = _EVAL_4608 & _EVAL_1414;
  assign _EVAL_3387 = _EVAL_4530[4];
  assign _EVAL_5222 = _EVAL_3387 == 1'h0;
  assign _EVAL_2925 = _EVAL_4530[2];
  assign _EVAL_2593 = _EVAL_5222 & _EVAL_2925;
  assign _EVAL_2358 = _EVAL_4530[3];
  assign _EVAL_2828 = _EVAL_2593 & _EVAL_2358;
  assign _EVAL_1587 = _EVAL_4530[0];
  assign _EVAL_3917 = _EVAL_1587 == 1'h0;
  assign _EVAL_981 = _EVAL_2828 & _EVAL_3917;
  assign _EVAL_2416 = _EVAL_2030[0];
  assign _EVAL_5261 = _EVAL_981 & _EVAL_2416;
  assign _EVAL_4152 = _EVAL_3922[2];
  assign _EVAL_1823 = _EVAL_5261 & _EVAL_4152;
  assign _EVAL_5034 = _EVAL_1823 & _EVAL_1319;
  assign _EVAL_977 = _EVAL_5324 | _EVAL_5034;
  assign _EVAL_781 = _EVAL_3568 & _EVAL_3360;
  assign _EVAL_1697 = _EVAL_16 & _EVAL_2369;
  assign _EVAL_2287 = _EVAL_214 & _EVAL_2219;
  assign _EVAL_1497 = _EVAL_1697 | _EVAL_2287;
  assign _EVAL_4937 = _EVAL_1497 & _EVAL_1180;
  assign _EVAL_3423 = _EVAL_268 & _EVAL_2219;
  assign _EVAL_3915 = _EVAL_627 | _EVAL_3423;
  assign _EVAL_796 = _EVAL_91 == _EVAL_3742;
  assign _EVAL_2654 = _EVAL_3915 & _EVAL_796;
  assign _EVAL_2551 = _EVAL_315 ? _EVAL_4937 : _EVAL_2654;
  assign _EVAL_1405 = _EVAL_3227 & _EVAL_2551;
  assign _EVAL_1742 = _EVAL_315 ? _EVAL_1405 : _EVAL_1405;
  assign _EVAL_478 = _EVAL_781 & _EVAL_1742;
  assign _EVAL_3825 = _EVAL_977 | _EVAL_478;
  assign _EVAL_3896 = _EVAL_315 ^ _EVAL_98;
  assign _EVAL_2231 = _EVAL_3896 ^ 1'h1;
  assign _EVAL_1776 = _EVAL_58 & _EVAL_39;
  assign _EVAL_1721 = _EVAL_268 & _EVAL_205;
  assign _EVAL_520 = _EVAL_1776 | _EVAL_1721;
  assign _EVAL_1444 = _EVAL_274 == _EVAL_91;
  assign _EVAL_2318 = _EVAL_520 & _EVAL_1444;
  assign _EVAL_2943 = _EVAL_58 & _EVAL_188;
  assign _EVAL_3202 = _EVAL_268 & _EVAL_250;
  assign _EVAL_2023 = _EVAL_2943 | _EVAL_3202;
  assign _EVAL_4816 = _EVAL_2023 & _EVAL_2144;
  assign _EVAL_4341 = _EVAL_2318 | _EVAL_4816;
  assign _EVAL_4521 = _EVAL_58 & _EVAL_260;
  assign _EVAL_2779 = _EVAL_3212 == _EVAL_91;
  assign _EVAL_384 = _EVAL_4521 & _EVAL_2779;
  assign _EVAL_1524 = _EVAL_4341 | _EVAL_384;
  assign _EVAL_1366 = _EVAL_16 & _EVAL_58;
  assign _EVAL_5026 = _EVAL_214 & _EVAL_268;
  assign _EVAL_4801 = _EVAL_1366 | _EVAL_5026;
  assign _EVAL_4741 = _EVAL_171 == _EVAL_91;
  assign _EVAL_347 = _EVAL_4801 & _EVAL_4741;
  assign _EVAL_415 = _EVAL_1524 | _EVAL_347;
  assign _EVAL_3100 = _EVAL_5289 == 1'h0;
  assign _EVAL_1759 = _EVAL_3226 & _EVAL_3100;
  assign _EVAL_400 = _EVAL_40 == 1'h0;
  assign _EVAL_1279 = _EVAL_153 == 3'h5;
  assign _EVAL_4171 = _EVAL_153 == 3'h6;
  assign _EVAL_2053 = _EVAL_1279 | _EVAL_4171;
  assign _EVAL_2547 = csr__EVAL_134 | _EVAL_2053;
  assign _EVAL_519 = _EVAL_153 == 3'h7;
  assign _EVAL_3843 = _EVAL_519 & _EVAL_1144;
  assign _EVAL_5423 = _EVAL_2547 | _EVAL_3843;
  assign _EVAL_4124 = _EVAL_3111 & _EVAL_5423;
  assign _EVAL_2274 = _EVAL_400 | _EVAL_4124;
  assign _EVAL_897 = _EVAL_154 != _EVAL_154;
  assign _EVAL_1564 = _EVAL_1 & _EVAL_897;
  assign _EVAL_836 = _EVAL_141 & _EVAL_1775;
  assign _EVAL_5158 = _EVAL_1564 | _EVAL_836;
  assign _EVAL_5143 = _EVAL_2274 | _EVAL_5158;
  assign _EVAL_4506 = _EVAL_1759 | _EVAL_5143;
  assign _EVAL_2528 = {_EVAL_32,_EVAL_172,_EVAL_212,_EVAL_165};
  assign _EVAL_1576 = _EVAL_2528 != 4'h0;
  assign _EVAL_3220 = _EVAL_4506 | _EVAL_1576;
  assign _EVAL_647 = _EVAL_3220 | _EVAL_184;
  assign _EVAL_1086 = _EVAL_415 | _EVAL_647;
  assign _EVAL_5395 = _EVAL_16 & _EVAL_148;
  assign _EVAL_1813 = _EVAL_214 & _EVAL_1;
  assign _EVAL_4641 = _EVAL_5395 | _EVAL_1813;
  assign _EVAL_4921 = _EVAL_154 == _EVAL_171;
  assign _EVAL_4456 = _EVAL_4641 & _EVAL_4921;
  assign _EVAL_3458 = _EVAL_16 & _EVAL_179;
  assign _EVAL_1635 = _EVAL_214 & _EVAL_141;
  assign _EVAL_3286 = _EVAL_3458 | _EVAL_1635;
  assign _EVAL_5192 = _EVAL_68 == _EVAL_171;
  assign _EVAL_1441 = _EVAL_3286 & _EVAL_5192;
  assign _EVAL_2166 = _EVAL_4456 | _EVAL_1441;
  assign _EVAL_2167 = _EVAL_16 & _EVAL_119;
  assign _EVAL_5164 = _EVAL_4127 == _EVAL_171;
  assign _EVAL_4687 = _EVAL_2167 & _EVAL_5164;
  assign _EVAL_1413 = _EVAL_2166 | _EVAL_4687;
  assign _EVAL_1651 = _EVAL_58 & _EVAL_16;
  assign _EVAL_2196 = _EVAL_268 & _EVAL_214;
  assign _EVAL_3215 = _EVAL_1651 | _EVAL_2196;
  assign _EVAL_4112 = _EVAL_91 == _EVAL_171;
  assign _EVAL_4795 = _EVAL_3215 & _EVAL_4112;
  assign _EVAL_1510 = _EVAL_1413 | _EVAL_4795;
  assign _EVAL_2976 = _EVAL_2908 == 1'h0;
  assign _EVAL_5302 = _EVAL_1661 & _EVAL_2976;
  assign _EVAL_2691 = _EVAL_59 == 1'h0;
  assign _EVAL_1310 = _EVAL_16 | _EVAL_39;
  assign _EVAL_464 = _EVAL_1310 | _EVAL_188;
  assign _EVAL_3103 = _EVAL_84 == 3'h5;
  assign _EVAL_5047 = _EVAL_84 == 3'h6;
  assign _EVAL_5002 = _EVAL_3103 | _EVAL_5047;
  assign _EVAL_3594 = csr__EVAL_134 | _EVAL_5002;
  assign _EVAL_552 = _EVAL_84 == 3'h7;
  assign _EVAL_4510 = _EVAL_552 & _EVAL_1144;
  assign _EVAL_2337 = _EVAL_3594 | _EVAL_4510;
  assign _EVAL_1869 = _EVAL_464 & _EVAL_2337;
  assign _EVAL_1424 = _EVAL_2691 | _EVAL_1869;
  assign _EVAL_2330 = _EVAL_274 != _EVAL_274;
  assign _EVAL_4100 = _EVAL_205 & _EVAL_2330;
  assign _EVAL_4864 = _EVAL_180 != _EVAL_180;
  assign _EVAL_1698 = _EVAL_250 & _EVAL_4864;
  assign _EVAL_1808 = _EVAL_4100 | _EVAL_1698;
  assign _EVAL_2461 = _EVAL_1424 | _EVAL_1808;
  assign _EVAL_5066 = _EVAL_5302 | _EVAL_2461;
  assign _EVAL_567 = {_EVAL_80,_EVAL_213,_EVAL_92,_EVAL_204};
  assign _EVAL_3174 = _EVAL_567 != 4'h0;
  assign _EVAL_1632 = _EVAL_5066 | _EVAL_3174;
  assign _EVAL_5355 = _EVAL_1632 | _EVAL_198;
  assign _EVAL_1640 = _EVAL_1510 | _EVAL_5355;
  assign _EVAL_3632 = _EVAL_315 ? _EVAL_1086 : _EVAL_1640;
  assign _EVAL_4247 = _EVAL_315 ? _EVAL_5355 : _EVAL_647;
  assign _EVAL_1646 = csr__EVAL_105 ? 1'h1 : _EVAL_4247;
  assign _EVAL_1547 = _EVAL_3632 | _EVAL_1646;
  assign _EVAL_518 = _EVAL_315 ? _EVAL_1661 : _EVAL_3226;
  assign _EVAL_3015 = _EVAL_1547 | _EVAL_518;
  assign _EVAL_324 = _EVAL_240[16];
  assign _EVAL_3951 = _EVAL_324 == 1'h0;
  assign _EVAL_1672 = _EVAL_3989 & _EVAL_3951;
  assign _EVAL_1979 = _EVAL_2317 | _EVAL_607;
  assign _EVAL_1894 = _EVAL_4517 & _EVAL_1979;
  assign _EVAL_5383 = _EVAL_607 | _EVAL_3356;
  assign _EVAL_4849 = _EVAL_3057 & _EVAL_5383;
  assign _EVAL_1451 = _EVAL_1894 | _EVAL_4849;
  assign _EVAL_1046 = _EVAL_1672 & _EVAL_1451;
  assign _EVAL_5319 = _EVAL_3015 | _EVAL_1046;
  assign _EVAL_538 = _EVAL_2231 & _EVAL_5319;
  assign _EVAL_4386 = _EVAL_3825 | _EVAL_538;
  assign _EVAL_2345 = _EVAL_4386 | _EVAL_601;
  assign _EVAL_3498 = _EVAL_3742 == _EVAL_1059;
  assign _EVAL_2734 = _EVAL_4721 & _EVAL_4736;
  assign _EVAL_2064 = _EVAL_4721 + _EVAL_2734;
  assign _EVAL_2003 = _EVAL_890 & _EVAL_1499;
  assign _EVAL_4751 = _EVAL_890 + _EVAL_2003;
  assign _EVAL_4776 = _EVAL_2064 + _EVAL_4751;
  assign _EVAL_2927 = _EVAL_4776[0];
  assign _EVAL_766 = _EVAL_2231 < 1'h1;
  assign _EVAL_626 = _EVAL_237 | _EVAL_766;
  assign _EVAL_3184 = _EVAL_1241 ? 5'h1f : 5'h0;
  assign _EVAL_2655 = _EVAL_269[11:10];
  assign _EVAL_3253 = _EVAL_269[4:3];
  assign _EVAL_1159 = {_EVAL_3184,_EVAL_3935,_EVAL_2243,_EVAL_2655,_EVAL_3253,1'h0};
  assign _EVAL_4702 = _EVAL_1159[12];
  assign _EVAL_453 = _EVAL_1159[10:5];
  assign _EVAL_2381 = _EVAL_1159[4:1];
  assign _EVAL_2949 = _EVAL_1159[11];
  assign _EVAL_814 = {_EVAL_4702,_EVAL_453,5'h0,2'h1,_EVAL_2725,3'h1,_EVAL_2381,_EVAL_2949,7'h63};
  assign _EVAL_3351 = {_EVAL_4702,_EVAL_453,5'h0,2'h1,_EVAL_2725,3'h0,_EVAL_2381,_EVAL_2949,7'h63};
  assign _EVAL_2071 = {_EVAL_2978,_EVAL_1285,_EVAL_4259,_EVAL_2173,5'h0,7'h6f};
  assign _EVAL_3131 = _EVAL_2655 == 2'h3;
  assign _EVAL_3655 = _EVAL_3972 == 3'h7;
  assign _EVAL_555 = _EVAL_3972 == 3'h6;
  assign _EVAL_4857 = _EVAL_3972 == 3'h5;
  assign _EVAL_4198 = _EVAL_3972 == 3'h4;
  assign _EVAL_3657 = _EVAL_3972 == 3'h3;
  assign _EVAL_975 = _EVAL_3657 ? 3'h7 : _EVAL_791;
  assign _EVAL_2684 = _EVAL_4198 ? 3'h0 : _EVAL_975;
  assign _EVAL_4037 = _EVAL_4857 ? 3'h0 : _EVAL_2684;
  assign _EVAL_1498 = _EVAL_555 ? 3'h2 : _EVAL_4037;
  assign _EVAL_1254 = _EVAL_3655 ? 3'h3 : _EVAL_1498;
  assign _EVAL_1391 = _EVAL_1241 ? 7'h3b : 7'h33;
  assign _EVAL_4487 = {2'h1,_EVAL_3643,2'h1,_EVAL_2725,_EVAL_1254,2'h1,_EVAL_2725,_EVAL_1391};
  assign _EVAL_5304 = {{6'd0}, _EVAL_4487};
  assign _EVAL_5125 = _EVAL_3935 == 2'h0;
  assign _EVAL_733 = {_EVAL_5125, 30'h0};
  assign _EVAL_2623 = _EVAL_5304 | _EVAL_733;
  assign _EVAL_1797 = _EVAL_2655 == 2'h2;
  assign _EVAL_1410 = _EVAL_1241 ? 7'h7f : 7'h0;
  assign _EVAL_2462 = {_EVAL_1410,_EVAL_5394,2'h1,_EVAL_2725,3'h7,2'h1,_EVAL_2725,7'h13};
  assign _EVAL_5359 = _EVAL_2655 == 2'h1;
  assign _EVAL_628 = {_EVAL_1241,_EVAL_5394,2'h1,_EVAL_2725,3'h5,2'h1,_EVAL_2725,7'h13};
  assign _EVAL_4619 = {{5'd0}, _EVAL_628};
  assign _EVAL_5308 = _EVAL_4619 | 31'h40000000;
  assign _EVAL_679 = _EVAL_5359 ? _EVAL_5308 : {{5'd0}, _EVAL_628};
  assign _EVAL_1317 = _EVAL_1797 ? _EVAL_2462 : {{1'd0}, _EVAL_679};
  assign _EVAL_795 = _EVAL_3131 ? {{1'd0}, _EVAL_2623} : _EVAL_1317;
  assign _EVAL_2324 = _EVAL_475 == 5'h2;
  assign _EVAL_4563 = {_EVAL_3511,_EVAL_3253,_EVAL_1112,_EVAL_2243,_EVAL_5194,4'h0,_EVAL_475,3'h0,_EVAL_475,7'h13};
  assign _EVAL_5365 = _EVAL_1241 ? 15'h7fff : 15'h0;
  assign _EVAL_1313 = {_EVAL_5365,_EVAL_5394,12'h0};
  assign _EVAL_2521 = _EVAL_1313[31:12];
  assign _EVAL_5078 = {_EVAL_2521,_EVAL_475,7'h37};
  assign _EVAL_1353 = _EVAL_2324 ? _EVAL_4563 : _EVAL_5078;
  assign _EVAL_2247 = {_EVAL_1410,_EVAL_5394,5'h0,3'h0,_EVAL_475,7'h13};
  assign _EVAL_2253 = {_EVAL_1410,_EVAL_5394,_EVAL_475,3'h0,_EVAL_475,7'h13};
  assign _EVAL_2204 = _EVAL_1897 ? _EVAL_1628 : _EVAL_2253;
  assign _EVAL_705 = _EVAL_654 ? _EVAL_2247 : _EVAL_2204;
  assign _EVAL_3257 = _EVAL_5161 ? _EVAL_1353 : _EVAL_705;
  assign _EVAL_3261 = _EVAL_4280 ? _EVAL_795 : _EVAL_3257;
  assign _EVAL_4584 = _EVAL_397 ? _EVAL_2071 : _EVAL_3261;
  assign _EVAL_4856 = _EVAL_4909 ? _EVAL_3351 : _EVAL_4584;
  assign _EVAL_1475 = _EVAL_3284 ? _EVAL_814 : _EVAL_4856;
  assign _EVAL_4855 = _EVAL_1475 & 32'h2024;
  assign _EVAL_1262 = _EVAL_4855 == 32'h24;
  assign _EVAL_2224 = _EVAL_3309 == 5'h1d;
  assign _EVAL_5291 = _EVAL_2224 ? _EVAL_1407 : _EVAL_3474;
  assign _EVAL_2964 = _EVAL_153[2];
  assign _EVAL_2619 = csr__EVAL_167;
  assign _EVAL_1244 = _EVAL_2619[2];
  assign _EVAL_1049 = _EVAL_21 | 32'h3;
  assign _EVAL_517 = _EVAL_1049 & 32'h30;
  assign _EVAL_4226 = _EVAL_3504 == 1'h0;
  assign _EVAL_2146 = _EVAL_3085 & _EVAL_4226;
  assign _EVAL_1555 = _EVAL_3229[6:2];
  assign _EVAL_5414 = _EVAL_1555 == 5'h0;
  assign _EVAL_346 = _EVAL_1555 == 5'h1;
  assign _EVAL_5393 = _EVAL_5414 | _EVAL_346;
  assign _EVAL_3372 = _EVAL_1555 == 5'h2;
  assign _EVAL_1426 = _EVAL_5393 | _EVAL_3372;
  assign _EVAL_3416 = _EVAL_1555 == 5'h3;
  assign _EVAL_5042 = _EVAL_1555 == 5'h7;
  assign _EVAL_2185 = _EVAL_3416 | _EVAL_5042;
  assign _EVAL_4568 = _EVAL_1555 == 5'hb;
  assign _EVAL_4793 = _EVAL_2185 | _EVAL_4568;
  assign _EVAL_3680 = _EVAL_1555 == 5'hf;
  assign _EVAL_2515 = _EVAL_4793 | _EVAL_3680;
  assign _EVAL_848 = _EVAL_1426 | _EVAL_2515;
  assign _EVAL_1015 = _EVAL_848 == 1'h0;
  assign _EVAL_1246 = _EVAL_2146 & _EVAL_1015;
  assign _EVAL_2110 = _EVAL_1913[22:0];
  assign _EVAL_3088 = _EVAL_315 ? _EVAL_188 : _EVAL_179;
  assign _EVAL_768 = _EVAL_315 ? _EVAL_3907 : _EVAL_5224;
  assign _EVAL_2449 = _EVAL_269[1:0];
  assign _EVAL_757 = _EVAL_2449 == 2'h3;
  assign _EVAL_3705 = _EVAL_269 | 32'h3;
  assign _EVAL_4869 = _EVAL_3705[19:15];
  assign _EVAL_544 = _EVAL_2449 == 2'h2;
  assign _EVAL_3171 = _EVAL_2522[19:15];
  assign _EVAL_2180 = _EVAL_2449 == 2'h1;
  assign _EVAL_2991 = _EVAL_1475[19:15];
  assign _EVAL_2074 = _EVAL_961[19:15];
  assign _EVAL_3806 = _EVAL_2180 ? _EVAL_2991 : _EVAL_2074;
  assign _EVAL_675 = _EVAL_544 ? _EVAL_3171 : _EVAL_3806;
  assign _EVAL_4252 = _EVAL_757 ? _EVAL_4869 : _EVAL_675;
  assign _EVAL_1206 = _EVAL_3176 == 1'h0;
  assign _EVAL_2763 = csr__EVAL_39;
  assign _EVAL_3149 = _EVAL_2763 == 1'h0;
  assign _EVAL_4688 = csr__EVAL_152;
  assign _EVAL_5378 = csr__EVAL_59;
  assign _EVAL_2012 = {_EVAL_4688,1'h0,1'h0,_EVAL_5378};
  assign _EVAL_5087 = _EVAL_2012 >> _EVAL_5168;
  assign _EVAL_1940 = _EVAL_5087[0];
  assign _EVAL_4215 = _EVAL_3149 & _EVAL_1940;
  assign _EVAL_2135 = csr__EVAL_3;
  assign _EVAL_4823 = _EVAL_4215 & _EVAL_2135;
  assign _EVAL_1139 = csr__EVAL_31;
  assign _EVAL_2134 = _EVAL_1139[1];
  assign _EVAL_3641 = _EVAL_4679;
  assign _EVAL_4885 = csr__EVAL_64;
  assign _EVAL_597 = _EVAL_3641 >= _EVAL_4885;
  assign _EVAL_4221 = _EVAL_1139[0];
  assign _EVAL_3210 = _EVAL_597 ^ _EVAL_4221;
  assign _EVAL_2867 = ~ _EVAL_3641;
  assign _EVAL_3930 = _EVAL_4885[0];
  assign _EVAL_1603 = _EVAL_4221 & _EVAL_3930;
  assign _EVAL_2940 = _EVAL_4885[1];
  assign _EVAL_5385 = _EVAL_1603 & _EVAL_2940;
  assign _EVAL_3075 = _EVAL_4885[2];
  assign _EVAL_641 = _EVAL_5385 & _EVAL_3075;
  assign _EVAL_331 = {_EVAL_641,_EVAL_5385,_EVAL_1603,_EVAL_4221};
  assign _EVAL_1079 = {{28'd0}, _EVAL_331};
  assign _EVAL_5297 = _EVAL_2867 | _EVAL_1079;
  assign _EVAL_2346 = ~ _EVAL_4885;
  assign _EVAL_1138 = _EVAL_2346 | _EVAL_1079;
  assign _EVAL_4085 = _EVAL_5297 == _EVAL_1138;
  assign _EVAL_2229 = _EVAL_2134 ? _EVAL_3210 : _EVAL_4085;
  assign _EVAL_2435 = _EVAL_4823 & _EVAL_2229;
  assign _EVAL_4624 = _EVAL_4530[4:2];
  assign _EVAL_2922 = _EVAL_4624 == 3'h7;
  assign _EVAL_3831 = _EVAL_3922[1:0];
  assign _EVAL_4163 = _EVAL_3831 != 2'h0;
  assign _EVAL_4044 = _EVAL_2922 & _EVAL_4163;
  assign _EVAL_5167 = _EVAL_4044 == 1'h0;
  assign _EVAL_5170 = _EVAL_3208 ? _EVAL_1024 : 3'h2;
  assign _EVAL_4699 = {{2'd0}, _EVAL_3188};
  assign _EVAL_1300 = _EVAL_5170 ^ _EVAL_4699;
  assign _EVAL_707 = _EVAL_1300[1];
  assign _EVAL_1100 = _EVAL_3401 | _EVAL_922;
  assign _EVAL_1487 = _EVAL_922 == 1'h0;
  assign _EVAL_1533 = _EVAL_1487 & _EVAL_340;
  assign _EVAL_3540 = _EVAL_4706 == _EVAL_1059;
  assign _EVAL_629 = _EVAL_1333 & _EVAL_3540;
  assign _EVAL_5183 = _EVAL_2506 & _EVAL_629;
  assign _EVAL_2869 = _EVAL_116 & _EVAL_159;
  assign _EVAL_702 = _EVAL_4162 == 3'h0;
  assign _EVAL_3037 = {_EVAL_330,_EVAL_1827,1'h1};
  assign _EVAL_2782 = _EVAL_3037 + _EVAL_4503;
  assign _EVAL_3892 = _EVAL_2782[32:1];
  assign _EVAL_5117 = _EVAL_702 ? _EVAL_3892 : 32'h0;
  assign _EVAL_1101 = _EVAL_4162[2:1];
  assign _EVAL_1941 = _EVAL_1101 == 2'h1;
  assign _EVAL_782 = _EVAL_1141[31];
  assign _EVAL_3938 = _EVAL_3901[31];
  assign _EVAL_2647 = _EVAL_782 ^ _EVAL_3938;
  assign _EVAL_1494 = _EVAL_3892[31];
  assign _EVAL_4413 = _EVAL_3938 == 1'h0;
  assign _EVAL_3031 = _EVAL_2723 ? _EVAL_4413 : _EVAL_782;
  assign _EVAL_5015 = _EVAL_2647 ? _EVAL_1494 : _EVAL_3031;
  assign _EVAL_696 = _EVAL_1941 & _EVAL_5015;
  assign _EVAL_2151 = {{31'd0}, _EVAL_696};
  assign _EVAL_1119 = _EVAL_5117 | _EVAL_2151;
  assign _EVAL_4585 = _EVAL_1119 | _EVAL_665;
  assign _EVAL_718 = _EVAL_4162 == 3'h5;
  assign _EVAL_676 = _EVAL_5412[31];
  assign _EVAL_681 = _EVAL_2282 & _EVAL_676;
  assign _EVAL_4668 = {_EVAL_681,_EVAL_5412};
  assign _EVAL_3186 = _EVAL_5412[31:16];
  assign _EVAL_4612 = {{16'd0}, _EVAL_3186};
  assign _EVAL_4211 = _EVAL_5412[15:0];
  assign _EVAL_2796 = {_EVAL_4211, 16'h0};
  assign _EVAL_744 = _EVAL_2796 & 32'hffff0000;
  assign _EVAL_4586 = _EVAL_4612 | _EVAL_744;
  assign _EVAL_562 = _EVAL_4586[31:8];
  assign _EVAL_4017 = {{8'd0}, _EVAL_562};
  assign _EVAL_4763 = _EVAL_4017 & 32'hff00ff;
  assign _EVAL_4861 = _EVAL_4586[23:0];
  assign _EVAL_1078 = {_EVAL_4861, 8'h0};
  assign _EVAL_2142 = _EVAL_1078 & 32'hff00ff00;
  assign _EVAL_1633 = _EVAL_4763 | _EVAL_2142;
  assign _EVAL_3905 = _EVAL_1633[31:4];
  assign _EVAL_1745 = {{4'd0}, _EVAL_3905};
  assign _EVAL_656 = _EVAL_1745 & 32'hf0f0f0f;
  assign _EVAL_1657 = _EVAL_1633[27:0];
  assign _EVAL_5333 = {_EVAL_1657, 4'h0};
  assign _EVAL_1898 = _EVAL_5333 & 32'hf0f0f0f0;
  assign _EVAL_3521 = _EVAL_656 | _EVAL_1898;
  assign _EVAL_1550 = _EVAL_3521[31:2];
  assign _EVAL_5038 = {{2'd0}, _EVAL_1550};
  assign _EVAL_1365 = _EVAL_5038 & 32'h33333333;
  assign _EVAL_3967 = _EVAL_3521[29:0];
  assign _EVAL_688 = {_EVAL_3967, 2'h0};
  assign _EVAL_4853 = _EVAL_688 & 32'hcccccccc;
  assign _EVAL_3446 = _EVAL_1365 | _EVAL_4853;
  assign _EVAL_1848 = _EVAL_3446[31:1];
  assign _EVAL_1197 = {{1'd0}, _EVAL_1848};
  assign _EVAL_2896 = _EVAL_1197 & 32'h55555555;
  assign _EVAL_3998 = _EVAL_3446[30:0];
  assign _EVAL_3251 = {_EVAL_3998, 1'h0};
  assign _EVAL_4408 = _EVAL_3251 & 32'haaaaaaaa;
  assign _EVAL_3547 = _EVAL_2896 | _EVAL_4408;
  assign _EVAL_3866 = _EVAL_2859 ? _EVAL_4668 : {{1'd0}, _EVAL_3547};
  assign _EVAL_303 = $signed(_EVAL_3866);
  assign _EVAL_3683 = _EVAL_1155[4:0];
  assign _EVAL_2894 = $signed(_EVAL_303) >>> _EVAL_3683;
  assign _EVAL_1866 = _EVAL_2894[31:0];
  assign _EVAL_5215 = _EVAL_718 ? _EVAL_1866 : 32'h0;
  assign _EVAL_1944 = _EVAL_4162 == 3'h1;
  assign _EVAL_5328 = _EVAL_1866[31:16];
  assign _EVAL_2264 = {{16'd0}, _EVAL_5328};
  assign _EVAL_3615 = _EVAL_1866[15:0];
  assign _EVAL_5124 = {_EVAL_3615, 16'h0};
  assign _EVAL_3601 = _EVAL_5124 & 32'hffff0000;
  assign _EVAL_4371 = _EVAL_2264 | _EVAL_3601;
  assign _EVAL_2516 = _EVAL_4371[31:8];
  assign _EVAL_4412 = {{8'd0}, _EVAL_2516};
  assign _EVAL_1331 = _EVAL_4412 & 32'hff00ff;
  assign _EVAL_2520 = _EVAL_4371[23:0];
  assign _EVAL_5336 = {_EVAL_2520, 8'h0};
  assign _EVAL_668 = _EVAL_5336 & 32'hff00ff00;
  assign _EVAL_3182 = _EVAL_1331 | _EVAL_668;
  assign _EVAL_5231 = _EVAL_3182[31:4];
  assign _EVAL_4958 = {{4'd0}, _EVAL_5231};
  assign _EVAL_3572 = _EVAL_4958 & 32'hf0f0f0f;
  assign _EVAL_642 = _EVAL_3182[27:0];
  assign _EVAL_1312 = {_EVAL_642, 4'h0};
  assign _EVAL_5033 = _EVAL_1312 & 32'hf0f0f0f0;
  assign _EVAL_3337 = _EVAL_3572 | _EVAL_5033;
  assign _EVAL_3564 = _EVAL_3337[31:2];
  assign _EVAL_4616 = {{2'd0}, _EVAL_3564};
  assign _EVAL_3833 = _EVAL_4616 & 32'h33333333;
  assign _EVAL_3189 = _EVAL_3337[29:0];
  assign _EVAL_658 = {_EVAL_3189, 2'h0};
  assign _EVAL_2663 = _EVAL_658 & 32'hcccccccc;
  assign _EVAL_4342 = _EVAL_3833 | _EVAL_2663;
  assign _EVAL_2984 = _EVAL_4342[31:1];
  assign _EVAL_3397 = {{1'd0}, _EVAL_2984};
  assign _EVAL_553 = _EVAL_3397 & 32'h55555555;
  assign _EVAL_2392 = _EVAL_4342[30:0];
  assign _EVAL_1265 = {_EVAL_2392, 1'h0};
  assign _EVAL_3891 = _EVAL_1265 & 32'haaaaaaaa;
  assign _EVAL_3749 = _EVAL_553 | _EVAL_3891;
  assign _EVAL_572 = _EVAL_1944 ? _EVAL_3749 : 32'h0;
  assign _EVAL_3726 = _EVAL_5215 | _EVAL_572;
  assign _EVAL_1495 = _EVAL_4585 | _EVAL_3726;
  assign _EVAL_2845 = _EVAL_1446 ? _EVAL_110 : _EVAL_1495;
  assign _EVAL_4399 = _EVAL_2869 ? _EVAL_234 : _EVAL_2845;
  assign _EVAL_924 = _EVAL_2219 & _EVAL_3498;
  assign _EVAL_1891 = _EVAL_3227 & _EVAL_924;
  assign _EVAL_3378 = _EVAL_4064 == 3'h0;
  assign _EVAL_4870 = {_EVAL_4659,_EVAL_2683,1'h1};
  assign _EVAL_1715 = {_EVAL_3977,_EVAL_1818};
  assign _EVAL_943 = _EVAL_4870 + _EVAL_1715;
  assign _EVAL_4330 = _EVAL_943[32:1];
  assign _EVAL_363 = _EVAL_3378 ? _EVAL_4330 : 32'h0;
  assign _EVAL_1784 = _EVAL_4064[2:1];
  assign _EVAL_986 = _EVAL_1784 == 2'h1;
  assign _EVAL_4946 = _EVAL_1102 ^ _EVAL_4572;
  assign _EVAL_3729 = _EVAL_4330[31];
  assign _EVAL_3756 = _EVAL_4946 ? _EVAL_3729 : _EVAL_354;
  assign _EVAL_1841 = _EVAL_986 & _EVAL_3756;
  assign _EVAL_2947 = {{31'd0}, _EVAL_1841};
  assign _EVAL_1489 = _EVAL_363 | _EVAL_2947;
  assign _EVAL_4717 = _EVAL_557 == 1'h0;
  assign _EVAL_4651 = _EVAL_358 & _EVAL_4717;
  assign _EVAL_2950 = _EVAL_1483 ^ _EVAL_3977;
  assign _EVAL_3447 = _EVAL_4651 ? _EVAL_2950 : 32'h0;
  assign _EVAL_1662 = _EVAL_4064 >= 3'h6;
  assign _EVAL_1791 = _EVAL_1483 & _EVAL_3977;
  assign _EVAL_2179 = _EVAL_1662 ? _EVAL_1791 : 32'h0;
  assign _EVAL_1833 = _EVAL_3447 | _EVAL_2179;
  assign _EVAL_2769 = _EVAL_1489 | _EVAL_1833;
  assign _EVAL_4694 = _EVAL_4064 == 3'h5;
  assign _EVAL_3487 = _EVAL_4694 ? _EVAL_1505 : 32'h0;
  assign _EVAL_698 = _EVAL_4064 == 3'h1;
  assign _EVAL_1720 = {{16'd0}, _EVAL_3885};
  assign _EVAL_571 = _EVAL_1505[15:0];
  assign _EVAL_3136 = {_EVAL_571, 16'h0};
  assign _EVAL_1295 = _EVAL_3136 & 32'hffff0000;
  assign _EVAL_484 = _EVAL_1720 | _EVAL_1295;
  assign _EVAL_2418 = _EVAL_484[31:8];
  assign _EVAL_5119 = {{8'd0}, _EVAL_2418};
  assign _EVAL_2713 = _EVAL_5119 & 32'hff00ff;
  assign _EVAL_1663 = _EVAL_484[23:0];
  assign _EVAL_4777 = {_EVAL_1663, 8'h0};
  assign _EVAL_4784 = _EVAL_4777 & 32'hff00ff00;
  assign _EVAL_385 = _EVAL_2713 | _EVAL_4784;
  assign _EVAL_638 = _EVAL_385[31:4];
  assign _EVAL_4331 = {{4'd0}, _EVAL_638};
  assign _EVAL_3206 = _EVAL_4331 & 32'hf0f0f0f;
  assign _EVAL_1554 = _EVAL_385[27:0];
  assign _EVAL_4315 = {_EVAL_1554, 4'h0};
  assign _EVAL_4529 = _EVAL_4315 & 32'hf0f0f0f0;
  assign _EVAL_2837 = _EVAL_3206 | _EVAL_4529;
  assign _EVAL_4868 = _EVAL_2837[31:2];
  assign _EVAL_2433 = {{2'd0}, _EVAL_4868};
  assign _EVAL_3773 = _EVAL_2433 & 32'h33333333;
  assign _EVAL_1058 = _EVAL_2837[29:0];
  assign _EVAL_825 = {_EVAL_1058, 2'h0};
  assign _EVAL_5005 = _EVAL_825 & 32'hcccccccc;
  assign _EVAL_3179 = _EVAL_3773 | _EVAL_5005;
  assign _EVAL_4922 = _EVAL_3179[31:1];
  assign _EVAL_4434 = {{1'd0}, _EVAL_4922};
  assign _EVAL_5028 = _EVAL_4434 & 32'h55555555;
  assign _EVAL_2755 = _EVAL_3179[30:0];
  assign _EVAL_4076 = {_EVAL_2755, 1'h0};
  assign _EVAL_3437 = _EVAL_4076 & 32'haaaaaaaa;
  assign _EVAL_2240 = _EVAL_5028 | _EVAL_3437;
  assign _EVAL_4258 = _EVAL_698 ? _EVAL_2240 : 32'h0;
  assign _EVAL_3595 = _EVAL_3487 | _EVAL_4258;
  assign _EVAL_3125 = _EVAL_2769 | _EVAL_3595;
  assign _EVAL_942 = _EVAL_3568 ? m__EVAL_2 : _EVAL_3125;
  assign _EVAL_3923 = _EVAL_854 ? csr__EVAL_84 : _EVAL_942;
  assign _EVAL_2039 = _EVAL_5099 == _EVAL_1059;
  assign _EVAL_932 = _EVAL_332 & _EVAL_2039;
  assign _EVAL_1961 = _EVAL_4774 & _EVAL_932;
  assign _EVAL_5350 = _EVAL_2812 == _EVAL_1059;
  assign _EVAL_5092 = _EVAL_5386 & _EVAL_5350;
  assign _EVAL_4599 = _EVAL_5252 & _EVAL_5092;
  assign _EVAL_3185 = _EVAL_4599 ? _EVAL_3187 : _EVAL_4679;
  assign _EVAL_1044 = _EVAL_1961 ? _EVAL_4863 : _EVAL_3185;
  assign _EVAL_2877 = _EVAL_1891 ? _EVAL_3923 : _EVAL_1044;
  assign _EVAL_3262 = _EVAL_5183 ? _EVAL_4399 : _EVAL_2877;
  assign _EVAL_2199 = _EVAL_1533 ? _EVAL_3262 : _EVAL_4679;
  assign _EVAL_2004 = _EVAL_4000 & _EVAL_3295;
  assign _EVAL_5323 = csr__EVAL_80[31:8];
  assign _EVAL_1803 = _EVAL_5323[0];
  assign _EVAL_450 = _EVAL_3624 & _EVAL_2145;
  assign _EVAL_3790 = _EVAL_4530[1:0];
  assign _EVAL_4114 = _EVAL_3790 == 2'h0;
  assign _EVAL_660 = _EVAL_2145 & _EVAL_4114;
  assign _EVAL_4426 = _EVAL_660 & _EVAL_3176;
  assign _EVAL_2871 = _EVAL_4426 == 1'h0;
  assign _EVAL_5263 = _EVAL_450 & _EVAL_2871;
  assign _EVAL_4235 = _EVAL_5263 == 1'h0;
  assign _EVAL_1549 = _EVAL_3105 & _EVAL_4235;
  assign _EVAL_2689 = _EVAL_4832[4];
  assign _EVAL_3811 = _EVAL_2689 == 1'h0;
  assign _EVAL_2829 = _EVAL_4832[2];
  assign _EVAL_4988 = _EVAL_3811 & _EVAL_2829;
  assign _EVAL_4661 = _EVAL_5283 == 1'h0;
  assign _EVAL_5409 = _EVAL_6[2];
  assign _EVAL_4117 = _EVAL_4661 & _EVAL_5409;
  assign _EVAL_4325 = _EVAL_6[3];
  assign _EVAL_3207 = _EVAL_4117 & _EVAL_4325;
  assign _EVAL_357 = _EVAL_6[0];
  assign _EVAL_2115 = _EVAL_357 == 1'h0;
  assign _EVAL_576 = _EVAL_3207 & _EVAL_2115;
  assign _EVAL_3349 = _EVAL_73[0];
  assign _EVAL_3807 = _EVAL_576 & _EVAL_3349;
  assign _EVAL_2616 = _EVAL_84[2];
  assign _EVAL_2438 = _EVAL_2616 == 1'h0;
  assign _EVAL_905 = _EVAL_3807 & _EVAL_2438;
  assign _EVAL_1821 = _EVAL_191[4];
  assign _EVAL_5419 = _EVAL_1821 == 1'h0;
  assign _EVAL_2850 = _EVAL_191[2];
  assign _EVAL_703 = _EVAL_5419 & _EVAL_2850;
  assign _EVAL_5417 = _EVAL_191[3];
  assign _EVAL_4023 = _EVAL_703 & _EVAL_5417;
  assign _EVAL_4078 = _EVAL_191[0];
  assign _EVAL_4209 = _EVAL_4078 == 1'h0;
  assign _EVAL_1061 = _EVAL_4023 & _EVAL_4209;
  assign _EVAL_3190 = _EVAL_121[0];
  assign _EVAL_3644 = _EVAL_1061 & _EVAL_3190;
  assign _EVAL_2233 = _EVAL_2964 == 1'h0;
  assign _EVAL_2403 = _EVAL_3644 & _EVAL_2233;
  assign _EVAL_2013 = _EVAL_315 ? _EVAL_905 : _EVAL_2403;
  assign _EVAL_5208 = _EVAL_4988 & _EVAL_3255;
  assign _EVAL_4141 = _EVAL_4832[0];
  assign _EVAL_5201 = _EVAL_4141 == 1'h0;
  assign _EVAL_1196 = _EVAL_5208 & _EVAL_5201;
  assign _EVAL_4449 = _EVAL_1196 & _EVAL_1762;
  assign _EVAL_5022 = _EVAL_315 ? _EVAL_84 : _EVAL_153;
  assign _EVAL_5107 = _EVAL_5022[2];
  assign _EVAL_2545 = _EVAL_4449 & _EVAL_5107;
  assign _EVAL_4826 = _EVAL_2013 | _EVAL_2545;
  assign _EVAL_1243 = _EVAL_4826 == 1'h0;
  assign _EVAL_3533 = _EVAL_4988 & _EVAL_1243;
  assign _EVAL_1267 = _EVAL_1549 | _EVAL_3533;
  assign _EVAL_2079 = _EVAL_205 == 1'h0;
  assign _EVAL_1273 = _EVAL_1379[1];
  assign _EVAL_3113 = _EVAL_1273 | _EVAL_4818;
  assign _EVAL_1490 = {_EVAL_3113,_EVAL_4322};
  assign _EVAL_2200 = $signed(_EVAL_1490);
  assign _EVAL_1165 = _EVAL_3880[31];
  assign _EVAL_2226 = _EVAL_1273 | _EVAL_1165;
  assign _EVAL_2174 = {_EVAL_2226,_EVAL_3880};
  assign _EVAL_5327 = $signed(_EVAL_2174);
  assign _EVAL_3979 = $signed(_EVAL_2200) < $signed(_EVAL_5327);
  assign _EVAL_3682 = _EVAL_3039[1:0];
  assign _EVAL_1330 = _EVAL_3682 == 2'h0;
  assign _EVAL_910 = _EVAL_946 & _EVAL_1330;
  assign _EVAL_4056 = _EVAL_910 & _EVAL_3588;
  assign _EVAL_838 = _EVAL_4240 & _EVAL_4056;
  assign _EVAL_3452 = _EVAL_3240 & _EVAL_2118;
  assign _EVAL_3658 = _EVAL_838 & _EVAL_3452;
  assign _EVAL_2270 = _EVAL_3658 ? _EVAL_1379 : 3'h2;
  assign _EVAL_664 = _EVAL_2270[0];
  assign _EVAL_2457 = _EVAL_2270[2];
  assign _EVAL_4680 = _EVAL_664 ^ _EVAL_2457;
  assign _EVAL_2434 = _EVAL_4322 == _EVAL_3880;
  assign _EVAL_1864 = _EVAL_2457 == 1'h0;
  assign _EVAL_2076 = _EVAL_2270[1];
  assign _EVAL_4170 = _EVAL_2076 == 1'h0;
  assign _EVAL_2480 = _EVAL_1864 & _EVAL_4170;
  assign _EVAL_1448 = _EVAL_664 ^ _EVAL_2480;
  assign _EVAL_5113 = _EVAL_2434 ? _EVAL_1448 : _EVAL_664;
  assign _EVAL_430 = _EVAL_3979 ? _EVAL_4680 : _EVAL_5113;
  assign _EVAL_4129 = _EVAL_430 ? 1'h0 : _EVAL_2118;
  assign _EVAL_815 = _EVAL_2579 == _EVAL_274;
  assign _EVAL_4069 = _EVAL_653 & _EVAL_815;
  assign _EVAL_3753 = _EVAL_4129 & _EVAL_4069;
  assign _EVAL_4789 = _EVAL_3117 == _EVAL_274;
  assign _EVAL_1887 = _EVAL_4043 & _EVAL_4789;
  assign _EVAL_3853 = _EVAL_2326 & _EVAL_1887;
  assign _EVAL_1430 = _EVAL_3670 == _EVAL_274;
  assign _EVAL_2649 = _EVAL_1724 & _EVAL_1430;
  assign _EVAL_581 = _EVAL_3624 & _EVAL_2649;
  assign _EVAL_1221 = _EVAL_581 ? _EVAL_3176 : 1'h1;
  assign _EVAL_4410 = _EVAL_3853 ? _EVAL_922 : _EVAL_1221;
  assign _EVAL_5354 = _EVAL_3231 ? _EVAL_3588 : _EVAL_4410;
  assign _EVAL_3689 = _EVAL_3753 ? _EVAL_1122 : _EVAL_5354;
  assign _EVAL_1543 = _EVAL_3227 & _EVAL_3085;
  assign _EVAL_3847 = _EVAL_3227 & _EVAL_1963;
  assign _EVAL_2635 = _EVAL_1543 & _EVAL_3847;
  assign _EVAL_4279 = _EVAL_2635 == 1'h0;
  assign _EVAL_2335 = _EVAL_3689 & _EVAL_4279;
  assign _EVAL_917 = _EVAL_2079 | _EVAL_2335;
  assign _EVAL_1726 = _EVAL_250 == 1'h0;
  assign _EVAL_4840 = _EVAL_2579 == _EVAL_180;
  assign _EVAL_2148 = _EVAL_653 & _EVAL_4840;
  assign _EVAL_4874 = _EVAL_4129 & _EVAL_2148;
  assign _EVAL_4846 = _EVAL_4135 == _EVAL_180;
  assign _EVAL_4159 = _EVAL_4692 & _EVAL_4846;
  assign _EVAL_2228 = _EVAL_4240 & _EVAL_4159;
  assign _EVAL_1530 = _EVAL_3117 == _EVAL_180;
  assign _EVAL_2844 = _EVAL_4043 & _EVAL_1530;
  assign _EVAL_1177 = _EVAL_2326 & _EVAL_2844;
  assign _EVAL_2773 = _EVAL_3670 == _EVAL_180;
  assign _EVAL_1515 = _EVAL_1724 & _EVAL_2773;
  assign _EVAL_853 = _EVAL_3624 & _EVAL_1515;
  assign _EVAL_5101 = _EVAL_853 ? _EVAL_3176 : 1'h1;
  assign _EVAL_4766 = _EVAL_1177 ? _EVAL_922 : _EVAL_5101;
  assign _EVAL_1388 = _EVAL_2228 ? _EVAL_3588 : _EVAL_4766;
  assign _EVAL_1718 = _EVAL_4874 ? _EVAL_1122 : _EVAL_1388;
  assign _EVAL_2341 = _EVAL_1543 & _EVAL_5055;
  assign _EVAL_1620 = _EVAL_2341 == 1'h0;
  assign _EVAL_3626 = _EVAL_1718 & _EVAL_1620;
  assign _EVAL_964 = _EVAL_1726 | _EVAL_3626;
  assign _EVAL_801 = _EVAL_917 & _EVAL_964;
  assign _EVAL_5141 = _EVAL_1 == 1'h0;
  assign _EVAL_4499 = _EVAL_2579 == _EVAL_154;
  assign _EVAL_1767 = _EVAL_653 & _EVAL_4499;
  assign _EVAL_2827 = _EVAL_4129 & _EVAL_1767;
  assign _EVAL_1183 = _EVAL_3117 == _EVAL_154;
  assign _EVAL_992 = _EVAL_4043 & _EVAL_1183;
  assign _EVAL_4654 = _EVAL_2326 & _EVAL_992;
  assign _EVAL_442 = _EVAL_3670 == _EVAL_154;
  assign _EVAL_875 = _EVAL_1724 & _EVAL_442;
  assign _EVAL_1858 = _EVAL_3624 & _EVAL_875;
  assign _EVAL_3408 = _EVAL_1858 ? _EVAL_3176 : 1'h1;
  assign _EVAL_4485 = _EVAL_4654 ? _EVAL_922 : _EVAL_3408;
  assign _EVAL_1315 = _EVAL_589 ? _EVAL_3588 : _EVAL_4485;
  assign _EVAL_1877 = _EVAL_2827 ? _EVAL_1122 : _EVAL_1315;
  assign _EVAL_5063 = _EVAL_3742 == _EVAL_154;
  assign _EVAL_1888 = _EVAL_2219 & _EVAL_5063;
  assign _EVAL_3527 = _EVAL_3227 & _EVAL_1888;
  assign _EVAL_467 = _EVAL_1543 & _EVAL_3527;
  assign _EVAL_5204 = _EVAL_467 == 1'h0;
  assign _EVAL_2007 = _EVAL_1877 & _EVAL_5204;
  assign _EVAL_2279 = _EVAL_5141 | _EVAL_2007;
  assign _EVAL_370 = _EVAL_141 == 1'h0;
  assign _EVAL_5347 = _EVAL_2579 == _EVAL_68;
  assign _EVAL_1594 = _EVAL_653 & _EVAL_5347;
  assign _EVAL_2986 = _EVAL_4129 & _EVAL_1594;
  assign _EVAL_4184 = _EVAL_4135 == _EVAL_68;
  assign _EVAL_3464 = _EVAL_4692 & _EVAL_4184;
  assign _EVAL_2468 = _EVAL_4240 & _EVAL_3464;
  assign _EVAL_4276 = _EVAL_3117 == _EVAL_68;
  assign _EVAL_2639 = _EVAL_4043 & _EVAL_4276;
  assign _EVAL_1693 = _EVAL_2326 & _EVAL_2639;
  assign _EVAL_1073 = _EVAL_3670 == _EVAL_68;
  assign _EVAL_4557 = _EVAL_1724 & _EVAL_1073;
  assign _EVAL_1440 = _EVAL_3624 & _EVAL_4557;
  assign _EVAL_503 = _EVAL_1440 ? _EVAL_3176 : 1'h1;
  assign _EVAL_438 = _EVAL_1693 ? _EVAL_922 : _EVAL_503;
  assign _EVAL_1229 = _EVAL_2468 ? _EVAL_3588 : _EVAL_438;
  assign _EVAL_2889 = _EVAL_2986 ? _EVAL_1122 : _EVAL_1229;
  assign _EVAL_4317 = _EVAL_3742 == _EVAL_68;
  assign _EVAL_1301 = _EVAL_2219 & _EVAL_4317;
  assign _EVAL_1993 = _EVAL_3227 & _EVAL_1301;
  assign _EVAL_1682 = _EVAL_1543 & _EVAL_1993;
  assign _EVAL_2618 = _EVAL_1682 == 1'h0;
  assign _EVAL_5103 = _EVAL_2889 & _EVAL_2618;
  assign _EVAL_699 = _EVAL_370 | _EVAL_5103;
  assign _EVAL_1980 = _EVAL_2279 & _EVAL_699;
  assign _EVAL_2482 = _EVAL_315 ? _EVAL_801 : _EVAL_1980;
  assign _EVAL_3139 = _EVAL_1267 & _EVAL_2482;
  assign _EVAL_3799 = _EVAL_725 | _EVAL_3139;
  assign _EVAL_3514 = _EVAL_315 ? _EVAL_3753 : _EVAL_2827;
  assign _EVAL_770 = _EVAL_313 == 3'h0;
  assign _EVAL_1839 = {_EVAL_929,_EVAL_3366,1'h1};
  assign _EVAL_3792 = _EVAL_5237 ? _EVAL_5102 : _EVAL_1560;
  assign _EVAL_1987 = {_EVAL_3792,_EVAL_5237};
  assign _EVAL_5199 = _EVAL_1839 + _EVAL_1987;
  assign _EVAL_3860 = _EVAL_5199[32:1];
  assign _EVAL_2830 = _EVAL_770 ? _EVAL_3860 : 32'h0;
  assign _EVAL_2211 = _EVAL_313[2:1];
  assign _EVAL_2432 = _EVAL_2211 == 2'h1;
  assign _EVAL_4366 = _EVAL_2983[31];
  assign _EVAL_3478 = _EVAL_3792[31];
  assign _EVAL_592 = _EVAL_4366 ^ _EVAL_3478;
  assign _EVAL_1986 = _EVAL_3860[31];
  assign _EVAL_491 = _EVAL_313[0];
  assign _EVAL_2010 = _EVAL_3478 == 1'h0;
  assign _EVAL_1092 = _EVAL_491 ? _EVAL_2010 : _EVAL_4366;
  assign _EVAL_3640 = _EVAL_592 ? _EVAL_1986 : _EVAL_1092;
  assign _EVAL_3058 = _EVAL_2432 & _EVAL_3640;
  assign _EVAL_3929 = {{31'd0}, _EVAL_3058};
  assign _EVAL_5137 = _EVAL_2830 | _EVAL_3929;
  assign _EVAL_3664 = _EVAL_491 == 1'h0;
  assign _EVAL_2610 = _EVAL_2538 & _EVAL_3664;
  assign _EVAL_4268 = _EVAL_2983 ^ _EVAL_3792;
  assign _EVAL_2988 = _EVAL_2610 ? _EVAL_4268 : 32'h0;
  assign _EVAL_1673 = _EVAL_313 >= 3'h6;
  assign _EVAL_2248 = _EVAL_2983 & _EVAL_3792;
  assign _EVAL_4739 = _EVAL_1673 ? _EVAL_2248 : 32'h0;
  assign _EVAL_1343 = _EVAL_2988 | _EVAL_4739;
  assign _EVAL_1739 = _EVAL_5137 | _EVAL_1343;
  assign _EVAL_1666 = _EVAL_313 == 3'h5;
  assign _EVAL_3468 = _EVAL_1666 ? _EVAL_1735 : 32'h0;
  assign _EVAL_4134 = _EVAL_313 == 3'h1;
  assign _EVAL_3916 = _EVAL_2336[31:2];
  assign _EVAL_2473 = {{2'd0}, _EVAL_3916};
  assign _EVAL_1217 = _EVAL_2473 & 32'h33333333;
  assign _EVAL_720 = _EVAL_1217 | _EVAL_3622;
  assign _EVAL_5080 = _EVAL_720[31:1];
  assign _EVAL_4323 = {{1'd0}, _EVAL_5080};
  assign _EVAL_3410 = _EVAL_4323 & 32'h55555555;
  assign _EVAL_2792 = _EVAL_720[30:0];
  assign _EVAL_2702 = {_EVAL_2792, 1'h0};
  assign _EVAL_381 = _EVAL_2702 & 32'haaaaaaaa;
  assign _EVAL_3411 = _EVAL_3410 | _EVAL_381;
  assign _EVAL_1512 = _EVAL_4134 ? _EVAL_3411 : 32'h0;
  assign _EVAL_5361 = _EVAL_3468 | _EVAL_1512;
  assign _EVAL_1572 = _EVAL_1739 | _EVAL_5361;
  assign _EVAL_2073 = _EVAL_315 ? _EVAL_3853 : _EVAL_4654;
  assign _EVAL_4207 = _EVAL_315 ? _EVAL_581 : _EVAL_1858;
  assign _EVAL_436 = _EVAL_4706 == _EVAL_274;
  assign _EVAL_1205 = _EVAL_1333 & _EVAL_436;
  assign _EVAL_4824 = _EVAL_2506 & _EVAL_1205;
  assign _EVAL_820 = _EVAL_4706 == _EVAL_154;
  assign _EVAL_5189 = _EVAL_1333 & _EVAL_820;
  assign _EVAL_2478 = _EVAL_2506 & _EVAL_5189;
  assign _EVAL_391 = _EVAL_315 ? _EVAL_4824 : _EVAL_2478;
  assign _EVAL_1129 = _EVAL_315 ? _EVAL_3847 : _EVAL_3527;
  assign _EVAL_4097 = _EVAL_5099 == _EVAL_274;
  assign _EVAL_2971 = _EVAL_332 & _EVAL_4097;
  assign _EVAL_1485 = _EVAL_4774 & _EVAL_2971;
  assign _EVAL_4810 = _EVAL_5099 == _EVAL_154;
  assign _EVAL_3801 = _EVAL_332 & _EVAL_4810;
  assign _EVAL_4977 = _EVAL_4774 & _EVAL_3801;
  assign _EVAL_4046 = _EVAL_315 ? _EVAL_1485 : _EVAL_4977;
  assign _EVAL_2464 = _EVAL_315 ? _EVAL_1228 : _EVAL_3364;
  assign _EVAL_1853 = _EVAL_708__EVAL_709_data;
  assign _EVAL_5376 = _EVAL_708__EVAL_711_data;
  assign _EVAL_5310 = _EVAL_315 ? _EVAL_1853 : _EVAL_5376;
  assign _EVAL_568 = _EVAL_2464 ? _EVAL_3187 : _EVAL_5310;
  assign _EVAL_4878 = _EVAL_4046 ? _EVAL_4863 : _EVAL_568;
  assign _EVAL_1457 = _EVAL_1129 ? _EVAL_3923 : _EVAL_4878;
  assign _EVAL_1974 = _EVAL_391 ? _EVAL_4399 : _EVAL_1457;
  assign _EVAL_1288 = _EVAL_4207 ? _EVAL_2919 : _EVAL_1974;
  assign _EVAL_1257 = _EVAL_2073 ? _EVAL_4679 : _EVAL_1288;
  assign _EVAL_886 = _EVAL_2668 ? _EVAL_1932 : _EVAL_1257;
  assign _EVAL_1431 = _EVAL_3514 ? _EVAL_1572 : _EVAL_886;
  assign _EVAL_3135 = _EVAL_1764 == 2'h1;
  assign _EVAL_4405 = _EVAL_1699 & _EVAL_3135;
  assign _EVAL_4292 = _EVAL_315 ? _EVAL_268 : _EVAL_214;
  assign _EVAL_3083 = _EVAL_315 ? _EVAL_58 : _EVAL_16;
  assign _EVAL_3426 = _EVAL_4292 | _EVAL_3083;
  assign _EVAL_5075 = _EVAL_2326 & _EVAL_3431;
  assign _EVAL_3723 = _EVAL_4803 & _EVAL_5075;
  assign _EVAL_2652 = _EVAL_2506 & _EVAL_4643;
  assign _EVAL_3581 = _EVAL_3723 & _EVAL_2652;
  assign _EVAL_4571 = _EVAL_3426 & _EVAL_3581;
  assign _EVAL_3870 = _EVAL_4571 & _EVAL_4360;
  assign _EVAL_4978 = _EVAL_405 | _EVAL_1588;
  assign _EVAL_2963 = _EVAL_55 & _EVAL_626;
  assign _EVAL_3028 = fpu__EVAL_10 > 3'h2;
  assign _EVAL_1020 = fpu__EVAL_20 & fpu__EVAL_16;
  assign _EVAL_2784 = fpu__EVAL_35;
  assign _EVAL_1114 = _EVAL_274 == _EVAL_2784;
  assign _EVAL_2414 = _EVAL_39 & _EVAL_1114;
  assign _EVAL_445 = _EVAL_180 == _EVAL_2784;
  assign _EVAL_3336 = _EVAL_188 & _EVAL_445;
  assign _EVAL_4554 = _EVAL_2414 | _EVAL_3336;
  assign _EVAL_1937 = _EVAL_3212 == _EVAL_2784;
  assign _EVAL_2598 = _EVAL_260 & _EVAL_1937;
  assign _EVAL_5317 = _EVAL_4554 | _EVAL_2598;
  assign _EVAL_765 = _EVAL_1020 & _EVAL_5317;
  assign _EVAL_3837 = _EVAL_154 == _EVAL_2784;
  assign _EVAL_1975 = _EVAL_148 & _EVAL_3837;
  assign _EVAL_5177 = _EVAL_68 == _EVAL_2784;
  assign _EVAL_2824 = _EVAL_179 & _EVAL_5177;
  assign _EVAL_1094 = _EVAL_1975 | _EVAL_2824;
  assign _EVAL_3442 = _EVAL_4127 == _EVAL_2784;
  assign _EVAL_1029 = _EVAL_119 & _EVAL_3442;
  assign _EVAL_5053 = _EVAL_1094 | _EVAL_1029;
  assign _EVAL_1089 = _EVAL_1020 & _EVAL_5053;
  assign _EVAL_2367 = _EVAL_315 ? _EVAL_765 : _EVAL_1089;
  assign _EVAL_3199 = _EVAL_3028 & _EVAL_2367;
  assign _EVAL_1406 = fpu__EVAL_39 > 3'h2;
  assign _EVAL_2273 = fpu__EVAL_22 & fpu__EVAL_56;
  assign _EVAL_4009 = fpu__EVAL_26;
  assign _EVAL_2276 = _EVAL_274 == _EVAL_4009;
  assign _EVAL_1873 = _EVAL_39 & _EVAL_2276;
  assign _EVAL_4438 = _EVAL_180 == _EVAL_4009;
  assign _EVAL_4502 = _EVAL_188 & _EVAL_4438;
  assign _EVAL_3612 = _EVAL_1873 | _EVAL_4502;
  assign _EVAL_3945 = _EVAL_3212 == _EVAL_4009;
  assign _EVAL_2993 = _EVAL_260 & _EVAL_3945;
  assign _EVAL_786 = _EVAL_3612 | _EVAL_2993;
  assign _EVAL_4293 = _EVAL_2273 & _EVAL_786;
  assign _EVAL_812 = _EVAL_154 == _EVAL_4009;
  assign _EVAL_2078 = _EVAL_148 & _EVAL_812;
  assign _EVAL_4012 = _EVAL_68 == _EVAL_4009;
  assign _EVAL_2334 = _EVAL_179 & _EVAL_4012;
  assign _EVAL_4990 = _EVAL_2078 | _EVAL_2334;
  assign _EVAL_3084 = _EVAL_4127 == _EVAL_4009;
  assign _EVAL_4511 = _EVAL_119 & _EVAL_3084;
  assign _EVAL_4681 = _EVAL_4990 | _EVAL_4511;
  assign _EVAL_4058 = _EVAL_2273 & _EVAL_4681;
  assign _EVAL_4263 = _EVAL_315 ? _EVAL_4293 : _EVAL_4058;
  assign _EVAL_4579 = _EVAL_1406 & _EVAL_4263;
  assign _EVAL_479 = _EVAL_3199 | _EVAL_4579;
  assign _EVAL_2672 = fpu__EVAL_34 > 3'h2;
  assign _EVAL_1892 = _EVAL_315 ? _EVAL_2025 : _EVAL_4623;
  assign _EVAL_4835 = _EVAL_2672 & _EVAL_1892;
  assign _EVAL_3698 = _EVAL_479 | _EVAL_4835;
  assign _EVAL_2411 = fpu__EVAL_51 > 3'h2;
  assign _EVAL_1686 = fpu__EVAL_48 & fpu__EVAL_42;
  assign _EVAL_521 = fpu__EVAL_25;
  assign _EVAL_4006 = _EVAL_274 == _EVAL_521;
  assign _EVAL_1872 = _EVAL_39 & _EVAL_4006;
  assign _EVAL_4775 = _EVAL_180 == _EVAL_521;
  assign _EVAL_745 = _EVAL_188 & _EVAL_4775;
  assign _EVAL_2385 = _EVAL_1872 | _EVAL_745;
  assign _EVAL_1945 = _EVAL_3212 == _EVAL_521;
  assign _EVAL_987 = _EVAL_260 & _EVAL_1945;
  assign _EVAL_5421 = _EVAL_2385 | _EVAL_987;
  assign _EVAL_1314 = _EVAL_1686 & _EVAL_5421;
  assign _EVAL_2293 = _EVAL_154 == _EVAL_521;
  assign _EVAL_1211 = _EVAL_148 & _EVAL_2293;
  assign _EVAL_3562 = _EVAL_68 == _EVAL_521;
  assign _EVAL_682 = _EVAL_179 & _EVAL_3562;
  assign _EVAL_1586 = _EVAL_1211 | _EVAL_682;
  assign _EVAL_4029 = _EVAL_4127 == _EVAL_521;
  assign _EVAL_4013 = _EVAL_119 & _EVAL_4029;
  assign _EVAL_2212 = _EVAL_1586 | _EVAL_4013;
  assign _EVAL_2288 = _EVAL_1686 & _EVAL_2212;
  assign _EVAL_4509 = _EVAL_315 ? _EVAL_1314 : _EVAL_2288;
  assign _EVAL_3654 = _EVAL_2411 & _EVAL_4509;
  assign _EVAL_5118 = _EVAL_3698 | _EVAL_3654;
  assign _EVAL_5322 = _EVAL_862 | _EVAL_5118;
  assign _EVAL_5402 = _EVAL_274 == _EVAL_5129;
  assign _EVAL_5415 = _EVAL_39 & _EVAL_5402;
  assign _EVAL_4369 = _EVAL_180 == _EVAL_5129;
  assign _EVAL_4265 = _EVAL_188 & _EVAL_4369;
  assign _EVAL_427 = _EVAL_5415 | _EVAL_4265;
  assign _EVAL_2580 = _EVAL_427 | _EVAL_2902;
  assign _EVAL_3970 = _EVAL_591 & _EVAL_2580;
  assign _EVAL_1371 = _EVAL_68 == _EVAL_5129;
  assign _EVAL_3129 = _EVAL_179 & _EVAL_1371;
  assign _EVAL_1669 = _EVAL_5373 | _EVAL_3129;
  assign _EVAL_805 = _EVAL_4127 == _EVAL_5129;
  assign _EVAL_3699 = _EVAL_119 & _EVAL_805;
  assign _EVAL_2492 = _EVAL_1669 | _EVAL_3699;
  assign _EVAL_3835 = _EVAL_591 & _EVAL_2492;
  assign _EVAL_2728 = _EVAL_315 ? _EVAL_3970 : _EVAL_3835;
  assign _EVAL_1743 = _EVAL_5322 | _EVAL_2728;
  assign _EVAL_4916 = _EVAL_1743 | _EVAL_2875;
  assign _EVAL_4111 = _EVAL_4299 & _EVAL_39;
  assign _EVAL_3303 = _EVAL_4692 & _EVAL_205;
  assign _EVAL_773 = _EVAL_4111 | _EVAL_3303;
  assign _EVAL_4187 = _EVAL_274 == _EVAL_4135;
  assign _EVAL_1900 = _EVAL_773 & _EVAL_4187;
  assign _EVAL_3348 = _EVAL_180 == _EVAL_4135;
  assign _EVAL_1252 = _EVAL_5187 & _EVAL_3348;
  assign _EVAL_1906 = _EVAL_1900 | _EVAL_1252;
  assign _EVAL_293 = _EVAL_4299 & _EVAL_260;
  assign _EVAL_2531 = _EVAL_3212 == _EVAL_4135;
  assign _EVAL_2170 = _EVAL_293 & _EVAL_2531;
  assign _EVAL_5346 = _EVAL_1906 | _EVAL_2170;
  assign _EVAL_435 = _EVAL_4299 & _EVAL_148;
  assign _EVAL_3343 = _EVAL_4692 & _EVAL_1;
  assign _EVAL_4042 = _EVAL_435 | _EVAL_3343;
  assign _EVAL_4071 = _EVAL_154 == _EVAL_4135;
  assign _EVAL_5040 = _EVAL_4042 & _EVAL_4071;
  assign _EVAL_4821 = _EVAL_4299 & _EVAL_179;
  assign _EVAL_3779 = _EVAL_4692 & _EVAL_141;
  assign _EVAL_2891 = _EVAL_4821 | _EVAL_3779;
  assign _EVAL_5116 = _EVAL_68 == _EVAL_4135;
  assign _EVAL_4381 = _EVAL_2891 & _EVAL_5116;
  assign _EVAL_4137 = _EVAL_5040 | _EVAL_4381;
  assign _EVAL_5098 = _EVAL_4137 | _EVAL_286;
  assign _EVAL_1131 = _EVAL_315 ? _EVAL_5346 : _EVAL_5098;
  assign _EVAL_3761 = _EVAL_4240 & _EVAL_1131;
  assign _EVAL_5147 = _EVAL_315 ? _EVAL_3761 : _EVAL_3761;
  assign _EVAL_2789 = _EVAL_4692 & _EVAL_2258;
  assign _EVAL_3589 = _EVAL_4299 | _EVAL_2789;
  assign _EVAL_4057 = _EVAL_5147 & _EVAL_3589;
  assign _EVAL_3895 = _EVAL_4916 | _EVAL_4057;
  assign _EVAL_4582 = _EVAL_315 ? _EVAL_650 : _EVAL_650;
  assign _EVAL_4286 = fpu__EVAL_0 > 3'h1;
  assign _EVAL_868 = fpu__EVAL_4 | _EVAL_4286;
  assign _EVAL_2182 = fpu__EVAL_49 & _EVAL_868;
  assign _EVAL_1584 = _EVAL_4582 & _EVAL_2182;
  assign _EVAL_4250 = _EVAL_3895 | _EVAL_1584;
  assign _EVAL_1422 = _EVAL_2369 & _EVAL_39;
  assign _EVAL_3213 = _EVAL_2219 & _EVAL_205;
  assign _EVAL_3264 = _EVAL_1422 | _EVAL_3213;
  assign _EVAL_2574 = _EVAL_274 == _EVAL_3742;
  assign _EVAL_4243 = _EVAL_3264 & _EVAL_2574;
  assign _EVAL_4852 = _EVAL_2369 & _EVAL_188;
  assign _EVAL_2585 = _EVAL_2219 & _EVAL_250;
  assign _EVAL_5287 = _EVAL_4852 | _EVAL_2585;
  assign _EVAL_1258 = _EVAL_180 == _EVAL_3742;
  assign _EVAL_3647 = _EVAL_5287 & _EVAL_1258;
  assign _EVAL_4742 = _EVAL_4243 | _EVAL_3647;
  assign _EVAL_3486 = _EVAL_2369 & _EVAL_260;
  assign _EVAL_1008 = _EVAL_3212 == _EVAL_3742;
  assign _EVAL_1667 = _EVAL_3486 & _EVAL_1008;
  assign _EVAL_4156 = _EVAL_4742 | _EVAL_1667;
  assign _EVAL_3234 = _EVAL_2369 & _EVAL_148;
  assign _EVAL_344 = _EVAL_2219 & _EVAL_1;
  assign _EVAL_2917 = _EVAL_3234 | _EVAL_344;
  assign _EVAL_4792 = _EVAL_154 == _EVAL_3742;
  assign _EVAL_5345 = _EVAL_2917 & _EVAL_4792;
  assign _EVAL_1799 = _EVAL_2369 & _EVAL_179;
  assign _EVAL_4500 = _EVAL_2219 & _EVAL_141;
  assign _EVAL_2597 = _EVAL_1799 | _EVAL_4500;
  assign _EVAL_4650 = _EVAL_68 == _EVAL_3742;
  assign _EVAL_594 = _EVAL_2597 & _EVAL_4650;
  assign _EVAL_3809 = _EVAL_5345 | _EVAL_594;
  assign _EVAL_966 = _EVAL_2369 & _EVAL_119;
  assign _EVAL_3501 = _EVAL_4127 == _EVAL_3742;
  assign _EVAL_3739 = _EVAL_966 & _EVAL_3501;
  assign _EVAL_2028 = _EVAL_3809 | _EVAL_3739;
  assign _EVAL_3290 = _EVAL_315 ? _EVAL_4156 : _EVAL_2028;
  assign _EVAL_4136 = _EVAL_3227 & _EVAL_3290;
  assign _EVAL_3541 = _EVAL_315 ? _EVAL_4136 : _EVAL_4136;
  assign _EVAL_4441 = _EVAL_3541 & _EVAL_3085;
  assign _EVAL_1234 = _EVAL_4441 & _EVAL_2219;
  assign _EVAL_2987 = _EVAL_4250 | _EVAL_1234;
  assign _EVAL_3812 = _EVAL_2963 & _EVAL_2987;
  assign _EVAL_4055 = _EVAL_2812 == _EVAL_2193;
  assign _EVAL_1011 = _EVAL_5386 & _EVAL_4055;
  assign _EVAL_2839 = _EVAL_3705[11:7];
  assign _EVAL_3158 = _EVAL_315 ? _EVAL_274 : _EVAL_154;
  assign _EVAL_4169 = {_EVAL_2400,_EVAL_4513,_EVAL_3158,_EVAL_5022};
  assign _EVAL_997 = $signed(_EVAL_4169);
  assign _EVAL_4665 = _EVAL_997[8];
  assign _EVAL_3928 = _EVAL_3309[2];
  assign _EVAL_1334 = _EVAL_4705 & _EVAL_3928;
  assign _EVAL_4467 = _EVAL_1334 & _EVAL_2923;
  assign _EVAL_4175 = _EVAL_873 == 1'h0;
  assign _EVAL_1519 = _EVAL_4467 & _EVAL_4175;
  assign _EVAL_1804 = _EVAL_4019[0];
  assign _EVAL_1278 = _EVAL_1519 & _EVAL_1804;
  assign _EVAL_2710 = _EVAL_1278 == 1'h0;
  assign _EVAL_856 = _EVAL_4776 > 3'h1;
  assign _EVAL_3659 = _EVAL_2812 == _EVAL_180;
  assign _EVAL_417 = _EVAL_5386 & _EVAL_3659;
  assign _EVAL_1556 = _EVAL_4468 ^ 32'h80000000;
  assign _EVAL_2936 = {1'b0,$signed(_EVAL_1556)};
  assign _EVAL_2262 = $signed(_EVAL_2936) & $signed(-33'sh20000);
  assign _EVAL_1385 = $signed(_EVAL_2262);
  assign _EVAL_476 = $signed(_EVAL_1385) == $signed(33'sh0);
  assign _EVAL_3043 = _EVAL_476 == 1'h0;
  assign _EVAL_5032 = _EVAL_545 & _EVAL_3043;
  assign _EVAL_1071 = _EVAL_315 ? _EVAL_5071 : _EVAL_2817;
  assign _EVAL_4716 = _EVAL_2118 & _EVAL_1071;
  assign _EVAL_3444 = _EVAL_315 ? _EVAL_4716 : _EVAL_4716;
  assign _EVAL_1998 = _EVAL_2118 & _EVAL_2847;
  assign _EVAL_2019 = _EVAL_315 ? _EVAL_1998 : _EVAL_1998;
  assign _EVAL_3191 = _EVAL_3444 | _EVAL_2019;
  assign _EVAL_3857 = _EVAL_5032 & _EVAL_3191;
  assign _EVAL_2163 = _EVAL_58 & _EVAL_3608;
  assign _EVAL_5303 = _EVAL_268 & _EVAL_4043;
  assign _EVAL_5255 = _EVAL_2163 | _EVAL_5303;
  assign _EVAL_4032 = _EVAL_91 == _EVAL_3117;
  assign _EVAL_1566 = _EVAL_5255 & _EVAL_4032;
  assign _EVAL_2340 = _EVAL_16 & _EVAL_3608;
  assign _EVAL_4930 = _EVAL_214 & _EVAL_4043;
  assign _EVAL_599 = _EVAL_2340 | _EVAL_4930;
  assign _EVAL_4867 = _EVAL_171 == _EVAL_3117;
  assign _EVAL_4677 = _EVAL_599 & _EVAL_4867;
  assign _EVAL_2882 = _EVAL_315 ? _EVAL_1566 : _EVAL_4677;
  assign _EVAL_395 = _EVAL_2326 & _EVAL_2882;
  assign _EVAL_4753 = _EVAL_315 ? _EVAL_395 : _EVAL_395;
  assign _EVAL_2069 = _EVAL_1349 | _EVAL_4753;
  assign _EVAL_940 = _EVAL_2138 & _EVAL_2069;
  assign _EVAL_2235 = _EVAL_3857 | _EVAL_940;
  assign _EVAL_3154 = _EVAL_4962 & _EVAL_148;
  assign _EVAL_4199 = _EVAL_1333 & _EVAL_1;
  assign _EVAL_2097 = _EVAL_3154 | _EVAL_4199;
  assign _EVAL_1565 = _EVAL_154 == _EVAL_4706;
  assign _EVAL_3061 = _EVAL_2097 & _EVAL_1565;
  assign _EVAL_3390 = _EVAL_4962 & _EVAL_179;
  assign _EVAL_5035 = _EVAL_1333 & _EVAL_141;
  assign _EVAL_804 = _EVAL_3390 | _EVAL_5035;
  assign _EVAL_3768 = _EVAL_68 == _EVAL_4706;
  assign _EVAL_691 = _EVAL_804 & _EVAL_3768;
  assign _EVAL_5174 = _EVAL_3061 | _EVAL_691;
  assign _EVAL_2972 = _EVAL_4962 & _EVAL_119;
  assign _EVAL_1700 = _EVAL_4127 == _EVAL_4706;
  assign _EVAL_958 = _EVAL_2972 & _EVAL_1700;
  assign _EVAL_4767 = _EVAL_5174 | _EVAL_958;
  assign _EVAL_2979 = _EVAL_4962 & _EVAL_39;
  assign _EVAL_842 = _EVAL_2979 | _EVAL_630;
  assign _EVAL_4893 = _EVAL_274 == _EVAL_4706;
  assign _EVAL_2704 = _EVAL_842 & _EVAL_4893;
  assign _EVAL_1170 = _EVAL_180 == _EVAL_4706;
  assign _EVAL_2771 = _EVAL_4724 & _EVAL_1170;
  assign _EVAL_4555 = _EVAL_2704 | _EVAL_2771;
  assign _EVAL_4691 = _EVAL_4962 & _EVAL_260;
  assign _EVAL_2210 = _EVAL_3212 == _EVAL_4706;
  assign _EVAL_4428 = _EVAL_4691 & _EVAL_2210;
  assign _EVAL_1437 = _EVAL_4555 | _EVAL_4428;
  assign _EVAL_570 = _EVAL_315 ? _EVAL_4767 : _EVAL_1437;
  assign _EVAL_3263 = _EVAL_2506 & _EVAL_570;
  assign _EVAL_4627 = _EVAL_315 ? _EVAL_3263 : _EVAL_3263;
  assign _EVAL_1946 = _EVAL_315 ? _EVAL_4714 : _EVAL_4714;
  assign _EVAL_3949 = _EVAL_4627 | _EVAL_1946;
  assign _EVAL_3059 = _EVAL_3404 & _EVAL_3949;
  assign _EVAL_3717 = _EVAL_2235 | _EVAL_3059;
  assign _EVAL_5273 = _EVAL_4362 & _EVAL_39;
  assign _EVAL_2177 = _EVAL_332 & _EVAL_205;
  assign _EVAL_2408 = _EVAL_5273 | _EVAL_2177;
  assign _EVAL_1935 = _EVAL_274 == _EVAL_5099;
  assign _EVAL_606 = _EVAL_2408 & _EVAL_1935;
  assign _EVAL_1851 = _EVAL_4362 & _EVAL_188;
  assign _EVAL_1800 = _EVAL_332 & _EVAL_250;
  assign _EVAL_4479 = _EVAL_1851 | _EVAL_1800;
  assign _EVAL_2045 = _EVAL_180 == _EVAL_5099;
  assign _EVAL_2855 = _EVAL_4479 & _EVAL_2045;
  assign _EVAL_3224 = _EVAL_606 | _EVAL_2855;
  assign _EVAL_334 = _EVAL_4362 & _EVAL_260;
  assign _EVAL_891 = _EVAL_3212 == _EVAL_5099;
  assign _EVAL_5375 = _EVAL_334 & _EVAL_891;
  assign _EVAL_1108 = _EVAL_3224 | _EVAL_5375;
  assign _EVAL_823 = _EVAL_315 ? _EVAL_5046 : _EVAL_1108;
  assign _EVAL_5234 = _EVAL_4000 & _EVAL_823;
  assign _EVAL_1977 = _EVAL_315 ? _EVAL_5234 : _EVAL_5234;
  assign _EVAL_4349 = _EVAL_58 & _EVAL_4362;
  assign _EVAL_2530 = _EVAL_268 & _EVAL_332;
  assign _EVAL_465 = _EVAL_4349 | _EVAL_2530;
  assign _EVAL_3996 = _EVAL_91 == _EVAL_5099;
  assign _EVAL_1346 = _EVAL_465 & _EVAL_3996;
  assign _EVAL_1595 = _EVAL_16 & _EVAL_4362;
  assign _EVAL_1861 = _EVAL_214 & _EVAL_332;
  assign _EVAL_3466 = _EVAL_1595 | _EVAL_1861;
  assign _EVAL_1925 = _EVAL_171 == _EVAL_5099;
  assign _EVAL_4281 = _EVAL_3466 & _EVAL_1925;
  assign _EVAL_3244 = _EVAL_315 ? _EVAL_1346 : _EVAL_4281;
  assign _EVAL_1725 = _EVAL_4000 & _EVAL_3244;
  assign _EVAL_1496 = _EVAL_315 ? _EVAL_1725 : _EVAL_1725;
  assign _EVAL_989 = _EVAL_1977 | _EVAL_1496;
  assign _EVAL_1989 = _EVAL_954 & _EVAL_989;
  assign _EVAL_2738 = _EVAL_3717 | _EVAL_1989;
  assign _EVAL_1363 = {_EVAL_1452,_EVAL_3117};
  assign _EVAL_4559 = $signed(_EVAL_1363);
  assign _EVAL_285 = {_EVAL_1452,_EVAL_2193};
  assign _EVAL_4338 = $signed(_EVAL_285);
  assign _EVAL_4202 = _EVAL_971 ? $signed(_EVAL_4559) : $signed(_EVAL_4338);
  assign _EVAL_3570 = $unsigned(_EVAL_4202);
  assign _EVAL_2576 = _EVAL_3570[11];
  assign _EVAL_5041 = _EVAL_4329 & 32'h90000010;
  assign _EVAL_5243 = _EVAL_1 & _EVAL_4071;
  assign _EVAL_4359 = _EVAL_4692 & _EVAL_5243;
  assign _EVAL_1329 = _EVAL_205 & _EVAL_4187;
  assign _EVAL_3450 = _EVAL_4692 & _EVAL_1329;
  assign _EVAL_878 = _EVAL_315 ? _EVAL_4359 : _EVAL_3450;
  assign _EVAL_3890 = _EVAL_4240 & _EVAL_878;
  assign _EVAL_2020 = _EVAL_1475 & 32'h30;
  assign _EVAL_1701 = {_EVAL_16,_EVAL_171};
  assign _EVAL_1161 = _EVAL_4160 >> _EVAL_1701;
  assign _EVAL_4772 = _EVAL_1161[0];
  assign _EVAL_4324 = _EVAL_2823 == _EVAL_1701;
  assign _EVAL_5216 = _EVAL_1535 & _EVAL_4324;
  assign _EVAL_2893 = _EVAL_4772 | _EVAL_5216;
  assign _EVAL_3237 = _EVAL_2617 == _EVAL_1701;
  assign _EVAL_3493 = divider__EVAL_2 & _EVAL_3237;
  assign _EVAL_4628 = _EVAL_2893 | _EVAL_3493;
  assign _EVAL_4542 = _EVAL_315 ? _EVAL_3763 : _EVAL_5360;
  assign _EVAL_972 = _EVAL_4240 & _EVAL_4542;
  assign _EVAL_4507 = _EVAL_315 ? _EVAL_972 : _EVAL_972;
  assign _EVAL_1173 = _EVAL_4608 & _EVAL_4507;
  assign _EVAL_3183 = _EVAL_315 ? _EVAL_4067 : _EVAL_1158;
  assign _EVAL_2809 = _EVAL_3624 & _EVAL_3183;
  assign _EVAL_4151 = _EVAL_315 ? _EVAL_2809 : _EVAL_2809;
  assign _EVAL_1650 = _EVAL_1823 & _EVAL_4151;
  assign _EVAL_4666 = _EVAL_1173 | _EVAL_1650;
  assign _EVAL_1135 = _EVAL_315 ? _EVAL_2654 : _EVAL_4937;
  assign _EVAL_282 = _EVAL_3227 & _EVAL_1135;
  assign _EVAL_3936 = _EVAL_315 ? _EVAL_282 : _EVAL_282;
  assign _EVAL_1592 = _EVAL_781 & _EVAL_3936;
  assign _EVAL_2136 = _EVAL_4666 | _EVAL_1592;
  assign _EVAL_5279 = _EVAL_315 ? _EVAL_1640 : _EVAL_1086;
  assign _EVAL_2861 = _EVAL_315 ? _EVAL_647 : _EVAL_5355;
  assign _EVAL_3722 = csr__EVAL_105 ? 1'h1 : _EVAL_2861;
  assign _EVAL_2622 = _EVAL_5279 | _EVAL_3722;
  assign _EVAL_3055 = _EVAL_2622 | _EVAL_327;
  assign _EVAL_1683 = _EVAL_3896 & _EVAL_3055;
  assign _EVAL_5369 = _EVAL_2136 | _EVAL_1683;
  assign _EVAL_1582 = _EVAL_5369 | _EVAL_601;
  assign _EVAL_2614 = _EVAL_1582 | _EVAL_1149;
  assign _EVAL_3130 = _EVAL_2614 | _EVAL_3528;
  assign _EVAL_3751 = _EVAL_2094 == 1'h0;
  assign _EVAL_3275 = _EVAL_4570 & _EVAL_3751;
  assign _EVAL_1239 = _EVAL_3275 & _EVAL_3119;
  assign _EVAL_2756 = _EVAL_3299 & _EVAL_1239;
  assign _EVAL_319 = _EVAL_2152 & _EVAL_4103;
  assign _EVAL_1287 = _EVAL_3299 & _EVAL_319;
  assign _EVAL_2535 = _EVAL_2756 | _EVAL_1287;
  assign _EVAL_5320 = _EVAL_3030 == 1'h0;
  assign _EVAL_2057 = _EVAL_2535 & _EVAL_5320;
  assign _EVAL_2687 = _EVAL_3269 | _EVAL_1910;
  assign _EVAL_434 = _EVAL_2118 & _EVAL_2687;
  assign _EVAL_4597 = _EVAL_190 == 1'h0;
  assign _EVAL_1695 = _EVAL_434 | _EVAL_4597;
  assign _EVAL_3341 = _EVAL_1695 | _EVAL_1997;
  assign _EVAL_1247 = _EVAL_2057 & _EVAL_3341;
  assign _EVAL_1209 = _EVAL_2198 & _EVAL_1247;
  assign _EVAL_5352 = _EVAL_107 == 1'h0;
  assign _EVAL_657 = _EVAL_434 & _EVAL_5352;
  assign _EVAL_3350 = _EVAL_29 == 1'h0;
  assign _EVAL_2795 = _EVAL_657 | _EVAL_3350;
  assign _EVAL_2188 = _EVAL_2057 & _EVAL_2795;
  assign _EVAL_1809 = _EVAL_1209 | _EVAL_2188;
  assign _EVAL_3339 = _EVAL_3130 | _EVAL_1809;
  assign _EVAL_3832 = _EVAL_3598 == 5'h3;
  assign _EVAL_2047 = _EVAL_315 ? _EVAL_153 : _EVAL_84;
  assign _EVAL_2277 = _EVAL_2047[0];
  assign _EVAL_3312 = _EVAL_3832 & _EVAL_2277;
  assign _EVAL_5076 = _EVAL_2277 == 1'h0;
  assign _EVAL_4900 = _EVAL_3832 & _EVAL_5076;
  assign _EVAL_3688 = _EVAL_315 ? _EVAL_68 : _EVAL_180;
  assign _EVAL_2338 = _EVAL_3688[3:2];
  assign _EVAL_4808 = _EVAL_416[2:1];
  assign _EVAL_1150 = _EVAL_2338 | _EVAL_4808;
  assign _EVAL_4718 = _EVAL_1150 != 2'h0;
  assign _EVAL_4205 = _EVAL_416[0];
  assign _EVAL_3889 = _EVAL_3688[4];
  assign _EVAL_3510 = _EVAL_4205 | _EVAL_3889;
  assign _EVAL_2842 = {{1'd0}, _EVAL_3510};
  assign _EVAL_5081 = _EVAL_3688[1:0];
  assign _EVAL_5286 = _EVAL_2842 | _EVAL_5081;
  assign _EVAL_2234 = _EVAL_5286 != 2'h0;
  assign _EVAL_3428 = _EVAL_4718 & _EVAL_2234;
  assign _EVAL_5019 = _EVAL_3428 | _EVAL_4718;
  assign _EVAL_1624 = _EVAL_5019 | _EVAL_2234;
  assign _EVAL_3663 = _EVAL_4900 & _EVAL_1624;
  assign _EVAL_1562 = _EVAL_3312 | _EVAL_3663;
  assign _EVAL_5088 = _EVAL_1287 & _EVAL_4205;
  assign _EVAL_976 = _EVAL_1562 | _EVAL_5088;
  assign _EVAL_1014 = _EVAL_1908 & _EVAL_3299;
  assign _EVAL_729 = _EVAL_976 | _EVAL_1014;
  assign _EVAL_2994 = _EVAL_1905 & _EVAL_729;
  assign _EVAL_3920 = _EVAL_3339 | _EVAL_2994;
  assign _EVAL_3918 = _EVAL_233 == 1'h0;
  assign _EVAL_4953 = _EVAL_2176 & _EVAL_3918;
  assign _EVAL_2930 = _EVAL_3299 & _EVAL_4953;
  assign _EVAL_5368 = _EVAL_3920 | _EVAL_2930;
  assign _EVAL_2206 = _EVAL_5368 | _EVAL_2738;
  assign _EVAL_3417 = _EVAL_2206 | _EVAL_3870;
  assign _EVAL_4140 = _EVAL_2798 == 1'h0;
  assign _EVAL_817 = _EVAL_3417 | _EVAL_4140;
  assign _EVAL_2561 = _EVAL_2118 & _EVAL_3747;
  assign _EVAL_4166 = _EVAL_327 & _EVAL_2561;
  assign _EVAL_3944 = _EVAL_817 | _EVAL_4166;
  assign _EVAL_816 = _EVAL_4299 | _EVAL_2258;
  assign _EVAL_4347 = _EVAL_4240 & _EVAL_816;
  assign _EVAL_881 = _EVAL_2573 | _EVAL_1854;
  assign _EVAL_4216 = _EVAL_3624 & _EVAL_881;
  assign _EVAL_1085 = _EVAL_4347 | _EVAL_4216;
  assign _EVAL_4845 = _EVAL_327 & _EVAL_1085;
  assign _EVAL_317 = _EVAL_3944 | _EVAL_4845;
  assign _EVAL_1520 = fpu__EVAL_20 | fpu__EVAL_22;
  assign _EVAL_1091 = fpu__EVAL_13 | _EVAL_1520;
  assign _EVAL_1455 = _EVAL_327 & _EVAL_1091;
  assign _EVAL_2888 = _EVAL_317 | _EVAL_1455;
  assign _EVAL_5366 = _EVAL_3452 == 1'h0;
  assign _EVAL_2022 = _EVAL_315 ? _EVAL_1440 : _EVAL_853;
  assign _EVAL_3222 = _EVAL_4706 == _EVAL_68;
  assign _EVAL_4015 = _EVAL_1333 & _EVAL_3222;
  assign _EVAL_389 = _EVAL_2506 & _EVAL_4015;
  assign _EVAL_2821 = _EVAL_4706 == _EVAL_180;
  assign _EVAL_4422 = _EVAL_1333 & _EVAL_2821;
  assign _EVAL_4463 = _EVAL_2506 & _EVAL_4422;
  assign _EVAL_2544 = _EVAL_315 ? _EVAL_389 : _EVAL_4463;
  assign _EVAL_1518 = _EVAL_315 ? _EVAL_1993 : _EVAL_5055;
  assign _EVAL_730 = _EVAL_5099 == _EVAL_68;
  assign _EVAL_5146 = _EVAL_332 & _EVAL_730;
  assign _EVAL_736 = _EVAL_4774 & _EVAL_5146;
  assign _EVAL_3001 = _EVAL_5099 == _EVAL_180;
  assign _EVAL_847 = _EVAL_332 & _EVAL_3001;
  assign _EVAL_2139 = _EVAL_4774 & _EVAL_847;
  assign _EVAL_4073 = _EVAL_315 ? _EVAL_736 : _EVAL_2139;
  assign _EVAL_1865 = _EVAL_2812 == _EVAL_68;
  assign _EVAL_4546 = _EVAL_5386 & _EVAL_1865;
  assign _EVAL_2825 = _EVAL_5252 & _EVAL_4546;
  assign _EVAL_3329 = _EVAL_5252 & _EVAL_417;
  assign _EVAL_3531 = _EVAL_315 ? _EVAL_2825 : _EVAL_3329;
  assign _EVAL_1214 = _EVAL_708__EVAL_712_data;
  assign _EVAL_4515 = _EVAL_708__EVAL_710_data;
  assign _EVAL_4770 = _EVAL_315 ? _EVAL_1214 : _EVAL_4515;
  assign _EVAL_872 = _EVAL_3531 ? _EVAL_3187 : _EVAL_4770;
  assign _EVAL_4561 = _EVAL_4073 ? _EVAL_4863 : _EVAL_872;
  assign _EVAL_2412 = _EVAL_1518 ? _EVAL_3923 : _EVAL_4561;
  assign _EVAL_1471 = _EVAL_2544 ? _EVAL_4399 : _EVAL_2412;
  assign _EVAL_422 = _EVAL_2022 ? _EVAL_2919 : _EVAL_1471;
  assign _EVAL_2363 = _EVAL_2667 == 1'h0;
  assign _EVAL_4316 = _EVAL_4721 & _EVAL_2363;
  assign _EVAL_2096 = _EVAL_993 == 1'h0;
  assign _EVAL_3867 = _EVAL_4721 & _EVAL_2096;
  assign _EVAL_4489 = _EVAL_3867 & _EVAL_4736;
  assign _EVAL_4287 = _EVAL_4316 + _EVAL_4489;
  assign _EVAL_906 = _EVAL_4947 == 1'h0;
  assign _EVAL_429 = _EVAL_4620 == 1'h0;
  assign _EVAL_5300 = _EVAL_906 & _EVAL_429;
  assign _EVAL_4453 = _EVAL_890 & _EVAL_5300;
  assign _EVAL_1486 = _EVAL_925 == 1'h0;
  assign _EVAL_3614 = _EVAL_3476 == 1'h0;
  assign _EVAL_2952 = _EVAL_1486 & _EVAL_3614;
  assign _EVAL_2453 = _EVAL_890 & _EVAL_2952;
  assign _EVAL_3602 = _EVAL_2453 & _EVAL_1499;
  assign _EVAL_307 = _EVAL_4453 + _EVAL_3602;
  assign _EVAL_3579 = _EVAL_4287 + _EVAL_307;
  assign _EVAL_2981 = _EVAL_3316 & _EVAL_3995;
  assign _EVAL_3677 = _EVAL_2981 ? _EVAL_1024 : 3'h2;
  assign _EVAL_1627 = _EVAL_3788 == 1'h0;
  assign _EVAL_634 = _EVAL_1049 & 32'h64;
  assign _EVAL_2227 = _EVAL_634 == 32'h0;
  assign _EVAL_2104 = _EVAL_1049 & 32'h50;
  assign _EVAL_2419 = _EVAL_2104 == 32'h10;
  assign _EVAL_3946 = _EVAL_2227 | _EVAL_2419;
  assign _EVAL_3836 = _EVAL_1049 & 32'h2024;
  assign _EVAL_2458 = _EVAL_3836 == 32'h24;
  assign _EVAL_4754 = _EVAL_3946 | _EVAL_2458;
  assign _EVAL_1684 = _EVAL_1049 & 32'h28;
  assign _EVAL_2553 = _EVAL_1684 == 32'h28;
  assign _EVAL_3323 = _EVAL_4754 | _EVAL_2553;
  assign _EVAL_5150 = _EVAL_517 == 32'h30;
  assign _EVAL_5214 = _EVAL_3323 | _EVAL_5150;
  assign _EVAL_3049 = _EVAL_1049 & 32'h90000010;
  assign _EVAL_502 = _EVAL_3049 == 32'h80000010;
  assign _EVAL_4352 = _EVAL_5214 | _EVAL_502;
  assign _EVAL_2980 = _EVAL_1049[11:7];
  assign _EVAL_4105 = _EVAL_2980 != 5'h0;
  assign _EVAL_1802 = _EVAL_4352 & _EVAL_4105;
  assign _EVAL_1502 = {{4'd0}, _EVAL_596};
  assign _EVAL_5372 = _EVAL_1502 ^ 9'h1ff;
  assign _EVAL_335 = _EVAL_2899 ? _EVAL_5372 : {{1'd0}, _EVAL_3894};
  assign _EVAL_3963 = _EVAL_335 + _EVAL_4547;
  assign _EVAL_1687 = {1'b0,$signed(_EVAL_3963)};
  assign _EVAL_2959 = _EVAL_1687[8:6];
  assign _EVAL_3926 = _EVAL_590 ? 3'h0 : _EVAL_2959;
  assign _EVAL_959 = csr__EVAL_150;
  assign _EVAL_965 = _EVAL_959 == 1'h0;
  assign _EVAL_721 = csr__EVAL_24;
  assign _EVAL_3937 = csr__EVAL_116;
  assign _EVAL_1553 = {_EVAL_721,1'h0,1'h0,_EVAL_3937};
  assign _EVAL_5132 = _EVAL_1553 >> _EVAL_5168;
  assign _EVAL_2155 = _EVAL_5132[0];
  assign _EVAL_1648 = _EVAL_3149 & _EVAL_2155;
  assign _EVAL_393 = csr__EVAL_133;
  assign _EVAL_3026 = _EVAL_1648 & _EVAL_393;
  assign _EVAL_2715 = csr__EVAL_35;
  assign _EVAL_471 = _EVAL_2715[1];
  assign _EVAL_3919 = csr__EVAL_132;
  assign _EVAL_3882 = _EVAL_3641 >= _EVAL_3919;
  assign _EVAL_3697 = _EVAL_2715[0];
  assign _EVAL_4233 = _EVAL_3882 ^ _EVAL_3697;
  assign _EVAL_1792 = _EVAL_3919[0];
  assign _EVAL_4964 = _EVAL_3697 & _EVAL_1792;
  assign _EVAL_3875 = _EVAL_3919[1];
  assign _EVAL_5169 = _EVAL_4964 & _EVAL_3875;
  assign _EVAL_2356 = _EVAL_3919[2];
  assign _EVAL_2272 = _EVAL_5169 & _EVAL_2356;
  assign _EVAL_2883 = {_EVAL_2272,_EVAL_5169,_EVAL_4964,_EVAL_3697};
  assign _EVAL_1798 = {{28'd0}, _EVAL_2883};
  assign _EVAL_3846 = _EVAL_2867 | _EVAL_1798;
  assign _EVAL_5027 = ~ _EVAL_3919;
  assign _EVAL_1418 = _EVAL_5027 | _EVAL_1798;
  assign _EVAL_4569 = _EVAL_3846 == _EVAL_1418;
  assign _EVAL_2105 = _EVAL_471 ? _EVAL_4233 : _EVAL_4569;
  assign _EVAL_1269 = _EVAL_3026 & _EVAL_2105;
  assign _EVAL_5229 = _EVAL_965 & _EVAL_1269;
  assign _EVAL_4782 = csr__EVAL_26;
  assign _EVAL_1009 = _EVAL_4782 == 1'h0;
  assign _EVAL_4261 = _EVAL_1009 | _EVAL_2435;
  assign _EVAL_3218 = _EVAL_5229 & _EVAL_4261;
  assign _EVAL_1817 = csr__EVAL_141;
  assign _EVAL_834 = _EVAL_1009 & _EVAL_2435;
  assign _EVAL_2100 = csr__EVAL_79;
  assign _EVAL_4459 = _EVAL_834 ? _EVAL_2100 : 1'h0;
  assign _EVAL_1967 = _EVAL_3218 ? _EVAL_1817 : _EVAL_4459;
  assign _EVAL_561 = _EVAL_315 ? _EVAL_5376 : _EVAL_1853;
  assign _EVAL_3278 = _EVAL_3742 == _EVAL_2495;
  assign _EVAL_472 = _EVAL_2219 & _EVAL_3278;
  assign _EVAL_1832 = _EVAL_3227 & _EVAL_472;
  assign _EVAL_2114 = _EVAL_332 & _EVAL_3512;
  assign _EVAL_418 = _EVAL_4774 & _EVAL_2114;
  assign _EVAL_3604 = _EVAL_2812 == _EVAL_2495;
  assign _EVAL_3007 = _EVAL_5386 & _EVAL_3604;
  assign _EVAL_948 = _EVAL_5252 & _EVAL_3007;
  assign _EVAL_1425 = _EVAL_948 ? _EVAL_3187 : _EVAL_1109;
  assign _EVAL_5313 = _EVAL_418 ? _EVAL_4863 : _EVAL_1425;
  assign _EVAL_3044 = _EVAL_1832 ? _EVAL_3923 : _EVAL_5313;
  assign _EVAL_4645 = _EVAL_4774 & _EVAL_4362;
  assign _EVAL_2611 = _EVAL_5099 == _EVAL_3711;
  assign _EVAL_3414 = _EVAL_4645 & _EVAL_2611;
  assign _EVAL_4190 = _EVAL_3444 & _EVAL_3747;
  assign _EVAL_995 = csr__EVAL_155 | csr__EVAL_89;
  assign _EVAL_3736 = _EVAL_315 ? _EVAL_1 : _EVAL_205;
  assign _EVAL_1597 = _EVAL_3736 == 1'h0;
  assign _EVAL_3047 = _EVAL_1597 & _EVAL_3751;
  assign _EVAL_4176 = _EVAL_316 & _EVAL_873;
  assign _EVAL_3496 = _EVAL_1446 & _EVAL_4176;
  assign _EVAL_3649 = csr__EVAL_12;
  assign _EVAL_4896 = _EVAL_3649[0];
  assign _EVAL_2996 = _EVAL_2619[0];
  assign _EVAL_4943 = _EVAL_4896 & _EVAL_2996;
  assign _EVAL_4389 = _EVAL_2619[1];
  assign _EVAL_3050 = _EVAL_4943 & _EVAL_4389;
  assign _EVAL_2676 = _EVAL_3050 & _EVAL_1244;
  assign _EVAL_1691 = _EVAL_2146 & _EVAL_2515;
  assign _EVAL_686 = _EVAL_3085 & _EVAL_3504;
  assign _EVAL_646 = _EVAL_2146 & _EVAL_3372;
  assign _EVAL_2557 = _EVAL_2146 & _EVAL_5393;
  assign _EVAL_1982 = _EVAL_3568 == 1'h0;
  assign _EVAL_4223 = _EVAL_2915 & _EVAL_1982;
  assign _EVAL_1889 = {_EVAL_4405,_EVAL_5120,_EVAL_5329,_EVAL_4223,_EVAL_854,4'h0};
  assign _EVAL_2065 = {_EVAL_1246,_EVAL_1691,_EVAL_686,_EVAL_646,_EVAL_2557,2'h0,_EVAL_781,_EVAL_4150,_EVAL_1889};
  assign _EVAL_2864 = {{6'd0}, _EVAL_2065};
  assign _EVAL_362 = _EVAL_5323 & _EVAL_2864;
  assign _EVAL_2605 = {_EVAL_188,_EVAL_180};
  assign _EVAL_3584 = _EVAL_4160 >> _EVAL_2605;
  assign _EVAL_1754 = _EVAL_3584[0];
  assign _EVAL_3542 = _EVAL_315 ? _EVAL_4463 : _EVAL_389;
  assign _EVAL_2697 = _EVAL_315 ? _EVAL_5055 : _EVAL_1993;
  assign _EVAL_2186 = _EVAL_315 ? _EVAL_2139 : _EVAL_736;
  assign _EVAL_4397 = _EVAL_315 ? _EVAL_3329 : _EVAL_2825;
  assign _EVAL_1793 = _EVAL_315 ? _EVAL_4515 : _EVAL_1214;
  assign _EVAL_2140 = _EVAL_4397 ? _EVAL_3187 : _EVAL_1793;
  assign _EVAL_2091 = _EVAL_2186 ? _EVAL_4863 : _EVAL_2140;
  assign _EVAL_3830 = _EVAL_2697 ? _EVAL_3923 : _EVAL_2091;
  assign _EVAL_3704 = _EVAL_3542 ? _EVAL_4399 : _EVAL_3830;
  assign _EVAL_907 = _EVAL_3922[2:1];
  assign _EVAL_4430 = {_EVAL_4019,_EVAL_1198,_EVAL_4715,_EVAL_4201,_EVAL_4706,_EVAL_3309,2'h3};
  assign _EVAL_1928 = _EVAL_3705 & 32'h64;
  assign _EVAL_348 = _EVAL_1928 == 32'h0;
  assign _EVAL_5067 = _EVAL_3705 & 32'h50;
  assign _EVAL_1755 = _EVAL_5067 == 32'h10;
  assign _EVAL_1807 = _EVAL_348 | _EVAL_1755;
  assign _EVAL_3435 = _EVAL_3705 & 32'h2024;
  assign _EVAL_4344 = _EVAL_3435 == 32'h24;
  assign _EVAL_1933 = _EVAL_1807 | _EVAL_4344;
  assign _EVAL_2005 = _EVAL_3705 & 32'h28;
  assign _EVAL_2714 = _EVAL_2005 == 32'h28;
  assign _EVAL_3254 = _EVAL_1933 | _EVAL_2714;
  assign _EVAL_4685 = _EVAL_3705 & 32'h30;
  assign _EVAL_3214 = _EVAL_4685 == 32'h30;
  assign _EVAL_2928 = _EVAL_3254 | _EVAL_3214;
  assign _EVAL_1226 = _EVAL_3705 & 32'h90000010;
  assign _EVAL_5396 = _EVAL_1226 == 32'h80000010;
  assign _EVAL_2736 = _EVAL_2928 | _EVAL_5396;
  assign _EVAL_2251 = _EVAL_2839 != 5'h0;
  assign _EVAL_1923 = _EVAL_2736 & _EVAL_2251;
  assign _EVAL_3014 = _EVAL_2522 & 32'h64;
  assign _EVAL_4340 = _EVAL_3014 == 32'h0;
  assign _EVAL_3096 = _EVAL_2522 & 32'h50;
  assign _EVAL_2323 = _EVAL_3096 == 32'h10;
  assign _EVAL_2083 = _EVAL_4340 | _EVAL_2323;
  assign _EVAL_1421 = _EVAL_2643 == 32'h24;
  assign _EVAL_5342 = _EVAL_2083 | _EVAL_1421;
  assign _EVAL_3762 = _EVAL_2522 & 32'h28;
  assign _EVAL_2294 = _EVAL_3762 == 32'h28;
  assign _EVAL_3554 = _EVAL_5342 | _EVAL_2294;
  assign _EVAL_4267 = _EVAL_2522 & 32'h30;
  assign _EVAL_2907 = _EVAL_4267 == 32'h30;
  assign _EVAL_536 = _EVAL_3554 | _EVAL_2907;
  assign _EVAL_835 = _EVAL_2522 & 32'h90000010;
  assign _EVAL_2267 = _EVAL_835 == 32'h80000010;
  assign _EVAL_785 = _EVAL_536 | _EVAL_2267;
  assign _EVAL_1332 = _EVAL_785 & _EVAL_4894;
  assign _EVAL_5331 = _EVAL_1475 & 32'h64;
  assign _EVAL_4304 = _EVAL_5331 == 32'h0;
  assign _EVAL_4275 = _EVAL_1475 & 32'h50;
  assign _EVAL_604 = _EVAL_4275 == 32'h10;
  assign _EVAL_410 = _EVAL_4304 | _EVAL_604;
  assign _EVAL_4128 = _EVAL_410 | _EVAL_1262;
  assign _EVAL_2957 = _EVAL_1475 & 32'h28;
  assign _EVAL_5294 = _EVAL_2957 == 32'h28;
  assign _EVAL_2444 = _EVAL_4128 | _EVAL_5294;
  assign _EVAL_3465 = _EVAL_2020 == 32'h30;
  assign _EVAL_3868 = _EVAL_2444 | _EVAL_3465;
  assign _EVAL_1419 = _EVAL_1475 & 32'h90000010;
  assign _EVAL_4081 = _EVAL_1419 == 32'h80000010;
  assign _EVAL_4647 = _EVAL_3868 | _EVAL_4081;
  assign _EVAL_3765 = _EVAL_1475[11:7];
  assign _EVAL_2754 = _EVAL_3765 != 5'h0;
  assign _EVAL_3744 = _EVAL_4647 & _EVAL_2754;
  assign _EVAL_1964 = _EVAL_961 & 32'h90000010;
  assign _EVAL_4610 = _EVAL_1964 == 32'h80000010;
  assign _EVAL_3721 = _EVAL_1679 | _EVAL_4610;
  assign _EVAL_5405 = _EVAL_961[11:7];
  assign _EVAL_3289 = _EVAL_5405 != 5'h0;
  assign _EVAL_2123 = _EVAL_3721 & _EVAL_3289;
  assign _EVAL_800 = _EVAL_2180 ? _EVAL_3744 : _EVAL_2123;
  assign _EVAL_1185 = _EVAL_544 ? _EVAL_1332 : _EVAL_800;
  assign _EVAL_692 = _EVAL_757 ? _EVAL_1923 : _EVAL_1185;
  assign _EVAL_3558 = _EVAL_2180 ? _EVAL_3765 : _EVAL_5405;
  assign _EVAL_5153 = _EVAL_544 ? _EVAL_2637 : _EVAL_3558;
  assign _EVAL_4611 = _EVAL_757 ? _EVAL_2839 : _EVAL_5153;
  assign _EVAL_4179 = _EVAL_692 ? _EVAL_4611 : 5'h0;
  assign _EVAL_1443 = _EVAL_4179;
  assign _EVAL_2366 = _EVAL_1588 & _EVAL_1922;
  assign _EVAL_4673 = _EVAL_884[12];
  assign _EVAL_1730 = _EVAL_4673 ? 19'h7ffff : 19'h0;
  assign _EVAL_5128 = {_EVAL_1730,_EVAL_884};
  assign _EVAL_2701 = _EVAL_2366 ? _EVAL_5128 : 32'h0;
  assign _EVAL_1736 = _EVAL_1588 & _EVAL_405;
  assign _EVAL_3969 = _EVAL_997[19];
  assign _EVAL_2489 = _EVAL_997[7:0];
  assign _EVAL_4425 = _EVAL_997[18:9];
  assign _EVAL_2641 = {_EVAL_3969,_EVAL_2489,_EVAL_4665,_EVAL_4425,1'h0};
  assign _EVAL_1991 = $signed(_EVAL_2641);
  assign _EVAL_1674 = $unsigned(_EVAL_1991);
  assign _EVAL_1688 = _EVAL_1674[20];
  assign _EVAL_1390 = _EVAL_1688 ? 11'h7ff : 11'h0;
  assign _EVAL_3981 = {_EVAL_1390,_EVAL_1674};
  assign _EVAL_672 = _EVAL_1736 ? _EVAL_3981 : 32'h0;
  assign _EVAL_407 = _EVAL_2701 | _EVAL_672;
  assign _EVAL_455 = _EVAL_1588 == 1'h0;
  assign _EVAL_2500 = _EVAL_455 & _EVAL_405;
  assign _EVAL_3288 = $unsigned(_EVAL_997);
  assign _EVAL_326 = {_EVAL_3288, 12'h0};
  assign _EVAL_3021 = _EVAL_2500 ? _EVAL_326 : 32'h0;
  assign _EVAL_3095 = _EVAL_407 | _EVAL_3021;
  assign _EVAL_4602 = _EVAL_1588 | _EVAL_4988;
  assign _EVAL_3080 = _EVAL_1922 == 1'h0;
  assign _EVAL_3583 = _EVAL_4602 & _EVAL_3080;
  assign _EVAL_583 = _EVAL_725 & _EVAL_3583;
  assign _EVAL_2048 = $unsigned(_EVAL_527);
  assign _EVAL_4800 = _EVAL_2048[11];
  assign _EVAL_1978 = _EVAL_4800 ? 20'hfffff : 20'h0;
  assign _EVAL_1765 = {_EVAL_1978,_EVAL_2048};
  assign _EVAL_4232 = _EVAL_583 ? _EVAL_1765 : 32'h0;
  assign _EVAL_1886 = _EVAL_3095 | _EVAL_4232;
  assign _EVAL_1344 = _EVAL_1922 & _EVAL_455;
  assign _EVAL_683 = _EVAL_315 ? _EVAL_4874 : _EVAL_2986;
  assign _EVAL_5179 = _EVAL_315 ? _EVAL_2228 : _EVAL_2468;
  assign _EVAL_3042 = _EVAL_315 ? _EVAL_1177 : _EVAL_1693;
  assign _EVAL_2081 = _EVAL_315 ? _EVAL_853 : _EVAL_1440;
  assign _EVAL_1464 = _EVAL_2081 ? _EVAL_2919 : _EVAL_3704;
  assign _EVAL_514 = _EVAL_3042 ? _EVAL_4679 : _EVAL_1464;
  assign _EVAL_4929 = _EVAL_5179 ? _EVAL_1932 : _EVAL_514;
  assign _EVAL_4744 = _EVAL_683 ? _EVAL_1572 : _EVAL_4929;
  assign _EVAL_2029 = _EVAL_1344 ? _EVAL_4744 : 32'h0;
  assign _EVAL_2194 = _EVAL_1886 | _EVAL_2029;
  assign _EVAL_4174 = _EVAL_315 ? _EVAL_1858 : _EVAL_581;
  assign _EVAL_3609 = _EVAL_315 ? _EVAL_2478 : _EVAL_4824;
  assign _EVAL_1656 = _EVAL_315 ? _EVAL_3527 : _EVAL_3847;
  assign _EVAL_4417 = _EVAL_315 ? _EVAL_4977 : _EVAL_1485;
  assign _EVAL_3197 = _EVAL_969 ? _EVAL_3187 : _EVAL_561;
  assign _EVAL_3695 = _EVAL_4417 ? _EVAL_4863 : _EVAL_3197;
  assign _EVAL_425 = _EVAL_1656 ? _EVAL_3923 : _EVAL_3695;
  assign _EVAL_481 = _EVAL_3609 ? _EVAL_4399 : _EVAL_425;
  assign _EVAL_2933 = _EVAL_4174 ? _EVAL_2919 : _EVAL_481;
  assign _EVAL_2425 = csr__EVAL_107;
  assign _EVAL_4734 = _EVAL_4215 & _EVAL_2425;
  assign _EVAL_3662 = _EVAL_4734 & _EVAL_2229;
  assign _EVAL_3074 = _EVAL_1009 & _EVAL_3662;
  assign _EVAL_2632 = _EVAL_3391 | _EVAL_1122;
  assign _EVAL_749 = _EVAL_4507 & _EVAL_4299;
  assign _EVAL_4709 = $signed(_EVAL_3432);
  assign _EVAL_3078 = _EVAL_214 | _EVAL_16;
  assign _EVAL_3630 = _EVAL_4158 == _EVAL_1701;
  assign _EVAL_1025 = _EVAL_1190 & _EVAL_3630;
  assign _EVAL_3345 = _EVAL_4628 | _EVAL_1025;
  assign _EVAL_2377 = _EVAL_3078 & _EVAL_3345;
  assign _EVAL_2184 = _EVAL_205 | _EVAL_39;
  assign _EVAL_5045 = {_EVAL_39,_EVAL_274};
  assign _EVAL_5403 = _EVAL_4160 >> _EVAL_5045;
  assign _EVAL_3921 = _EVAL_5403[0];
  assign _EVAL_4337 = _EVAL_2823 == _EVAL_5045;
  assign _EVAL_4310 = _EVAL_1535 & _EVAL_4337;
  assign _EVAL_2292 = _EVAL_3921 | _EVAL_4310;
  assign _EVAL_337 = _EVAL_2617 == _EVAL_5045;
  assign _EVAL_1459 = divider__EVAL_2 & _EVAL_337;
  assign _EVAL_1199 = _EVAL_2292 | _EVAL_1459;
  assign _EVAL_1056 = _EVAL_4158 == _EVAL_5045;
  assign _EVAL_4657 = _EVAL_1190 & _EVAL_1056;
  assign _EVAL_1395 = _EVAL_1199 | _EVAL_4657;
  assign _EVAL_3576 = _EVAL_2184 & _EVAL_1395;
  assign _EVAL_2165 = _EVAL_2377 | _EVAL_3576;
  assign _EVAL_3287 = _EVAL_250 | _EVAL_188;
  assign _EVAL_2311 = _EVAL_2823 == _EVAL_2605;
  assign _EVAL_2410 = _EVAL_1535 & _EVAL_2311;
  assign _EVAL_3152 = _EVAL_1754 | _EVAL_2410;
  assign _EVAL_4478 = _EVAL_2617 == _EVAL_2605;
  assign _EVAL_3097 = divider__EVAL_2 & _EVAL_4478;
  assign _EVAL_4346 = _EVAL_3152 | _EVAL_3097;
  assign _EVAL_3267 = _EVAL_4158 == _EVAL_2605;
  assign _EVAL_2398 = _EVAL_1190 & _EVAL_3267;
  assign _EVAL_2539 = _EVAL_4346 | _EVAL_2398;
  assign _EVAL_3235 = _EVAL_3287 & _EVAL_2539;
  assign _EVAL_5160 = _EVAL_2165 | _EVAL_3235;
  assign _EVAL_1204 = _EVAL_5160 | _EVAL_532;
  assign _EVAL_1176 = _EVAL_315 ? _EVAL_1204 : _EVAL_3256;
  assign _EVAL_2402 = _EVAL_2963 & _EVAL_1176;
  assign _EVAL_950 = _EVAL_3616 == 2'h1;
  assign _EVAL_2017 = _EVAL_1588 & _EVAL_950;
  assign _EVAL_2168 = _EVAL_2017 | _EVAL_2013;
  assign _EVAL_1360 = _EVAL_2168 | _EVAL_2545;
  assign _EVAL_824 = _EVAL_1122 == 1'h0;
  assign _EVAL_1846 = _EVAL_449 & _EVAL_824;
  assign _EVAL_2479 = _EVAL_3588 == 1'h0;
  assign _EVAL_4285 = _EVAL_5147 & _EVAL_2479;
  assign _EVAL_5251 = _EVAL_1846 | _EVAL_4285;
  assign _EVAL_2905 = _EVAL_315 ? _EVAL_3033 : _EVAL_1714;
  assign _EVAL_3380 = _EVAL_2326 & _EVAL_2905;
  assign _EVAL_2708 = _EVAL_315 ? _EVAL_3380 : _EVAL_3380;
  assign _EVAL_3013 = _EVAL_2708 & _EVAL_1487;
  assign _EVAL_4815 = _EVAL_5251 | _EVAL_3013;
  assign _EVAL_855 = _EVAL_4582 & _EVAL_1206;
  assign _EVAL_2881 = _EVAL_4815 | _EVAL_855;
  assign _EVAL_1118 = _EVAL_1360 & _EVAL_2881;
  assign _EVAL_1115 = _EVAL_2963 & _EVAL_1118;
  assign _EVAL_2117 = {1'h0,_EVAL_95,1'h0,_EVAL_2402,_EVAL_1115};
  assign _EVAL_4074 = _EVAL_649 == 5'h3;
  assign _EVAL_5008 = _EVAL_4607[0];
  assign _EVAL_1055 = _EVAL_4074 & _EVAL_5008;
  assign _EVAL_1664 = _EVAL_2583 & _EVAL_3624;
  assign _EVAL_2154 = _EVAL_2765 ? 2'h2 : 2'h0;
  assign _EVAL_4913 = _EVAL_2542 ? 3'h4 : 3'h6;
  assign _EVAL_1045 = _EVAL_2542 ? 4'h6 : 4'h8;
  assign _EVAL_3826 = _EVAL_1521 ? {{1'd0}, _EVAL_4913} : _EVAL_1045;
  assign _EVAL_4603 = _EVAL_2542 ? 3'h2 : 3'h4;
  assign _EVAL_1202 = _EVAL_2753 ? _EVAL_3826 : {{1'd0}, _EVAL_4603};
  assign _EVAL_3543 = _EVAL_5226 ? {{2'd0}, _EVAL_2154} : _EVAL_1202;
  assign _EVAL_4642 = {{28'd0}, _EVAL_3543};
  assign _EVAL_1834 = _EVAL_3132 + _EVAL_4642;
  assign _EVAL_5306 = _EVAL_1834 != _EVAL_4157;
  assign _EVAL_2681 = _EVAL_1664 & _EVAL_5306;
  assign _EVAL_2342 = _EVAL_1055 | _EVAL_2681;
  assign _EVAL_506 = _EVAL_2342 ? 1'h1 : _EVAL_937;
  assign _EVAL_2040 = _EVAL_3624 ? 1'h1 : _EVAL_506;
  assign _EVAL_5154 = csr__EVAL_20;
  assign _EVAL_2709 = _EVAL_315 ? _EVAL_2028 : _EVAL_4156;
  assign _EVAL_5239 = _EVAL_3227 & _EVAL_2709;
  assign _EVAL_5133 = _EVAL_315 ? _EVAL_5239 : _EVAL_5239;
  assign _EVAL_2122 = _EVAL_5133 & _EVAL_3085;
  assign _EVAL_716 = _EVAL_2122 & _EVAL_2219;
  assign _EVAL_4435 = _EVAL_4000 & _EVAL_490;
  assign _EVAL_3052 = _EVAL_1664 == 1'h0;
  assign _EVAL_3520 = _EVAL_881 | _EVAL_3176;
  assign _EVAL_5341 = {_EVAL_2030,_EVAL_2495};
  assign _EVAL_1462 = $signed(_EVAL_5341);
  assign _EVAL_2450 = $unsigned(_EVAL_1462);
  assign _EVAL_5050 = _EVAL_2450[11];
  assign _EVAL_833 = _EVAL_5050 ? 20'hfffff : 20'h0;
  assign _EVAL_4472 = {_EVAL_833,_EVAL_2450};
  assign _EVAL_4333 = _EVAL_2499 ? _EVAL_4472 : 32'h0;
  assign _EVAL_4960 = _EVAL_4706 == _EVAL_2495;
  assign _EVAL_3434 = _EVAL_1333 & _EVAL_4960;
  assign _EVAL_4882 = _EVAL_2506 & _EVAL_3434;
  assign _EVAL_2153 = _EVAL_4882 ? _EVAL_4399 : _EVAL_3044;
  assign _EVAL_1152 = _EVAL_2989 ? _EVAL_2153 : 32'h0;
  assign _EVAL_4041 = _EVAL_4333 | _EVAL_1152;
  assign _EVAL_2351 = _EVAL_2145 ? {{28'd0}, _EVAL_3515} : _EVAL_4041;
  assign _EVAL_944 = _EVAL_3520 ? 32'h0 : _EVAL_2351;
  assign _EVAL_4967 = _EVAL_3624 ? _EVAL_944 : {{27'd0}, _EVAL_3370};
  assign _EVAL_2546 = _EVAL_1557[6:0];
  assign _EVAL_297 = 128'h1 << _EVAL_2546;
  assign _EVAL_5349 = _EVAL_3019 | _EVAL_297;
  assign _EVAL_1943 = _EVAL_1588 ? _EVAL_3080 : 1'h1;
  assign _EVAL_1248 = _EVAL_725 & _EVAL_1943;
  assign _EVAL_3319 = _EVAL_315 ? _EVAL_1980 : _EVAL_801;
  assign _EVAL_3073 = _EVAL_315 ? _EVAL_4281 : _EVAL_1346;
  assign _EVAL_4079 = _EVAL_4000 & _EVAL_3073;
  assign _EVAL_4106 = csr__EVAL_60;
  assign _EVAL_3259 = csr__EVAL_161;
  assign _EVAL_985 = {_EVAL_4106,1'h0,1'h0,_EVAL_3259};
  assign _EVAL_1466 = _EVAL_985 >> _EVAL_5168;
  assign _EVAL_655 = _EVAL_1466[0];
  assign _EVAL_3571 = _EVAL_3149 & _EVAL_655;
  assign _EVAL_1411 = csr__EVAL_67;
  assign _EVAL_4217 = _EVAL_3571 & _EVAL_1411;
  assign _EVAL_497 = _EVAL_3649[1];
  assign _EVAL_3844 = _EVAL_3641 >= _EVAL_2619;
  assign _EVAL_4689 = _EVAL_3844 ^ _EVAL_4896;
  assign _EVAL_2852 = {_EVAL_2676,_EVAL_3050,_EVAL_4943,_EVAL_4896};
  assign _EVAL_420 = {{28'd0}, _EVAL_2852};
  assign _EVAL_368 = _EVAL_2867 | _EVAL_420;
  assign _EVAL_4533 = ~ _EVAL_2619;
  assign _EVAL_1368 = _EVAL_4533 | _EVAL_420;
  assign _EVAL_2082 = _EVAL_368 == _EVAL_1368;
  assign _EVAL_2036 = _EVAL_497 ? _EVAL_4689 : _EVAL_2082;
  assign _EVAL_2575 = _EVAL_4217 & _EVAL_2036;
  assign _EVAL_1222 = _EVAL_2912[31];
  assign _EVAL_2879 = _EVAL_3963[8:7];
  assign _EVAL_5259 = _EVAL_2879 == 2'h3;
  assign _EVAL_394 = _EVAL_299 == 1'h0;
  assign _EVAL_947 = _EVAL_5259 & _EVAL_394;
  assign _EVAL_1038 = {{2'd0}, _EVAL_947};
  assign _EVAL_4291 = _EVAL_3926 | _EVAL_1038;
  assign _EVAL_4075 = _EVAL_1687[5:0];
  assign _EVAL_3606 = _EVAL_2353[22:0];
  assign _EVAL_1004 = {_EVAL_1222,_EVAL_4291,_EVAL_4075,_EVAL_3606};
  assign _EVAL_3732 = _EVAL_448 | _EVAL_4008;
  assign _EVAL_625 = {{2'd0}, _EVAL_3732};
  assign _EVAL_2035 = _EVAL_3677 ^ _EVAL_625;
  assign _EVAL_2661 = _EVAL_2035[0];
  assign _EVAL_2787 = _EVAL_2035[2];
  assign _EVAL_5173 = _EVAL_2787 == 1'h0;
  assign _EVAL_2286 = _EVAL_2035[1];
  assign _EVAL_5384 = _EVAL_2286 == 1'h0;
  assign _EVAL_4932 = _EVAL_5173 & _EVAL_5384;
  assign _EVAL_1153 = _EVAL_2661 ^ _EVAL_4932;
  assign _EVAL_1238 = _EVAL_1973 ? _EVAL_1153 : _EVAL_2661;
  assign _EVAL_2841 = csr__EVAL_123[12:0];
  assign _EVAL_1883 = csr__EVAL_29;
  assign _EVAL_1602 = _EVAL_1883[0];
  assign _EVAL_3795 = _EVAL_3399[0];
  assign _EVAL_4133 = _EVAL_1602 & _EVAL_3795;
  assign _EVAL_2445 = _EVAL_3399[1];
  assign _EVAL_4356 = _EVAL_4133 & _EVAL_2445;
  assign _EVAL_4132 = _EVAL_3399[2];
  assign _EVAL_1579 = _EVAL_4356 & _EVAL_4132;
  assign _EVAL_4700 = {_EVAL_1579,_EVAL_4356,_EVAL_4133,_EVAL_1602};
  assign _EVAL_5136 = _EVAL_4531 == 1'h0;
  assign _EVAL_3693 = _EVAL_5136 ? _EVAL_2331 : _EVAL_3845;
  assign _EVAL_4601 = _EVAL_3693;
  assign _EVAL_5388 = _EVAL_3742 == _EVAL_4460;
  assign _EVAL_5171 = _EVAL_2219 & _EVAL_5388;
  assign _EVAL_4236 = _EVAL_3227 & _EVAL_5171;
  assign _EVAL_3032 = _EVAL_612 == 1'h0;
  assign _EVAL_1454 = _EVAL_5114 & 32'h64;
  assign _EVAL_292 = _EVAL_1454 == 32'h0;
  assign _EVAL_414 = _EVAL_292 | _EVAL_3271;
  assign _EVAL_4165 = _EVAL_414 | _EVAL_2990;
  assign _EVAL_1316 = _EVAL_5114 & 32'h28;
  assign _EVAL_1907 = _EVAL_1316 == 32'h28;
  assign _EVAL_2232 = _EVAL_4165 | _EVAL_1907;
  assign _EVAL_1738 = _EVAL_5114 & 32'h30;
  assign _EVAL_4314 = _EVAL_1738 == 32'h30;
  assign _EVAL_5109 = _EVAL_2232 | _EVAL_4314;
  assign _EVAL_2043 = _EVAL_5114 & 32'h90000010;
  assign _EVAL_1622 = _EVAL_2043 == 32'h80000010;
  assign _EVAL_3553 = _EVAL_5109 | _EVAL_1622;
  assign _EVAL_3433 = _EVAL_3943 != 5'h0;
  assign _EVAL_582 = _EVAL_3553 & _EVAL_3433;
  assign _EVAL_4884 = _EVAL_2302 & 32'h64;
  assign _EVAL_2760 = _EVAL_4884 == 32'h0;
  assign _EVAL_3332 = _EVAL_2302 & 32'h50;
  assign _EVAL_4253 = _EVAL_3332 == 32'h10;
  assign _EVAL_4332 = _EVAL_2760 | _EVAL_4253;
  assign _EVAL_3479 = _EVAL_2302 & 32'h2024;
  assign _EVAL_3388 = _EVAL_3479 == 32'h24;
  assign _EVAL_2312 = _EVAL_4332 | _EVAL_3388;
  assign _EVAL_1456 = _EVAL_2302 & 32'h28;
  assign _EVAL_3563 = _EVAL_1456 == 32'h28;
  assign _EVAL_1814 = _EVAL_2312 | _EVAL_3563;
  assign _EVAL_371 = _EVAL_2302 & 32'h30;
  assign _EVAL_1689 = _EVAL_371 == 32'h30;
  assign _EVAL_3371 = _EVAL_1814 | _EVAL_1689;
  assign _EVAL_2024 = _EVAL_2302 & 32'h90000010;
  assign _EVAL_4096 = _EVAL_2024 == 32'h80000010;
  assign _EVAL_5014 = _EVAL_3371 | _EVAL_4096;
  assign _EVAL_1538 = _EVAL_504 != 5'h0;
  assign _EVAL_1867 = _EVAL_5014 & _EVAL_1538;
  assign _EVAL_4797 = _EVAL_4329 & 32'h64;
  assign _EVAL_4107 = _EVAL_4797 == 32'h0;
  assign _EVAL_4631 = _EVAL_4329 & 32'h50;
  assign _EVAL_4738 = _EVAL_4631 == 32'h10;
  assign _EVAL_4618 = _EVAL_4107 | _EVAL_4738;
  assign _EVAL_860 = _EVAL_4329 & 32'h2024;
  assign _EVAL_1195 = _EVAL_860 == 32'h24;
  assign _EVAL_549 = _EVAL_4618 | _EVAL_1195;
  assign _EVAL_892 = _EVAL_841 == 32'h28;
  assign _EVAL_4652 = _EVAL_549 | _EVAL_892;
  assign _EVAL_4090 = _EVAL_4329 & 32'h30;
  assign _EVAL_5149 = _EVAL_4090 == 32'h30;
  assign _EVAL_2220 = _EVAL_4652 | _EVAL_5149;
  assign _EVAL_1359 = _EVAL_5041 == 32'h80000010;
  assign _EVAL_916 = _EVAL_2220 | _EVAL_1359;
  assign _EVAL_2465 = _EVAL_5382 != 5'h0;
  assign _EVAL_5371 = _EVAL_916 & _EVAL_2465;
  assign _EVAL_3611 = _EVAL_1926 ? _EVAL_1867 : _EVAL_5371;
  assign _EVAL_1207 = _EVAL_2164 ? _EVAL_582 : _EVAL_3611;
  assign _EVAL_1942 = _EVAL_1535 | _EVAL_2869;
  assign _EVAL_4002 = _EVAL_2345 | _EVAL_1149;
  assign _EVAL_5404 = _EVAL_3149 & _EVAL_451;
  assign _EVAL_1051 = csr__EVAL_34;
  assign _EVAL_2370 = _EVAL_5404 & _EVAL_1051;
  assign _EVAL_2496 = _EVAL_1883[1];
  assign _EVAL_1871 = _EVAL_3641 >= _EVAL_3399;
  assign _EVAL_2291 = _EVAL_1871 ^ _EVAL_1602;
  assign _EVAL_4956 = {{28'd0}, _EVAL_4700};
  assign _EVAL_1087 = _EVAL_2867 | _EVAL_4956;
  assign _EVAL_3449 = ~ _EVAL_3399;
  assign _EVAL_5001 = _EVAL_3449 | _EVAL_4956;
  assign _EVAL_1829 = _EVAL_1087 == _EVAL_5001;
  assign _EVAL_2269 = _EVAL_2496 ? _EVAL_2291 : _EVAL_1829;
  assign _EVAL_1277 = _EVAL_2370 & _EVAL_2269;
  assign _EVAL_2112 = _EVAL_3672 == 1'h0;
  assign _EVAL_2352 = _EVAL_416[6:4];
  assign _EVAL_3219 = {{1'd0}, _EVAL_2352};
  assign _EVAL_3819 = _EVAL_315 ? _EVAL_1437 : _EVAL_4767;
  assign _EVAL_1463 = _EVAL_2506 & _EVAL_3819;
  assign _EVAL_4436 = _EVAL_3309[4:2];
  assign _EVAL_3958 = _EVAL_2100 == 1'h0;
  assign _EVAL_2711 = _EVAL_3884 ? _EVAL_5412 : 32'h0;
  assign _EVAL_534 = _EVAL_3496 == 1'h0;
  assign _EVAL_3592 = _EVAL_4480 & _EVAL_534;
  assign _EVAL_2767 = _EVAL_2326 & _EVAL_4842;
  assign _EVAL_728 = _EVAL_5022[1:0];
  assign _EVAL_3445 = _EVAL_728 == 2'h1;
  assign _EVAL_3398 = _EVAL_707 == 1'h0;
  assign _EVAL_2067 = _EVAL_1118 | _EVAL_1176;
  assign _EVAL_372 = _EVAL_3688[3:0];
  assign _EVAL_1904 = _EVAL_372 == 4'h0;
  assign _EVAL_4955 = _EVAL_4900 & _EVAL_1904;
  assign _EVAL_2974 = _EVAL_1476 ? 3'h4 : 3'h6;
  assign _EVAL_3002 = _EVAL_1476 ? 4'h6 : 4'h8;
  assign _EVAL_5406 = _EVAL_1187 ? {{1'd0}, _EVAL_2974} : _EVAL_3002;
  assign _EVAL_1453 = _EVAL_1476 ? 3'h2 : 3'h4;
  assign _EVAL_3794 = _EVAL_2329 ? _EVAL_5406 : {{1'd0}, _EVAL_1453};
  assign _EVAL_2690 = $signed(_EVAL_3794);
  assign _EVAL_2862 = _EVAL_3170 ? $signed({{9{_EVAL_2690[3]}},_EVAL_2690}) : $signed(_EVAL_3159);
  assign _EVAL_3022 = fpu__EVAL_41 == 1'h0;
  assign _EVAL_4130 = fpu__EVAL_49 & _EVAL_3022;
  assign _EVAL_1216 = _EVAL_4130 ? 1'h1 : _EVAL_1097;
  assign _EVAL_3260 = _EVAL_854 & _EVAL_5185;
  assign _EVAL_1157 = _EVAL_5363 == 5'h0;
  assign _EVAL_3459 = _EVAL_3260 & _EVAL_1157;
  assign _EVAL_1398 = _EVAL_3459 == 1'h0;
  assign _EVAL_3009 = _EVAL_4987 & _EVAL_1398;
  assign _EVAL_5230 = {_EVAL_4075,_EVAL_3606};
  assign _EVAL_1601 = _EVAL_1009 | _EVAL_3662;
  assign _EVAL_996 = _EVAL_416[5];
  assign _EVAL_3818 = _EVAL_2756 | _EVAL_2203;
  assign _EVAL_3597 = _EVAL_3598[2];
  assign _EVAL_3361 = _EVAL_4570 & _EVAL_3597;
  assign _EVAL_2740 = _EVAL_315 ? _EVAL_141 : _EVAL_250;
  assign _EVAL_1380 = _EVAL_2740 == 1'h0;
  assign _EVAL_486 = _EVAL_3361 & _EVAL_1380;
  assign _EVAL_2945 = _EVAL_3818 | _EVAL_486;
  assign _EVAL_4944 = _EVAL_3736 & _EVAL_2945;
  assign _EVAL_1504 = _EVAL_98 != _EVAL_315;
  assign _EVAL_1181 = _EVAL_2084 & _EVAL_1504;
  assign _EVAL_325 = _EVAL_315 ? _EVAL_4654 : _EVAL_3853;
  assign _EVAL_2921 = csr__EVAL_93;
  assign _EVAL_839 = _EVAL_3571 & _EVAL_2921;
  assign _EVAL_5068 = _EVAL_839 & _EVAL_2036;
  assign _EVAL_359 = _EVAL_4607[1:0];
  assign _EVAL_5260 = _EVAL_359 != 2'h0;
  assign _EVAL_3517 = fpu__EVAL_29 == _EVAL_4400;
  assign _EVAL_4475 = _EVAL_4729 & _EVAL_3517;
  assign _EVAL_4365 = csr__EVAL_128;
  assign _EVAL_5275 = _EVAL_4365 == 1'h0;
  assign _EVAL_283 = _EVAL_5275 & _EVAL_5068;
  assign _EVAL_4270 = _EVAL_965 | _EVAL_1269;
  assign _EVAL_4025 = _EVAL_283 & _EVAL_4270;
  assign _EVAL_4534 = _EVAL_3624 == 1'h0;
  assign _EVAL_5175 = _EVAL_1895 & _EVAL_4534;
  assign _EVAL_1705 = _EVAL_3227 == 1'h0;
  assign _EVAL_565 = _EVAL_1591 & _EVAL_1705;
  assign _EVAL_569 = _EVAL_5175 | _EVAL_565;
  assign _EVAL_5123 = _EVAL_3309 == 5'h1f;
  assign _EVAL_1589 = _EVAL_3309 == 5'h1e;
  assign _EVAL_1526 = _EVAL_1589 ? _EVAL_1407 : _EVAL_5291;
  assign _EVAL_477 = _EVAL_5123 ? _EVAL_1407 : _EVAL_1526;
  assign _EVAL_4256 = _EVAL_1042 ? {{16'd0}, _EVAL_477} : _EVAL_4430;
  assign _EVAL_1860 = _EVAL_111[5];
  assign _EVAL_3301 = _EVAL_1860 == 1'h0;
  assign _EVAL_1082 = _EVAL_649[0];
  assign _EVAL_4301 = _EVAL_1082 == 1'h0;
  assign _EVAL_1326 = _EVAL_3227 & _EVAL_4405;
  assign _EVAL_1536 = _EVAL_2506 & _EVAL_3746;
  assign _EVAL_934 = fpu__EVAL_0 > 3'h0;
  assign _EVAL_2250 = fpu__EVAL_4 | _EVAL_934;
  assign _EVAL_4118 = _EVAL_1300[0];
  assign _EVAL_5152 = _EVAL_1300[2];
  assign _EVAL_3297 = _EVAL_4118 ^ _EVAL_5152;
  assign _EVAL_2466 = _EVAL_5152 == 1'h0;
  assign _EVAL_3513 = _EVAL_2466 & _EVAL_3398;
  assign _EVAL_1561 = _EVAL_4118 ^ _EVAL_3513;
  assign _EVAL_2664 = _EVAL_1973 ? _EVAL_1561 : _EVAL_4118;
  assign _EVAL_4560 = _EVAL_1225 ? _EVAL_3297 : _EVAL_2664;
  assign _EVAL_3285 = _EVAL_4560 | _EVAL_1511;
  assign _EVAL_4409 = _EVAL_2326 & _EVAL_3052;
  assign _EVAL_2566 = _EVAL_4114 == 1'h0;
  assign _EVAL_1788 = _EVAL_2624 ^ _EVAL_2911;
  assign _EVAL_3011 = _EVAL_2566 | _EVAL_1788;
  assign _EVAL_4393 = _EVAL_2145 & _EVAL_3011;
  assign _EVAL_2092 = _EVAL_4393 ? _EVAL_4461 : _EVAL_4238;
  assign _EVAL_5358 = _EVAL_267;
  assign _EVAL_2999 = _EVAL_2067 | _EVAL_2987;
  assign _EVAL_2451 = divider__EVAL_2 | _EVAL_296;
  assign _EVAL_3153 = _EVAL_2545 & _EVAL_2451;
  assign _EVAL_3675 = _EVAL_2999 | _EVAL_3153;
  assign _EVAL_2534 = _EVAL_2118 & _EVAL_768;
  assign _EVAL_1389 = _EVAL_315 ? _EVAL_2534 : _EVAL_2534;
  assign _EVAL_2147 = _EVAL_449 | _EVAL_1389;
  assign _EVAL_5155 = _EVAL_5032 & _EVAL_2147;
  assign _EVAL_670 = _EVAL_315 ? _EVAL_4677 : _EVAL_1566;
  assign _EVAL_3582 = _EVAL_2326 & _EVAL_670;
  assign _EVAL_3903 = _EVAL_315 ? _EVAL_3582 : _EVAL_3582;
  assign _EVAL_4928 = _EVAL_2708 | _EVAL_3903;
  assign _EVAL_734 = _EVAL_2138 & _EVAL_4928;
  assign _EVAL_2011 = _EVAL_5155 | _EVAL_734;
  assign _EVAL_1137 = _EVAL_315 ? _EVAL_1463 : _EVAL_1463;
  assign _EVAL_3491 = _EVAL_315 ? _EVAL_4227 : _EVAL_2733;
  assign _EVAL_1585 = _EVAL_2506 & _EVAL_3491;
  assign _EVAL_4875 = _EVAL_315 ? _EVAL_1585 : _EVAL_1585;
  assign _EVAL_399 = _EVAL_1137 | _EVAL_4875;
  assign _EVAL_756 = _EVAL_3404 & _EVAL_399;
  assign _EVAL_1461 = _EVAL_2011 | _EVAL_756;
  assign _EVAL_3757 = _EVAL_315 ? _EVAL_1108 : _EVAL_5046;
  assign _EVAL_3121 = _EVAL_4000 & _EVAL_3757;
  assign _EVAL_4980 = _EVAL_315 ? _EVAL_3121 : _EVAL_3121;
  assign _EVAL_697 = _EVAL_315 ? _EVAL_4079 : _EVAL_4079;
  assign _EVAL_1750 = _EVAL_4980 | _EVAL_697;
  assign _EVAL_2205 = _EVAL_954 & _EVAL_1750;
  assign _EVAL_3539 = _EVAL_1461 | _EVAL_2205;
  assign _EVAL_1612 = _EVAL_4002 | _EVAL_3539;
  assign _EVAL_3292 = _EVAL_315 ? _EVAL_90 : _EVAL_247;
  assign _EVAL_3863 = _EVAL_3292 == 1'h0;
  assign _EVAL_1381 = _EVAL_1612 | _EVAL_3863;
  assign _EVAL_1249 = _EVAL_518 & _EVAL_2561;
  assign _EVAL_329 = _EVAL_1381 | _EVAL_1249;
  assign _EVAL_3815 = _EVAL_518 & _EVAL_1085;
  assign _EVAL_1309 = _EVAL_329 | _EVAL_3815;
  assign _EVAL_1539 = _EVAL_518 & _EVAL_1091;
  assign _EVAL_4194 = _EVAL_1309 | _EVAL_1539;
  assign _EVAL_2299 = _EVAL_3675 | _EVAL_4194;
  assign _EVAL_2379 = _EVAL_2299 == 1'h0;
  assign _EVAL_4225 = _EVAL_612 & _EVAL_2443;
  assign _EVAL_2510 = _EVAL_3896 < 1'h1;
  assign _EVAL_4573 = _EVAL_237 | _EVAL_2510;
  assign _EVAL_4788 = _EVAL_55 & _EVAL_4573;
  assign _EVAL_539 = _EVAL_315 ? _EVAL_3256 : _EVAL_1204;
  assign _EVAL_2001 = _EVAL_4788 & _EVAL_539;
  assign _EVAL_2508 = _EVAL_205 & _EVAL_3377;
  assign _EVAL_1013 = _EVAL_3497 | _EVAL_4000;
  assign _EVAL_4827 = _EVAL_1013 | _EVAL_612;
  assign _EVAL_3587 = _EVAL_240[2];
  assign _EVAL_2239 = _EVAL_4827 | _EVAL_3587;
  assign _EVAL_1124 = _EVAL_5099 == _EVAL_2193;
  assign _EVAL_4701 = _EVAL_332 & _EVAL_1124;
  assign _EVAL_1770 = _EVAL_4774 & _EVAL_4701;
  assign _EVAL_3725 = _EVAL_315 ? _EVAL_2288 : _EVAL_1314;
  assign _EVAL_3201 = _EVAL_2302[24:20];
  assign _EVAL_5277 = _EVAL_4329[24:20];
  assign _EVAL_3321 = _EVAL_1926 ? _EVAL_3201 : _EVAL_5277;
  assign _EVAL_3070 = {1'h0,_EVAL_24,_EVAL_156,_EVAL_174,_EVAL_246,_EVAL_36};
  assign _EVAL_701 = {{18'd0}, _EVAL_3070};
  assign _EVAL_2354 = _EVAL_5111 | _EVAL_3520;
  assign _EVAL_3112 = _EVAL_3705[24:20];
  assign _EVAL_3873 = _EVAL_1334 & _EVAL_2710;
  assign _EVAL_4671 = _EVAL_4436 == 3'h7;
  assign _EVAL_4005 = _EVAL_1988 & _EVAL_1400;
  assign _EVAL_1840 = _EVAL_1446 & _EVAL_4005;
  assign _EVAL_3973 = {3'h0,_EVAL_3873,_EVAL_4671,_EVAL_1840,_EVAL_4072,_EVAL_3592,1'h0};
  assign _EVAL_1734 = csr__EVAL_57;
  assign _EVAL_4300 = _EVAL_5404 & _EVAL_1734;
  assign _EVAL_1862 = _EVAL_4300 & _EVAL_2269;
  assign _EVAL_4491 = _EVAL_5275 | _EVAL_2575;
  assign _EVAL_4908 = _EVAL_1862 & _EVAL_4491;
  assign _EVAL_3216 = _EVAL_5154 == 1'h0;
  assign _EVAL_3731 = _EVAL_5275 & _EVAL_2575;
  assign _EVAL_5311 = csr__EVAL_62;
  assign _EVAL_4639 = _EVAL_1648 & _EVAL_5311;
  assign _EVAL_810 = _EVAL_4639 & _EVAL_2105;
  assign _EVAL_4902 = _EVAL_965 | _EVAL_810;
  assign _EVAL_635 = _EVAL_3731 & _EVAL_4902;
  assign _EVAL_2967 = csr__EVAL_65;
  assign _EVAL_4297 = _EVAL_2967 == 1'h0;
  assign _EVAL_2913 = _EVAL_965 & _EVAL_810;
  assign _EVAL_609 = _EVAL_2913 & _EVAL_1601;
  assign _EVAL_402 = _EVAL_1817 == 1'h0;
  assign _EVAL_4831 = _EVAL_3074 ? _EVAL_3958 : 1'h0;
  assign _EVAL_1392 = _EVAL_609 ? _EVAL_402 : _EVAL_4831;
  assign _EVAL_2507 = _EVAL_635 ? _EVAL_4297 : _EVAL_1392;
  assign _EVAL_1460 = _EVAL_4908 ? _EVAL_3216 : _EVAL_2507;
  assign _EVAL_1747 = _EVAL_1446 & _EVAL_81;
  assign _EVAL_5399 = _EVAL_1747 == 1'h0;
  assign _EVAL_4372 = _EVAL_4643 & _EVAL_5399;
  assign _EVAL_4914 = _EVAL_4372 | _EVAL_5104;
  assign _EVAL_559 = _EVAL_1702 | _EVAL_3939;
  assign _EVAL_4272 = _EVAL_3223 == 2'h3;
  assign _EVAL_1402 = _EVAL_4272 ? _EVAL_1802 : _EVAL_1207;
  assign _EVAL_2343 = _EVAL_4272 ? _EVAL_2980 : _EVAL_1847;
  assign _EVAL_3333 = _EVAL_1402 ? _EVAL_2343 : 5'h0;
  assign _EVAL_5278 = _EVAL_1146[1:0];
  assign _EVAL_2840 = _EVAL_5278 == 2'h1;
  assign _EVAL_4802 = _EVAL_5226 == 1'h0;
  assign _EVAL_1610 = _EVAL_4252;
  assign _EVAL_4783 = _EVAL_315 ? _EVAL_2468 : _EVAL_2228;
  assign _EVAL_1052 = _EVAL_315 ? _EVAL_1693 : _EVAL_1177;
  assign _EVAL_4690 = _EVAL_1052 ? _EVAL_4679 : _EVAL_422;
  assign _EVAL_1223 = _EVAL_4783 ? _EVAL_1932 : _EVAL_4690;
  assign _EVAL_2275 = _EVAL_416[3];
  assign _EVAL_1874 = _EVAL_416[2];
  assign _EVAL_5418 = _EVAL_1874 ? 3'h7 : 3'h6;
  assign _EVAL_953 = 4'h8 | _EVAL_3219;
  assign _EVAL_4743 = _EVAL_1874 ? 4'h4 : _EVAL_953;
  assign _EVAL_2189 = _EVAL_2275 ? {{1'd0}, _EVAL_5418} : _EVAL_4743;
  assign _EVAL_2493 = _EVAL_3119 ? 4'h1 : _EVAL_2189;
  assign _EVAL_3313 = fpu__EVAL_25 == _EVAL_4400;
  assign _EVAL_4011 = _EVAL_1686 & _EVAL_3313;
  assign _EVAL_5084 = _EVAL_1475[24:20];
  assign _EVAL_3955 = _EVAL_4151 & _EVAL_2573;
  assign _EVAL_3900 = _EVAL_749 | _EVAL_3955;
  assign _EVAL_4959 = _EVAL_315 ? _EVAL_4260 : _EVAL_821;
  assign _EVAL_5059 = _EVAL_3900 | _EVAL_4959;
  assign _EVAL_893 = _EVAL_1020 & _EVAL_58;
  assign _EVAL_1763 = _EVAL_91 == fpu__EVAL_35;
  assign _EVAL_617 = _EVAL_893 & _EVAL_1763;
  assign _EVAL_3784 = _EVAL_1020 & _EVAL_16;
  assign _EVAL_3020 = _EVAL_171 == fpu__EVAL_35;
  assign _EVAL_1522 = _EVAL_3784 & _EVAL_3020;
  assign _EVAL_2428 = _EVAL_315 ? _EVAL_617 : _EVAL_1522;
  assign _EVAL_1200 = _EVAL_5059 | _EVAL_2428;
  assign _EVAL_1191 = fpu__EVAL_10 > 3'h1;
  assign _EVAL_2591 = _EVAL_315 ? _EVAL_1089 : _EVAL_765;
  assign _EVAL_526 = _EVAL_1191 & _EVAL_2591;
  assign _EVAL_2975 = fpu__EVAL_39 > 3'h1;
  assign _EVAL_3367 = _EVAL_315 ? _EVAL_4058 : _EVAL_4293;
  assign _EVAL_4387 = _EVAL_2975 & _EVAL_3367;
  assign _EVAL_1976 = _EVAL_526 | _EVAL_4387;
  assign _EVAL_2706 = _EVAL_1976 | _EVAL_3808;
  assign _EVAL_3620 = fpu__EVAL_51 > 3'h1;
  assign _EVAL_4540 = _EVAL_3620 & _EVAL_3725;
  assign _EVAL_1947 = _EVAL_2706 | _EVAL_4540;
  assign _EVAL_4414 = _EVAL_1200 | _EVAL_1947;
  assign _EVAL_3392 = _EVAL_315 ? _EVAL_3835 : _EVAL_3970;
  assign _EVAL_3933 = _EVAL_4414 | _EVAL_3392;
  assign _EVAL_398 = _EVAL_1349 & _EVAL_3608;
  assign _EVAL_885 = _EVAL_3933 | _EVAL_398;
  assign _EVAL_2469 = _EVAL_315 ? _EVAL_3304 : _EVAL_3353;
  assign _EVAL_1629 = _EVAL_3624 & _EVAL_2469;
  assign _EVAL_1341 = _EVAL_315 ? _EVAL_1629 : _EVAL_1629;
  assign _EVAL_3764 = _EVAL_1341 & fpu__EVAL_49;
  assign _EVAL_3242 = _EVAL_885 | _EVAL_3764;
  assign _EVAL_2511 = _EVAL_3242 | _EVAL_4190;
  assign _EVAL_3376 = _EVAL_315 ? _EVAL_5098 : _EVAL_5346;
  assign _EVAL_726 = _EVAL_4240 & _EVAL_3376;
  assign _EVAL_406 = _EVAL_315 ? _EVAL_726 : _EVAL_726;
  assign _EVAL_973 = _EVAL_406 & _EVAL_3589;
  assign _EVAL_4242 = _EVAL_2511 | _EVAL_973;
  assign _EVAL_1261 = fpu__EVAL_49 & _EVAL_2250;
  assign _EVAL_2308 = _EVAL_1341 & _EVAL_1261;
  assign _EVAL_1259 = _EVAL_4242 | _EVAL_2308;
  assign _EVAL_1189 = _EVAL_1259 | _EVAL_716;
  assign _EVAL_4189 = _EVAL_4788 & _EVAL_1189;
  assign _EVAL_4415 = _EVAL_315 ? _EVAL_148 : _EVAL_39;
  assign _EVAL_4125 = _EVAL_1278 & _EVAL_3788;
  assign _EVAL_2541 = _EVAL_1278 & _EVAL_1627;
  assign _EVAL_5070 = {5'h0,_EVAL_1162,_EVAL_3496,_EVAL_4125,_EVAL_2541,_EVAL_3973};
  assign _EVAL_5422 = _EVAL_838 & _EVAL_5366;
  assign _EVAL_318 = _EVAL_5422 ? _EVAL_1379 : 3'h2;
  assign _EVAL_1340 = _EVAL_318[0];
  assign _EVAL_2851 = _EVAL_318[2];
  assign _EVAL_454 = _EVAL_1340 ^ _EVAL_2851;
  assign _EVAL_1305 = _EVAL_3232[8:7];
  assign _EVAL_401 = _EVAL_1305 == 2'h3;
  assign _EVAL_4653 = _EVAL_3232[6];
  assign _EVAL_4851 = _EVAL_401 & _EVAL_4653;
  assign _EVAL_1236 = _EVAL_4653 == 1'h0;
  assign _EVAL_4931 = _EVAL_401 & _EVAL_1236;
  assign _EVAL_753 = _EVAL_4851 | _EVAL_4931;
  assign _EVAL_1660 = _EVAL_3255 | _EVAL_3445;
  assign _EVAL_4465 = _EVAL_4788 & _EVAL_3299;
  assign _EVAL_2604 = _EVAL_4465 & _EVAL_4953;
  assign _EVAL_2415 = _EVAL_315 ? _EVAL_4527 : _EVAL_2283;
  assign _EVAL_3610 = _EVAL_5206 & 12'h444;
  assign _EVAL_1948 = _EVAL_3610 == 12'h40;
  assign _EVAL_1370 = _EVAL_5206 & 12'h412;
  assign _EVAL_2087 = _EVAL_1370 == 12'h412;
  assign _EVAL_2543 = _EVAL_1948 | _EVAL_2087;
  assign _EVAL_4926 = _EVAL_2415 & _EVAL_2543;
  assign _EVAL_3023 = csr__EVAL_123[4:0];
  assign _EVAL_1531 = _EVAL_3023 == 5'h0;
  assign _EVAL_2581 = _EVAL_1531 | _EVAL_174;
  assign _EVAL_2554 = _EVAL_3285 | _EVAL_4474;
  assign _EVAL_487 = _EVAL_5422 & _EVAL_3170;
  assign _EVAL_3325 = {{2'd0}, _EVAL_487};
  assign _EVAL_3931 = _EVAL_318 ^ _EVAL_3325;
  assign _EVAL_1794 = _EVAL_3931[0];
  assign _EVAL_595 = _EVAL_3931[2];
  assign _EVAL_2805 = _EVAL_1794 ^ _EVAL_595;
  assign _EVAL_687 = _EVAL_595 == 1'h0;
  assign _EVAL_843 = _EVAL_3931[1];
  assign _EVAL_3502 = _EVAL_843 == 1'h0;
  assign _EVAL_4825 = _EVAL_687 & _EVAL_3502;
  assign _EVAL_543 = _EVAL_1794 ^ _EVAL_4825;
  assign _EVAL_788 = _EVAL_2434 ? _EVAL_543 : _EVAL_1794;
  assign _EVAL_1508 = _EVAL_3979 ? _EVAL_2805 : _EVAL_788;
  assign _EVAL_1548 = _EVAL_2554 | _EVAL_1508;
  assign _EVAL_5221 = _EVAL_2581 | _EVAL_1548;
  assign _EVAL_888 = _EVAL_5221 == 1'h0;
  assign _EVAL_5060 = _EVAL_2661 ^ _EVAL_2787;
  assign _EVAL_4905 = divider__EVAL_2 & _EVAL_296;
  assign _EVAL_2088 = _EVAL_3997 == 1'h0;
  assign _EVAL_3305 = _EVAL_2118 & _EVAL_2088;
  assign _EVAL_1074 = _EVAL_3305 == 1'h0;
  assign _EVAL_3076 = _EVAL_838 & _EVAL_1074;
  assign _EVAL_4146 = _EVAL_3076 ? _EVAL_1379 : 3'h2;
  assign _EVAL_3334 = _EVAL_487 & _EVAL_1074;
  assign _EVAL_1953 = {{2'd0}, _EVAL_3334};
  assign _EVAL_2536 = _EVAL_4146 ^ _EVAL_1953;
  assign _EVAL_4532 = _EVAL_2536[0];
  assign _EVAL_2555 = _EVAL_2536[2];
  assign _EVAL_4670 = _EVAL_4532 ^ _EVAL_2555;
  assign _EVAL_5188 = _EVAL_2679[0];
  assign _EVAL_1282 = _EVAL_2679[1];
  assign _EVAL_4575 = _EVAL_1282 == 1'h0;
  assign _EVAL_2722 = _EVAL_1568 & _EVAL_4575;
  assign _EVAL_2062 = _EVAL_5188 ^ _EVAL_2722;
  assign _EVAL_3975 = _EVAL_3401 == 1'h0;
  assign _EVAL_3984 = _EVAL_3975 | _EVAL_4596;
  assign _EVAL_5270 = _EVAL_5275 | _EVAL_5068;
  assign _EVAL_1470 = _EVAL_1277 & _EVAL_5270;
  assign _EVAL_541 = _EVAL_834 ? _EVAL_3958 : 1'h0;
  assign _EVAL_4345 = _EVAL_3218 ? _EVAL_402 : _EVAL_541;
  assign _EVAL_3382 = _EVAL_4025 ? _EVAL_4297 : _EVAL_4345;
  assign _EVAL_912 = _EVAL_1470 ? _EVAL_3216 : _EVAL_3382;
  assign _EVAL_4363 = _EVAL_4605 == 1'h0;
  assign _EVAL_883 = _EVAL_1536 & _EVAL_5031;
  assign _EVAL_3358 = _EVAL_779 == 1'h0;
  assign _EVAL_2187 = _EVAL_3440 & _EVAL_3358;
  assign _EVAL_2941 = _EVAL_2187 & _EVAL_4376;
  assign _EVAL_360 = _EVAL_4596 & _EVAL_2941;
  assign _EVAL_1210 = _EVAL_4007 & _EVAL_1849;
  assign _EVAL_2171 = _EVAL_4596 & _EVAL_1210;
  assign _EVAL_4143 = _EVAL_360 | _EVAL_2171;
  assign _EVAL_3369 = _EVAL_1460 & _EVAL_4143;
  assign _EVAL_3488 = _EVAL_4596 & _EVAL_1215;
  assign _EVAL_2589 = _EVAL_3488 | _EVAL_2171;
  assign _EVAL_846 = _EVAL_912 & _EVAL_2589;
  assign _EVAL_4077 = _EVAL_846 ? 4'h3 : 4'he;
  assign _EVAL_2375 = _EVAL_3369 ? 4'h3 : _EVAL_4077;
  assign _EVAL_4246 = _EVAL_4607[2:1];
  assign _EVAL_4860 = _EVAL_5188 ^ _EVAL_5127;
  assign _EVAL_1757 = _EVAL_1973 ? _EVAL_2062 : _EVAL_5188;
  assign _EVAL_4979 = _EVAL_1225 ? _EVAL_4860 : _EVAL_1757;
  assign _EVAL_2559 = _EVAL_240[1];
  assign _EVAL_2961 = _EVAL_2963 & _EVAL_1588;
  assign _EVAL_4378 = _EVAL_2961 & _EVAL_2379;
  assign _EVAL_3194 = _EVAL_2559 | _EVAL_4378;
  assign _EVAL_4379 = {{63'd0}, _EVAL_1535};
  assign _EVAL_3127 = _EVAL_4379 << _EVAL_2823;
  assign _EVAL_4149 = _EVAL_612 & _EVAL_4512;
  assign _EVAL_5121 = _EVAL_545 == 1'h0;
  assign _EVAL_3400 = {_EVAL_416,_EVAL_3688};
  assign _EVAL_2849 = _EVAL_3208 ? _EVAL_356 : _EVAL_4968;
  assign _EVAL_3829 = _EVAL_2400[5];
  assign _EVAL_2698 = _EVAL_3598[0];
  assign _EVAL_5416 = _EVAL_2698 == 1'h0;
  assign _EVAL_2870 = _EVAL_4706 == _EVAL_4460;
  assign _EVAL_4523 = _EVAL_1333 & _EVAL_2870;
  assign _EVAL_1493 = _EVAL_2506 & _EVAL_4523;
  assign _EVAL_1076 = _EVAL_4236 ? _EVAL_3923 : _EVAL_579;
  assign _EVAL_4482 = _EVAL_1493 ? _EVAL_4399 : _EVAL_1076;
  assign _EVAL_4444 = _EVAL_1206 ? _EVAL_4482 : _EVAL_2919;
  assign _EVAL_955 = _EVAL_2145 ? _EVAL_4157 : _EVAL_4444;
  assign _EVAL_4906 = fpu__EVAL_26 == _EVAL_1480;
  assign _EVAL_1037 = _EVAL_1187 ? _EVAL_1453 : _EVAL_2974;
  assign _EVAL_3692 = _EVAL_1476 ? 2'h0 : 2'h2;
  assign _EVAL_509 = _EVAL_2329 ? _EVAL_1037 : {{1'd0}, _EVAL_3692};
  assign _EVAL_566 = _EVAL_315 ? _EVAL_2908 : _EVAL_5289;
  assign _EVAL_333 = _EVAL_566 | _EVAL_4926;
  assign _EVAL_4188 = _EVAL_333 == 1'h0;
  assign _EVAL_2909 = _EVAL_518 & _EVAL_4188;
  assign _EVAL_5400 = _EVAL_838 ? _EVAL_1379 : 3'h2;
  assign _EVAL_4837 = _EVAL_5400 ^ _EVAL_3325;
  assign _EVAL_4145 = _EVAL_4837[0];
  assign _EVAL_3685 = _EVAL_4837[2];
  assign _EVAL_4213 = _EVAL_3685 == 1'h0;
  assign _EVAL_5296 = _EVAL_4837[1];
  assign _EVAL_1438 = _EVAL_5296 == 1'h0;
  assign _EVAL_2396 = _EVAL_4213 & _EVAL_1438;
  assign _EVAL_1771 = _EVAL_4145 ^ _EVAL_2396;
  assign _EVAL_1637 = _EVAL_1913[32];
  assign _EVAL_3427 = $signed(_EVAL_618) < $signed(10'sh82);
  assign _EVAL_2470 = _EVAL_3427 ? 8'h0 : _EVAL_2577;
  assign _EVAL_4785 = _EVAL_753 ? 8'hff : 8'h0;
  assign _EVAL_5139 = _EVAL_2470 | _EVAL_4785;
  assign _EVAL_1043 = {1'h0,_EVAL_3258,_EVAL_2110};
  assign _EVAL_466 = _EVAL_1043[24:1];
  assign _EVAL_3770 = _EVAL_618[4:0];
  assign _EVAL_5343 = 5'h1 - _EVAL_3770;
  assign _EVAL_4501 = _EVAL_466 >> _EVAL_5343;
  assign _EVAL_2675 = _EVAL_4501[22:0];
  assign _EVAL_1796 = _EVAL_1043[22:0];
  assign _EVAL_1751 = _EVAL_4931 ? 23'h0 : _EVAL_1796;
  assign _EVAL_3899 = _EVAL_3427 ? _EVAL_2675 : _EVAL_1751;
  assign _EVAL_4035 = {_EVAL_1637,_EVAL_5139,_EVAL_3899};
  assign _EVAL_3791 = _EVAL_5099 == _EVAL_4400;
  assign _EVAL_1072 = _EVAL_4645 & _EVAL_3791;
  assign _EVAL_5357 = 1'h1;
  assign _EVAL_4094 = fpu__EVAL_26 == _EVAL_4400;
  assign _EVAL_1394 = _EVAL_1024[1:0];
  assign _EVAL_306 = _EVAL_1394 != 2'h0;
  assign _EVAL_2834 = _EVAL_854 & _EVAL_306;
  assign _EVAL_4830 = _EVAL_951 | _EVAL_1352;
  assign _EVAL_1151 = _EVAL_2834 == 1'h0;
  assign _EVAL_3861 = _EVAL_854 & _EVAL_1151;
  assign _EVAL_3018 = _EVAL_4830 | _EVAL_3861;
  assign _EVAL_4704 = _EVAL_3227 & _EVAL_3018;
  assign _EVAL_1289 = _EVAL_3194 | _EVAL_2327;
  assign _EVAL_2304 = csr__EVAL_80[1:0];
  assign _EVAL_1361 = _EVAL_1 & _EVAL_4368;
  assign _EVAL_4556 = _EVAL_653 & _EVAL_1361;
  assign _EVAL_2169 = _EVAL_653 & _EVAL_2508;
  assign _EVAL_3816 = _EVAL_315 ? _EVAL_4556 : _EVAL_2169;
  assign _EVAL_4108 = _EVAL_2118 & _EVAL_3816;
  assign _EVAL_1284 = _EVAL_315 ? _EVAL_4108 : _EVAL_4108;
  assign _EVAL_939 = _EVAL_1284 & _EVAL_824;
  assign _EVAL_4102 = _EVAL_315 ? _EVAL_3890 : _EVAL_3890;
  assign _EVAL_3469 = _EVAL_4102 & _EVAL_2479;
  assign _EVAL_3006 = _EVAL_939 | _EVAL_3469;
  assign _EVAL_3690 = _EVAL_2326 & _EVAL_5097;
  assign _EVAL_2887 = _EVAL_315 ? _EVAL_3690 : _EVAL_3690;
  assign _EVAL_4997 = _EVAL_2887 & _EVAL_1487;
  assign _EVAL_5096 = _EVAL_3006 | _EVAL_4997;
  assign _EVAL_2191 = _EVAL_1 & _EVAL_4970;
  assign _EVAL_999 = _EVAL_1724 & _EVAL_2191;
  assign _EVAL_3280 = _EVAL_1724 & _EVAL_1741;
  assign _EVAL_493 = _EVAL_315 ? _EVAL_999 : _EVAL_3280;
  assign _EVAL_3824 = _EVAL_3624 & _EVAL_493;
  assign _EVAL_3306 = _EVAL_315 ? _EVAL_3824 : _EVAL_3824;
  assign _EVAL_4940 = _EVAL_3306 & _EVAL_1206;
  assign _EVAL_5012 = _EVAL_5096 | _EVAL_4940;
  assign _EVAL_4296 = _EVAL_3299 & _EVAL_5012;
  assign _EVAL_328 = _EVAL_4296 | _EVAL_539;
  assign _EVAL_5280 = _EVAL_328 | _EVAL_1189;
  assign _EVAL_802 = _EVAL_5280 | _EVAL_2888;
  assign _EVAL_3098 = _EVAL_3896 ? _EVAL_2299 : _EVAL_802;
  assign _EVAL_2093 = _EVAL_1049[19:15];
  assign _EVAL_3320 = _EVAL_5114[19:15];
  assign _EVAL_2729 = _EVAL_2302[19:15];
  assign _EVAL_3067 = _EVAL_4329[19:15];
  assign _EVAL_1339 = _EVAL_1926 ? _EVAL_2729 : _EVAL_3067;
  assign _EVAL_4635 = _EVAL_2164 ? _EVAL_3320 : _EVAL_1339;
  assign _EVAL_5228 = _EVAL_4272 ? _EVAL_2093 : _EVAL_4635;
  assign _EVAL_3110 = _EVAL_5228;
  assign _EVAL_3489 = _EVAL_3361 & _EVAL_3319;
  assign _EVAL_684 = _EVAL_3736 | _EVAL_3489;
  assign _EVAL_4629 = _EVAL_4160 | _EVAL_3127;
  assign _EVAL_2223 = $signed(_EVAL_3400);
  assign _EVAL_1435 = _EVAL_2203 ? $signed(_EVAL_3911) : $signed(_EVAL_2223);
  assign _EVAL_4762 = csr__EVAL_70 | _EVAL_5226;
  assign _EVAL_2300 = _EVAL_4762 | _EVAL_3369;
  assign _EVAL_3537 = _EVAL_719 == 1'h0;
  assign _EVAL_1050 = _EVAL_4596 & _EVAL_4802;
  assign _EVAL_3483 = _EVAL_678 == 1'h0;
  assign _EVAL_1506 = _EVAL_1050 & _EVAL_3483;
  assign _EVAL_4950 = _EVAL_1506 ? 1'h1 : _EVAL_4842;
  assign _EVAL_5410 = _EVAL_1815 ? _EVAL_3537 : _EVAL_4950;
  assign _EVAL_5037 = _EVAL_1699 == 1'h0;
  assign _EVAL_288 = fpu__EVAL_29 == _EVAL_3711;
  assign _EVAL_3735 = _EVAL_4721 & _EVAL_3712;
  assign _EVAL_4508 = _EVAL_1803 ? _EVAL_1647 : _EVAL_3735;
  assign _EVAL_4740 = _EVAL_2273 & _EVAL_5082;
  assign _EVAL_2218 = fpu__EVAL_57 == _EVAL_4745;
  assign _EVAL_3429 = _EVAL_351 & _EVAL_2218;
  assign _EVAL_1820 = fpu__EVAL_25 == _EVAL_4745;
  assign _EVAL_3407 = _EVAL_1686 & _EVAL_1820;
  assign _EVAL_3560 = _EVAL_3407 ? fpu__EVAL_2 : _EVAL_4208;
  assign _EVAL_1148 = _EVAL_3429 ? fpu__EVAL_30 : _EVAL_3560;
  assign _EVAL_2570 = _EVAL_4740 ? fpu__EVAL_60 : _EVAL_1148;
  assign _EVAL_2590 = _EVAL_315 ? _EVAL_2986 : _EVAL_4874;
  assign _EVAL_4083 = _EVAL_2590 ? _EVAL_1572 : _EVAL_1223;
  assign _EVAL_1955 = _EVAL_3299 == 1'h0;
  assign _EVAL_4484 = _EVAL_2555 == 1'h0;
  assign _EVAL_3914 = _EVAL_2536[1];
  assign _EVAL_353 = _EVAL_3914 == 1'h0;
  assign _EVAL_921 = _EVAL_4484 & _EVAL_353;
  assign _EVAL_4010 = _EVAL_4532 ^ _EVAL_921;
  assign _EVAL_2086 = _EVAL_2434 ? _EVAL_4010 : _EVAL_4532;
  assign _EVAL_4667 = _EVAL_3979 ? _EVAL_4670 : _EVAL_2086;
  assign _EVAL_2181 = _EVAL_4667 ? 1'h0 : _EVAL_2118;
  assign _EVAL_4606 = _EVAL_4192[6:2];
  assign _EVAL_4703 = _EVAL_649[4:2];
  assign _EVAL_4080 = _EVAL_4703 == 3'h7;
  assign _EVAL_5235 = _EVAL_359 == 2'h0;
  assign _EVAL_3793 = _EVAL_4240 & _EVAL_4608;
  assign _EVAL_2426 = _EVAL_5252 & _EVAL_1011;
  assign _EVAL_4589 = _EVAL_2426 ? _EVAL_3187 : _EVAL_5367;
  assign _EVAL_3848 = _EVAL_1770 ? _EVAL_4863 : _EVAL_4589;
  assign _EVAL_2982 = _EVAL_3790 == 2'h1;
  assign _EVAL_915 = _EVAL_2145 & _EVAL_2982;
  assign _EVAL_1760 = _EVAL_3074 ? _EVAL_2100 : 1'h0;
  assign _EVAL_433 = _EVAL_609 ? _EVAL_1817 : _EVAL_1760;
  assign _EVAL_3307 = _EVAL_635 ? _EVAL_2967 : _EVAL_433;
  assign _EVAL_4519 = _EVAL_4908 ? _EVAL_5154 : _EVAL_3307;
  assign _EVAL_4219 = _EVAL_2806 ? 3'h7 : 3'h5;
  assign _EVAL_3569 = _EVAL_1127 ? 4'hd : {{1'd0}, _EVAL_4219};
  assign _EVAL_3418 = _EVAL_525 ? 4'hf : _EVAL_3569;
  assign _EVAL_1080 = _EVAL_5037 | _EVAL_1250;
  assign _EVAL_5029 = _EVAL_4203 ? 4'h6 : 4'h8;
  assign _EVAL_378 = _EVAL_2060 ? {{1'd0}, _EVAL_4439} : _EVAL_5029;
  assign _EVAL_4385 = _EVAL_2603 ? _EVAL_378 : {{1'd0}, _EVAL_2157};
  assign _EVAL_4053 = {{28'd0}, _EVAL_4385};
  assign _EVAL_341 = _EVAL_5043 + _EVAL_4053;
  assign _EVAL_1026 = _EVAL_1080 ? _EVAL_341 : _EVAL_1104;
  assign _EVAL_4761 = {{19{_EVAL_2862[12]}},_EVAL_2862};
  assign _EVAL_4548 = $signed(_EVAL_4709) + $signed(_EVAL_4761);
  assign _EVAL_3024 = $unsigned(_EVAL_4548);
  assign _EVAL_3625 = _EVAL_3208 ? {{1'd0}, _EVAL_1026} : _EVAL_3024;
  assign _EVAL_5397 = _EVAL_3047 ? _EVAL_2799 : 32'h0;
  assign _EVAL_3342 = _EVAL_315 ? _EVAL_2827 : _EVAL_3753;
  assign _EVAL_4829 = _EVAL_315 ? _EVAL_589 : _EVAL_3231;
  assign _EVAL_1175 = _EVAL_325 ? _EVAL_4679 : _EVAL_2933;
  assign _EVAL_5000 = _EVAL_4829 ? _EVAL_1932 : _EVAL_1175;
  assign _EVAL_489 = _EVAL_3342 ? _EVAL_1572 : _EVAL_5000;
  assign _EVAL_4733 = _EVAL_3736 ? _EVAL_489 : 32'h0;
  assign _EVAL_5364 = _EVAL_5397 | _EVAL_4733;
  assign _EVAL_379 = _EVAL_2583 == 1'h0;
  assign _EVAL_2503 = _EVAL_379 & _EVAL_2326;
  assign _EVAL_2307 = _EVAL_2092 != _EVAL_3132;
  assign _EVAL_5105 = _EVAL_2503 & _EVAL_2307;
  assign _EVAL_832 = _EVAL_2886 == 1'h0;
  assign _EVAL_3236 = _EVAL_832 | csr__EVAL_39;
  assign _EVAL_2860 = _EVAL_915 & _EVAL_3236;
  assign _EVAL_1384 = _EVAL_5105 | _EVAL_2860;
  assign _EVAL_4308 = _EVAL_1384 ? 1'h1 : _EVAL_980;
  assign _EVAL_680 = _EVAL_1216 | _EVAL_4308;
  assign _EVAL_4725 = _EVAL_2583 & _EVAL_680;
  assign _EVAL_2107 = _EVAL_4725 ? _EVAL_2040 : _EVAL_506;
  assign _EVAL_1482 = _EVAL_5410 | _EVAL_2107;
  assign _EVAL_4462 = {_EVAL_416,_EVAL_3688,_EVAL_2059,_EVAL_2047};
  assign _EVAL_1787 = $signed(_EVAL_4462);
  assign _EVAL_5312 = _EVAL_47 == 1'h0;
  assign _EVAL_1779 = _EVAL_2273 & _EVAL_4094;
  assign _EVAL_4858 = _EVAL_2843 | _EVAL_233;
  assign _EVAL_1107 = $unsigned(_EVAL_1435);
  assign _EVAL_3877 = _EVAL_1107[11];
  assign _EVAL_3472 = _EVAL_3877 ? 20'hfffff : 20'h0;
  assign _EVAL_1121 = {_EVAL_3472,_EVAL_1107};
  assign _EVAL_2533 = _EVAL_4944 ? _EVAL_1121 : 32'h0;
  assign _EVAL_1852 = _EVAL_1508 | _EVAL_4560;
  assign _EVAL_5108 = _EVAL_55 & _EVAL_129;
  assign _EVAL_2820 = _EVAL_237 & _EVAL_254;
  assign _EVAL_573 = _EVAL_2084 ? 1'h0 : _EVAL_3896;
  assign _EVAL_4773 = _EVAL_573 < 1'h1;
  assign _EVAL_845 = _EVAL_2820 | _EVAL_4773;
  assign _EVAL_2800 = _EVAL_5108 & _EVAL_845;
  assign _EVAL_5272 = _EVAL_956 | _EVAL_2800;
  assign _EVAL_957 = _EVAL_802 == 1'h0;
  assign _EVAL_460 = _EVAL_4788 & _EVAL_957;
  assign _EVAL_4543 = _EVAL_956 | _EVAL_460;
  assign _EVAL_2486 = _EVAL_2851 == 1'h0;
  assign _EVAL_819 = _EVAL_318[1];
  assign _EVAL_4693 = _EVAL_819 == 1'h0;
  assign _EVAL_5249 = _EVAL_2486 & _EVAL_4693;
  assign _EVAL_1034 = _EVAL_5271 | _EVAL_1384;
  assign _EVAL_4638 = _EVAL_4788 & _EVAL_4296;
  assign _EVAL_4070 = {_EVAL_2604,_EVAL_95,1'h0,_EVAL_2001,_EVAL_4638};
  assign _EVAL_2613 = {_EVAL_4189,1'h0,_EVAL_4435,_EVAL_2004,_EVAL_1034,_EVAL_1852,_EVAL_4070};
  assign _EVAL_2645 = {{13'd0}, _EVAL_2613};
  assign _EVAL_437 = fpu__EVAL_29 == _EVAL_1480;
  assign _EVAL_1744 = _EVAL_4729 & _EVAL_437;
  assign _EVAL_3536 = _EVAL_1744 ? fpu__EVAL_21 : _EVAL_2741__EVAL_2748_data;
  assign _EVAL_2835 = fpu__EVAL_57 == _EVAL_3711;
  assign _EVAL_1321 = _EVAL_351 & _EVAL_2835;
  assign _EVAL_3375 = _EVAL_416[1];
  assign _EVAL_4062 = _EVAL_1287 & _EVAL_3375;
  assign _EVAL_4375 = _EVAL_4706 == _EVAL_2193;
  assign _EVAL_1613 = _EVAL_1333 & _EVAL_4375;
  assign _EVAL_2103 = _EVAL_2506 & _EVAL_1613;
  assign _EVAL_510 = _EVAL_3227 & _EVAL_5093;
  assign _EVAL_3805 = _EVAL_510 ? _EVAL_3923 : _EVAL_3848;
  assign _EVAL_4290 = _EVAL_2103 ? _EVAL_4399 : _EVAL_3805;
  assign _EVAL_1931 = {{31'd0}, _EVAL_127};
  assign _EVAL_535 = _EVAL_3333;
  assign _EVAL_2776 = _EVAL_3299 ? _EVAL_5340 : _EVAL_4415;
  assign _EVAL_3249 = _EVAL_5136 ? _EVAL_4319 : _EVAL_3196;
  assign _EVAL_3748 = _EVAL_3405 == 32'h2;
  assign _EVAL_1403 = _EVAL_3421 & _EVAL_3748;
  assign _EVAL_4022 = _EVAL_359 == 2'h1;
  assign _EVAL_4919 = _EVAL_779 | _EVAL_4022;
  assign _EVAL_4440 = _EVAL_1452[5];
  assign _EVAL_1786 = _EVAL_4919 & _EVAL_4440;
  assign _EVAL_5011 = _EVAL_3751 ? 4'h0 : _EVAL_2493;
  assign _EVAL_1163 = _EVAL_2963 & _EVAL_3153;
  assign _EVAL_1845 = _EVAL_1957 ? 2'h1 : 2'h2;
  assign _EVAL_4975 = _EVAL_663 ? 4'hc : {{2'd0}, _EVAL_1845};
  assign _EVAL_5211 = _EVAL_1593 ? 4'h3 : _EVAL_4975;
  assign _EVAL_1903 = _EVAL_3035 ? 4'he : _EVAL_5211;
  assign _EVAL_651 = _EVAL_3227 & _EVAL_951;
  assign _EVAL_4027 = _EVAL_3227 & _EVAL_1352;
  assign _EVAL_5100 = _EVAL_5031 & _EVAL_5104;
  assign _EVAL_3090 = $unsigned(_EVAL_1787);
  assign _EVAL_4224 = {_EVAL_3090, 12'h0};
  assign _EVAL_5073 = _EVAL_1597 ? _EVAL_4224 : 32'h0;
  assign _EVAL_831 = _EVAL_5073 | _EVAL_2533;
  assign _EVAL_2175 = _EVAL_2740 & _EVAL_1955;
  assign _EVAL_829 = _EVAL_2175 ? _EVAL_4083 : 32'h0;
  assign _EVAL_1938 = _EVAL_831 | _EVAL_829;
  assign _EVAL_4442 = _EVAL_4543 ? _EVAL_1938 : {{27'd0}, _EVAL_350};
  assign _EVAL_528 = _EVAL_2869 & _EVAL_1860;
  assign _EVAL_3708 = _EVAL_1049[24:20];
  assign _EVAL_2178 = _EVAL_2164 ? _EVAL_4536 : _EVAL_3321;
  assign _EVAL_3574 = _EVAL_4272 ? _EVAL_3708 : _EVAL_2178;
  assign _EVAL_4370 = _EVAL_3574;
  assign _EVAL_990 = _EVAL_315 ? _EVAL_260 : _EVAL_119;
  assign _EVAL_1095 = _EVAL_2400[6:2];
  assign _EVAL_4354 = _EVAL_2820 | _EVAL_766;
  assign _EVAL_3821 = _EVAL_5108 & _EVAL_4354;
  assign _EVAL_5253 = _EVAL_5022[2:1];
  assign _EVAL_4367 = _EVAL_5253 == 2'h1;
  assign _EVAL_5276 = _EVAL_2963 & _EVAL_2379;
  assign _EVAL_4994 = _EVAL_5099 == _EVAL_4745;
  assign _EVAL_392 = _EVAL_4645 & _EVAL_4994;
  assign _EVAL_1716 = _EVAL_5363[2];
  assign _EVAL_4553 = _EVAL_3742[2];
  assign _EVAL_5074 = _EVAL_1716 == _EVAL_4553;
  assign _EVAL_674 = _EVAL_2047[1:0];
  assign _EVAL_1826 = _EVAL_674 == 2'h1;
  assign _EVAL_1678 = _EVAL_2094 | _EVAL_1826;
  assign _EVAL_2962 = _EVAL_2239 | _EVAL_296;
  assign _EVAL_1433 = _EVAL_2962 | _EVAL_896;
  assign _EVAL_1733 = _EVAL_1433 | _EVAL_159;
  assign _EVAL_1169 = _EVAL_2424 & _EVAL_2840;
  assign _EVAL_4003 = _EVAL_890 & _EVAL_1169;
  assign _EVAL_3548 = _EVAL_4645 & _EVAL_4809;
  assign _EVAL_4251 = _EVAL_4437 ? _EVAL_4290 : 32'h0;
  assign _EVAL_516 = _EVAL_2304 == 2'h1;
  assign _EVAL_2098 = _EVAL_890 & _EVAL_3362;
  assign _EVAL_3425 = _EVAL_1803 ? 1'h0 : _EVAL_2098;
  assign _EVAL_3395 = _EVAL_4508 + _EVAL_3425;
  assign _EVAL_2572 = _EVAL_516 ? {{1'd0}, _EVAL_559} : _EVAL_3395;
  assign _EVAL_2832 = _EVAL_2841 == 13'h0;
  assign _EVAL_530 = {{6'd0}, _EVAL_5070};
  assign _EVAL_511 = _EVAL_379 & _EVAL_680;
  assign _EVAL_4269 = _EVAL_511 ? 1'h0 : _EVAL_2326;
  assign _EVAL_5207 = _EVAL_1815 ? 1'h1 : _EVAL_4269;
  assign _EVAL_4735 = _EVAL_2554 ? 1'h0 : _EVAL_5207;
  assign _EVAL_3775 = _EVAL_5136 ? _EVAL_4863 : _EVAL_3727;
  assign _EVAL_3169 = _EVAL_3775;
  assign _EVAL_4581 = _EVAL_5170[2];
  assign _EVAL_3865 = _EVAL_4581 == 1'h0;
  assign _EVAL_669 = _EVAL_2506 & _EVAL_4962;
  assign _EVAL_2563 = _EVAL_669 | _EVAL_528;
  assign _EVAL_1268 = fpu__EVAL_57 == _EVAL_1480;
  assign _EVAL_3987 = _EVAL_351 & _EVAL_1268;
  assign _EVAL_1875 = _EVAL_5344 | _EVAL_3176;
  assign _EVAL_2405 = _EVAL_2593 & _EVAL_3917;
  assign _EVAL_447 = _EVAL_1671 ? 3'h4 : 3'h6;
  assign _EVAL_1918 = _EVAL_1671 ? 4'h6 : 4'h8;
  assign _EVAL_4277 = _EVAL_3276 ? {{1'd0}, _EVAL_447} : _EVAL_1918;
  assign _EVAL_867 = _EVAL_1671 ? 3'h2 : 3'h4;
  assign _EVAL_1959 = _EVAL_4736 ? _EVAL_4277 : {{1'd0}, _EVAL_867};
  assign _EVAL_4142 = _EVAL_3588 & _EVAL_4692;
  assign _EVAL_928 = _EVAL_4142 == 1'h0;
  assign _EVAL_619 = _EVAL_3831 == 2'h1;
  assign _EVAL_2050 = _EVAL_2358 | _EVAL_619;
  assign _EVAL_5209 = _EVAL_2030[5];
  assign _EVAL_1423 = _EVAL_2050 & _EVAL_5209;
  assign _EVAL_4836 = _EVAL_2522[24:20];
  assign _EVAL_894 = _EVAL_961[24:20];
  assign _EVAL_919 = _EVAL_2180 ? _EVAL_5084 : _EVAL_894;
  assign _EVAL_2836 = _EVAL_544 ? _EVAL_4836 : _EVAL_919;
  assign _EVAL_3225 = _EVAL_757 ? _EVAL_3112 : _EVAL_2836;
  assign _EVAL_908 = _EVAL_2059 != 5'h0;
  assign _EVAL_456 = _EVAL_1335 == 2'h3;
  assign _EVAL_3477 = _EVAL_1248 ? _EVAL_1431 : 32'h0;
  assign _EVAL_383 = _EVAL_1780 & _EVAL_5031;
  assign _EVAL_4343 = _EVAL_5170[0];
  assign _EVAL_931 = _EVAL_3587 | _EVAL_159;
  assign _EVAL_2384 = _EVAL_3688 != 5'h0;
  assign _EVAL_4063 = {_EVAL_2384,_EVAL_908};
  assign _EVAL_1201 = _EVAL_5363 & 5'h1b;
  assign _EVAL_301 = 5'h1 == _EVAL_1201;
  assign _EVAL_4148 = _EVAL_301 == 1'h0;
  assign _EVAL_365 = _EVAL_1815 ? 1'h0 : _EVAL_639;
  assign _EVAL_2658 = _EVAL_2231 ? _EVAL_2299 : _EVAL_802;
  assign _EVAL_4759 = _EVAL_612 & _EVAL_4844;
  assign _EVAL_3518 = _EVAL_150 == 1'h0;
  assign _EVAL_3925 = _EVAL_60 & _EVAL_3518;
  assign _EVAL_2297 = _EVAL_3925;
  assign _EVAL_859 = _EVAL_951 == 1'h0;
  assign _EVAL_1939 = _EVAL_4519 & _EVAL_4143;
  assign _EVAL_1174 = _EVAL_990 ? 1'h1 : _EVAL_3088;
  assign _EVAL_1186 = _EVAL_4729 & _EVAL_288;
  assign _EVAL_339 = _EVAL_5323 & _EVAL_530;
  assign _EVAL_1130 = _EVAL_931 | _EVAL_669;
  assign _EVAL_1574 = {1'h0,_EVAL_4399};
  assign _EVAL_2772 = _EVAL_1574[31:0];
  assign _EVAL_5285 = _EVAL_2922 & _EVAL_5167;
  assign _EVAL_673 = _EVAL_2273 & _EVAL_4906;
  assign _EVAL_439 = fpu__EVAL_25 == _EVAL_1480;
  assign _EVAL_1835 = _EVAL_1686 & _EVAL_439;
  assign _EVAL_1773 = _EVAL_1835 ? fpu__EVAL_2 : _EVAL_3536;
  assign _EVAL_3122 = _EVAL_3987 ? fpu__EVAL_30 : _EVAL_1773;
  assign _EVAL_4758 = _EVAL_673 ? fpu__EVAL_60 : _EVAL_3122;
  assign _EVAL_1876 = fpu__EVAL_57 == _EVAL_4400;
  assign _EVAL_5051 = _EVAL_351 & _EVAL_1876;
  assign _EVAL_633 = fpu__EVAL_25 == _EVAL_3711;
  assign _EVAL_767 = _EVAL_1686 & _EVAL_633;
  assign _EVAL_3706 = _EVAL_3752[0];
  assign _EVAL_4883 = _EVAL_4988 & _EVAL_5201;
  assign _EVAL_4636 = _EVAL_4080 & _EVAL_5260;
  assign _EVAL_1652 = _EVAL_63;
  assign _EVAL_1732 = _EVAL_4382 & _EVAL_164;
  assign _EVAL_3621 = _EVAL_4145 ^ _EVAL_3685;
  assign _EVAL_4567 = _EVAL_365 == 1'h0;
  assign _EVAL_2548 = _EVAL_3971 & _EVAL_215;
  assign _EVAL_3994 = _EVAL_63;
  assign _EVAL_4732 = _EVAL_1083 & _EVAL_340;
  assign _EVAL_3045 = _EVAL_4732 | _EVAL_922;
  assign _EVAL_5057 = _EVAL_4636 == 1'h0;
  assign _EVAL_4402 = _EVAL_3165 == 1'h0;
  assign _EVAL_2494 = _EVAL_545 & _EVAL_4402;
  assign _EVAL_4355 = _EVAL_5312 & _EVAL_2494;
  assign _EVAL_1028 = _EVAL_3624 ? _EVAL_955 : {{27'd0}, _EVAL_2683};
  assign _EVAL_2296 = {{63'd0}, _EVAL_2869};
  assign _EVAL_5089 = _EVAL_2296 << _EVAL_111;
  assign _EVAL_3272 = ~ _EVAL_5089;
  assign _EVAL_2556 = _EVAL_2300 | _EVAL_846;
  assign _EVAL_789 = _EVAL_2556 | _EVAL_1939;
  assign _EVAL_515 = _EVAL_4025 ? _EVAL_2967 : _EVAL_1967;
  assign _EVAL_2537 = _EVAL_1470 ? _EVAL_5154 : _EVAL_515;
  assign _EVAL_1070 = _EVAL_2537 & _EVAL_2589;
  assign _EVAL_874 = _EVAL_789 | _EVAL_1070;
  assign _EVAL_3365 = _EVAL_1482 | _EVAL_874;
  assign _EVAL_2325 = _EVAL_1186 ? fpu__EVAL_21 : _EVAL_2741__EVAL_2750_data;
  assign _EVAL_4731 = _EVAL_3694 == 1'h0;
  assign _EVAL_5268 = _EVAL_649[2];
  assign _EVAL_3453 = _EVAL_4704 & _EVAL_4405;
  assign _EVAL_4173 = _EVAL_1749 | _EVAL_301;
  assign _EVAL_3041 = _EVAL_3453 & _EVAL_4173;
  assign _EVAL_4452 = _EVAL_1749 & _EVAL_5074;
  assign _EVAL_722 = {{29'd0}, _EVAL_509};
  assign _EVAL_4059 = _EVAL_1733 | _EVAL_1732;
  assign _EVAL_1099 = _EVAL_1597 | _EVAL_3299;
  assign _EVAL_3906 = _EVAL_3208 ? _EVAL_2399 : _EVAL_2371;
  assign _EVAL_2699 = 1'h1;
  assign _EVAL_3769 = _EVAL_111[4:0];
  assign _EVAL_2631 = _EVAL_3769 != 5'h0;
  assign _EVAL_4640 = _EVAL_3360 ? _EVAL_5363 : 5'h0;
  assign _EVAL_4457 = {{27'd0}, _EVAL_4640};
  assign _EVAL_3785 = _EVAL_2576 ? 20'hfffff : 20'h0;
  assign _EVAL_3354 = {_EVAL_3785,_EVAL_3570};
  assign _EVAL_1680 = _EVAL_4698 ? _EVAL_3354 : 32'h0;
  assign _EVAL_3822 = _EVAL_1680 | _EVAL_4251;
  assign _EVAL_1468 = _EVAL_3045 ? 32'h0 : _EVAL_3822;
  assign _EVAL_693 = _EVAL_1558 ? _EVAL_1468 : {{27'd0}, _EVAL_1415};
  assign _EVAL_3338 = _EVAL_1130 | _EVAL_4347;
  assign _EVAL_4336 = _EVAL_2506 & _EVAL_4914;
  assign _EVAL_3241 = _EVAL_4336 == 1'h0;
  assign _EVAL_1838 = _EVAL_1122 & _EVAL_653;
  assign _EVAL_1709 = 64'h0 << _EVAL_25;
  assign _EVAL_4750 = 64'h1 | _EVAL_1709;
  assign _EVAL_2630 = ~ _EVAL_4750;
  assign _EVAL_3104 = _EVAL_4629 & _EVAL_2630;
  assign _EVAL_2504 = _EVAL_3104 & _EVAL_3272;
  assign _EVAL_3003 = _EVAL_3538 & _EVAL_2864;
  assign _EVAL_3559 = _EVAL_5170[1];
  assign _EVAL_4204 = _EVAL_3559 == 1'h0;
  assign _EVAL_2497 = _EVAL_3865 & _EVAL_4204;
  assign _EVAL_5077 = _EVAL_4595[2:0];
  assign _EVAL_4274 = _EVAL_3841 == 5'h3;
  assign _EVAL_3988 = _EVAL_4274 & _EVAL_3706;
  assign _EVAL_4443 = _EVAL_4721 & _EVAL_3988;
  assign _EVAL_1062 = _EVAL_3624 & _EVAL_2922;
  assign _EVAL_4945 = _EVAL_1335 == 2'h2;
  assign _EVAL_2161 = _EVAL_4945 ? {{1'd0}, _EVAL_1740} : _EVAL_5069;
  assign _EVAL_4804 = {_EVAL_3747,_EVAL_2579};
  assign _EVAL_5202 = _EVAL_444 ? 4'h4 : _EVAL_3418;
  assign _EVAL_4030 = _EVAL_3301 & _EVAL_2631;
  assign _EVAL_797 = _EVAL_531 ? _EVAL_4035 : _EVAL_4290;
  assign _EVAL_4404 = _EVAL_797[15:0];
  assign _EVAL_382 = {_EVAL_4404,_EVAL_4404};
  assign _EVAL_2322 = _EVAL_4022 ? _EVAL_382 : _EVAL_797;
  assign _EVAL_3211 = ~ _EVAL_1230;
  assign _EVAL_1748 = _EVAL_3211 | 32'h1;
  assign _EVAL_2621 = ~ _EVAL_1748;
  assign _EVAL_2056 = _EVAL_1253 ? _EVAL_2443 : _EVAL_490;
  assign _EVAL_5135 = _EVAL_4343 ^ _EVAL_4581;
  assign _EVAL_851 = _EVAL_4343 ^ _EVAL_2497;
  assign _EVAL_4676 = _EVAL_1973 ? _EVAL_851 : _EVAL_4343;
  assign _EVAL_4917 = _EVAL_1225 ? _EVAL_5135 : _EVAL_4676;
  assign _EVAL_3310 = _EVAL_2554 ? 1'h0 : _EVAL_2181;
  assign _EVAL_4871 = _EVAL_142 == 1'h0;
  assign _EVAL_1399 = _EVAL_4858 | _EVAL_4871;
  assign _EVAL_1465 = _EVAL_2767 | _EVAL_1965;
  assign _EVAL_904 = _EVAL_2047[2:1];
  assign _EVAL_882 = _EVAL_1253 | _EVAL_1647;
  assign _EVAL_5131 = _EVAL_882 | _EVAL_490;
  assign _EVAL_1614 = _EVAL_5131 ? 4'h0 : _EVAL_1959;
  assign _EVAL_2997 = {{28'd0}, _EVAL_1614};
  assign _EVAL_1782 = _EVAL_1660 & _EVAL_3829;
  assign _EVAL_4834 = _EVAL_1782 | _EVAL_4367;
  assign _EVAL_3181 = _EVAL_4883 & _EVAL_4834;
  assign _EVAL_4052 = _EVAL_4776 > 3'h0;
  assign _EVAL_2195 = _EVAL_2922 & _EVAL_4152;
  assign _EVAL_2132 = _EVAL_907 == 2'h1;
  assign _EVAL_2514 = _EVAL_1423 | _EVAL_2132;
  assign _EVAL_624 = _EVAL_1838 == 1'h0;
  assign _EVAL_2238 = _EVAL_624 & _EVAL_5121;
  assign _EVAL_2063 = _EVAL_3361 & _EVAL_5416;
  assign _EVAL_605 = _EVAL_1678 & _EVAL_996;
  assign _EVAL_5049 = _EVAL_904 == 2'h1;
  assign _EVAL_637 = _EVAL_605 | _EVAL_5049;
  assign _EVAL_4756 = _EVAL_2063 & _EVAL_637;
  assign _EVAL_586 = _EVAL_797[7:0];
  assign _EVAL_1338 = {_EVAL_586,_EVAL_586,_EVAL_586,_EVAL_586};
  assign _EVAL_1971 = _EVAL_3728 + _EVAL_2997;
  assign _EVAL_2584 = _EVAL_1511 ? {{1'd0}, _EVAL_1971} : _EVAL_3625;
  assign _EVAL_1790 = _EVAL_4595[3];
  assign _EVAL_2873 = _EVAL_1790 ? _EVAL_341 : _EVAL_5043;
  assign _EVAL_2386 = _EVAL_2873[31:3];
  assign _EVAL_2924 = _EVAL_2583 & _EVAL_3365;
  assign _EVAL_5145 = ~ _EVAL_270;
  assign _EVAL_3403 = _EVAL_5145 | 32'h1;
  assign _EVAL_994 = _EVAL_2304 == 2'h3;
  assign _EVAL_1328 = _EVAL_3009 & _EVAL_859;
  assign _EVAL_3603 = csr__EVAL_148 | _EVAL_87;
  assign _EVAL_4390 = _EVAL_3922 >= 3'h6;
  assign _EVAL_403 = _EVAL_4148 | _EVAL_4452;
  assign _EVAL_2863 = _EVAL_3338 | _EVAL_4216;
  assign _EVAL_5348 = _EVAL_5136 ? _EVAL_3196 : _EVAL_4319;
  assign _EVAL_2838 = _EVAL_5348;
  assign _EVAL_936 = _EVAL_1416 | _EVAL_1281;
  assign _EVAL_2355 = _EVAL_2506 | _EVAL_3227;
  assign _EVAL_4212 = fpu__EVAL_26 == _EVAL_3711;
  assign _EVAL_4590 = _EVAL_2304 == 2'h2;
  assign _EVAL_3106 = {{28'd0}, _EVAL_1903};
  assign _EVAL_4178 = {_EVAL_3812,_EVAL_1163,_EVAL_4225,_EVAL_4149,_EVAL_1034,_EVAL_1852,_EVAL_2117};
  assign _EVAL_2031 = {{13'd0}, _EVAL_4178};
  assign _EVAL_2446 = _EVAL_5323 & _EVAL_2031;
  assign _EVAL_723 = ~ _EVAL_3403;
  assign _EVAL_3016 = csr__EVAL_123;
  assign _EVAL_1822 = _EVAL_3016;
  assign _EVAL_1260 = _EVAL_416[6:2];
  assign _EVAL_2592 = _EVAL_1340 ^ _EVAL_5249;
  assign _EVAL_5227 = _EVAL_2434 ? _EVAL_2592 : _EVAL_1340;
  assign _EVAL_2455 = _EVAL_3432 + _EVAL_722;
  assign _EVAL_4669 = _EVAL_3208 ? _EVAL_3384 : _EVAL_4481;
  assign _EVAL_1605 = _EVAL_1149 & _EVAL_888;
  assign _EVAL_3108 = _EVAL_5136 ? _EVAL_3727 : _EVAL_4863;
  assign _EVAL_1166 = _EVAL_3108;
  assign _EVAL_2517 = _EVAL_21;
  assign _EVAL_3754 = _EVAL_4246 == 2'h1;
  assign _EVAL_4985 = _EVAL_5323 & _EVAL_701;
  assign _EVAL_4021 = _EVAL_2927 == 1'h0;
  assign _EVAL_4220 = _EVAL_266;
  assign _EVAL_2051 = _EVAL_4080 & _EVAL_5057;
  assign _EVAL_2890 = _EVAL_2051 & _EVAL_4872;
  assign _EVAL_1994 = _EVAL_3029 == 1'h0;
  assign _EVAL_1619 = _EVAL_1558 ? _EVAL_2199 : {{27'd0}, _EVAL_1827};
  assign _EVAL_777 = _EVAL_2853 ? _EVAL_4035 : _EVAL_1619;
  assign _EVAL_4576 = _EVAL_2326 ? _EVAL_777 : _EVAL_1619;
  assign _EVAL_4427 = _EVAL_1452[2];
  assign _EVAL_1902 = _EVAL_4427 == 1'h0;
  assign _EVAL_2068 = _EVAL_2890 & _EVAL_1902;
  assign _EVAL_3311 = _EVAL_4590 ? {{1'd0}, _EVAL_3637} : _EVAL_2572;
  assign _EVAL_443 = _EVAL_2273 & _EVAL_4212;
  assign _EVAL_2906 = _EVAL_3440 & _EVAL_5268;
  assign _EVAL_2281 = _EVAL_2906 & _EVAL_4301;
  assign _EVAL_3198 = _EVAL_1786 | _EVAL_3754;
  assign _EVAL_4038 = _EVAL_2281 & _EVAL_3198;
  assign _EVAL_3385 = _EVAL_3663 | _EVAL_4062;
  assign _EVAL_3381 = _EVAL_4543 ? _EVAL_5364 : {{27'd0}, _EVAL_3366};
  assign _EVAL_2305 = _EVAL_4539[2];
  assign _EVAL_3109 = {_EVAL_4962,_EVAL_4706};
  assign _EVAL_4764 = _EVAL_3984 | _EVAL_3045;
  assign _EVAL_758 = _EVAL_767 ? fpu__EVAL_2 : _EVAL_2325;
  assign _EVAL_4918 = _EVAL_1321 ? fpu__EVAL_30 : _EVAL_758;
  assign _EVAL_3855 = _EVAL_443 ? fpu__EVAL_60 : _EVAL_4918;
  assign _EVAL_4723 = _EVAL_3016;
  assign _EVAL_1583 = _EVAL_3979 ? _EVAL_454 : _EVAL_5227;
  assign _EVAL_5356 = _EVAL_2803 ? 4'h6 : _EVAL_5202;
  assign _EVAL_3383 = _EVAL_3413 ? 1'h1 : _EVAL_2244;
  assign _EVAL_3200 = _EVAL_1420 | _EVAL_3477;
  assign _EVAL_1007 = _EVAL_5276 ? _EVAL_3200 : {{27'd0}, _EVAL_483};
  assign _EVAL_4889 = _EVAL_98 ? _EVAL_121 : _EVAL_73;
  assign _EVAL_4806 = _EVAL_4003 & csr__EVAL_39;
  assign _EVAL_3115 = {_EVAL_1222,_EVAL_4291};
  assign _EVAL_1634 = _EVAL_2405 & _EVAL_2514;
  assign _EVAL_4131 = _EVAL_3538 & _EVAL_701;
  assign _EVAL_2245 = _EVAL_3208 ? _EVAL_1250 : _EVAL_3170;
  assign _EVAL_3803 = _EVAL_5323 & _EVAL_2645;
  assign _EVAL_661 = _EVAL_3538 & _EVAL_530;
  assign _EVAL_3473 = _EVAL_126;
  assign _EVAL_3247 = _EVAL_3249;
  assign _EVAL_4887 = {_EVAL_2386,_EVAL_5077};
  assign _EVAL_5004 = _EVAL_660 & _EVAL_2871;
  assign _EVAL_5362 = _EVAL_5136 ? _EVAL_3845 : _EVAL_2331;
  assign _EVAL_537 = _EVAL_5362;
  assign _EVAL_4004 = _EVAL_3538 & _EVAL_2645;
  assign _EVAL_1027 = _EVAL_267;
  assign _EVAL_4924 = _EVAL_3538 & _EVAL_2031;
  assign _EVAL_1325 = _EVAL_5276 ? _EVAL_2194 : {{27'd0}, _EVAL_498};
  assign _EVAL_2804 = _EVAL_3225;
  assign _EVAL_3138 = _EVAL_811 & _EVAL_3032;
  assign _EVAL_5269 = _EVAL_269;
  assign csr__EVAL_49 = _EVAL_456 ? 2'h0 : _EVAL_2161;
  assign _EVAL_136 = csr__EVAL_103;
  assign csr__EVAL_87 = _EVAL_2758 | _EVAL_4457;
  assign bullet_clock_gate_in = _EVAL_267;
  assign _EVAL_41 = _EVAL_1511 == 1'h0;
  assign divider__EVAL_5 = _EVAL_4135;
  assign _EVAL_28 = csr__EVAL_131;
  assign _EVAL_187 = csr__EVAL_64;
  assign fpu__EVAL_11 = _EVAL_3670;
  assign _EVAL_173 = csr__EVAL_15;
  assign _EVAL_178 = csr__EVAL_82;
  assign _EVAL_181 = csr__EVAL_33;
  assign _EVAL_238 = _EVAL_3208 ? _EVAL_4887 : _EVAL_2455;
  assign _EVAL_94 = _EVAL_930 ? _EVAL_4804 : 6'h0;
  assign _EVAL_144 = csr__EVAL_150;
  assign csr__EVAL_74 = _EVAL_4721 & _EVAL_4362;
  assign divider__EVAL_1 = _EVAL_3880;
  assign _EVAL_0 = csr__EVAL_67;
  assign _EVAL_67 = csr__EVAL_110;
  assign _EVAL_193 = _EVAL_4917 | _EVAL_1583;
  assign csr__EVAL_86 = _EVAL_127;
  assign _EVAL_253 = csr__EVAL_106;
  assign _EVAL_230 = csr__EVAL_37;
  assign _EVAL_75 = _EVAL_3208 ? _EVAL_3178 : _EVAL_3291;
  assign fpu__EVAL_6 = _EVAL_3548 ? _EVAL_1004 : _EVAL_4758;
  assign _EVAL_52 = csr__EVAL_5;
  assign _EVAL_243 = csr__EVAL_108;
  assign _EVAL_157 = csr__EVAL_57;
  assign divider__EVAL_9 = _EVAL_569 | _EVAL_3138;
  assign _EVAL_218 = _EVAL_3208 ? _EVAL_1469 : _EVAL_5039;
  assign _EVAL_189 = csr__EVAL_145;
  assign _EVAL_17 = csr__EVAL_29;
  assign _EVAL_120 = csr__EVAL_161;
  assign _EVAL_275 = _EVAL_3208 ? _EVAL_3645 : _EVAL_5213;
  assign m__EVAL_0 = _EVAL_1994 ? 32'h0 : divider__EVAL_6;
  assign _EVAL_139 = csr__EVAL_56;
  assign _EVAL_10 = csr__EVAL_158;
  assign _EVAL_177 = _EVAL_1511 == 1'h0;
  assign _EVAL_93 = _EVAL_3208 ? _EVAL_706 : _EVAL_3934;
  assign _EVAL_257 = csr__EVAL_16;
  assign _EVAL_211 = csr__EVAL_55;
  assign _EVAL_60 = _EVAL_856 | _EVAL_150;
  assign _EVAL_209 = _EVAL_1104;
  assign _EVAL_195 = csr__EVAL_166;
  assign _EVAL_271 = csr__EVAL_104;
  assign _EVAL_124 = csr__EVAL_28;
  assign csr__EVAL_53 = bullet_clock_gate_out;
  assign fpu__EVAL_36 = _EVAL_2573;
  assign _EVAL_62 = _EVAL_5199[32:1];
  assign _EVAL_143 = csr__EVAL_45;
  assign csr__EVAL_23 = {_EVAL_1328,_EVAL_1972};
  assign _EVAL_279 = csr__EVAL_32;
  assign divider__EVAL_2 = _EVAL_3793 & _EVAL_4692;
  assign _EVAL_244 = _EVAL_3208 ? _EVAL_1000 : _EVAL_366;
  assign _EVAL_245 = 1'h0;
  assign csr__EVAL_117 = _EVAL_1403 ? _EVAL_4256 : _EVAL_2711;
  assign _EVAL_79 = _EVAL_883 & _EVAL_4819;
  assign _EVAL_3 = csr__EVAL_129;
  assign _EVAL_199 = csr__EVAL_96;
  assign _EVAL_112 = csr__EVAL_157;
  assign _EVAL_5 = 32'h0;
  assign fpu__EVAL_27 = _EVAL_1206 ? _EVAL_4482 : _EVAL_2919;
  assign _EVAL_83 = csr__EVAL_17;
  assign _EVAL_269 = _EVAL_5136 ? _EVAL_3025 : _EVAL_2656;
  assign _EVAL_240 = csr__EVAL_51;
  assign m__EVAL_5 = bullet_clock_gate_out;
  assign fpu__EVAL_38 = _EVAL_1491;
  assign _EVAL_109 = _EVAL_2305 == 1'h0;
  assign _EVAL_21 = _EVAL_5136 ? _EVAL_2656 : _EVAL_3025;
  assign _EVAL_155 = csr__EVAL_39;
  assign _EVAL_231 = csr__EVAL_133;
  assign csr__EVAL_6 = _EVAL_4;
  assign _EVAL_113 = csr__EVAL_19;
  assign _EVAL_74 = csr__EVAL_141;
  assign _EVAL_13 = _EVAL_3208 ? _EVAL_2587 : _EVAL_4088;
  assign _EVAL_38 = _EVAL_3077;
  assign _EVAL_53 = csr__EVAL_10;
  assign _EVAL_70 = csr__EVAL_128;
  assign _EVAL_273 = csr__EVAL_160;
  assign fpu_clock_gate_in = _EVAL_267;
  assign _EVAL_123 = _EVAL_4052 | _EVAL_49;
  assign _EVAL_266 = _EVAL_5136 ? _EVAL_4600 : _EVAL_3142;
  assign csr__EVAL_41 = _EVAL_994 ? 2'h0 : _EVAL_3311;
  assign _EVAL_125 = csr__EVAL_98;
  assign _EVAL_65 = _EVAL_1896;
  assign _EVAL_50 = _EVAL_4788 & _EVAL_3299;
  assign _EVAL_101 = csr__EVAL_3;
  assign fpu__EVAL_28 = _EVAL_2495;
  assign _EVAL_197 = csr__EVAL_7;
  assign _EVAL_8 = csr__EVAL_62;
  assign _EVAL_161 = csr__EVAL_159;
  assign _EVAL_89 = csr__EVAL_66;
  assign fpu__EVAL_1 = _EVAL_890 == 1'h0;
  assign _EVAL_150 = _EVAL_2927 & _EVAL_1647;
  assign _EVAL_201 = _EVAL_2245 == 1'h0;
  assign fpu__EVAL = fpu_clock_gate_out;
  assign _EVAL_192 = _EVAL_3208 | _EVAL_838;
  assign _EVAL_9 = csr__EVAL_126;
  assign m__EVAL_3 = divider__EVAL_4;
  assign fpu__EVAL_58 = _EVAL_5095;
  assign fpu__EVAL_5 = _EVAL_4530;
  assign fpu__EVAL_32 = _EVAL_392 ? _EVAL_1004 : _EVAL_2570;
  assign _EVAL_99 = _EVAL_1511 ? _EVAL_3270 : _EVAL_2849;
  assign _EVAL_254 = _EVAL_2658 == 1'h0;
  assign fpu__EVAL_31 = _EVAL_4390 ? csr__EVAL_99 : _EVAL_3922;
  assign m__EVAL_4 = _EVAL_1994 ? 32'h0 : divider__EVAL_1;
  assign _EVAL_258 = _EVAL_3208 ? _EVAL_1250 : _EVAL_3170;
  assign _EVAL_152 = csr__EVAL_93;
  assign _EVAL_129 = _EVAL_3098 == 1'h0;
  assign divider__EVAL_7 = bullet_clock_gate_out;
  assign _EVAL_167 = _EVAL_1225 ? _EVAL_5060 : _EVAL_1238;
  assign fpu_clock_gate_en = _EVAL_896;
  assign _EVAL_166 = csr__EVAL_167;
  assign divider__EVAL_10 = _EVAL_63;
  assign _EVAL_256 = csr__EVAL_121;
  assign csr__EVAL_165 = _EVAL_134;
  assign csr__EVAL_155 = _EVAL_3565 & _EVAL_4583;
  assign _EVAL_117 = _EVAL_1511 & _EVAL_3393;
  assign _EVAL_114 = _EVAL_3208 ? _EVAL_5025 : _EVAL_3730;
  assign _EVAL_248 = _EVAL_3573;
  assign _EVAL_130 = csr__EVAL_125;
  assign _EVAL_37 = csr__EVAL_156;
  assign csr__EVAL_1 = _EVAL_3579[1:0];
  assign m__EVAL_1 = _EVAL_4240 & _EVAL_3029;
  assign divider__EVAL_4 = {{1'd0}, _EVAL_1379};
  assign _EVAL_27 = csr__EVAL_59;
  assign _EVAL_223 = csr__EVAL_13;
  assign _EVAL_162 = csr__EVAL_132;
  assign _EVAL_219 = csr__EVAL_34;
  assign _EVAL_12 = csr__EVAL_153;
  assign _EVAL_145 = csr__EVAL_97;
  assign _EVAL_194 = csr__EVAL_113;
  assign csr__EVAL_146 = _EVAL_63;
  assign _EVAL_128 = csr__EVAL_152;
  assign _EVAL_11 = csr__EVAL_151;
  assign _EVAL_30 = csr__EVAL_20;
  assign csr__EVAL_102 = _EVAL_4218;
  assign _EVAL_100 = csr__EVAL_39;
  assign _EVAL_49 = _EVAL_4021 & _EVAL_1647;
  assign _EVAL_241 = csr__EVAL_35;
  assign _EVAL_14 = csr__EVAL_100;
  assign _EVAL_221 = csr__EVAL_31;
  assign _EVAL_118 = _EVAL_2118 & _EVAL_2494;
  assign _EVAL_210 = csr__EVAL_11;
  assign bullet_clock_gate_en = _EVAL_3448 | _EVAL_1732;
  assign _EVAL_7 = csr__EVAL_76;
  assign csr__EVAL_18 = {_EVAL_4889,_EVAL_4305};
  assign _EVAL_116 = _EVAL_3241 & _EVAL_3448;
  assign _EVAL_19 = csr__EVAL_65;
  assign _EVAL_185 = _EVAL_3208 ? _EVAL_3384 : _EVAL_4481;
  assign _EVAL_126 = _EVAL_5136 ? _EVAL_3142 : _EVAL_4600;
  assign _EVAL_151 = {_EVAL_2386,_EVAL_5077};
  assign _EVAL_262 = csr__EVAL_43;
  assign fpu__EVAL_15 = _EVAL_1854;
  assign divider__EVAL_6 = _EVAL_4322;
  assign fpu__EVAL_33 = _EVAL_5344;
  assign _EVAL_131 = csr__EVAL_9;
  assign _EVAL_42 = csr__EVAL_116;
  assign _EVAL_85 = _EVAL_5235 ? _EVAL_1338 : _EVAL_2322;
  assign _EVAL_200 = csr__EVAL_136;
  assign fpu__EVAL_50 = _EVAL_2030;
  assign csr__EVAL = _EVAL_5009;
  assign _EVAL_217 = csr__EVAL_12;
  assign _EVAL_61 = csr__EVAL_0;
  assign m__EVAL = _EVAL_63;
  assign _EVAL_77 = csr__EVAL_147;
  assign _EVAL_227 = csr__EVAL_60;
  assign fpu__EVAL_19 = _EVAL_3414 ? _EVAL_1004 : _EVAL_3855;
  assign _EVAL_264 = csr__EVAL_101;
  assign _EVAL_182 = _EVAL_79;
  assign _EVAL_239 = csr__EVAL_24;
  assign _EVAL_18 = _EVAL_1511 ? _EVAL_4550 : _EVAL_4669;
  assign divider__EVAL_0 = _EVAL_4759 == 1'h0;
  assign _EVAL_252 = csr__EVAL_112;
  assign _EVAL_69 = 1'h0;
  assign _EVAL_132 = csr__EVAL_76;
  assign _EVAL_46 = csr__EVAL_54;
  assign csr__EVAL_50 = _EVAL_267;
  assign _EVAL_228 = csr__EVAL_38;
  assign _EVAL_33 = _EVAL_3208 ? _EVAL_899 : _EVAL_2955;
  assign _EVAL_54 = _EVAL_1326 & _EVAL_403;
  assign _EVAL_149 = csr__EVAL_81;
  assign _EVAL_26 = csr__EVAL_79;
  assign _EVAL_229 = _EVAL_1511 ? _EVAL_2948 : _EVAL_3906;
  assign csr__EVAL_47 = fpu__EVAL_12;
  assign _EVAL_207 = csr__EVAL_26;
  assign _EVAL_140 = csr__EVAL_119;
  assign fpu__EVAL_49 = _EVAL_3624 & _EVAL_881;
  assign fpu__EVAL_46 = _EVAL_63;
  assign _EVAL_135 = csr__EVAL_21;
  assign _EVAL_56 = _EVAL_3208 ? _EVAL_2969 : _EVAL_4812;
  assign _EVAL_34 = _EVAL_2326 == 1'h0;
  assign csr__EVAL_109 = _EVAL_277;
  assign _EVAL_276 = _EVAL_1508 | _EVAL_3285;
  assign _EVAL_48 = csr__EVAL_58;
  assign _EVAL_72 = csr__EVAL_114;
  assign _EVAL_86 = csr__EVAL_137;
  assign _EVAL_88 = csr__EVAL_162;
  assign _EVAL_43 = _EVAL_1511 & _EVAL_2056;
  assign _EVAL_225 = _EVAL_4806 | _EVAL_4443;
  assign _EVAL_82 = csr__EVAL_107;
  assign _EVAL_66 = csr__EVAL_142;
  assign csr__EVAL_144 = fpu__EVAL_47;
  assign csr__EVAL_78 = _EVAL_3421 ? _EVAL_3405 : {{28'd0}, _EVAL_5356};
  assign _EVAL = csr__EVAL_154;
  assign _EVAL_103 = csr__EVAL_149;
  assign _EVAL_235 = csr__EVAL_164;
  assign _EVAL_160 = csr__EVAL_75;
  assign _EVAL_263 = _EVAL_2584[31:0];
  assign _EVAL_44 = csr__EVAL_2;
  assign csr__EVAL_77 = _EVAL_105;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    _EVAL_708[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    _EVAL_2741[initvar] = _RAND_1[32:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_284 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_313 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_332 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_350 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_356 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_366 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_375 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_380 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_396 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_483 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_490 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_494 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_498 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_531 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_545 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_601 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_612 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_623 = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_639 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_649 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_653 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_666 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_678 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_690 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_706 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_780 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_792 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_811 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_861 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_869 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_896 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_899 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_922 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_925 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_935 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_937 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_946 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_949 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_951 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_952 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_954 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_971 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_980 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_983 = _RAND_45[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_993 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_1000 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_1024 = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_1042 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1059 = _RAND_50[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1097 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1103 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1104 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1109 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1122 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1134 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1146 = _RAND_57[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1149 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1187 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1198 = _RAND_60[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1250 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1253 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1294 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1333 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1347 = _RAND_65[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1352 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1356 = _RAND_67[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1379 = _RAND_68[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1415 = _RAND_69[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1446 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1452 = _RAND_71[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1469 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1476 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1480 = _RAND_74[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1491 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1499 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1511 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1521 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1591 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1617 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1641 = _RAND_81[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1647 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1654 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1671 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1699 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1702 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1724 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {4{`RANDOM}};
  _EVAL_1727 = _RAND_88[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1737 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1740 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1795 = _RAND_91[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1818 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1827 = _RAND_93[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1828 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1854 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1895 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1896 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1908 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  _EVAL_1913 = _RAND_99[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1915 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1921 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1965 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1968 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1972 = _RAND_104[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_2030 = _RAND_105[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_2060 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_2089 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_2118 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_2138 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_2145 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_2172 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_2176 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_2193 = _RAND_113[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _EVAL_2219 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_2244 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_2258 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_2268 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {4{`RANDOM}};
  _EVAL_2278 = _RAND_118[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_2280 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_2282 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_2320 = _RAND_121[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_2326 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_2329 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_2331 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_2369 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_2371 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_2383 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_2397 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_2399 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_2409 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_2423 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_2424 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_2443 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_2495 = _RAND_134[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_2499 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_2506 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_2542 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_2573 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_2579 = _RAND_139[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_2583 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_2587 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _EVAL_2596 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2603 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _EVAL_2624 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _EVAL_2644 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2656 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _EVAL_2667 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _EVAL_2683 = _RAND_148[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _EVAL_2686 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _EVAL_2753 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _EVAL_2758 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _EVAL_2765 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _EVAL_2794 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _EVAL_2823 = _RAND_154[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _EVAL_2843 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _EVAL_2853 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _EVAL_2880 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _EVAL_2886 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _EVAL_2911 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _EVAL_2912 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _EVAL_2919 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _EVAL_2948 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _EVAL_2955 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _EVAL_2969 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _EVAL_2989 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _EVAL_3000 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {4{`RANDOM}};
  _EVAL_3019 = _RAND_167[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _EVAL_3025 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _EVAL_3029 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _EVAL_3039 = _RAND_170[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _EVAL_3053 = _RAND_171[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _EVAL_3064 = _RAND_172[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _EVAL_3077 = _RAND_173[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _EVAL_3085 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _EVAL_3094 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _EVAL_3102 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _EVAL_3117 = _RAND_177[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _EVAL_3132 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _EVAL_3134 = _RAND_179[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _EVAL_3142 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _EVAL_3165 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _EVAL_3170 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _EVAL_3176 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _EVAL_3178 = _RAND_184[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _EVAL_3196 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _EVAL_3204 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _EVAL_3217 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _EVAL_3227 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _EVAL_3229 = _RAND_189[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _EVAL_3240 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _EVAL_3270 = _RAND_191[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _EVAL_3276 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _EVAL_3291 = _RAND_193[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _EVAL_3295 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _EVAL_3302 = _RAND_195[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _EVAL_3309 = _RAND_196[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _EVAL_3355 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _EVAL_3362 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _EVAL_3366 = _RAND_199[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _EVAL_3370 = _RAND_200[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {4{`RANDOM}};
  _EVAL_3384 = _RAND_201[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _EVAL_3386 = _RAND_202[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _EVAL_3391 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _EVAL_3393 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _EVAL_3401 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _EVAL_3404 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _EVAL_3405 = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _EVAL_3413 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _EVAL_3415 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _EVAL_3421 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _EVAL_3432 = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _EVAL_3448 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _EVAL_3476 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _EVAL_3481 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _EVAL_3494 = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _EVAL_3523 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _EVAL_3573 = _RAND_217[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _EVAL_3588 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _EVAL_3608 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _EVAL_3624 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _EVAL_3629 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _EVAL_3637 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _EVAL_3645 = _RAND_223[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _EVAL_3670 = _RAND_224[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _EVAL_3694 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _EVAL_3711 = _RAND_226[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _EVAL_3712 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _EVAL_3727 = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _EVAL_3728 = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _EVAL_3730 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _EVAL_3742 = _RAND_231[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _EVAL_3747 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _EVAL_3750 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _EVAL_3752 = _RAND_234[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _EVAL_3771 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _EVAL_3798 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _EVAL_3814 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _EVAL_3840 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _EVAL_3841 = _RAND_239[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _EVAL_3845 = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _EVAL_3851 = _RAND_241[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _EVAL_3858 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _EVAL_3880 = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _EVAL_3888 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _EVAL_3902 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _EVAL_3922 = _RAND_246[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _EVAL_3934 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _EVAL_3939 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _EVAL_3940 = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _EVAL_3974 = _RAND_250[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _EVAL_3986 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _EVAL_3997 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _EVAL_4000 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _EVAL_4014 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _EVAL_4019 = _RAND_255[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _EVAL_4043 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _EVAL_4064 = _RAND_257[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _EVAL_4088 = _RAND_258[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _EVAL_4092 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _EVAL_4095 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _EVAL_4115 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _EVAL_4135 = _RAND_262[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {4{`RANDOM}};
  _EVAL_4154 = _RAND_263[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _EVAL_4157 = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {2{`RANDOM}};
  _EVAL_4160 = _RAND_265[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _EVAL_4162 = _RAND_266[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _EVAL_4167 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _EVAL_4168 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _EVAL_4192 = _RAND_269[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _EVAL_4195 = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _EVAL_4201 = _RAND_271[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _EVAL_4203 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _EVAL_4218 = _RAND_273[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _EVAL_4240 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _EVAL_4299 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _EVAL_4319 = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _EVAL_4322 = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _EVAL_4360 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _EVAL_4362 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _EVAL_4373 = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _EVAL_4400 = _RAND_281[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _EVAL_4423 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _EVAL_4437 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _EVAL_4460 = _RAND_284[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _EVAL_4461 = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _EVAL_4468 = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {4{`RANDOM}};
  _EVAL_4481 = _RAND_287[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _EVAL_4512 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _EVAL_4530 = _RAND_289[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _EVAL_4531 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _EVAL_4535 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _EVAL_4539 = _RAND_292[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {4{`RANDOM}};
  _EVAL_4550 = _RAND_293[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _EVAL_4562 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _EVAL_4596 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _EVAL_4600 = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _EVAL_4607 = _RAND_297[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _EVAL_4614 = _RAND_298[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _EVAL_4620 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _EVAL_4632 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _EVAL_4633 = _RAND_301[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _EVAL_4649 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _EVAL_4656 = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _EVAL_4679 = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _EVAL_4684 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _EVAL_4692 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _EVAL_4698 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _EVAL_4706 = _RAND_308[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _EVAL_4715 = _RAND_309[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _EVAL_4736 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _EVAL_4745 = _RAND_311[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _EVAL_4748 = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _EVAL_4790 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _EVAL_4796 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _EVAL_4805 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _EVAL_4812 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _EVAL_4819 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _EVAL_4842 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _EVAL_4844 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _EVAL_4863 = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {4{`RANDOM}};
  _EVAL_4915 = _RAND_321[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _EVAL_4927 = _RAND_322[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _EVAL_4936 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _EVAL_4939 = _RAND_324[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _EVAL_4947 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _EVAL_4962 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _EVAL_4968 = _RAND_327[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _EVAL_5009 = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _EVAL_5017 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _EVAL_5025 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _EVAL_5039 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _EVAL_5043 = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _EVAL_5052 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _EVAL_5095 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _EVAL_5099 = _RAND_335[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _EVAL_5178 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _EVAL_5213 = _RAND_337[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _EVAL_5226 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _EVAL_5233 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _EVAL_5237 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _EVAL_5265 = _RAND_341[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _EVAL_5335 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _EVAL_5344 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _EVAL_5363 = _RAND_344[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _EVAL_5367 = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _EVAL_5412 = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge bullet_clock_gate_out) begin
    if(_EVAL_708__EVAL_713_en & _EVAL_708__EVAL_713_mask) begin
      _EVAL_708[_EVAL_708__EVAL_713_addr] <= _EVAL_708__EVAL_713_data;
    end
    if(_EVAL_708__EVAL_714_en & _EVAL_708__EVAL_714_mask) begin
      _EVAL_708[_EVAL_708__EVAL_714_addr] <= _EVAL_708__EVAL_714_data;
    end
    if(_EVAL_708__EVAL_715_en & _EVAL_708__EVAL_715_mask) begin
      _EVAL_708[_EVAL_708__EVAL_715_addr] <= _EVAL_708__EVAL_715_data;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_284 <= _EVAL_39;
        end else begin
          _EVAL_284 <= _EVAL_148;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_284 <= _EVAL_148;
        end else begin
          _EVAL_284 <= _EVAL_39;
        end
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_1099) begin
        _EVAL_313 <= 3'h0;
      end else begin
        if (_EVAL_315) begin
          _EVAL_313 <= _EVAL_153;
        end else begin
          _EVAL_313 <= _EVAL_84;
        end
      end
    end
    if (_EVAL_2869) begin
      _EVAL_332 <= _EVAL_4030;
    end else begin
      if (_EVAL_2506) begin
        _EVAL_332 <= _EVAL_1333;
      end
    end
    _EVAL_350 <= _EVAL_4442[4:0];
    if (_EVAL_3624) begin
      _EVAL_356 <= _EVAL_3302;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_366 <= _EVAL_76;
      end else begin
        _EVAL_366 <= _EVAL_224;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_3088) begin
        if (_EVAL_315) begin
          _EVAL_375 <= _EVAL_180;
        end else begin
          _EVAL_375 <= _EVAL_68;
        end
      end
    end
    if (_EVAL_3624) begin
      if (_EVAL_2145) begin
        _EVAL_380 <= 1'h0;
      end else begin
        _EVAL_380 <= _EVAL_2499;
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_396 <= _EVAL_106;
        end else begin
          _EVAL_396 <= _EVAL_71;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_396 <= _EVAL_71;
        end else begin
          _EVAL_396 <= _EVAL_106;
        end
      end
    end
    _EVAL_483 <= _EVAL_1007[4:0];
    if (_EVAL_2506) begin
      if (_EVAL_147) begin
        if (_EVAL_3995) begin
          _EVAL_490 <= 1'h1;
        end else begin
          _EVAL_490 <= _EVAL_2268;
        end
      end else begin
        _EVAL_490 <= _EVAL_2268;
      end
    end
    if (_EVAL_5276) begin
      _EVAL_494 <= _EVAL_1344;
    end
    _EVAL_498 <= _EVAL_1325[4:0];
    if (_EVAL_2118) begin
      _EVAL_531 <= _EVAL_2596;
    end
    if (_EVAL_4543) begin
      if (_EVAL_315) begin
        _EVAL_545 <= _EVAL_170;
      end else begin
        _EVAL_545 <= _EVAL_242;
      end
    end
    _EVAL_612 <= _EVAL_1281 & _EVAL_859;
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_623 <= _EVAL_180;
      end else begin
        _EVAL_623 <= _EVAL_68;
      end
    end
    if (_EVAL_2118) begin
      _EVAL_639 <= _EVAL_3997;
    end
    if (_EVAL_2118) begin
      _EVAL_649 <= _EVAL_4633;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_653 <= _EVAL_214;
        end else begin
          _EVAL_653 <= _EVAL_268;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_653 <= _EVAL_268;
        end else begin
          _EVAL_653 <= _EVAL_214;
        end
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_666 <= _EVAL_250;
        end else begin
          _EVAL_666 <= _EVAL_141;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_666 <= _EVAL_141;
        end else begin
          _EVAL_666 <= _EVAL_250;
        end
      end
    end
    _EVAL_678 <= _EVAL_47;
    if (_EVAL_2118) begin
      _EVAL_690 <= _EVAL_666;
    end
    if (_EVAL_3624) begin
      _EVAL_706 <= _EVAL_3217;
    end
    if (_EVAL_5276) begin
      if (_EVAL_4978) begin
        _EVAL_780 <= 3'h0;
      end else begin
        if (_EVAL_315) begin
          _EVAL_780 <= _EVAL_84;
        end else begin
          _EVAL_780 <= _EVAL_153;
        end
      end
    end
    if (_EVAL_4543) begin
      _EVAL_792 <= _EVAL_4944;
    end
    _EVAL_811 <= _EVAL_1591;
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_861 <= _EVAL_108;
      end else begin
        _EVAL_861 <= _EVAL_220;
      end
    end
    if (_EVAL_63) begin
      _EVAL_869 <= 1'h0;
    end else begin
      _EVAL_869 <= 1'h1;
    end
    if (_EVAL_3624) begin
      _EVAL_899 <= _EVAL_5335;
    end
    if (_EVAL_2118) begin
      _EVAL_922 <= _EVAL_1122;
    end
    _EVAL_925 <= csr__EVAL_39;
    if (_EVAL_4543) begin
      if (_EVAL_315) begin
        _EVAL_935 <= _EVAL_265;
      end else begin
        _EVAL_935 <= _EVAL_137;
      end
    end
    if (_EVAL_2118) begin
      _EVAL_937 <= _EVAL_3000;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_946 <= _EVAL_4047;
      end else begin
        _EVAL_946 <= _EVAL_469;
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_2740) begin
        if (_EVAL_2590) begin
          _EVAL_949 <= _EVAL_1572;
        end else begin
          if (_EVAL_4783) begin
            _EVAL_949 <= _EVAL_1932;
          end else begin
            if (_EVAL_1052) begin
              _EVAL_949 <= _EVAL_4679;
            end else begin
              if (_EVAL_2022) begin
                _EVAL_949 <= _EVAL_2919;
              end else begin
                if (_EVAL_2544) begin
                  if (_EVAL_2869) begin
                    _EVAL_949 <= _EVAL_234;
                  end else begin
                    if (_EVAL_1446) begin
                      _EVAL_949 <= _EVAL_110;
                    end else begin
                      _EVAL_949 <= _EVAL_1495;
                    end
                  end
                end else begin
                  if (_EVAL_1518) begin
                    if (_EVAL_854) begin
                      _EVAL_949 <= csr__EVAL_84;
                    end else begin
                      if (_EVAL_3568) begin
                        _EVAL_949 <= m__EVAL_2;
                      end else begin
                        _EVAL_949 <= _EVAL_3125;
                      end
                    end
                  end else begin
                    if (_EVAL_4073) begin
                      _EVAL_949 <= _EVAL_4863;
                    end else begin
                      if (_EVAL_3531) begin
                        if (_EVAL_2257) begin
                          _EVAL_949 <= divider__EVAL_8;
                        end else begin
                          if (_EVAL_3629) begin
                            _EVAL_949 <= fpu__EVAL_9;
                          end else begin
                            _EVAL_949 <= _EVAL_3727;
                          end
                        end
                      end else begin
                        if (_EVAL_315) begin
                          _EVAL_949 <= _EVAL_1214;
                        end else begin
                          _EVAL_949 <= _EVAL_4515;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_3624) begin
      if (_EVAL_4130) begin
        _EVAL_951 <= 1'h1;
      end else begin
        _EVAL_951 <= _EVAL_1097;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_3514) begin
        _EVAL_952 <= _EVAL_1572;
      end else begin
        if (_EVAL_2668) begin
          _EVAL_952 <= _EVAL_1932;
        end else begin
          if (_EVAL_2073) begin
            _EVAL_952 <= _EVAL_4679;
          end else begin
            if (_EVAL_4207) begin
              _EVAL_952 <= _EVAL_2919;
            end else begin
              if (_EVAL_391) begin
                if (_EVAL_2869) begin
                  _EVAL_952 <= _EVAL_234;
                end else begin
                  if (_EVAL_1446) begin
                    _EVAL_952 <= _EVAL_110;
                  end else begin
                    _EVAL_952 <= _EVAL_1495;
                  end
                end
              end else begin
                if (_EVAL_1129) begin
                  if (_EVAL_854) begin
                    _EVAL_952 <= csr__EVAL_84;
                  end else begin
                    if (_EVAL_3568) begin
                      _EVAL_952 <= m__EVAL_2;
                    end else begin
                      _EVAL_952 <= _EVAL_3125;
                    end
                  end
                end else begin
                  if (_EVAL_4046) begin
                    _EVAL_952 <= _EVAL_4863;
                  end else begin
                    if (_EVAL_2464) begin
                      if (_EVAL_2257) begin
                        _EVAL_952 <= divider__EVAL_8;
                      end else begin
                        if (_EVAL_3629) begin
                          _EVAL_952 <= fpu__EVAL_9;
                        end else begin
                          _EVAL_952 <= _EVAL_3727;
                        end
                      end
                    end else begin
                      if (_EVAL_315) begin
                        _EVAL_952 <= _EVAL_1853;
                      end else begin
                        _EVAL_952 <= _EVAL_5376;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_2506) begin
      _EVAL_954 <= _EVAL_3404;
    end
    if (_EVAL_2118) begin
      _EVAL_971 <= _EVAL_2686;
    end
    if (_EVAL_4240) begin
      _EVAL_980 <= _EVAL_2280;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_983 <= _EVAL_73;
        end else begin
          _EVAL_983 <= _EVAL_121;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_983 <= _EVAL_121;
        end else begin
          _EVAL_983 <= _EVAL_73;
        end
      end
    end
    _EVAL_993 <= csr__EVAL_39;
    if (_EVAL_3624) begin
      _EVAL_1000 <= _EVAL_3204;
    end
    if (_EVAL_3624) begin
      _EVAL_1024 <= _EVAL_3922;
    end
    if (_EVAL_1558) begin
      _EVAL_1042 <= _EVAL_2542;
    end
    if (_EVAL_2118) begin
      _EVAL_1059 <= _EVAL_3134;
    end
    if (_EVAL_4240) begin
      if (_EVAL_4905) begin
        _EVAL_1097 <= 1'h1;
      end else begin
        _EVAL_1097 <= _EVAL_4936;
      end
    end
    _EVAL_1103 <= _EVAL_163;
    if (_EVAL_450) begin
      _EVAL_1104 <= _EVAL_4461;
    end
    if (_EVAL_4240) begin
      if (_EVAL_3750) begin
        _EVAL_1109 <= _EVAL_3880;
      end
    end
    if (_EVAL_4543) begin
      _EVAL_1122 <= _EVAL_3489;
    end
    _EVAL_1134 <= _EVAL_661 != 24'h0;
    if (_EVAL_3227) begin
      _EVAL_1146 <= _EVAL_4614;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_1187 <= _EVAL_106;
      end else begin
        _EVAL_1187 <= _EVAL_71;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_1198 <= _EVAL_2193;
    end
    if (_EVAL_3624) begin
      _EVAL_1250 <= _EVAL_2911;
    end
    if (_EVAL_2355) begin
      _EVAL_1253 <= _EVAL_4704;
    end
    if (_EVAL_2118) begin
      _EVAL_1294 <= _EVAL_4195;
    end
    if (_EVAL_1558) begin
      _EVAL_1333 <= _EVAL_4043;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_1347 <= _EVAL_180;
        end else begin
          _EVAL_1347 <= _EVAL_68;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_1347 <= _EVAL_68;
        end else begin
          _EVAL_1347 <= _EVAL_180;
        end
      end
    end
    if (_EVAL_3624) begin
      if (_EVAL_1384) begin
        _EVAL_1352 <= 1'h1;
      end else begin
        _EVAL_1352 <= _EVAL_980;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_1174) begin
        if (_EVAL_990) begin
          _EVAL_1356 <= _EVAL_1095;
        end else begin
          if (_EVAL_315) begin
            _EVAL_1356 <= _EVAL_180;
          end else begin
            _EVAL_1356 <= _EVAL_68;
          end
        end
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_1379 <= _EVAL_84;
      end else begin
        _EVAL_1379 <= _EVAL_153;
      end
    end
    _EVAL_1415 <= _EVAL_693[4:0];
    if (_EVAL_1558) begin
      _EVAL_1446 <= _EVAL_4596;
    end
    if (_EVAL_2118) begin
      _EVAL_1452 <= _EVAL_983;
    end
    if (_EVAL_3624) begin
      _EVAL_1469 <= _EVAL_2089;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_1476 <= _EVAL_186;
      end else begin
        _EVAL_1476 <= _EVAL_78;
      end
    end
    if (_EVAL_4240) begin
      if (_EVAL_2258) begin
        _EVAL_1480 <= _EVAL_3053;
      end
    end
    if (_EVAL_4240) begin
      _EVAL_1491 <= _EVAL_2244;
    end
    if (_EVAL_3227) begin
      _EVAL_1499 <= _EVAL_2603;
    end
    _EVAL_1511 <= _EVAL_995 | _EVAL_4139;
    if (_EVAL_2118) begin
      _EVAL_1521 <= _EVAL_396;
    end
    _EVAL_1591 <= _EVAL_1895;
    if (_EVAL_4543) begin
      _EVAL_1617 <= _EVAL_3047;
    end
    if (_EVAL_3624) begin
      _EVAL_1641 <= _EVAL_2495;
    end
    if (_EVAL_352) begin
      _EVAL_1647 <= 1'h1;
    end else begin
      _EVAL_1647 <= csr__EVAL_155;
    end
    if (_EVAL_4240) begin
      _EVAL_1654 <= _EVAL_3750;
    end
    if (_EVAL_2506) begin
      _EVAL_1671 <= _EVAL_1042;
    end
    if (_EVAL_3624) begin
      _EVAL_1699 <= _EVAL_2145;
    end
    _EVAL_1702 <= _EVAL_3803 != 24'h0;
    if (_EVAL_4240) begin
      _EVAL_1724 <= _EVAL_4692;
    end
    if (_EVAL_2118) begin
      _EVAL_1727 <= _EVAL_2278;
    end
    if (_EVAL_5276) begin
      _EVAL_1737 <= _EVAL_1248;
    end
    _EVAL_1740 <= _EVAL_4131 != 24'h0;
    if (_EVAL_4543) begin
      if (_EVAL_5340) begin
        if (_EVAL_315) begin
          _EVAL_1795 <= _EVAL_68;
        end else begin
          _EVAL_1795 <= _EVAL_180;
        end
      end
    end
    if (_EVAL_3624) begin
      _EVAL_1818 <= _EVAL_1634;
    end
    _EVAL_1827 <= _EVAL_4576[4:0];
    if (_EVAL_4240) begin
      _EVAL_1828 <= _EVAL_4812;
    end
    if (_EVAL_4240) begin
      _EVAL_1854 <= _EVAL_2258;
    end
    _EVAL_1895 <= divider__EVAL & divider__EVAL_2;
    if (_EVAL_4543) begin
      if (_EVAL_3385) begin
        _EVAL_1908 <= 1'h1;
      end else begin
        if (_EVAL_1002) begin
          _EVAL_1908 <= 1'h0;
        end
      end
    end else begin
      if (_EVAL_1002) begin
        _EVAL_1908 <= 1'h0;
      end
    end
    if (_EVAL_2118) begin
      if (_EVAL_1072) begin
        _EVAL_1913 <= _EVAL_1004;
      end else begin
        if (_EVAL_1779) begin
          _EVAL_1913 <= fpu__EVAL_60;
        end else begin
          if (_EVAL_5051) begin
            _EVAL_1913 <= fpu__EVAL_30;
          end else begin
            if (_EVAL_4011) begin
              _EVAL_1913 <= fpu__EVAL_2;
            end else begin
              if (_EVAL_4475) begin
                _EVAL_1913 <= fpu__EVAL_21;
              end else begin
                _EVAL_1913 <= _EVAL_2741__EVAL_2742_data;
              end
            end
          end
        end
      end
    end
    if (_EVAL_5276) begin
      _EVAL_1915 <= _EVAL_1736;
    end
    if (_EVAL_4543) begin
      _EVAL_1921 <= _EVAL_3106;
    end
    _EVAL_1965 <= _EVAL_147;
    if (_EVAL_5276) begin
      _EVAL_1968 <= _EVAL_4065;
    end
    if (_EVAL_1062) begin
      _EVAL_1972 <= _EVAL_3831;
    end
    if (_EVAL_4240) begin
      _EVAL_2030 <= _EVAL_4192;
    end
    if (_EVAL_3624) begin
      _EVAL_2060 <= _EVAL_5233;
    end
    if (_EVAL_4240) begin
      _EVAL_2089 <= _EVAL_5039;
    end
    if (_EVAL_1548) begin
      _EVAL_2118 <= 1'h0;
    end else begin
      _EVAL_2118 <= _EVAL_5272;
    end
    if (_EVAL_2118) begin
      _EVAL_2138 <= _EVAL_5032;
    end
    if (_EVAL_4240) begin
      _EVAL_2145 <= _EVAL_946;
    end
    if (_EVAL_4240) begin
      _EVAL_2172 <= _EVAL_4088;
    end
    if (_EVAL_1399) begin
      _EVAL_2176 <= 1'h0;
    end else begin
      if (_EVAL_1465) begin
        _EVAL_2176 <= 1'h1;
      end
    end
    if (_EVAL_2118) begin
      _EVAL_2193 <= _EVAL_1347;
    end
    if (_EVAL_3624) begin
      _EVAL_2219 <= _EVAL_1724;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_2244 <= _EVAL_188;
      end else begin
        _EVAL_2244 <= _EVAL_179;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_2258 <= _EVAL_39;
      end else begin
        _EVAL_2258 <= _EVAL_148;
      end
    end
    if (_EVAL_1558) begin
      if (_EVAL_1815) begin
        _EVAL_2268 <= _EVAL_3537;
      end else begin
        if (_EVAL_1506) begin
          _EVAL_2268 <= 1'h1;
        end else begin
          _EVAL_2268 <= _EVAL_4842;
        end
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_315) begin
        _EVAL_2278 <= _EVAL_23;
      end else begin
        _EVAL_2278 <= _EVAL_97;
      end
    end
    if (_EVAL_5276) begin
      if (csr__EVAL_105) begin
        _EVAL_2280 <= 1'h1;
      end else begin
        _EVAL_2280 <= _EVAL_2909;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_2282 <= _EVAL_4038;
    end
    if (_EVAL_5276) begin
      if (_EVAL_3671) begin
        if (_EVAL_315) begin
          _EVAL_2320 <= _EVAL_274;
        end else begin
          _EVAL_2320 <= _EVAL_154;
        end
      end
    end
    if (_EVAL_2554) begin
      _EVAL_2326 <= 1'h0;
    end else begin
      if (_EVAL_4667) begin
        _EVAL_2326 <= 1'h0;
      end else begin
        _EVAL_2326 <= _EVAL_2118;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_2329 <= _EVAL_115;
      end else begin
        _EVAL_2329 <= _EVAL_251;
      end
    end
    if (_EVAL_3227) begin
      _EVAL_2331 <= _EVAL_4373;
    end
    if (_EVAL_3624) begin
      _EVAL_2369 <= _EVAL_2573;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_2371 <= _EVAL_137;
      end else begin
        _EVAL_2371 <= _EVAL_265;
      end
    end
    if (_EVAL_3624) begin
      if (_EVAL_1493) begin
        if (_EVAL_2869) begin
          _EVAL_2383 <= _EVAL_234;
        end else begin
          if (_EVAL_1446) begin
            _EVAL_2383 <= _EVAL_110;
          end else begin
            _EVAL_2383 <= _EVAL_1495;
          end
        end
      end else begin
        if (_EVAL_4236) begin
          if (_EVAL_854) begin
            _EVAL_2383 <= csr__EVAL_84;
          end else begin
            if (_EVAL_3568) begin
              _EVAL_2383 <= m__EVAL_2;
            end else begin
              _EVAL_2383 <= _EVAL_3125;
            end
          end
        end else begin
          if (_EVAL_3876) begin
            _EVAL_2383 <= _EVAL_4863;
          end else begin
            if (_EVAL_3273) begin
              if (_EVAL_2257) begin
                _EVAL_2383 <= divider__EVAL_8;
              end else begin
                if (_EVAL_3629) begin
                  _EVAL_2383 <= fpu__EVAL_9;
                end else begin
                  _EVAL_2383 <= _EVAL_3727;
                end
              end
            end else begin
              _EVAL_2383 <= _EVAL_3494;
            end
          end
        end
      end
    end
    if (_EVAL_2118) begin
      _EVAL_2397 <= _EVAL_1921;
    end
    if (_EVAL_3624) begin
      _EVAL_2399 <= _EVAL_4649;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_2409 <= _EVAL_115;
        end else begin
          _EVAL_2409 <= _EVAL_251;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_2409 <= _EVAL_251;
        end else begin
          _EVAL_2409 <= _EVAL_115;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2423 <= _EVAL_723;
    end else begin
      if (_EVAL_3285) begin
        _EVAL_2423 <= _EVAL_263;
      end else begin
        if (_EVAL_2327) begin
          if (_EVAL_4409) begin
            _EVAL_2423 <= _EVAL_1834;
          end else begin
            if (_EVAL_4393) begin
              _EVAL_2423 <= _EVAL_4461;
            end else begin
              _EVAL_2423 <= _EVAL_4238;
            end
          end
        end
      end
    end
    if (_EVAL_3227) begin
      _EVAL_2424 <= _EVAL_1699;
    end
    if (_EVAL_3227) begin
      _EVAL_2443 <= _EVAL_951;
    end
    if (_EVAL_4240) begin
      _EVAL_2495 <= _EVAL_623;
    end
    if (_EVAL_4240) begin
      _EVAL_2499 <= _EVAL_2794;
    end
    if (_EVAL_2554) begin
      _EVAL_2506 <= 1'h0;
    end else begin
      if (_EVAL_1815) begin
        _EVAL_2506 <= 1'h1;
      end else begin
        if (_EVAL_511) begin
          _EVAL_2506 <= 1'h0;
        end else begin
          _EVAL_2506 <= _EVAL_2326;
        end
      end
    end
    if (_EVAL_2118) begin
      _EVAL_2542 <= _EVAL_4115;
    end
    if (_EVAL_4240) begin
      _EVAL_2573 <= _EVAL_4299;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_2579 <= _EVAL_171;
        end else begin
          _EVAL_2579 <= _EVAL_91;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_2579 <= _EVAL_91;
        end else begin
          _EVAL_2579 <= _EVAL_171;
        end
      end
    end
    _EVAL_2583 <= _EVAL_3310 & _EVAL_2088;
    if (_EVAL_3624) begin
      _EVAL_2587 <= _EVAL_2172;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_2596 <= _EVAL_188;
        end else begin
          _EVAL_2596 <= _EVAL_179;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_2596 <= _EVAL_179;
        end else begin
          _EVAL_2596 <= _EVAL_188;
        end
      end
    end
    if (_EVAL_3624) begin
      _EVAL_2603 <= _EVAL_4423;
    end
    if (_EVAL_4240) begin
      if (_EVAL_3979) begin
        _EVAL_2624 <= _EVAL_3621;
      end else begin
        if (_EVAL_2434) begin
          _EVAL_2624 <= _EVAL_1771;
        end else begin
          _EVAL_2624 <= _EVAL_4145;
        end
      end
    end
    _EVAL_2644 <= _EVAL_4735 & _EVAL_4567;
    if (_EVAL_936) begin
      if (_EVAL_4203) begin
        _EVAL_2656 <= {{16'd0}, _EVAL_1032};
      end else begin
        _EVAL_2656 <= _EVAL_4961;
      end
    end
    _EVAL_2667 <= csr__EVAL_39;
    _EVAL_2683 <= _EVAL_1028[4:0];
    if (_EVAL_4543) begin
      _EVAL_2686 <= _EVAL_2203;
    end
    if (_EVAL_2118) begin
      _EVAL_2753 <= _EVAL_2409;
    end
    if (_EVAL_3624) begin
      if (_EVAL_2195) begin
        _EVAL_2758 <= 32'h0;
      end else begin
        if (_EVAL_3624) begin
          if (_EVAL_1875) begin
            if (_EVAL_1206) begin
              if (_EVAL_1493) begin
                if (_EVAL_2869) begin
                  _EVAL_2758 <= _EVAL_234;
                end else begin
                  if (_EVAL_1446) begin
                    _EVAL_2758 <= _EVAL_110;
                  end else begin
                    _EVAL_2758 <= _EVAL_1495;
                  end
                end
              end else begin
                if (_EVAL_4236) begin
                  if (_EVAL_854) begin
                    _EVAL_2758 <= csr__EVAL_84;
                  end else begin
                    if (_EVAL_3568) begin
                      _EVAL_2758 <= m__EVAL_2;
                    end else begin
                      _EVAL_2758 <= _EVAL_3125;
                    end
                  end
                end else begin
                  if (_EVAL_3876) begin
                    _EVAL_2758 <= _EVAL_4863;
                  end else begin
                    if (_EVAL_3273) begin
                      if (_EVAL_2257) begin
                        _EVAL_2758 <= divider__EVAL_8;
                      end else begin
                        if (_EVAL_3629) begin
                          _EVAL_2758 <= fpu__EVAL_9;
                        end else begin
                          _EVAL_2758 <= _EVAL_3727;
                        end
                      end
                    end else begin
                      _EVAL_2758 <= _EVAL_2919;
                    end
                  end
                end
              end
            end else begin
              _EVAL_2758 <= _EVAL_2919;
            end
          end
        end
      end
    end else begin
      if (_EVAL_3624) begin
        if (_EVAL_1875) begin
          if (_EVAL_1206) begin
            if (_EVAL_1493) begin
              _EVAL_2758 <= _EVAL_4399;
            end else begin
              if (_EVAL_4236) begin
                _EVAL_2758 <= _EVAL_3923;
              end else begin
                if (_EVAL_3876) begin
                  _EVAL_2758 <= _EVAL_4863;
                end else begin
                  if (_EVAL_3273) begin
                    _EVAL_2758 <= _EVAL_3187;
                  end else begin
                    _EVAL_2758 <= _EVAL_2919;
                  end
                end
              end
            end
          end else begin
            _EVAL_2758 <= _EVAL_2919;
          end
        end
      end
    end
    if (_EVAL_2118) begin
      _EVAL_2765 <= _EVAL_3355;
    end
    if (_EVAL_5276) begin
      _EVAL_2794 <= _EVAL_583;
    end
    if (_EVAL_3971) begin
      _EVAL_2823 <= _EVAL_3109;
    end
    _EVAL_2843 <= _EVAL_47;
    if (_EVAL_2118) begin
      _EVAL_2853 <= _EVAL_284;
    end
    if (_EVAL_2548) begin
      _EVAL_2880 <= _EVAL_5009;
    end
    if (_EVAL_4240) begin
      _EVAL_2886 <= _EVAL_861;
    end
    if (_EVAL_4240) begin
      _EVAL_2911 <= _EVAL_3170;
    end
    if (_EVAL_2563) begin
      _EVAL_2912 <= _EVAL_2772;
    end
    if (_EVAL_4240) begin
      if (_EVAL_928) begin
        _EVAL_2919 <= _EVAL_4322;
      end else begin
        if (_EVAL_2717) begin
          _EVAL_2919 <= _EVAL_1932;
        end
      end
    end
    if (_EVAL_2355) begin
      if (_EVAL_4704) begin
        _EVAL_2948 <= _EVAL_2399;
      end else begin
        _EVAL_2948 <= _EVAL_4535;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_2955 <= _EVAL_35;
      end else begin
        _EVAL_2955 <= _EVAL_168;
      end
    end
    if (_EVAL_3624) begin
      _EVAL_2969 <= _EVAL_1828;
    end
    if (_EVAL_4240) begin
      _EVAL_2989 <= _EVAL_494;
    end
    if (_EVAL_4543) begin
      if (csr__EVAL_105) begin
        _EVAL_3000 <= 1'h1;
      end else begin
        if (_EVAL_315) begin
          _EVAL_3000 <= _EVAL_3226;
        end else begin
          _EVAL_3000 <= _EVAL_1661;
        end
      end
    end
    if (_EVAL_2832) begin
      _EVAL_3019 <= 128'h0;
    end else begin
      if (_EVAL_3102) begin
        _EVAL_3019 <= _EVAL_5349;
      end
    end
    if (_EVAL_936) begin
      if (_EVAL_1042) begin
        _EVAL_3025 <= {{16'd0}, _EVAL_477};
      end else begin
        _EVAL_3025 <= _EVAL_4430;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3029 <= _EVAL_905;
      end else begin
        _EVAL_3029 <= _EVAL_2403;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3039 <= _EVAL_6;
      end else begin
        _EVAL_3039 <= _EVAL_191;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3053 <= _EVAL_274;
      end else begin
        _EVAL_3053 <= _EVAL_154;
      end
    end
    if (_EVAL_4240) begin
      _EVAL_3064 <= _EVAL_3291;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1768) begin
        _EVAL_3077 <= _EVAL_4063;
      end else begin
        _EVAL_3077 <= _EVAL_674;
      end
    end
    if (_EVAL_3624) begin
      _EVAL_3085 <= _EVAL_1854;
    end
    _EVAL_3094 <= _EVAL_116 & _EVAL_159;
    _EVAL_3102 <= _EVAL_3971 & _EVAL_215;
    if (_EVAL_2118) begin
      _EVAL_3117 <= _EVAL_2579;
    end
    if (_EVAL_2118) begin
      _EVAL_3132 <= _EVAL_3940;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_3134 <= _EVAL_274;
        end else begin
          _EVAL_3134 <= _EVAL_154;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_3134 <= _EVAL_154;
        end else begin
          _EVAL_3134 <= _EVAL_274;
        end
      end
    end
    if (_EVAL_2506) begin
      _EVAL_3142 <= _EVAL_5009;
    end
    if (_EVAL_4543) begin
      _EVAL_3165 <= _EVAL_2084;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3170 <= _EVAL_57;
      end else begin
        _EVAL_3170 <= _EVAL_20;
      end
    end
    if (_EVAL_4240) begin
      _EVAL_3176 <= _EVAL_3588;
    end
    if (_EVAL_3624) begin
      _EVAL_3178 <= _EVAL_3064;
    end
    if (_EVAL_2506) begin
      _EVAL_3196 <= _EVAL_4656;
    end
    if (_EVAL_4240) begin
      _EVAL_3204 <= _EVAL_366;
    end
    if (_EVAL_4240) begin
      _EVAL_3217 <= _EVAL_3934;
    end
    if (_EVAL_2554) begin
      _EVAL_3227 <= 1'h0;
    end else begin
      if (_EVAL_2924) begin
        _EVAL_3227 <= 1'h0;
      end else begin
        if (_EVAL_1815) begin
          _EVAL_3227 <= 1'h0;
        end else begin
          if (_EVAL_4725) begin
            _EVAL_3227 <= 1'h0;
          end else begin
            _EVAL_3227 <= _EVAL_3624;
          end
        end
      end
    end
    if (_EVAL_3624) begin
      _EVAL_3229 <= _EVAL_2030;
    end
    if (_EVAL_5276) begin
      if (_EVAL_2693) begin
        _EVAL_3240 <= 1'h0;
      end else begin
        _EVAL_3240 <= _EVAL_1046;
      end
    end
    if (_EVAL_2355) begin
      if (_EVAL_4704) begin
        _EVAL_3270 <= _EVAL_356;
      end else begin
        _EVAL_3270 <= _EVAL_3974;
      end
    end
    if (_EVAL_2506) begin
      _EVAL_3276 <= _EVAL_4796;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3291 <= _EVAL_158;
      end else begin
        _EVAL_3291 <= _EVAL_222;
      end
    end
    if (_EVAL_2506) begin
      if (_EVAL_1523) begin
        _EVAL_3295 <= 1'h1;
      end else begin
        _EVAL_3295 <= _EVAL_3888;
      end
    end
    if (_EVAL_4240) begin
      _EVAL_3302 <= _EVAL_4968;
    end
    if (_EVAL_1558) begin
      _EVAL_3309 <= _EVAL_649;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_3355 <= _EVAL_206;
        end else begin
          _EVAL_3355 <= _EVAL_278;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_3355 <= _EVAL_278;
        end else begin
          _EVAL_3355 <= _EVAL_206;
        end
      end
    end
    _EVAL_3362 <= _EVAL_362 != 24'h0;
    _EVAL_3366 <= _EVAL_3381[4:0];
    _EVAL_3370 <= _EVAL_4967[4:0];
    if (_EVAL_3624) begin
      _EVAL_3384 <= _EVAL_4915;
    end
    if (_EVAL_4240) begin
      _EVAL_3386 <= _EVAL_5213;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_3391 <= _EVAL_205;
        end else begin
          _EVAL_3391 <= _EVAL_1;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_3391 <= _EVAL_1;
        end else begin
          _EVAL_3391 <= _EVAL_205;
        end
      end
    end
    if (_EVAL_2355) begin
      _EVAL_3393 <= _EVAL_3041;
    end
    if (_EVAL_2118) begin
      _EVAL_3401 <= _EVAL_3391;
    end
    if (_EVAL_1558) begin
      _EVAL_3404 <= _EVAL_2138;
    end
    if (_EVAL_1558) begin
      if (csr__EVAL_70) begin
        _EVAL_3405 <= csr__EVAL_44;
      end else begin
        if (_EVAL_5226) begin
          _EVAL_3405 <= _EVAL_2397;
        end else begin
          _EVAL_3405 <= {{28'd0}, _EVAL_2375};
        end
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3413 <= _EVAL_260;
      end else begin
        _EVAL_3413 <= _EVAL_119;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_3415 <= _EVAL_4437;
    end
    if (_EVAL_1558) begin
      _EVAL_3421 <= _EVAL_874;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3432 <= _EVAL_2;
      end else begin
        _EVAL_3432 <= _EVAL_138;
      end
    end
    _EVAL_3476 <= csr__EVAL_83[2];
    if (_EVAL_4543) begin
      _EVAL_3481 <= _EVAL_2175;
    end
    if (_EVAL_4240) begin
      _EVAL_3494 <= _EVAL_952;
    end
    _EVAL_3523 <= _EVAL_3003 != 24'h0;
    if (_EVAL_4543) begin
      if (_EVAL_1768) begin
        _EVAL_3573 <= 5'h5;
      end else begin
        _EVAL_3573 <= {{1'd0}, _EVAL_5011};
      end
    end
    if (_EVAL_5276) begin
      _EVAL_3588 <= _EVAL_3139;
    end
    if (_EVAL_2118) begin
      _EVAL_3608 <= _EVAL_3747;
    end
    if (_EVAL_2554) begin
      _EVAL_3624 <= 1'h0;
    end else begin
      _EVAL_3624 <= _EVAL_4240;
    end
    if (_EVAL_3227) begin
      _EVAL_3629 <= _EVAL_3085;
    end
    _EVAL_3637 <= _EVAL_4985 != 24'h0;
    if (_EVAL_3624) begin
      _EVAL_3645 <= _EVAL_3386;
    end
    if (_EVAL_4240) begin
      _EVAL_3670 <= _EVAL_4135;
    end
    if (_EVAL_1558) begin
      if (_EVAL_1815) begin
        _EVAL_3694 <= 1'h0;
      end else begin
        _EVAL_3694 <= _EVAL_639;
      end
    end
    if (_EVAL_4240) begin
      if (_EVAL_3383) begin
        if (_EVAL_3413) begin
          _EVAL_3711 <= _EVAL_4606;
        end else begin
          _EVAL_3711 <= _EVAL_623;
        end
      end
    end
    _EVAL_3712 <= _EVAL_339 != 24'h0;
    if (_EVAL_3227) begin
      _EVAL_3727 <= _EVAL_3923;
    end
    if (_EVAL_2355) begin
      if (_EVAL_651) begin
        _EVAL_3728 <= _EVAL_5043;
      end else begin
        if (csr__EVAL_89) begin
          _EVAL_3728 <= csr__EVAL_40;
        end else begin
          if (_EVAL_4027) begin
            if (_EVAL_4979) begin
              _EVAL_3728 <= _EVAL_1104;
            end else begin
              _EVAL_3728 <= _EVAL_341;
            end
          end else begin
            if (_EVAL_5100) begin
              _EVAL_3728 <= csr__EVAL_40;
            end else begin
              _EVAL_3728 <= _EVAL_5009;
            end
          end
        end
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3730 <= _EVAL_226;
      end else begin
        _EVAL_3730 <= _EVAL_31;
      end
    end
    if (_EVAL_3624) begin
      _EVAL_3742 <= _EVAL_3670;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_3747 <= _EVAL_16;
        end else begin
          _EVAL_3747 <= _EVAL_58;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_3747 <= _EVAL_58;
        end else begin
          _EVAL_3747 <= _EVAL_16;
        end
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3750 <= _EVAL_250;
      end else begin
        _EVAL_3750 <= _EVAL_141;
      end
    end
    if (_EVAL_2506) begin
      _EVAL_3752 <= _EVAL_4201;
    end
    _EVAL_3771 <= _EVAL_167;
    if (_EVAL_2118) begin
      _EVAL_3798 <= _EVAL_935;
    end
    _EVAL_3814 <= _EVAL_383 & _EVAL_2112;
    if (_EVAL_4543) begin
      _EVAL_3840 <= _EVAL_1597;
    end
    if (_EVAL_2506) begin
      _EVAL_3841 <= _EVAL_3309;
    end
    if (_EVAL_2506) begin
      _EVAL_3845 <= _EVAL_4748;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1843) begin
        if (_EVAL_1030) begin
          _EVAL_3851 <= _EVAL_1260;
        end else begin
          if (_EVAL_315) begin
            _EVAL_3851 <= _EVAL_68;
          end else begin
            _EVAL_3851 <= _EVAL_180;
          end
        end
      end
    end
    if (_EVAL_1558) begin
      _EVAL_3858 <= _EVAL_971;
    end
    if (_EVAL_5276) begin
      if (_EVAL_1922) begin
        if (_EVAL_683) begin
          _EVAL_3880 <= _EVAL_1572;
        end else begin
          if (_EVAL_5179) begin
            _EVAL_3880 <= _EVAL_1932;
          end else begin
            if (_EVAL_3042) begin
              _EVAL_3880 <= _EVAL_4679;
            end else begin
              if (_EVAL_2081) begin
                _EVAL_3880 <= _EVAL_2919;
              end else begin
                if (_EVAL_3542) begin
                  _EVAL_3880 <= _EVAL_4399;
                end else begin
                  if (_EVAL_2697) begin
                    _EVAL_3880 <= _EVAL_3923;
                  end else begin
                    if (_EVAL_2186) begin
                      _EVAL_3880 <= _EVAL_4863;
                    end else begin
                      if (_EVAL_4397) begin
                        _EVAL_3880 <= _EVAL_3187;
                      end else begin
                        if (_EVAL_315) begin
                          _EVAL_3880 <= _EVAL_4515;
                        end else begin
                          _EVAL_3880 <= _EVAL_1214;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_1558) begin
      if (_EVAL_4725) begin
        if (_EVAL_3624) begin
          _EVAL_3888 <= 1'h1;
        end else begin
          if (_EVAL_2342) begin
            _EVAL_3888 <= 1'h1;
          end else begin
            _EVAL_3888 <= _EVAL_937;
          end
        end
      end else begin
        if (_EVAL_2342) begin
          _EVAL_3888 <= 1'h1;
        end else begin
          _EVAL_3888 <= _EVAL_937;
        end
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_3902 <= _EVAL_198;
        end else begin
          _EVAL_3902 <= _EVAL_184;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_3902 <= _EVAL_184;
        end else begin
          _EVAL_3902 <= _EVAL_198;
        end
      end
    end
    if (_EVAL_4240) begin
      _EVAL_3922 <= _EVAL_1379;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_3934 <= _EVAL_272;
      end else begin
        _EVAL_3934 <= _EVAL_169;
      end
    end
    _EVAL_3939 <= _EVAL_2446 != 24'h0;
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_3940 <= _EVAL_2;
        end else begin
          _EVAL_3940 <= _EVAL_138;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_3940 <= _EVAL_138;
        end else begin
          _EVAL_3940 <= _EVAL_2;
        end
      end
    end
    if (_EVAL_1558) begin
      _EVAL_3974 <= _EVAL_4927;
    end
    if (_EVAL_4240) begin
      _EVAL_3986 <= _EVAL_3730;
    end
    if (_EVAL_4543) begin
      if (_EVAL_2084) begin
        _EVAL_3997 <= 1'h0;
      end else begin
        _EVAL_3997 <= _EVAL_3896;
      end
    end
    _EVAL_4000 <= _EVAL_1416 & _EVAL_4363;
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4014 <= _EVAL_205;
      end else begin
        _EVAL_4014 <= _EVAL_1;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_4019 <= _EVAL_1452;
    end
    if (_EVAL_2118) begin
      _EVAL_4043 <= _EVAL_653;
    end
    if (_EVAL_3624) begin
      if (_EVAL_2354) begin
        _EVAL_4064 <= {{2'd0}, _EVAL_3520};
      end else begin
        _EVAL_4064 <= _EVAL_3922;
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4088 <= _EVAL_202;
      end else begin
        _EVAL_4088 <= _EVAL_96;
      end
    end
    if (_EVAL_5276) begin
      _EVAL_4092 <= _EVAL_2366;
    end
    if (_EVAL_4543) begin
      if (_EVAL_315) begin
        _EVAL_4095 <= _EVAL_1;
      end else begin
        _EVAL_4095 <= _EVAL_205;
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_4115 <= _EVAL_186;
        end else begin
          _EVAL_4115 <= _EVAL_78;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_4115 <= _EVAL_78;
        end else begin
          _EVAL_4115 <= _EVAL_186;
        end
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4135 <= _EVAL_171;
      end else begin
        _EVAL_4135 <= _EVAL_91;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_4154 <= _EVAL_1727;
    end
    if (_EVAL_4240) begin
      _EVAL_4157 <= _EVAL_3432;
    end
    if (_EVAL_63) begin
      _EVAL_4160 <= 64'h0;
    end else begin
      if (_EVAL_1942) begin
        _EVAL_4160 <= _EVAL_2504;
      end
    end
    if (_EVAL_1558) begin
      if (_EVAL_4764) begin
        _EVAL_4162 <= {{2'd0}, _EVAL_3045};
      end else begin
        _EVAL_4162 <= _EVAL_4607;
      end
    end
    _EVAL_4167 <= _EVAL_4004 != 24'h0;
    _EVAL_4168 <= _EVAL_4924 != 24'h0;
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4192 <= _EVAL_73;
      end else begin
        _EVAL_4192 <= _EVAL_121;
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_3342) begin
        _EVAL_4195 <= _EVAL_1572;
      end else begin
        if (_EVAL_4829) begin
          _EVAL_4195 <= _EVAL_1932;
        end else begin
          if (_EVAL_325) begin
            _EVAL_4195 <= _EVAL_4679;
          end else begin
            if (_EVAL_4174) begin
              _EVAL_4195 <= _EVAL_2919;
            end else begin
              if (_EVAL_3609) begin
                _EVAL_4195 <= _EVAL_4399;
              end else begin
                if (_EVAL_1656) begin
                  _EVAL_4195 <= _EVAL_3923;
                end else begin
                  if (_EVAL_4417) begin
                    _EVAL_4195 <= _EVAL_4863;
                  end else begin
                    if (_EVAL_969) begin
                      _EVAL_4195 <= _EVAL_3187;
                    end else begin
                      if (_EVAL_315) begin
                        _EVAL_4195 <= _EVAL_5376;
                      end else begin
                        _EVAL_4195 <= _EVAL_1853;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_1558) begin
      _EVAL_4201 <= _EVAL_4607;
    end
    if (_EVAL_3624) begin
      _EVAL_4203 <= _EVAL_4562;
    end
    if (_EVAL_1062) begin
      _EVAL_4218 <= _EVAL_5341;
    end
    if (_EVAL_1548) begin
      _EVAL_4240 <= 1'h0;
    end else begin
      _EVAL_4240 <= _EVAL_3821;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4299 <= _EVAL_16;
      end else begin
        _EVAL_4299 <= _EVAL_58;
      end
    end
    if (_EVAL_3227) begin
      _EVAL_4319 <= _EVAL_2383;
    end
    if (_EVAL_5276) begin
      if (_EVAL_3799) begin
        if (_EVAL_3514) begin
          _EVAL_4322 <= _EVAL_1572;
        end else begin
          if (_EVAL_2668) begin
            _EVAL_4322 <= _EVAL_1932;
          end else begin
            if (_EVAL_2073) begin
              _EVAL_4322 <= _EVAL_4679;
            end else begin
              if (_EVAL_4207) begin
                _EVAL_4322 <= _EVAL_2919;
              end else begin
                if (_EVAL_391) begin
                  _EVAL_4322 <= _EVAL_4399;
                end else begin
                  if (_EVAL_1129) begin
                    _EVAL_4322 <= _EVAL_3923;
                  end else begin
                    if (_EVAL_4046) begin
                      _EVAL_4322 <= _EVAL_4863;
                    end else begin
                      if (_EVAL_2464) begin
                        _EVAL_4322 <= _EVAL_3187;
                      end else begin
                        if (_EVAL_315) begin
                          _EVAL_4322 <= _EVAL_1853;
                        end else begin
                          _EVAL_4322 <= _EVAL_5376;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    _EVAL_4360 <= _EVAL_159 & _EVAL_3128;
    if (_EVAL_2869) begin
      _EVAL_4362 <= _EVAL_1860;
    end else begin
      if (_EVAL_2506) begin
        _EVAL_4362 <= _EVAL_4962;
      end
    end
    if (_EVAL_3624) begin
      if (_EVAL_1654) begin
        if (_EVAL_4882) begin
          _EVAL_4373 <= _EVAL_4399;
        end else begin
          if (_EVAL_1832) begin
            _EVAL_4373 <= _EVAL_3923;
          end else begin
            if (_EVAL_418) begin
              _EVAL_4373 <= _EVAL_4863;
            end else begin
              if (_EVAL_948) begin
                _EVAL_4373 <= _EVAL_3187;
              end else begin
                _EVAL_4373 <= _EVAL_1109;
              end
            end
          end
        end
      end
    end
    if (_EVAL_4543) begin
      if (_EVAL_2776) begin
        if (_EVAL_3299) begin
          if (_EVAL_315) begin
            _EVAL_4400 <= _EVAL_68;
          end else begin
            _EVAL_4400 <= _EVAL_180;
          end
        end else begin
          if (_EVAL_315) begin
            _EVAL_4400 <= _EVAL_154;
          end else begin
            _EVAL_4400 <= _EVAL_274;
          end
        end
      end
    end
    if (_EVAL_4240) begin
      _EVAL_4423 <= _EVAL_2329;
    end
    if (_EVAL_2118) begin
      _EVAL_4437 <= _EVAL_3481;
    end
    if (_EVAL_4240) begin
      _EVAL_4460 <= _EVAL_3053;
    end
    if (_EVAL_4580) begin
      _EVAL_4461 <= _EVAL_2621;
    end
    if (_EVAL_4543) begin
      if (_EVAL_684) begin
        if (_EVAL_3342) begin
          _EVAL_4468 <= _EVAL_1572;
        end else begin
          if (_EVAL_4829) begin
            _EVAL_4468 <= _EVAL_1932;
          end else begin
            if (_EVAL_325) begin
              _EVAL_4468 <= _EVAL_4679;
            end else begin
              if (_EVAL_4174) begin
                _EVAL_4468 <= _EVAL_2919;
              end else begin
                if (_EVAL_3609) begin
                  _EVAL_4468 <= _EVAL_4399;
                end else begin
                  if (_EVAL_1656) begin
                    _EVAL_4468 <= _EVAL_3923;
                  end else begin
                    if (_EVAL_4417) begin
                      _EVAL_4468 <= _EVAL_4863;
                    end else begin
                      if (_EVAL_969) begin
                        _EVAL_4468 <= _EVAL_3187;
                      end else begin
                        if (_EVAL_315) begin
                          _EVAL_4468 <= _EVAL_5376;
                        end else begin
                          _EVAL_4468 <= _EVAL_1853;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4481 <= _EVAL_97;
      end else begin
        _EVAL_4481 <= _EVAL_23;
      end
    end
    if (_EVAL_3227) begin
      _EVAL_4512 <= _EVAL_1352;
    end
    if (_EVAL_4240) begin
      _EVAL_4530 <= _EVAL_3039;
    end
    _EVAL_4531 <= _EVAL_1416 & _EVAL_4731;
    if (_EVAL_1558) begin
      _EVAL_4535 <= _EVAL_3798;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_4539 <= _EVAL_84;
        end else begin
          _EVAL_4539 <= _EVAL_153;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_4539 <= _EVAL_153;
        end else begin
          _EVAL_4539 <= _EVAL_84;
        end
      end
    end
    if (_EVAL_2355) begin
      if (_EVAL_4704) begin
        _EVAL_4550 <= _EVAL_3384;
      end else begin
        _EVAL_4550 <= _EVAL_4154;
      end
    end
    if (_EVAL_4240) begin
      _EVAL_4562 <= _EVAL_1476;
    end
    if (_EVAL_2118) begin
      _EVAL_4596 <= _EVAL_545;
    end
    if (_EVAL_3227) begin
      _EVAL_4600 <= _EVAL_5043;
    end
    if (_EVAL_2118) begin
      _EVAL_4607 <= _EVAL_4539;
    end
    if (_EVAL_3624) begin
      _EVAL_4614 <= _EVAL_4530;
    end
    _EVAL_4620 <= csr__EVAL_83[2];
    if (_EVAL_5276) begin
      _EVAL_4632 <= _EVAL_3181;
    end
    if (_EVAL_4543) begin
      if (_EVAL_1181) begin
        if (_EVAL_315) begin
          _EVAL_4633 <= _EVAL_6;
        end else begin
          _EVAL_4633 <= _EVAL_191;
        end
      end else begin
        if (_EVAL_315) begin
          _EVAL_4633 <= _EVAL_191;
        end else begin
          _EVAL_4633 <= _EVAL_6;
        end
      end
    end
    if (_EVAL_4240) begin
      _EVAL_4649 <= _EVAL_2371;
    end
    if (_EVAL_1558) begin
      if (_EVAL_5183) begin
        _EVAL_4656 <= _EVAL_4399;
      end else begin
        if (_EVAL_1891) begin
          _EVAL_4656 <= _EVAL_3923;
        end else begin
          if (_EVAL_1961) begin
            _EVAL_4656 <= _EVAL_4863;
          end else begin
            if (_EVAL_4599) begin
              _EVAL_4656 <= _EVAL_3187;
            end else begin
              _EVAL_4656 <= _EVAL_1294;
            end
          end
        end
      end
    end
    if (_EVAL_2118) begin
      if (_EVAL_2238) begin
        _EVAL_4679 <= _EVAL_4468;
      end else begin
        if (_EVAL_2632) begin
          _EVAL_4679 <= _EVAL_1572;
        end
      end
    end
    if (_EVAL_5276) begin
      _EVAL_4684 <= _EVAL_2500;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4692 <= _EVAL_214;
      end else begin
        _EVAL_4692 <= _EVAL_268;
      end
    end
    if (_EVAL_2118) begin
      _EVAL_4698 <= _EVAL_792;
    end
    if (_EVAL_1558) begin
      _EVAL_4706 <= _EVAL_3117;
    end
    if (_EVAL_1558) begin
      _EVAL_4715 <= _EVAL_1059;
    end
    if (_EVAL_2506) begin
      _EVAL_4736 <= _EVAL_5178;
    end
    if (_EVAL_4240) begin
      if (_EVAL_2244) begin
        _EVAL_4745 <= _EVAL_623;
      end
    end
    if (_EVAL_1558) begin
      if (_EVAL_690) begin
        if (_EVAL_2103) begin
          _EVAL_4748 <= _EVAL_4399;
        end else begin
          if (_EVAL_510) begin
            _EVAL_4748 <= _EVAL_3923;
          end else begin
            if (_EVAL_1770) begin
              _EVAL_4748 <= _EVAL_4863;
            end else begin
              if (_EVAL_2426) begin
                _EVAL_4748 <= _EVAL_3187;
              end else begin
                _EVAL_4748 <= _EVAL_5367;
              end
            end
          end
        end
      end
    end
    if (_EVAL_3624) begin
      _EVAL_4790 <= _EVAL_2989;
    end
    if (_EVAL_1558) begin
      _EVAL_4796 <= _EVAL_1521;
    end
    _EVAL_4805 <= _EVAL_147;
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4812 <= _EVAL_232;
      end else begin
        _EVAL_4812 <= _EVAL_102;
      end
    end
    if (_EVAL_2326) begin
      _EVAL_4819 <= _EVAL_2068;
    end
    if (_EVAL_2118) begin
      if (_EVAL_4355) begin
        _EVAL_4842 <= 1'h1;
      end else begin
        _EVAL_4842 <= _EVAL_3902;
      end
    end
    if (_EVAL_3227) begin
      _EVAL_4844 <= _EVAL_2219;
    end
    if (_EVAL_2869) begin
      _EVAL_4863 <= _EVAL_4399;
    end else begin
      if (_EVAL_3672) begin
        _EVAL_4863 <= _EVAL_5412;
      end else begin
        if (_EVAL_2506) begin
          _EVAL_4863 <= _EVAL_4399;
        end
      end
    end
    if (_EVAL_4240) begin
      _EVAL_4915 <= _EVAL_4481;
    end
    if (_EVAL_2118) begin
      _EVAL_4927 <= _EVAL_5265;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4936 <= _EVAL_198;
      end else begin
        _EVAL_4936 <= _EVAL_184;
      end
    end
    if (_EVAL_3227) begin
      _EVAL_4939 <= _EVAL_3742;
    end
    _EVAL_4947 <= csr__EVAL_39;
    if (_EVAL_1558) begin
      _EVAL_4962 <= _EVAL_3608;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_4968 <= _EVAL_183;
      end else begin
        _EVAL_4968 <= _EVAL_208;
      end
    end
    if (_EVAL_3624) begin
      if (_EVAL_5285) begin
        _EVAL_5009 <= _EVAL_2423;
      end else begin
        if (_EVAL_1558) begin
          if (_EVAL_1815) begin
            _EVAL_5009 <= _EVAL_2423;
          end else begin
            _EVAL_5009 <= _EVAL_3132;
          end
        end
      end
    end else begin
      if (_EVAL_1558) begin
        if (_EVAL_1815) begin
          _EVAL_5009 <= _EVAL_2423;
        end else begin
          _EVAL_5009 <= _EVAL_3132;
        end
      end
    end
    if (_EVAL_1558) begin
      _EVAL_5017 <= _EVAL_4698;
    end
    if (_EVAL_3624) begin
      _EVAL_5025 <= _EVAL_3986;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_5039 <= _EVAL_45;
      end else begin
        _EVAL_5039 <= _EVAL_104;
      end
    end
    if (_EVAL_3624) begin
      _EVAL_5043 <= _EVAL_4157;
    end
    if (_EVAL_3624) begin
      _EVAL_5052 <= _EVAL_5004;
    end
    if (_EVAL_4240) begin
      _EVAL_5095 <= _EVAL_3413;
    end
    if (_EVAL_2869) begin
      _EVAL_5099 <= _EVAL_3769;
    end else begin
      if (_EVAL_2506) begin
        _EVAL_5099 <= _EVAL_4706;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_5178 <= _EVAL_2753;
    end
    if (_EVAL_5276) begin
      if (_EVAL_315) begin
        _EVAL_5213 <= _EVAL_51;
      end else begin
        _EVAL_5213 <= _EVAL_64;
      end
    end
    if (_EVAL_2118) begin
      _EVAL_5226 <= _EVAL_3165;
    end
    if (_EVAL_4240) begin
      _EVAL_5233 <= _EVAL_1187;
    end
    if (_EVAL_4543) begin
      _EVAL_5237 <= _EVAL_4756;
    end
    if (_EVAL_4543) begin
      if (_EVAL_315) begin
        _EVAL_5265 <= _EVAL_208;
      end else begin
        _EVAL_5265 <= _EVAL_183;
      end
    end
    if (_EVAL_4240) begin
      _EVAL_5335 <= _EVAL_2955;
    end
    if (_EVAL_4240) begin
      _EVAL_5344 <= _EVAL_4014;
    end
    if (_EVAL_3624) begin
      _EVAL_5363 <= _EVAL_4460;
    end
    if (_EVAL_2118) begin
      if (_EVAL_666) begin
        _EVAL_5367 <= _EVAL_949;
      end
    end
    if (_EVAL_2326) begin
      if (_EVAL_5226) begin
        _EVAL_5412 <= _EVAL_1834;
      end else begin
        if (_EVAL_2853) begin
          _EVAL_5412 <= _EVAL_4035;
        end else begin
          if (_EVAL_1558) begin
            if (_EVAL_1100) begin
              if (_EVAL_1533) begin
                if (_EVAL_5183) begin
                  _EVAL_5412 <= _EVAL_4399;
                end else begin
                  if (_EVAL_1891) begin
                    _EVAL_5412 <= _EVAL_3923;
                  end else begin
                    if (_EVAL_1961) begin
                      _EVAL_5412 <= _EVAL_4863;
                    end else begin
                      if (_EVAL_4599) begin
                        _EVAL_5412 <= _EVAL_3187;
                      end else begin
                        _EVAL_5412 <= _EVAL_4679;
                      end
                    end
                  end
                end
              end else begin
                _EVAL_5412 <= _EVAL_4679;
              end
            end
          end
        end
      end
    end else begin
      if (_EVAL_1558) begin
        if (_EVAL_1100) begin
          if (_EVAL_1533) begin
            if (_EVAL_5183) begin
              _EVAL_5412 <= _EVAL_4399;
            end else begin
              if (_EVAL_1891) begin
                _EVAL_5412 <= _EVAL_3923;
              end else begin
                if (_EVAL_1961) begin
                  _EVAL_5412 <= _EVAL_4863;
                end else begin
                  if (_EVAL_4599) begin
                    _EVAL_5412 <= _EVAL_3187;
                  end else begin
                    _EVAL_5412 <= _EVAL_4679;
                  end
                end
              end
            end
          end else begin
            _EVAL_5412 <= _EVAL_4679;
          end
        end
      end
    end
  end
  always @(posedge fpu_clock_gate_out) begin
    if(_EVAL_2741__EVAL_2751_en & _EVAL_2741__EVAL_2751_mask) begin
      _EVAL_2741[_EVAL_2741__EVAL_2751_addr] <= _EVAL_2741__EVAL_2751_data;
    end
    if(_EVAL_2741__EVAL_2752_en & _EVAL_2741__EVAL_2752_mask) begin
      _EVAL_2741[_EVAL_2741__EVAL_2752_addr] <= _EVAL_2741__EVAL_2752_data;
    end
  end
  always @(posedge _EVAL_267) begin
    _EVAL_601 <= _EVAL_3603 | _EVAL_1605;
    _EVAL_896 <= _EVAL_2863 | fpu__EVAL_40;
    if (_EVAL_5221) begin
      _EVAL_1149 <= 1'h0;
    end else begin
      if (_EVAL_4543) begin
        if (_EVAL_4955) begin
          _EVAL_1149 <= 1'h1;
        end
      end
    end
    _EVAL_1896 <= _EVAL_1289 | _EVAL_2355;
    if (_EVAL_63) begin
      _EVAL_3448 <= 1'h1;
    end else begin
      _EVAL_3448 <= _EVAL_4059;
    end
  end
endmodule
