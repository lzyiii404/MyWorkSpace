//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_241_assert(
  input  [1:0]  _EVAL,
  input         _EVAL_0,
  input  [12:0] _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [24:0] _EVAL_9,
  input  [12:0] _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_45;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_48;
  reg [31:0] _RAND_1;
  reg  _EVAL_54;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_70;
  reg [31:0] _RAND_3;
  reg  _EVAL_82;
  reg [31:0] _RAND_4;
  reg [12:0] _EVAL_88;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_95;
  reg [31:0] _RAND_6;
  reg  _EVAL_149;
  reg [31:0] _RAND_7;
  reg [31:0] _EVAL_200;
  reg [31:0] _RAND_8;
  reg [24:0] _EVAL_201;
  reg [31:0] _RAND_9;
  reg  _EVAL_208;
  reg [31:0] _RAND_10;
  reg [12:0] _EVAL_210;
  reg [31:0] _RAND_11;
  reg [4351:0] _EVAL_230;
  reg [4351:0] _RAND_12;
  reg [1:0] _EVAL_233;
  reg [31:0] _RAND_13;
  wire  _EVAL_237;
  wire  _EVAL_65;
  wire  _EVAL_157;
  wire  _EVAL_206;
  wire  _EVAL_183;
  wire  _EVAL_224;
  wire  _EVAL_232;
  wire  _EVAL_188;
  wire  _EVAL_115;
  wire  _EVAL_20;
  wire  _EVAL_41;
  wire [8191:0] _EVAL_156;
  wire [8191:0] _EVAL_218;
  wire [4351:0] _EVAL_192;
  wire [4351:0] _EVAL_17;
  wire  _EVAL_166;
  wire  _EVAL_209;
  wire  _EVAL_78;
  wire  _EVAL_83;
  wire  _EVAL_121;
  wire  _EVAL_91;
  wire  _EVAL_57;
  wire  _EVAL_76;
  wire  _EVAL_175;
  wire [1:0] _EVAL_215;
  wire [1:0] _EVAL_59;
  wire  _EVAL_51;
  wire  _EVAL_29;
  wire  _EVAL_21;
  wire  _EVAL_164;
  wire  _EVAL_180;
  wire  _EVAL_18;
  wire  _EVAL_184;
  wire  _EVAL_72;
  wire  _EVAL_163;
  wire  _EVAL_26;
  wire  _EVAL_142;
  wire  _EVAL_173;
  wire  _EVAL_99;
  wire  _EVAL_211;
  wire  _EVAL_225;
  wire  _EVAL_158;
  wire  _EVAL_205;
  wire  _EVAL_178;
  wire  _EVAL_81;
  wire  _EVAL_126;
  wire  _EVAL_73;
  wire  _EVAL_235;
  wire [3:0] _EVAL_222;
  wire  _EVAL_122;
  wire  _EVAL_189;
  wire  _EVAL_140;
  wire  _EVAL_105;
  wire  _EVAL_216;
  wire  _EVAL_66;
  wire  _EVAL_96;
  wire  _EVAL_236;
  wire  _EVAL_103;
  wire  _EVAL_125;
  wire  _EVAL_19;
  wire  _EVAL_234;
  wire  _EVAL_134;
  wire  _EVAL_85;
  wire  _EVAL_151;
  wire  _EVAL_132;
  wire  _EVAL_116;
  wire  _EVAL_84;
  wire  _EVAL_231;
  wire  _EVAL_100;
  wire  _EVAL_75;
  wire [4:0] _EVAL_160;
  wire [3:0] _EVAL_33;
  wire [3:0] _EVAL_87;
  wire  _EVAL_30;
  wire  _EVAL_214;
  wire  _EVAL_162;
  wire  _EVAL_109;
  wire  _EVAL_101;
  wire  _EVAL_168;
  wire [1:0] _EVAL_141;
  wire [1:0] _EVAL_50;
  wire [24:0] _EVAL_68;
  wire [24:0] _EVAL_191;
  wire  _EVAL_169;
  wire  _EVAL_71;
  wire  _EVAL_220;
  wire  _EVAL_27;
  wire  _EVAL_171;
  wire [31:0] _EVAL_170;
  wire  _EVAL_152;
  wire  _EVAL_46;
  wire  _EVAL_15;
  wire  _EVAL_161;
  wire  _EVAL_60;
  wire  _EVAL_147;
  wire  _EVAL_52;
  wire  _EVAL_118;
  wire  _EVAL_67;
  wire  _EVAL_194;
  wire  _EVAL_106;
  wire [8191:0] _EVAL_24;
  wire [8191:0] _EVAL_136;
  wire [4351:0] _EVAL_227;
  wire [4351:0] _EVAL_56;
  wire [4351:0] _EVAL_22;
  wire  _EVAL_174;
  wire  _EVAL_150;
  wire  _EVAL_64;
  wire  _EVAL_53;
  wire  _EVAL_120;
  wire  _EVAL_176;
  wire  _EVAL_42;
  wire  _EVAL_137;
  wire  _EVAL_238;
  wire  _EVAL_127;
  wire  _EVAL_228;
  wire  _EVAL_190;
  wire  _EVAL_155;
  wire  _EVAL_159;
  wire  _EVAL_61;
  wire [24:0] _EVAL_36;
  wire [25:0] _EVAL_112;
  wire  _EVAL_165;
  wire  _EVAL_108;
  wire  _EVAL_199;
  wire  _EVAL_223;
  wire  _EVAL_177;
  wire [4351:0] _EVAL_63;
  wire  _EVAL_102;
  wire  _EVAL_124;
  wire  _EVAL_203;
  wire  _EVAL_148;
  wire  _EVAL_145;
  wire  _EVAL_138;
  wire  _EVAL_213;
  wire  _EVAL_217;
  wire  _EVAL_212;
  wire  _EVAL_154;
  wire  _EVAL_86;
  wire  _EVAL_167;
  wire  _EVAL_226;
  wire  _EVAL_181;
  wire  _EVAL_16;
  wire [3:0] _EVAL_62;
  wire  _EVAL_186;
  wire [4351:0] _EVAL_117;
  wire [4351:0] _EVAL_79;
  wire  _EVAL_28;
  wire  _EVAL_135;
  wire  _EVAL_94;
  wire  _EVAL_196;
  wire  _EVAL_49;
  wire  _EVAL_107;
  wire  _EVAL_40;
  wire  _EVAL_207;
  wire  _EVAL_119;
  wire  _EVAL_38;
  wire  _EVAL_131;
  wire  _EVAL_37;
  wire  _EVAL_34;
  wire  _EVAL_153;
  wire  _EVAL_113;
  wire  _EVAL_55;
  wire  _EVAL_31;
  wire  _EVAL_182;
  wire  _EVAL_97;
  wire  _EVAL_110;
  wire  _EVAL_143;
  wire  _EVAL_43;
  wire  _EVAL_114;
  wire  _EVAL_229;
  wire  _EVAL_187;
  wire [25:0] _EVAL_130;
  wire [25:0] _EVAL_221;
  wire  _EVAL_139;
  wire  _EVAL_133;
  wire  _EVAL_172;
  wire  _EVAL_98;
  wire  _EVAL_44;
  wire  _EVAL_90;
  wire  _EVAL_202;
  wire  _EVAL_47;
  wire  _EVAL_25;
  wire  _EVAL_123;
  wire  _EVAL_198;
  wire  _EVAL_89;
  wire  _EVAL_193;
  wire  _EVAL_195;
  wire  _EVAL_39;
  wire  _EVAL_32;
  wire  _EVAL_179;
  wire  _EVAL_69;
  wire  _EVAL_93;
  wire  _EVAL_77;
  wire  _EVAL_144;
  wire  _EVAL_58;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_237 = _EVAL_9 == _EVAL_201;
  assign _EVAL_65 = _EVAL_237 | _EVAL_0;
  assign _EVAL_157 = _EVAL_65 == 1'h0;
  assign _EVAL_206 = _EVAL_13 == _EVAL_48;
  assign _EVAL_183 = _EVAL_206 | _EVAL_0;
  assign _EVAL_224 = _EVAL_3 & _EVAL_12;
  assign _EVAL_232 = _EVAL_149 == 1'h0;
  assign _EVAL_188 = _EVAL_224 & _EVAL_232;
  assign _EVAL_115 = _EVAL_6 == 3'h6;
  assign _EVAL_20 = _EVAL_115 == 1'h0;
  assign _EVAL_41 = _EVAL_188 & _EVAL_20;
  assign _EVAL_156 = 8192'h1 << _EVAL_1;
  assign _EVAL_218 = _EVAL_41 ? _EVAL_156 : 8192'h0;
  assign _EVAL_192 = _EVAL_218[4351:0];
  assign _EVAL_17 = ~ _EVAL_192;
  assign _EVAL_166 = _EVAL_2 == 3'h0;
  assign _EVAL_209 = _EVAL_166 | _EVAL_0;
  assign _EVAL_78 = _EVAL_209 == 1'h0;
  assign _EVAL_83 = _EVAL_10 <= 13'h10ff;
  assign _EVAL_121 = _EVAL_83 | _EVAL_0;
  assign _EVAL_91 = _EVAL_121 == 1'h0;
  assign _EVAL_57 = _EVAL_2 <= 3'h4;
  assign _EVAL_76 = _EVAL >= 2'h2;
  assign _EVAL_175 = _EVAL[0];
  assign _EVAL_215 = 2'h1 << _EVAL_175;
  assign _EVAL_59 = _EVAL_215 | 2'h1;
  assign _EVAL_51 = _EVAL_59[1];
  assign _EVAL_29 = _EVAL_9[1];
  assign _EVAL_21 = _EVAL_51 & _EVAL_29;
  assign _EVAL_164 = _EVAL_76 | _EVAL_21;
  assign _EVAL_180 = _EVAL_59[0];
  assign _EVAL_18 = _EVAL_9[0];
  assign _EVAL_184 = _EVAL_29 & _EVAL_18;
  assign _EVAL_72 = _EVAL_180 & _EVAL_184;
  assign _EVAL_163 = _EVAL_164 | _EVAL_72;
  assign _EVAL_26 = _EVAL_18 == 1'h0;
  assign _EVAL_142 = _EVAL_29 & _EVAL_26;
  assign _EVAL_173 = _EVAL_180 & _EVAL_142;
  assign _EVAL_99 = _EVAL_164 | _EVAL_173;
  assign _EVAL_211 = _EVAL_29 == 1'h0;
  assign _EVAL_225 = _EVAL_51 & _EVAL_211;
  assign _EVAL_158 = _EVAL_76 | _EVAL_225;
  assign _EVAL_205 = _EVAL_211 & _EVAL_18;
  assign _EVAL_178 = _EVAL_180 & _EVAL_205;
  assign _EVAL_81 = _EVAL_158 | _EVAL_178;
  assign _EVAL_126 = _EVAL_211 & _EVAL_26;
  assign _EVAL_73 = _EVAL_180 & _EVAL_126;
  assign _EVAL_235 = _EVAL_158 | _EVAL_73;
  assign _EVAL_222 = {_EVAL_163,_EVAL_99,_EVAL_81,_EVAL_235};
  assign _EVAL_122 = _EVAL_8 == _EVAL_222;
  assign _EVAL_189 = _EVAL_57 | _EVAL_0;
  assign _EVAL_140 = _EVAL_230 != 4352'h0;
  assign _EVAL_105 = _EVAL_140 == 1'h0;
  assign _EVAL_216 = plusarg_reader_out == 32'h0;
  assign _EVAL_66 = _EVAL_105 | _EVAL_216;
  assign _EVAL_96 = _EVAL_200 < plusarg_reader_out;
  assign _EVAL_236 = _EVAL_66 | _EVAL_96;
  assign _EVAL_103 = _EVAL_13 == 3'h5;
  assign _EVAL_125 = _EVAL_11 & _EVAL_103;
  assign _EVAL_19 = _EVAL_6 == 3'h5;
  assign _EVAL_234 = _EVAL_76 | _EVAL_0;
  assign _EVAL_134 = _EVAL_234 == 1'h0;
  assign _EVAL_85 = _EVAL_1 <= 13'h10ff;
  assign _EVAL_151 = _EVAL_85 | _EVAL_0;
  assign _EVAL_132 = _EVAL_151 == 1'h0;
  assign _EVAL_116 = _EVAL_2 != 3'h0;
  assign _EVAL_84 = _EVAL_6 == _EVAL_95;
  assign _EVAL_231 = _EVAL_84 | _EVAL_0;
  assign _EVAL_100 = _EVAL_231 == 1'h0;
  assign _EVAL_75 = _EVAL_13 == 3'h0;
  assign _EVAL_160 = 5'h3 << _EVAL;
  assign _EVAL_33 = ~ _EVAL_222;
  assign _EVAL_87 = _EVAL_8 & _EVAL_33;
  assign _EVAL_30 = _EVAL_87 == 4'h0;
  assign _EVAL_214 = _EVAL_30 | _EVAL_0;
  assign _EVAL_162 = _EVAL_5 == 1'h0;
  assign _EVAL_109 = _EVAL_6 == 3'h4;
  assign _EVAL_101 = _EVAL_12 & _EVAL_109;
  assign _EVAL_168 = _EVAL_6 == 3'h1;
  assign _EVAL_141 = _EVAL_160[1:0];
  assign _EVAL_50 = ~ _EVAL_141;
  assign _EVAL_68 = {{23'd0}, _EVAL_50};
  assign _EVAL_191 = _EVAL_9 & _EVAL_68;
  assign _EVAL_169 = _EVAL_191 == 25'h0;
  assign _EVAL_71 = _EVAL_169 | _EVAL_0;
  assign _EVAL_220 = _EVAL_7 == _EVAL_233;
  assign _EVAL_27 = _EVAL_14 & _EVAL_11;
  assign _EVAL_171 = _EVAL_27 | _EVAL_224;
  assign _EVAL_170 = _EVAL_200 + 32'h1;
  assign _EVAL_152 = _EVAL_162 | _EVAL_0;
  assign _EVAL_46 = _EVAL_152 == 1'h0;
  assign _EVAL_15 = _EVAL_2 <= 3'h3;
  assign _EVAL_161 = _EVAL_15 | _EVAL_0;
  assign _EVAL_60 = _EVAL_6 == 3'h2;
  assign _EVAL_147 = _EVAL_10 == _EVAL_88;
  assign _EVAL_52 = _EVAL_12 & _EVAL_60;
  assign _EVAL_118 = _EVAL_0 == 1'h0;
  assign _EVAL_67 = _EVAL <= 2'h2;
  assign _EVAL_194 = _EVAL_82 == 1'h0;
  assign _EVAL_106 = _EVAL_27 & _EVAL_194;
  assign _EVAL_24 = 8192'h1 << _EVAL_10;
  assign _EVAL_136 = _EVAL_106 ? _EVAL_24 : 8192'h0;
  assign _EVAL_227 = _EVAL_136[4351:0];
  assign _EVAL_56 = _EVAL_227 | _EVAL_230;
  assign _EVAL_22 = _EVAL_56 >> _EVAL_1;
  assign _EVAL_174 = _EVAL_13 == 3'h6;
  assign _EVAL_150 = _EVAL_11 & _EVAL_174;
  assign _EVAL_64 = _EVAL_54 == 1'h0;
  assign _EVAL_53 = _EVAL_64 == 1'h0;
  assign _EVAL_120 = _EVAL_12 & _EVAL_53;
  assign _EVAL_176 = _EVAL_22[0];
  assign _EVAL_42 = _EVAL_7 >= 2'h2;
  assign _EVAL_137 = _EVAL_42 | _EVAL_0;
  assign _EVAL_238 = _EVAL_137 == 1'h0;
  assign _EVAL_127 = _EVAL_183 == 1'h0;
  assign _EVAL_228 = _EVAL_149 - 1'h1;
  assign _EVAL_190 = _EVAL_13 == 3'h2;
  assign _EVAL_155 = _EVAL_11 & _EVAL_190;
  assign _EVAL_159 = _EVAL_13 == 3'h7;
  assign _EVAL_61 = _EVAL_2 <= 3'h2;
  assign _EVAL_36 = _EVAL_9 ^ 25'h1900000;
  assign _EVAL_112 = {1'b0,$signed(_EVAL_36)};
  assign _EVAL_165 = _EVAL_61 | _EVAL_0;
  assign _EVAL_108 = _EVAL_54 - 1'h1;
  assign _EVAL_199 = _EVAL_6 <= 3'h6;
  assign _EVAL_223 = _EVAL_199 | _EVAL_0;
  assign _EVAL_177 = _EVAL_223 == 1'h0;
  assign _EVAL_63 = _EVAL_230 >> _EVAL_10;
  assign _EVAL_102 = _EVAL_63[0];
  assign _EVAL_124 = _EVAL_102 == 1'h0;
  assign _EVAL_203 = _EVAL_124 | _EVAL_0;
  assign _EVAL_148 = _EVAL_208 == 1'h0;
  assign _EVAL_145 = _EVAL_27 & _EVAL_148;
  assign _EVAL_138 = _EVAL_1 == _EVAL_210;
  assign _EVAL_213 = _EVAL_13 == 3'h1;
  assign _EVAL_217 = _EVAL_148 == 1'h0;
  assign _EVAL_212 = _EVAL_11 & _EVAL_217;
  assign _EVAL_154 = _EVAL_82 - 1'h1;
  assign _EVAL_86 = _EVAL_6 == 3'h0;
  assign _EVAL_167 = _EVAL_224 & _EVAL_64;
  assign _EVAL_226 = _EVAL_236 | _EVAL_0;
  assign _EVAL_181 = _EVAL_226 == 1'h0;
  assign _EVAL_16 = _EVAL_176 | _EVAL_0;
  assign _EVAL_62 = ~ _EVAL_8;
  assign _EVAL_186 = _EVAL_62 == 4'h0;
  assign _EVAL_117 = _EVAL_230 | _EVAL_227;
  assign _EVAL_79 = _EVAL_117 & _EVAL_17;
  assign _EVAL_28 = _EVAL_12 & _EVAL_19;
  assign _EVAL_135 = _EVAL_186 | _EVAL_0;
  assign _EVAL_94 = _EVAL_135 == 1'h0;
  assign _EVAL_196 = _EVAL_147 | _EVAL_0;
  assign _EVAL_49 = _EVAL_196 == 1'h0;
  assign _EVAL_107 = _EVAL_165 == 1'h0;
  assign _EVAL_40 = _EVAL_227 != _EVAL_192;
  assign _EVAL_207 = _EVAL_227 != 4352'h0;
  assign _EVAL_119 = _EVAL_207 == 1'h0;
  assign _EVAL_38 = _EVAL_40 | _EVAL_119;
  assign _EVAL_131 = _EVAL_38 | _EVAL_0;
  assign _EVAL_37 = _EVAL_131 == 1'h0;
  assign _EVAL_34 = _EVAL_116 | _EVAL_0;
  assign _EVAL_153 = _EVAL_12 & _EVAL_115;
  assign _EVAL_113 = _EVAL == _EVAL_70;
  assign _EVAL_55 = _EVAL_113 | _EVAL_0;
  assign _EVAL_31 = _EVAL_55 == 1'h0;
  assign _EVAL_182 = _EVAL_214 == 1'h0;
  assign _EVAL_97 = _EVAL_138 | _EVAL_0;
  assign _EVAL_110 = _EVAL_189 == 1'h0;
  assign _EVAL_143 = _EVAL_220 | _EVAL_0;
  assign _EVAL_43 = _EVAL_11 & _EVAL_159;
  assign _EVAL_114 = _EVAL_12 & _EVAL_168;
  assign _EVAL_229 = _EVAL_2 == _EVAL_45;
  assign _EVAL_187 = _EVAL_13 == 3'h4;
  assign _EVAL_130 = $signed(_EVAL_112) & $signed(-26'sh2000);
  assign _EVAL_221 = $signed(_EVAL_130);
  assign _EVAL_139 = _EVAL_13 == 3'h3;
  assign _EVAL_133 = _EVAL_11 & _EVAL_139;
  assign _EVAL_172 = _EVAL_143 == 1'h0;
  assign _EVAL_98 = _EVAL_229 | _EVAL_0;
  assign _EVAL_44 = _EVAL_208 - 1'h1;
  assign _EVAL_90 = _EVAL_161 == 1'h0;
  assign _EVAL_202 = $signed(_EVAL_221) == $signed(26'sh0);
  assign _EVAL_47 = _EVAL_67 & _EVAL_202;
  assign _EVAL_25 = _EVAL_34 == 1'h0;
  assign _EVAL_123 = _EVAL_11 & _EVAL_187;
  assign _EVAL_198 = _EVAL_47 | _EVAL_0;
  assign _EVAL_89 = _EVAL_198 == 1'h0;
  assign _EVAL_193 = _EVAL_98 == 1'h0;
  assign _EVAL_195 = _EVAL_11 & _EVAL_213;
  assign _EVAL_39 = _EVAL_71 == 1'h0;
  assign _EVAL_32 = _EVAL_122 | _EVAL_0;
  assign _EVAL_179 = _EVAL_32 == 1'h0;
  assign _EVAL_69 = _EVAL_12 & _EVAL_86;
  assign _EVAL_93 = _EVAL_11 & _EVAL_75;
  assign _EVAL_77 = _EVAL_97 == 1'h0;
  assign _EVAL_144 = _EVAL_16 == 1'h0;
  assign _EVAL_58 = _EVAL_203 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_45 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_48 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_54 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_70 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_82 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_88 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_95 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_149 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_200 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_201 = _RAND_9[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_208 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_210 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {136{`RANDOM}};
  _EVAL_230 = _RAND_12[4351:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_233 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_145) begin
      _EVAL_45 <= _EVAL_2;
    end
    if (_EVAL_145) begin
      _EVAL_48 <= _EVAL_13;
    end
    if (_EVAL_0) begin
      _EVAL_54 <= 1'h0;
    end else begin
      if (_EVAL_224) begin
        if (_EVAL_64) begin
          _EVAL_54 <= 1'h0;
        end else begin
          _EVAL_54 <= _EVAL_108;
        end
      end
    end
    if (_EVAL_145) begin
      _EVAL_70 <= _EVAL;
    end
    if (_EVAL_0) begin
      _EVAL_82 <= 1'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_194) begin
          _EVAL_82 <= 1'h0;
        end else begin
          _EVAL_82 <= _EVAL_154;
        end
      end
    end
    if (_EVAL_145) begin
      _EVAL_88 <= _EVAL_10;
    end
    if (_EVAL_167) begin
      _EVAL_95 <= _EVAL_6;
    end
    if (_EVAL_0) begin
      _EVAL_149 <= 1'h0;
    end else begin
      if (_EVAL_224) begin
        if (_EVAL_232) begin
          _EVAL_149 <= 1'h0;
        end else begin
          _EVAL_149 <= _EVAL_228;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_200 <= 32'h0;
    end else begin
      if (_EVAL_171) begin
        _EVAL_200 <= 32'h0;
      end else begin
        _EVAL_200 <= _EVAL_170;
      end
    end
    if (_EVAL_145) begin
      _EVAL_201 <= _EVAL_9;
    end
    if (_EVAL_0) begin
      _EVAL_208 <= 1'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_148) begin
          _EVAL_208 <= 1'h0;
        end else begin
          _EVAL_208 <= _EVAL_44;
        end
      end
    end
    if (_EVAL_167) begin
      _EVAL_210 <= _EVAL_1;
    end
    if (_EVAL_0) begin
      _EVAL_230 <= 4352'h0;
    end else begin
      _EVAL_230 <= _EVAL_79;
    end
    if (_EVAL_167) begin
      _EVAL_233 <= _EVAL_7;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c90cfc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec016fa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11d9541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0505c93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85e19fdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcabb8fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90baf95e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1fccef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83bad5e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28d036e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b86af47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f72f3dd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4abfdd60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(963ba72e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52375a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb5097d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84464999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(699db296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9735f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f24fc19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2bc7242)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef71a0f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0aa0ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ef3f450)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ee5306)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61bdb6fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95168fff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffb18b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c39b515b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87b16cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cc0e4c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2449ba4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86f8d6e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b008805)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e0cb892)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94bdbe9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddc81708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e749f7ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e254fe65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5659fbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39e02354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2768722)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26a5d75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67251080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(550779d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f7e004b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc26366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f401985)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c4de0d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfe13d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba41293e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(273aba98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffe33829)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65aebf6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7fc4143)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4ab71f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6adeff0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd5308a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(976132ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588d7d0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ee4470)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6658e10c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(758bba49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c80c1df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea886a22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27b700d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80bac186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d2dd058)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c11c6f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f88923f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6e28fc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3e6aad0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
