//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_304_assert(
  input  [1:0]  _EVAL_1,
  input  [2:0]  _EVAL_23,
  input         _EVAL_53,
  input  [11:0] _EVAL_102,
  input         _EVAL_146,
  input         _EVAL_155,
  input  [1:0]  _EVAL_252,
  input         _EVAL_1073,
  input         _EVAL_352,
  input         _EVAL_2099,
  input         _EVAL_1186,
  input         _EVAL_1014,
  input         _EVAL_1722,
  input         _EVAL_1310,
  input         _EVAL_898,
  input         _EVAL_1902,
  input         _EVAL_739,
  input         _EVAL_1937,
  input  [31:0] _EVAL_579,
  input         _EVAL_2017,
  input         _EVAL_826,
  input         _EVAL_283,
  input         _EVAL_1767,
  input         _EVAL_755,
  input         _EVAL_569,
  input         _EVAL_1031,
  input         _EVAL_1752,
  input         _EVAL_1291,
  input         _EVAL_2208,
  input         _EVAL_262,
  input         _EVAL_1833,
  input         _EVAL_1297,
  input         _EVAL_2143,
  input         _EVAL_1713,
  input         _EVAL_772,
  input         _EVAL_531,
  input         _EVAL_1559,
  input         _EVAL_1746,
  input         _EVAL_484,
  input         _EVAL_666,
  input         _EVAL_1358,
  input         _EVAL_2066,
  input         _EVAL_1374,
  input         _EVAL_800,
  input         _EVAL_1617,
  input         _EVAL_1437,
  input         _EVAL_316,
  input         _EVAL_1386,
  input         _EVAL_1560,
  input         _EVAL_677,
  input         _EVAL_425,
  input         _EVAL_323,
  input         _EVAL_1657,
  input         _EVAL_1872,
  input         _EVAL_596,
  input         _EVAL_212,
  input         _EVAL_1213,
  input         _EVAL_1396,
  input         _EVAL_237,
  input         _EVAL_780,
  input         _EVAL_539,
  input         _EVAL_1647,
  input         _EVAL_1418,
  input         _EVAL_1285,
  input         _EVAL_1864,
  input         _EVAL_747,
  input         _EVAL_2155,
  input         _EVAL_1500,
  input         _EVAL_843,
  input         _EVAL_1394
);
  wire  _EVAL_1971;
  wire  _EVAL_1868;
  wire  _EVAL_712;
  wire  _EVAL_1726;
  wire  _EVAL_1214;
  wire  _EVAL_1727;
  wire  _EVAL_1537;
  wire  _EVAL_1846;
  wire  _EVAL_2096;
  wire  _EVAL_291;
  wire  _EVAL_2020;
  wire  _EVAL_1546;
  wire  _EVAL_2233;
  wire  _EVAL_875;
  wire  _EVAL_382;
  wire  _EVAL_685;
  wire  _EVAL_1250;
  wire  _EVAL_2189;
  wire  _EVAL_1314;
  wire  _EVAL_1119;
  wire  _EVAL_398;
  wire  _EVAL_1309;
  wire  _EVAL_1205;
  wire  _EVAL_640;
  wire  _EVAL_1002;
  wire  _EVAL_696;
  wire  _EVAL_429;
  wire  _EVAL_1434;
  wire  _EVAL_301;
  wire  _EVAL_671;
  wire  _EVAL_1070;
  wire  _EVAL_1918;
  wire  _EVAL_1841;
  wire  _EVAL_2212;
  wire  _EVAL_1911;
  wire  _EVAL_1477;
  wire  _EVAL_2040;
  wire  _EVAL_200;
  wire  _EVAL_880;
  wire  _EVAL_983;
  wire  _EVAL_1460;
  wire  _EVAL_1267;
  wire  _EVAL_1599;
  wire  _EVAL_1787;
  wire  _EVAL_921;
  wire  _EVAL_493;
  wire  _EVAL_1703;
  wire  _EVAL_966;
  wire  _EVAL_1409;
  wire  _EVAL_1341;
  wire  _EVAL_623;
  wire  _EVAL_335;
  wire  _EVAL_1301;
  wire  _EVAL_191;
  wire  _EVAL_841;
  wire  _EVAL_444;
  wire  _EVAL_758;
  wire  _EVAL_2178;
  wire  _EVAL_1037;
  wire  _EVAL_1987;
  wire  _EVAL_1116;
  wire  _EVAL_629;
  wire  _EVAL_515;
  wire  _EVAL_1036;
  wire  _EVAL_454;
  wire  _EVAL_668;
  wire  _EVAL_272;
  wire  _EVAL_618;
  wire  _EVAL_1510;
  wire  _EVAL_1653;
  wire  _EVAL_1768;
  wire  _EVAL_1802;
  wire  _EVAL_1897;
  wire  _EVAL_1435;
  wire  _EVAL_748;
  wire  _EVAL_1511;
  wire  _EVAL_1574;
  wire  _EVAL_1169;
  wire  _EVAL_1604;
  wire  _EVAL_1542;
  wire  _EVAL_1175;
  wire  _EVAL_590;
  wire  _EVAL_1089;
  wire  _EVAL_588;
  wire  _EVAL_2022;
  wire  _EVAL_1313;
  wire  _EVAL_2166;
  wire  _EVAL_560;
  wire  _EVAL_1870;
  wire  _EVAL_1690;
  wire  _EVAL_1337;
  wire  _EVAL_2055;
  wire  _EVAL_319;
  wire  _EVAL_1319;
  wire  _EVAL_633;
  wire  _EVAL_2037;
  wire  _EVAL_423;
  wire  _EVAL_1206;
  wire  _EVAL_1252;
  wire  _EVAL_234;
  wire  _EVAL_1462;
  wire [1:0] _EVAL_536;
  wire [1:0] _EVAL_754;
  wire [2:0] _EVAL_1224;
  wire  _EVAL_1614;
  wire  _EVAL_1637;
  wire  _EVAL_1268;
  wire  _EVAL_788;
  wire  _EVAL_1187;
  wire  _EVAL_833;
  wire  _EVAL_1699;
  wire  _EVAL_2060;
  wire  _EVAL_2083;
  wire  _EVAL_734;
  wire  _EVAL_2045;
  wire  _EVAL_1227;
  wire  _EVAL_1766;
  wire  _EVAL_468;
  wire  _EVAL_1303;
  wire  _EVAL_1513;
  wire  _EVAL_1221;
  wire  _EVAL_1375;
  wire  _EVAL_1894;
  wire  _EVAL_1197;
  wire  _EVAL_553;
  wire  _EVAL_1209;
  wire  _EVAL_355;
  wire  _EVAL_2206;
  wire  _EVAL_1215;
  wire  _EVAL_727;
  wire  _EVAL_915;
  wire  _EVAL_1996;
  wire  _EVAL_701;
  wire  _EVAL_1778;
  wire  _EVAL_218;
  wire  _EVAL_469;
  wire  _EVAL_1755;
  wire  _EVAL_834;
  wire  _EVAL_1069;
  wire  _EVAL_472;
  wire  _EVAL_1530;
  wire  _EVAL_1179;
  wire  _EVAL_840;
  wire  _EVAL_1066;
  wire  _EVAL_1113;
  wire  _EVAL_613;
  wire  _EVAL_1057;
  wire  _EVAL_1230;
  wire  _EVAL_938;
  wire  _EVAL_933;
  wire  _EVAL_332;
  wire  _EVAL_1867;
  wire  _EVAL_911;
  wire  _EVAL_791;
  wire  _EVAL_585;
  wire  _EVAL_1154;
  wire  _EVAL_690;
  wire  _EVAL_1998;
  wire  _EVAL_1378;
  wire  _EVAL_568;
  wire  _EVAL_406;
  wire  _EVAL_614;
  wire  _EVAL_1299;
  wire  _EVAL_2134;
  wire  _EVAL_563;
  wire  _EVAL_723;
  wire  _EVAL_202;
  wire  _EVAL_1370;
  wire  _EVAL_433;
  wire  _EVAL_480;
  wire  _EVAL_2053;
  wire  _EVAL_288;
  wire  _EVAL_757;
  wire  _EVAL_1360;
  wire  _EVAL_1549;
  wire  _EVAL_600;
  wire  _EVAL_764;
  wire  _EVAL_524;
  wire  _EVAL_1760;
  wire  _EVAL_582;
  wire  _EVAL_837;
  wire  _EVAL_1933;
  wire  _EVAL_1716;
  wire  _EVAL_1944;
  wire  _EVAL_1192;
  wire  _EVAL_1195;
  wire  _EVAL_2051;
  wire  _EVAL_410;
  wire  _EVAL_774;
  wire  _EVAL_575;
  wire  _EVAL_1744;
  wire  _EVAL_1000;
  wire  _EVAL_1274;
  wire  _EVAL_1892;
  wire  _EVAL_2014;
  wire  _EVAL_1612;
  wire  _EVAL_839;
  wire  _EVAL_1263;
  wire  _EVAL_598;
  wire  _EVAL_2119;
  wire  _EVAL_586;
  wire  _EVAL_2109;
  wire  _EVAL_1857;
  wire  _EVAL_372;
  wire  _EVAL_637;
  wire  _EVAL_2196;
  wire  _EVAL_1039;
  wire  _EVAL_894;
  wire  _EVAL_1006;
  wire  _EVAL_1173;
  wire  _EVAL_501;
  wire  _EVAL_687;
  wire  _EVAL_2034;
  wire  _EVAL_2198;
  wire  _EVAL_1806;
  wire  _EVAL_235;
  wire  _EVAL_1290;
  wire  _EVAL_1706;
  wire  _EVAL_1280;
  wire  _EVAL_2093;
  wire  _EVAL_2231;
  wire  _EVAL_1860;
  wire  _EVAL_1701;
  wire  _EVAL_366;
  wire  _EVAL_2128;
  wire  _EVAL_1327;
  wire  _EVAL_1429;
  wire  _EVAL_1821;
  wire  _EVAL_1622;
  wire  _EVAL_1738;
  wire  _EVAL_498;
  wire  _EVAL_627;
  wire  _EVAL_879;
  wire  _EVAL_1858;
  wire  _EVAL_1817;
  wire  _EVAL_1670;
  wire  _EVAL_245;
  wire  _EVAL_172;
  wire  _EVAL_1109;
  wire  _EVAL_2075;
  wire  _EVAL_1304;
  wire  _EVAL_818;
  wire  _EVAL_2107;
  wire  _EVAL_766;
  wire  _EVAL_1325;
  wire  _EVAL_2026;
  wire  _EVAL_1810;
  wire  _EVAL_2016;
  wire  _EVAL_562;
  wire  _EVAL_1596;
  wire  _EVAL_413;
  wire  _EVAL_917;
  wire  _EVAL_1198;
  wire  _EVAL_1140;
  wire  _EVAL_1450;
  wire  _EVAL_1527;
  wire  _EVAL_1686;
  wire  _EVAL_1265;
  wire  _EVAL_721;
  wire  _EVAL_1654;
  wire  _EVAL_453;
  wire  _EVAL_1687;
  wire  _EVAL_695;
  wire  _EVAL_1776;
  wire  _EVAL_241;
  wire  _EVAL_554;
  wire  _EVAL_226;
  wire  _EVAL_1643;
  wire  _EVAL_1528;
  wire  _EVAL_1962;
  wire  _EVAL_610;
  wire  _EVAL_1829;
  wire  _EVAL_420;
  wire  _EVAL_789;
  wire  _EVAL_1915;
  wire  _EVAL_401;
  wire  _EVAL_1258;
  wire  _EVAL_593;
  wire  _EVAL_1323;
  wire  _EVAL_934;
  wire  _EVAL_1240;
  wire  _EVAL_1335;
  wire  _EVAL_1257;
  wire  _EVAL_1581;
  wire  _EVAL_927;
  wire  _EVAL_1412;
  wire  _EVAL_393;
  wire  _EVAL_1013;
  wire  _EVAL_1665;
  wire  _EVAL_447;
  wire  _EVAL_664;
  wire  _EVAL_2088;
  wire  _EVAL_1992;
  wire  _EVAL_1316;
  wire  _EVAL_628;
  wire  _EVAL_929;
  wire  _EVAL_1185;
  wire  _EVAL_1270;
  wire  _EVAL_1758;
  wire  _EVAL_481;
  wire  _EVAL_1990;
  wire  _EVAL_2111;
  wire  _EVAL_603;
  wire  _EVAL_544;
  wire  _EVAL_1682;
  wire  _EVAL_1222;
  wire  _EVAL_2242;
  wire  _EVAL_1753;
  wire  _EVAL_943;
  wire  _EVAL_1415;
  wire  _EVAL_1218;
  wire  _EVAL_1705;
  wire  _EVAL_2072;
  wire  _EVAL_945;
  wire  _EVAL_1041;
  wire  _EVAL_1237;
  wire  _EVAL_1839;
  wire  _EVAL_1958;
  wire  _EVAL_238;
  wire  _EVAL_1422;
  wire  _EVAL_1204;
  wire  _EVAL_2171;
  wire  _EVAL_661;
  wire  _EVAL_856;
  wire  _EVAL_1749;
  wire  _EVAL_1728;
  wire  _EVAL_1844;
  wire  _EVAL_1522;
  wire  _EVAL_1333;
  wire  _EVAL_768;
  wire  _EVAL_1245;
  wire  _EVAL_2000;
  wire  _EVAL_989;
  wire  _EVAL_1834;
  wire  _EVAL_972;
  wire  _EVAL_1798;
  wire  _EVAL_642;
  wire  _EVAL_799;
  wire  _EVAL_179;
  wire  _EVAL_704;
  wire  _EVAL_1675;
  wire  _EVAL_725;
  wire  _EVAL_1485;
  wire  _EVAL_2061;
  wire  _EVAL_2148;
  wire  _EVAL_965;
  wire  _EVAL_1660;
  wire  _EVAL_815;
  wire  _EVAL_1284;
  wire  _EVAL_1572;
  wire  _EVAL_1497;
  wire  _EVAL_1071;
  wire  _EVAL_617;
  wire  _EVAL_494;
  wire  _EVAL_183;
  wire  _EVAL_1591;
  wire  _EVAL_2052;
  wire  _EVAL_1399;
  wire  _EVAL_1611;
  wire  _EVAL_1148;
  wire  _EVAL_289;
  wire  _EVAL_1812;
  wire  _EVAL_414;
  wire  _EVAL_1757;
  wire  _EVAL_367;
  wire  _EVAL_221;
  wire  _EVAL_391;
  wire  _EVAL_1732;
  wire  _EVAL_1351;
  wire  _EVAL_986;
  wire  _EVAL_1080;
  wire  _EVAL_1007;
  wire  _EVAL_853;
  wire  _EVAL_1975;
  wire  _EVAL_1397;
  wire  _EVAL_1677;
  wire  _EVAL_706;
  wire  _EVAL_1935;
  wire  _EVAL_838;
  wire  _EVAL_1243;
  wire  _EVAL_698;
  wire  _EVAL_1903;
  wire  _EVAL_1480;
  wire  _EVAL_1135;
  wire  _EVAL_2098;
  wire  _EVAL_1916;
  wire  _EVAL_499;
  wire  _EVAL_519;
  wire  _EVAL_1413;
  wire  _EVAL_1883;
  assign _EVAL_1971 = _EVAL_352 | _EVAL_2099;
  assign _EVAL_1868 = _EVAL_1971 | _EVAL_1186;
  assign _EVAL_712 = _EVAL_1868 & _EVAL_1014;
  assign _EVAL_1726 = _EVAL_102 == 12'hb13;
  assign _EVAL_1214 = _EVAL_102 == 12'h329;
  assign _EVAL_1727 = _EVAL_102 == 12'h337;
  assign _EVAL_1537 = _EVAL_102 == 12'hc13;
  assign _EVAL_1846 = _EVAL_23 == 3'h2;
  assign _EVAL_2096 = _EVAL_102 == 12'hc18;
  assign _EVAL_291 = _EVAL_1846 & _EVAL_2096;
  assign _EVAL_2020 = _EVAL_1868 & _EVAL_531;
  assign _EVAL_1546 = _EVAL_102 == 12'hb9c;
  assign _EVAL_2233 = _EVAL_102 == 12'hc06;
  assign _EVAL_875 = _EVAL_1846 & _EVAL_2233;
  assign _EVAL_382 = _EVAL_102 == 12'hb9d;
  assign _EVAL_685 = _EVAL_102 == 12'hc9a;
  assign _EVAL_1250 = _EVAL_1846 & _EVAL_685;
  assign _EVAL_2189 = _EVAL_102 == 12'h339;
  assign _EVAL_1314 = _EVAL_102 == 12'hc08;
  assign _EVAL_1119 = _EVAL_579 == 32'h80000007;
  assign _EVAL_398 = _EVAL_102 == 12'h333;
  assign _EVAL_1309 = _EVAL_1868 & _EVAL_398;
  assign _EVAL_1205 = _EVAL_102 == 12'hc9d;
  assign _EVAL_640 = _EVAL_102 == 12'hc10;
  assign _EVAL_1002 = _EVAL_1846 & _EVAL_640;
  assign _EVAL_696 = _EVAL_1868 & _EVAL_2208;
  assign _EVAL_429 = _EVAL_1868 & _EVAL_2017;
  assign _EVAL_1434 = _EVAL_1846 & _EVAL_1205;
  assign _EVAL_301 = _EVAL_102 == 12'hc0f;
  assign _EVAL_671 = _EVAL_1846 & _EVAL_301;
  assign _EVAL_1070 = _EVAL_102 == 12'hb92;
  assign _EVAL_1918 = _EVAL_1868 & _EVAL_1070;
  assign _EVAL_1841 = _EVAL_102 == 12'hb8a;
  assign _EVAL_2212 = _EVAL_1868 & _EVAL_1841;
  assign _EVAL_1911 = _EVAL_102 == 12'hc86;
  assign _EVAL_1477 = _EVAL_102 == 12'hb8f;
  assign _EVAL_2040 = _EVAL_102 == 12'hc0c;
  assign _EVAL_200 = _EVAL_102 == 12'hb88;
  assign _EVAL_880 = _EVAL_1868 & _EVAL_200;
  assign _EVAL_983 = _EVAL_102 == 12'h3bf;
  assign _EVAL_1460 = _EVAL_1868 & _EVAL_983;
  assign _EVAL_1267 = _EVAL_102 == 12'hb0f;
  assign _EVAL_1599 = _EVAL_102 == 12'hc17;
  assign _EVAL_1787 = _EVAL_1846 & _EVAL_1599;
  assign _EVAL_921 = _EVAL_102 == 12'hb14;
  assign _EVAL_493 = _EVAL_1868 & _EVAL_921;
  assign _EVAL_1703 = _EVAL_102 == 12'h332;
  assign _EVAL_966 = _EVAL_102 == 12'hb0e;
  assign _EVAL_1409 = _EVAL_1868 & _EVAL_966;
  assign _EVAL_1341 = _EVAL_579 == 32'h2;
  assign _EVAL_623 = _EVAL_1937 & _EVAL_1341;
  assign _EVAL_335 = _EVAL_102 == 12'h331;
  assign _EVAL_1301 = _EVAL_102 == 12'hc92;
  assign _EVAL_191 = _EVAL_102 == 12'hc9e;
  assign _EVAL_841 = _EVAL_579 == 32'h3;
  assign _EVAL_444 = _EVAL_1868 & _EVAL_1833;
  assign _EVAL_758 = _EVAL_102 == 12'hc98;
  assign _EVAL_2178 = _EVAL_1846 & _EVAL_758;
  assign _EVAL_1037 = _EVAL_102 == 12'hc9c;
  assign _EVAL_1987 = _EVAL_579 == 32'h4;
  assign _EVAL_1116 = _EVAL_1937 & _EVAL_1987;
  assign _EVAL_629 = _EVAL_102 == 12'hb94;
  assign _EVAL_515 = _EVAL_1868 & _EVAL_629;
  assign _EVAL_1036 = _EVAL_102 == 12'hb9a;
  assign _EVAL_454 = _EVAL_1868 & _EVAL_1036;
  assign _EVAL_668 = _EVAL_102 == 12'hb85;
  assign _EVAL_272 = _EVAL_1868 & _EVAL_668;
  assign _EVAL_618 = _EVAL_102 == 12'h32b;
  assign _EVAL_1510 = _EVAL_1868 & _EVAL_618;
  assign _EVAL_1653 = _EVAL_102 == 12'hb91;
  assign _EVAL_1768 = _EVAL_102 == 12'hc0a;
  assign _EVAL_1802 = _EVAL_102 == 12'hb16;
  assign _EVAL_1897 = _EVAL_1868 & _EVAL_1802;
  assign _EVAL_1435 = _EVAL_102 == 12'hc8d;
  assign _EVAL_748 = _EVAL_102 == 12'hb0c;
  assign _EVAL_1511 = _EVAL_1868 & _EVAL_748;
  assign _EVAL_1574 = _EVAL_252 > 2'h0;
  assign _EVAL_1169 = _EVAL_1574 | _EVAL_146;
  assign _EVAL_1604 = _EVAL_102 == 12'h33a;
  assign _EVAL_1542 = _EVAL_102 == 12'hc09;
  assign _EVAL_1175 = _EVAL_102 == 12'hc96;
  assign _EVAL_590 = _EVAL_1846 & _EVAL_1175;
  assign _EVAL_1089 = _EVAL_102 == 12'hc93;
  assign _EVAL_588 = _EVAL_1846 & _EVAL_1089;
  assign _EVAL_2022 = _EVAL_579 == 32'h7;
  assign _EVAL_1313 = _EVAL_102 == 12'h335;
  assign _EVAL_2166 = _EVAL_1868 & _EVAL_1313;
  assign _EVAL_560 = _EVAL_1868 & _EVAL_1477;
  assign _EVAL_1870 = _EVAL_102 == 12'hc89;
  assign _EVAL_1690 = _EVAL_1846 & _EVAL_1870;
  assign _EVAL_1337 = _EVAL_102 == 12'hc8f;
  assign _EVAL_2055 = _EVAL_579 == 32'h8000000b;
  assign _EVAL_319 = _EVAL_1937 & _EVAL_2055;
  assign _EVAL_1319 = _EVAL_102 == 12'hc88;
  assign _EVAL_633 = _EVAL_1868 & _EVAL_1285;
  assign _EVAL_2037 = _EVAL_102 == 12'h336;
  assign _EVAL_423 = _EVAL_1868 & _EVAL_2037;
  assign _EVAL_1206 = _EVAL_102 == 12'hb05;
  assign _EVAL_1252 = _EVAL_1868 & _EVAL_1206;
  assign _EVAL_234 = _EVAL_102 == 12'h33c;
  assign _EVAL_1462 = _EVAL_1868 & _EVAL_234;
  assign _EVAL_536 = _EVAL_898 + _EVAL_1902;
  assign _EVAL_754 = _EVAL_739 + _EVAL_155;
  assign _EVAL_1224 = _EVAL_536 + _EVAL_754;
  assign _EVAL_1614 = _EVAL_1224 <= 3'h1;
  assign _EVAL_1637 = _EVAL_1614 | _EVAL_146;
  assign _EVAL_1268 = _EVAL_102 == 12'h326;
  assign _EVAL_788 = _EVAL_1868 & _EVAL_1268;
  assign _EVAL_1187 = _EVAL_102 == 12'hb0d;
  assign _EVAL_833 = _EVAL_1868 & _EVAL_1437;
  assign _EVAL_1699 = _EVAL_102 == 12'hb87;
  assign _EVAL_2060 = _EVAL_1868 & _EVAL_1699;
  assign _EVAL_2083 = _EVAL_102 == 12'hb95;
  assign _EVAL_734 = _EVAL_102 == 12'hb1b;
  assign _EVAL_2045 = _EVAL_1868 & _EVAL_734;
  assign _EVAL_1227 = _EVAL_102 == 12'hb98;
  assign _EVAL_1766 = _EVAL_1868 & _EVAL_1227;
  assign _EVAL_468 = _EVAL_1868 & _EVAL_1267;
  assign _EVAL_1303 = _EVAL_102 == 12'hc95;
  assign _EVAL_1513 = _EVAL_1846 & _EVAL_1303;
  assign _EVAL_1221 = _EVAL_102 == 12'h3b8;
  assign _EVAL_1375 = _EVAL_102 == 12'h33e;
  assign _EVAL_1894 = _EVAL_1868 & _EVAL_1375;
  assign _EVAL_1197 = _EVAL_102 == 12'hc1c;
  assign _EVAL_553 = _EVAL_1846 & _EVAL_1197;
  assign _EVAL_1209 = _EVAL_102 == 12'hc8e;
  assign _EVAL_355 = _EVAL_1868 & _EVAL_2143;
  assign _EVAL_2206 = _EVAL_102 == 12'hb17;
  assign _EVAL_1215 = _EVAL_102 == 12'hb0a;
  assign _EVAL_727 = _EVAL_102 == 12'hb99;
  assign _EVAL_915 = _EVAL_1868 & _EVAL_755;
  assign _EVAL_1996 = _EVAL_102 == 12'hc19;
  assign _EVAL_701 = _EVAL_1846 & _EVAL_1996;
  assign _EVAL_1778 = _EVAL_102 == 12'hb07;
  assign _EVAL_218 = _EVAL_1868 & _EVAL_1778;
  assign _EVAL_469 = _EVAL_102 == 12'hc9f;
  assign _EVAL_1755 = _EVAL_102 == 12'h32c;
  assign _EVAL_834 = _EVAL_102 == 12'h334;
  assign _EVAL_1069 = _EVAL_1169 == 1'h0;
  assign _EVAL_472 = _EVAL_102 == 12'hb93;
  assign _EVAL_1530 = _EVAL_1868 & _EVAL_472;
  assign _EVAL_1179 = _EVAL_1868 & _EVAL_727;
  assign _EVAL_840 = _EVAL_102 == 12'h3a2;
  assign _EVAL_1066 = _EVAL_1868 & _EVAL_840;
  assign _EVAL_1113 = _EVAL_102 == 12'hc8c;
  assign _EVAL_613 = _EVAL_1846 & _EVAL_1113;
  assign _EVAL_1057 = _EVAL_1 <= 2'h1;
  assign _EVAL_1230 = _EVAL_1394 | _EVAL_1057;
  assign _EVAL_938 = _EVAL_102 == 12'hc14;
  assign _EVAL_933 = _EVAL_1637 == 1'h0;
  assign _EVAL_332 = _EVAL_102 == 12'hc91;
  assign _EVAL_1867 = _EVAL_1846 & _EVAL_332;
  assign _EVAL_911 = _EVAL_102 == 12'hc1f;
  assign _EVAL_791 = _EVAL_1846 & _EVAL_911;
  assign _EVAL_585 = _EVAL_102 == 12'hb08;
  assign _EVAL_1154 = _EVAL_1868 & _EVAL_585;
  assign _EVAL_690 = _EVAL_102 == 12'h33f;
  assign _EVAL_1998 = _EVAL_102 == 12'h32f;
  assign _EVAL_1378 = _EVAL_102 == 12'hb96;
  assign _EVAL_568 = _EVAL_102 == 12'h328;
  assign _EVAL_406 = _EVAL_1868 & _EVAL_568;
  assign _EVAL_614 = _EVAL_1868 & _EVAL_1386;
  assign _EVAL_1299 = _EVAL_1868 & _EVAL_1767;
  assign _EVAL_2134 = _EVAL_1868 & _EVAL_1998;
  assign _EVAL_563 = _EVAL_102 == 12'hc1a;
  assign _EVAL_723 = _EVAL_102 == 12'h325;
  assign _EVAL_202 = _EVAL_1868 & _EVAL_723;
  assign _EVAL_1370 = _EVAL_1846 & _EVAL_1542;
  assign _EVAL_433 = _EVAL_102 == 12'h338;
  assign _EVAL_480 = _EVAL_1868 & _EVAL_433;
  assign _EVAL_2053 = _EVAL_102 == 12'h32d;
  assign _EVAL_288 = _EVAL_1868 & _EVAL_2053;
  assign _EVAL_757 = _EVAL_1868 & _EVAL_677;
  assign _EVAL_1360 = _EVAL_102 == 12'hc99;
  assign _EVAL_1549 = _EVAL_579 == 32'h5;
  assign _EVAL_600 = _EVAL_1937 & _EVAL_1549;
  assign _EVAL_764 = _EVAL_1846 & _EVAL_191;
  assign _EVAL_524 = _EVAL_102 == 12'hb0b;
  assign _EVAL_1760 = _EVAL_1868 & _EVAL_524;
  assign _EVAL_582 = _EVAL_1868 & _EVAL_1653;
  assign _EVAL_837 = _EVAL_1937 & _EVAL_841;
  assign _EVAL_1933 = _EVAL_102 == 12'hb15;
  assign _EVAL_1716 = _EVAL_1868 & _EVAL_1933;
  assign _EVAL_1944 = _EVAL_102 == 12'hffc;
  assign _EVAL_1192 = _EVAL_102 == 12'hc85;
  assign _EVAL_1195 = _EVAL_1846 & _EVAL_1192;
  assign _EVAL_2051 = _EVAL_1868 & _EVAL_2189;
  assign _EVAL_410 = _EVAL_1868 & _EVAL_1291;
  assign _EVAL_774 = _EVAL_1937 & _EVAL_1119;
  assign _EVAL_575 = _EVAL_102 == 12'hb8c;
  assign _EVAL_1744 = _EVAL_102 == 12'hb89;
  assign _EVAL_1000 = _EVAL_102 == 12'hc8b;
  assign _EVAL_1274 = _EVAL_1846 & _EVAL_1000;
  assign _EVAL_1892 = _EVAL_102 == 12'hc94;
  assign _EVAL_2014 = _EVAL_1846 & _EVAL_1892;
  assign _EVAL_1612 = _EVAL_102 == 12'hb1d;
  assign _EVAL_839 = _EVAL_1846 & _EVAL_1560;
  assign _EVAL_1263 = _EVAL_102 == 12'hb90;
  assign _EVAL_598 = _EVAL_102 == 12'hc97;
  assign _EVAL_2119 = _EVAL_1846 & _EVAL_598;
  assign _EVAL_586 = _EVAL_1868 & _EVAL_1617;
  assign _EVAL_2109 = _EVAL_102 == 12'hb18;
  assign _EVAL_1857 = _EVAL_579 == 32'hb;
  assign _EVAL_372 = _EVAL_1937 & _EVAL_1857;
  assign _EVAL_637 = _EVAL_1868 & _EVAL_1187;
  assign _EVAL_2196 = _EVAL_1868 & _EVAL_1727;
  assign _EVAL_1039 = _EVAL_1868 & _EVAL_1310;
  assign _EVAL_894 = _EVAL_102 == 12'hb97;
  assign _EVAL_1006 = _EVAL_1868 & _EVAL_894;
  assign _EVAL_1173 = _EVAL_1868 & _EVAL_1358;
  assign _EVAL_501 = _EVAL_102 == 12'h3be;
  assign _EVAL_687 = _EVAL_102 == 12'h327;
  assign _EVAL_2034 = _EVAL_102 == 12'h3bb;
  assign _EVAL_2198 = _EVAL_102 == 12'hc05;
  assign _EVAL_1806 = _EVAL_1 == 2'h0;
  assign _EVAL_235 = _EVAL_102 == 12'hc87;
  assign _EVAL_1290 = _EVAL_102 == 12'hc9b;
  assign _EVAL_1706 = _EVAL_1868 & _EVAL_1559;
  assign _EVAL_1280 = _EVAL_1868 & _EVAL_1546;
  assign _EVAL_2093 = _EVAL_1868 & _EVAL_539;
  assign _EVAL_2231 = _EVAL_1846 & _EVAL_1435;
  assign _EVAL_1860 = _EVAL_1868 & _EVAL_1213;
  assign _EVAL_1701 = _EVAL_102 == 12'hc12;
  assign _EVAL_366 = _EVAL_1846 & _EVAL_1701;
  assign _EVAL_2128 = _EVAL_102 == 12'h3ba;
  assign _EVAL_1327 = _EVAL_1868 & _EVAL_2128;
  assign _EVAL_1429 = _EVAL_1868 & _EVAL_834;
  assign _EVAL_1821 = _EVAL_102 == 12'hc15;
  assign _EVAL_1622 = _EVAL_1846 & _EVAL_1821;
  assign _EVAL_1738 = _EVAL_1868 & _EVAL_1755;
  assign _EVAL_498 = _EVAL_1846 & _EVAL_747;
  assign _EVAL_627 = _EVAL_1868 & _EVAL_1263;
  assign _EVAL_879 = _EVAL_102 == 12'hb9e;
  assign _EVAL_1858 = _EVAL_1868 & _EVAL_1221;
  assign _EVAL_1817 = _EVAL_1846 & _EVAL_2066;
  assign _EVAL_1670 = _EVAL_102 == 12'h3a3;
  assign _EVAL_245 = _EVAL_1868 & _EVAL_1670;
  assign _EVAL_172 = _EVAL_1868 & _EVAL_666;
  assign _EVAL_1109 = _EVAL_1846 & _EVAL_235;
  assign _EVAL_2075 = _EVAL_102 == 12'h330;
  assign _EVAL_1304 = _EVAL_1868 & _EVAL_2075;
  assign _EVAL_818 = _EVAL_1868 & _EVAL_1215;
  assign _EVAL_2107 = _EVAL_1846 & _EVAL_1944;
  assign _EVAL_766 = _EVAL_1846 & _EVAL_2040;
  assign _EVAL_1325 = _EVAL_102 == 12'h3bd;
  assign _EVAL_2026 = _EVAL_102 == 12'hb11;
  assign _EVAL_1810 = _EVAL_1868 & _EVAL_2026;
  assign _EVAL_2016 = _EVAL_1846 & _EVAL_212;
  assign _EVAL_562 = _EVAL_1868 & _EVAL_1325;
  assign _EVAL_1596 = _EVAL_1868 & _EVAL_1396;
  assign _EVAL_413 = _EVAL_1846 & _EVAL_323;
  assign _EVAL_917 = _EVAL_1868 & _EVAL_501;
  assign _EVAL_1198 = _EVAL_102 == 12'hb06;
  assign _EVAL_1140 = _EVAL_1868 & _EVAL_1647;
  assign _EVAL_1450 = _EVAL_102 == 12'hb9f;
  assign _EVAL_1527 = _EVAL_1868 & _EVAL_1450;
  assign _EVAL_1686 = _EVAL_579 == 32'h6;
  assign _EVAL_1265 = _EVAL_1937 & _EVAL_1686;
  assign _EVAL_721 = _EVAL_1846 & _EVAL_1768;
  assign _EVAL_1654 = _EVAL_1868 & _EVAL_1872;
  assign _EVAL_453 = _EVAL_1868 & _EVAL_826;
  assign _EVAL_1687 = _EVAL_102 == 12'hc07;
  assign _EVAL_695 = _EVAL_102 == 12'hb8b;
  assign _EVAL_1776 = _EVAL_1073 == 1'h0;
  assign _EVAL_241 = _EVAL_1846 & _EVAL_596;
  assign _EVAL_554 = _EVAL_102 == 12'hc0b;
  assign _EVAL_226 = _EVAL_102 == 12'hb86;
  assign _EVAL_1643 = _EVAL_102 == 12'hb19;
  assign _EVAL_1528 = _EVAL_1868 & _EVAL_1643;
  assign _EVAL_1962 = _EVAL_1868 & _EVAL_1864;
  assign _EVAL_610 = _EVAL_1846 & _EVAL_800;
  assign _EVAL_1829 = _EVAL_102 == 12'hb8e;
  assign _EVAL_420 = _EVAL_1868 & _EVAL_1829;
  assign _EVAL_789 = _EVAL_102 == 12'h3bc;
  assign _EVAL_1915 = _EVAL_1846 & _EVAL_2198;
  assign _EVAL_401 = _EVAL_1868 & _EVAL_1604;
  assign _EVAL_1258 = _EVAL_1846 & _EVAL_1314;
  assign _EVAL_593 = _EVAL_1868 & _EVAL_772;
  assign _EVAL_1323 = _EVAL_102 == 12'hc1d;
  assign _EVAL_934 = _EVAL_1846 & _EVAL_1323;
  assign _EVAL_1240 = _EVAL_1846 & _EVAL_1290;
  assign _EVAL_1335 = _EVAL_1846 & _EVAL_2155;
  assign _EVAL_1257 = _EVAL_102 == 12'h32a;
  assign _EVAL_1581 = _EVAL_1868 & _EVAL_1257;
  assign _EVAL_927 = _EVAL_579 == 32'h80000003;
  assign _EVAL_1412 = _EVAL_1937 & _EVAL_927;
  assign _EVAL_393 = _EVAL_1868 & _EVAL_1703;
  assign _EVAL_1013 = _EVAL_1868 & _EVAL_1713;
  assign _EVAL_1665 = _EVAL_102 == 12'hc1e;
  assign _EVAL_447 = _EVAL_1846 & _EVAL_1665;
  assign _EVAL_664 = _EVAL_102 == 12'hb1f;
  assign _EVAL_2088 = _EVAL_102 == 12'hc0e;
  assign _EVAL_1992 = _EVAL_1868 & _EVAL_687;
  assign _EVAL_1316 = _EVAL_1868 & _EVAL_1214;
  assign _EVAL_628 = _EVAL_102 == 12'hc16;
  assign _EVAL_929 = _EVAL_1868 & _EVAL_1418;
  assign _EVAL_1185 = _EVAL_102 == 12'hb1e;
  assign _EVAL_1270 = _EVAL_1868 & _EVAL_1185;
  assign _EVAL_1758 = _EVAL_102 == 12'hb8d;
  assign _EVAL_481 = _EVAL_1846 & _EVAL_628;
  assign _EVAL_1990 = _EVAL_1846 & _EVAL_1319;
  assign _EVAL_2111 = _EVAL_1846 & _EVAL_938;
  assign _EVAL_603 = _EVAL_1868 & _EVAL_2083;
  assign _EVAL_544 = _EVAL_1868 & _EVAL_1722;
  assign _EVAL_1682 = _EVAL_1868 & _EVAL_1378;
  assign _EVAL_1222 = _EVAL_102 == 12'hb12;
  assign _EVAL_2242 = _EVAL_1868 & _EVAL_664;
  assign _EVAL_1753 = _EVAL_102 == 12'hb9b;
  assign _EVAL_943 = _EVAL_1868 & _EVAL_1753;
  assign _EVAL_1415 = _EVAL_102 == 12'h33d;
  assign _EVAL_1218 = _EVAL_102 == 12'hc1b;
  assign _EVAL_1705 = _EVAL_1846 & _EVAL_1218;
  assign _EVAL_2072 = _EVAL_102 == 12'hc90;
  assign _EVAL_945 = _EVAL_1868 & _EVAL_1297;
  assign _EVAL_1041 = _EVAL_102 == 12'hb09;
  assign _EVAL_1237 = _EVAL_1868 & _EVAL_1041;
  assign _EVAL_1839 = _EVAL_1846 & _EVAL_1209;
  assign _EVAL_1958 = _EVAL_579 == 32'h8;
  assign _EVAL_238 = _EVAL_1846 & _EVAL_2072;
  assign _EVAL_1422 = _EVAL_1846 & _EVAL_469;
  assign _EVAL_1204 = _EVAL_1868 & _EVAL_1198;
  assign _EVAL_2171 = _EVAL_1846 & _EVAL_563;
  assign _EVAL_661 = _EVAL_1868 & _EVAL_226;
  assign _EVAL_856 = _EVAL_102 == 12'h33b;
  assign _EVAL_1749 = _EVAL_1846 & _EVAL_554;
  assign _EVAL_1728 = _EVAL_1868 & _EVAL_695;
  assign _EVAL_1844 = _EVAL_102 == 12'h32e;
  assign _EVAL_1522 = _EVAL_1868 & _EVAL_1844;
  assign _EVAL_1333 = _EVAL_1776 | _EVAL_1806;
  assign _EVAL_768 = _EVAL_1868 & _EVAL_1744;
  assign _EVAL_1245 = _EVAL_1846 & _EVAL_1337;
  assign _EVAL_2000 = _EVAL_1868 & _EVAL_1746;
  assign _EVAL_989 = _EVAL_1846 & _EVAL_2088;
  assign _EVAL_1834 = _EVAL_1868 & _EVAL_484;
  assign _EVAL_972 = _EVAL_1868 & _EVAL_1415;
  assign _EVAL_1798 = _EVAL_102 == 12'hb1a;
  assign _EVAL_642 = _EVAL_1868 & _EVAL_2206;
  assign _EVAL_799 = _EVAL_1846 & _EVAL_1911;
  assign _EVAL_179 = _EVAL_1230 | _EVAL_146;
  assign _EVAL_704 = _EVAL_1868 & _EVAL_1031;
  assign _EVAL_1675 = _EVAL_1868 & _EVAL_690;
  assign _EVAL_725 = _EVAL_1868 & _EVAL_789;
  assign _EVAL_1485 = _EVAL_1868 & _EVAL_1752;
  assign _EVAL_2061 = _EVAL_1868 & _EVAL_2034;
  assign _EVAL_2148 = _EVAL_102 == 12'hc8a;
  assign _EVAL_965 = _EVAL_1846 & _EVAL_2148;
  assign _EVAL_1660 = _EVAL_1937 & _EVAL_1958;
  assign _EVAL_815 = _EVAL_1333 | _EVAL_146;
  assign _EVAL_1284 = _EVAL_1868 & _EVAL_1726;
  assign _EVAL_1572 = _EVAL_1868 & _EVAL_575;
  assign _EVAL_1497 = _EVAL_815 == 1'h0;
  assign _EVAL_1071 = _EVAL_102 == 12'hb1c;
  assign _EVAL_617 = _EVAL_1868 & _EVAL_1071;
  assign _EVAL_494 = _EVAL_1868 & _EVAL_1374;
  assign _EVAL_183 = _EVAL_1846 & _EVAL_1687;
  assign _EVAL_1591 = _EVAL_1846 & _EVAL_1360;
  assign _EVAL_2052 = _EVAL_1846 & _EVAL_316;
  assign _EVAL_1399 = _EVAL_1868 & _EVAL_335;
  assign _EVAL_1611 = _EVAL_1846 & _EVAL_1037;
  assign _EVAL_1148 = _EVAL_102 == 12'hc11;
  assign _EVAL_289 = _EVAL_1868 & _EVAL_1657;
  assign _EVAL_1812 = _EVAL_102 == 12'hb10;
  assign _EVAL_414 = _EVAL_1868 & _EVAL_2109;
  assign _EVAL_1757 = _EVAL_1868 & _EVAL_1222;
  assign _EVAL_367 = _EVAL_1846 & _EVAL_1301;
  assign _EVAL_221 = _EVAL_1868 & _EVAL_1812;
  assign _EVAL_391 = _EVAL_579 == 32'h1;
  assign _EVAL_1732 = _EVAL_1937 & _EVAL_391;
  assign _EVAL_1351 = _EVAL_179 == 1'h0;
  assign _EVAL_986 = _EVAL_102 == 12'h3b9;
  assign _EVAL_1080 = _EVAL_1868 & _EVAL_283;
  assign _EVAL_1007 = _EVAL_1846 & _EVAL_1148;
  assign _EVAL_853 = _EVAL_1868 & _EVAL_780;
  assign _EVAL_1975 = _EVAL_1868 & _EVAL_1798;
  assign _EVAL_1397 = _EVAL_1868 & _EVAL_1612;
  assign _EVAL_1677 = _EVAL_146 == 1'h0;
  assign _EVAL_706 = _EVAL_1868 & _EVAL_986;
  assign _EVAL_1935 = _EVAL_1868 & _EVAL_382;
  assign _EVAL_838 = _EVAL_1868 & _EVAL_856;
  assign _EVAL_1243 = _EVAL_1937 & _EVAL_2022;
  assign _EVAL_698 = _EVAL_102 == 12'hc0d;
  assign _EVAL_1903 = _EVAL_1846 & _EVAL_698;
  assign _EVAL_1480 = _EVAL_1868 & _EVAL_879;
  assign _EVAL_1135 = _EVAL_1846 & _EVAL_425;
  assign _EVAL_2098 = _EVAL_1846 & _EVAL_262;
  assign _EVAL_1916 = _EVAL_1846 & _EVAL_1500;
  assign _EVAL_499 = _EVAL_1868 & _EVAL_1758;
  assign _EVAL_519 = _EVAL_1868 & _EVAL_569;
  assign _EVAL_1413 = _EVAL_1868 & _EVAL_237;
  assign _EVAL_1883 = _EVAL_1846 & _EVAL_1537;
  always @(posedge _EVAL_53) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_627 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d827667c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34f665a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1732 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a7710b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1675 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1979a4e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1528 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffc83ec3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1299 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1afc0c8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_875 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69e4eb1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1135 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bf5c93a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_696 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddae5c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b800bec2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1660 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dec2b15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57df8ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_444 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ef0dba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1622 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c5e1b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1270 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(709038fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62de7888)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_915 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5151e92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1b88849)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1867 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9140a01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_642 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d179cba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1513 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf524e88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4604cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c120a34d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1903 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73d26e76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_933) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ecc008b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_768 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5336a167)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1265 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ac5e10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2045 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e2d1a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1990 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e952cf90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d3039d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1327 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e08ed3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a304701d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2061 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c6fd14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1510 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0fc4cb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3724fa22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1530 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aac14fe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_406 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5140c8f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1243 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f8c394c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_706 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41b77a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_671 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8f5c06f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6c96807)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1839 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e91f362)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1309 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7065364d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7143e86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2119 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c42e5d56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1109 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(147b80ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(463ed6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_481 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e04d2695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2014 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b07498a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_1069) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1962 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fae31a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2093 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9a56d8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1154 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a0ac939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1918 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cb95be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1250 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cc9d2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_818 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e032baf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_603 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a142eda5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc90e737)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1749 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcd53ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1460 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c619dcc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1611 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8db1015)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2178 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cb0080e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1274 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b36978b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1581 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d559ce60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1654 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e859743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1706 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9234956)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_943 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7917c50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f3f686)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_480 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63ebfe4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_593 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7213b13c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46a57442)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_833 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92407d32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1370 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb9eba6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1787 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17d1b182)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_366 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9433624)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_519 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1388d1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_582 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df1a9bcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1817 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c1fd84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_1069) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45253f03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1497) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1351) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a20d37ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1690 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b5e2ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_468 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c76424e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1335 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e9e93b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_610 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(970d61b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_933) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_917 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c69e2e00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1002 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9ea90c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_637 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16b2d249)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1116 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(544185fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53adff8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2134 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5c21e99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1258 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ebd9a27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1397 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b26fe7cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e1e88f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1858 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c77008b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65a3fb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24c69aa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1039 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(505aa10d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_590 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbad1a53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1316 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4b14e8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_560 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4b5bd24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_454 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca3be4bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1284 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ea20bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472e0b84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1006 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d922385)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1304 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2587ae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_453 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be095eb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e57e40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2000 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77537ed0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1766 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52bccae6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1860 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6eda505)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2196 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5df7d9db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1179 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd41584a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_429 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb4e8e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1522 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(838b6f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_493 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d17c8454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1195 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a914dcae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1591 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e071ebd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2020 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4653d4ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5664abe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1894 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(628f60c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1399 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8feb6756)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1883 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de0ceb89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_788 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(919b36b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d08409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(569ee470)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1705 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29b2cb3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f2b3670)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1252 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9011f9d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74299daf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1511 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(473223f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1245 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab6d014)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2107 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10aed55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2212 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7078d693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61b253d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1738 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72ebe2ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2052 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86a80eb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_704 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18751c65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_623 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c29a370f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70ccb2f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82454e04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55322d80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_945 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73f57b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1760 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c92b2953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_965 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18417fb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2242 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39ce339a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_721 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1703bd0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e9b7bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1897 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6dfe87a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83f36b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2051 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fbbc11d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_757 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1fdf073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_372 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3e267e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1351) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_839 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f590cf0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d20bd19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_774 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c51dd02d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2166 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2415c13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1485 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673179da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1080 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e540c721)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1527 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f530aedd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_600 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97a3c410)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bf16920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_393 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b603caee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4cf085f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_420 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f2af1f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80b0126)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_972 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb74efe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_838 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc511b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_880 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3bf2af1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1975 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebfddb6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2231 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d68bebc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1240 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8a728dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1497) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e824304d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_791 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f7c81f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1682 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecc4ba18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2016 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ffc2af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_553 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(921da9bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5248ef45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_712 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab3d4f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1572 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6af25338)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1915 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(153de2ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1173 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4e99312)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(247f3e88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_799 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(461ae642)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_701 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e0a2541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1462 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12bb3b96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e378fef2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1429 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c235df54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(267887ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1140 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df8e699d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1422 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d4717cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1204 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(260e0482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_929 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed1dcc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1480 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b7e83a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1007 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8137bb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1935 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc35ff40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1434 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51eb07d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_989 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bed4288)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_498 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39a37740)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(575a7150)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1237 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea0a1dec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ca84ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2171 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75bcb192)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_633 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb780c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2111 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e942de0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5120e2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1596 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(801dc077)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1716 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44e48d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2060 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c96ff8bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(578058f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2098 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8317592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1992 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8781154)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_410 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a1fb9af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(617ce01c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1013 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74f5fcfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_934 & _EVAL_1677) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d117df60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
