//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_304(
  input  [31:0] _EVAL,
  output [29:0] _EVAL_0,
  input  [1:0]  _EVAL_1,
  output [31:0] _EVAL_2,
  output        _EVAL_3,
  output [7:0]  _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  output [7:0]  _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  output [1:0]  _EVAL_12,
  output        _EVAL_13,
  output [31:0] _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input  [11:0] _EVAL_18,
  output        _EVAL_19,
  output        _EVAL_20,
  output [1:0]  _EVAL_21,
  output [1:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  output [1:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  output [1:0]  _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  output [1:0]  _EVAL_35,
  output        _EVAL_36,
  output [29:0] _EVAL_37,
  output        _EVAL_38,
  output        _EVAL_39,
  output [31:0] _EVAL_40,
  input  [1:0]  _EVAL_41,
  output        _EVAL_42,
  output [1:0]  _EVAL_43,
  output [31:0] _EVAL_44,
  output [1:0]  _EVAL_45,
  output        _EVAL_46,
  input         _EVAL_47,
  output        _EVAL_48,
  input  [1:0]  _EVAL_49,
  input         _EVAL_50,
  output [31:0] _EVAL_51,
  output        _EVAL_52,
  input         _EVAL_53,
  output [29:0] _EVAL_54,
  output [1:0]  _EVAL_55,
  output        _EVAL_56,
  output        _EVAL_57,
  output        _EVAL_58,
  output        _EVAL_59,
  output        _EVAL_60,
  output        _EVAL_61,
  output        _EVAL_62,
  output        _EVAL_63,
  output [31:0] _EVAL_64,
  output        _EVAL_65,
  output [29:0] _EVAL_66,
  output        _EVAL_67,
  output [1:0]  _EVAL_68,
  output        _EVAL_69,
  output        _EVAL_70,
  output        _EVAL_71,
  output        _EVAL_72,
  output [1:0]  _EVAL_73,
  input         _EVAL_74,
  output        _EVAL_75,
  output [1:0]  _EVAL_76,
  input         _EVAL_77,
  input  [31:0] _EVAL_78,
  output        _EVAL_79,
  output [31:0] _EVAL_80,
  output        _EVAL_81,
  output [1:0]  _EVAL_82,
  output [31:0] _EVAL_83,
  output [31:0] _EVAL_84,
  output        _EVAL_85,
  input         _EVAL_86,
  input  [31:0] _EVAL_87,
  output [2:0]  _EVAL_88,
  output        _EVAL_89,
  output        _EVAL_90,
  output        _EVAL_91,
  output        _EVAL_92,
  output        _EVAL_93,
  output        _EVAL_94,
  output        _EVAL_95,
  output [31:0] _EVAL_96,
  output        _EVAL_97,
  output        _EVAL_98,
  output [2:0]  _EVAL_99,
  output [1:0]  _EVAL_100,
  output [29:0] _EVAL_101,
  input  [11:0] _EVAL_102,
  output        _EVAL_103,
  output        _EVAL_104,
  output        _EVAL_105,
  output        _EVAL_106,
  output        _EVAL_107,
  output        _EVAL_108,
  input         _EVAL_109,
  output        _EVAL_110,
  output        _EVAL_111,
  output        _EVAL_112,
  output [31:0] _EVAL_113,
  output        _EVAL_114,
  output [7:0]  _EVAL_115,
  output        _EVAL_116,
  input  [31:0] _EVAL_117,
  output [31:0] _EVAL_118,
  output        _EVAL_119,
  output [1:0]  _EVAL_120,
  output [1:0]  _EVAL_121,
  output        _EVAL_122,
  output [31:0] _EVAL_123,
  output        _EVAL_124,
  output        _EVAL_125,
  output [31:0] _EVAL_126,
  output [26:0] _EVAL_127,
  output        _EVAL_128,
  output        _EVAL_129,
  output        _EVAL_130,
  output        _EVAL_131,
  output [31:0] _EVAL_132,
  output        _EVAL_133,
  output        _EVAL_134,
  output [1:0]  _EVAL_135,
  output [31:0] _EVAL_136,
  output        _EVAL_137,
  output [1:0]  _EVAL_138,
  output        _EVAL_139,
  output        _EVAL_140,
  output        _EVAL_141,
  output [29:0] _EVAL_142,
  output        _EVAL_143,
  input  [4:0]  _EVAL_144,
  output [31:0] _EVAL_145,
  input         _EVAL_146,
  output        _EVAL_147,
  output        _EVAL_148,
  output        _EVAL_149,
  output        _EVAL_150,
  output [1:0]  _EVAL_151,
  output        _EVAL_152,
  output        _EVAL_153,
  output        _EVAL_154,
  input         _EVAL_155,
  output [29:0] _EVAL_156,
  output        _EVAL_157,
  output [31:0] _EVAL_158,
  output [1:0]  _EVAL_159,
  output [31:0] _EVAL_160,
  output        _EVAL_161,
  output [29:0] _EVAL_162,
  output        _EVAL_163,
  output        _EVAL_164,
  input         _EVAL_165,
  output [31:0] _EVAL_166,
  output [31:0] _EVAL_167
);
  reg [33:0] _EVAL_171;
  reg [63:0] _RAND_0;
  reg  _EVAL_178;
  reg [31:0] _RAND_1;
  reg  _EVAL_181;
  reg [31:0] _RAND_2;
  reg [29:0] _EVAL_182;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_194;
  reg [31:0] _RAND_4;
  reg  _EVAL_203;
  reg [31:0] _RAND_5;
  reg  _EVAL_207;
  reg [31:0] _RAND_6;
  reg [1:0] _EVAL_252;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_267;
  reg [31:0] _RAND_8;
  reg [29:0] _EVAL_286;
  reg [31:0] _RAND_9;
  reg  _EVAL_297;
  reg [31:0] _RAND_10;
  reg [5:0] _EVAL_305;
  reg [31:0] _RAND_11;
  reg [1:0] _EVAL_317;
  reg [31:0] _RAND_12;
  reg  _EVAL_333;
  reg [31:0] _RAND_13;
  reg  _EVAL_334;
  reg [31:0] _RAND_14;
  reg  _EVAL_346;
  reg [31:0] _RAND_15;
  reg  _EVAL_361;
  reg [31:0] _RAND_16;
  reg  _EVAL_381;
  reg [31:0] _RAND_17;
  reg [31:0] _EVAL_422;
  reg [31:0] _RAND_18;
  reg  _EVAL_436;
  reg [31:0] _RAND_19;
  reg  _EVAL_442;
  reg [31:0] _RAND_20;
  reg [7:0] _EVAL_463;
  reg [31:0] _RAND_21;
  reg [1:0] _EVAL_491;
  reg [31:0] _RAND_22;
  reg  _EVAL_523;
  reg [31:0] _RAND_23;
  reg  _EVAL_528;
  reg [31:0] _RAND_24;
  reg [31:0] _EVAL_537;
  reg [31:0] _RAND_25;
  reg  _EVAL_551;
  reg [31:0] _RAND_26;
  reg [4:0] _EVAL_584;
  reg [31:0] _RAND_27;
  reg  _EVAL_594;
  reg [31:0] _RAND_28;
  reg [2:0] _EVAL_597;
  reg [31:0] _RAND_29;
  reg  _EVAL_609;
  reg [31:0] _RAND_30;
  reg  _EVAL_611;
  reg [31:0] _RAND_31;
  reg [1:0] _EVAL_631;
  reg [31:0] _RAND_32;
  reg  _EVAL_645;
  reg [31:0] _RAND_33;
  reg  _EVAL_692;
  reg [31:0] _RAND_34;
  reg  _EVAL_710;
  reg [31:0] _RAND_35;
  reg [1:0] _EVAL_715;
  reg [31:0] _RAND_36;
  reg  _EVAL_726;
  reg [31:0] _RAND_37;
  reg [31:0] _EVAL_745;
  reg [31:0] _RAND_38;
  reg [57:0] _EVAL_751;
  reg [63:0] _RAND_39;
  reg [1:0] _EVAL_759;
  reg [31:0] _RAND_40;
  reg [1:0] _EVAL_760;
  reg [31:0] _RAND_41;
  reg  _EVAL_762;
  reg [31:0] _RAND_42;
  reg  _EVAL_795;
  reg [31:0] _RAND_43;
  reg [29:0] _EVAL_842;
  reg [31:0] _RAND_44;
  reg [31:0] _EVAL_900;
  reg [31:0] _RAND_45;
  reg  _EVAL_926;
  reg [31:0] _RAND_46;
  reg  _EVAL_941;
  reg [31:0] _RAND_47;
  reg  _EVAL_944;
  reg [31:0] _RAND_48;
  reg  _EVAL_958;
  reg [31:0] _RAND_49;
  reg [31:0] _EVAL_978;
  reg [31:0] _RAND_50;
  reg  _EVAL_990;
  reg [31:0] _RAND_51;
  reg  _EVAL_992;
  reg [31:0] _RAND_52;
  reg [1:0] _EVAL_1011;
  reg [31:0] _RAND_53;
  reg  _EVAL_1022;
  reg [31:0] _RAND_54;
  reg [31:0] _EVAL_1048;
  reg [31:0] _RAND_55;
  reg  _EVAL_1062;
  reg [31:0] _RAND_56;
  reg [31:0] _EVAL_1063;
  reg [31:0] _RAND_57;
  reg  _EVAL_1073;
  reg [31:0] _RAND_58;
  reg [26:0] _EVAL_1078;
  reg [31:0] _RAND_59;
  reg  _EVAL_1138;
  reg [31:0] _RAND_60;
  reg  _EVAL_1162;
  reg [31:0] _RAND_61;
  reg  _EVAL_1167;
  reg [31:0] _RAND_62;
  reg  _EVAL_1168;
  reg [31:0] _RAND_63;
  reg  _EVAL_1178;
  reg [31:0] _RAND_64;
  reg  _EVAL_1193;
  reg [31:0] _RAND_65;
  reg [57:0] _EVAL_1212;
  reg [63:0] _RAND_66;
  reg [31:0] _EVAL_1223;
  reg [31:0] _RAND_67;
  reg [31:0] _EVAL_1239;
  reg [31:0] _RAND_68;
  reg  _EVAL_1241;
  reg [31:0] _RAND_69;
  reg [5:0] _EVAL_1249;
  reg [31:0] _RAND_70;
  reg  _EVAL_1261;
  reg [31:0] _RAND_71;
  reg [31:0] _EVAL_1282;
  reg [31:0] _RAND_72;
  reg [1:0] _EVAL_1344;
  reg [31:0] _RAND_73;
  reg  _EVAL_1354;
  reg [31:0] _RAND_74;
  reg  _EVAL_1366;
  reg [31:0] _RAND_75;
  reg  _EVAL_1376;
  reg [31:0] _RAND_76;
  reg  _EVAL_1381;
  reg [31:0] _RAND_77;
  reg  _EVAL_1385;
  reg [31:0] _RAND_78;
  reg [31:0] _EVAL_1392;
  reg [31:0] _RAND_79;
  reg [5:0] _EVAL_1419;
  reg [31:0] _RAND_80;
  reg  _EVAL_1421;
  reg [31:0] _RAND_81;
  reg [1:0] _EVAL_1424;
  reg [31:0] _RAND_82;
  reg [1:0] _EVAL_1425;
  reg [31:0] _RAND_83;
  reg [1:0] _EVAL_1440;
  reg [31:0] _RAND_84;
  reg [2:0] _EVAL_1458;
  reg [31:0] _RAND_85;
  reg [1:0] _EVAL_1466;
  reg [31:0] _RAND_86;
  reg [1:0] _EVAL_1479;
  reg [31:0] _RAND_87;
  reg [1:0] _EVAL_1494;
  reg [31:0] _RAND_88;
  reg  _EVAL_1499;
  reg [31:0] _RAND_89;
  reg [31:0] _EVAL_1532;
  reg [31:0] _RAND_90;
  reg [1:0] _EVAL_1545;
  reg [31:0] _RAND_91;
  reg  _EVAL_1555;
  reg [31:0] _RAND_92;
  reg  _EVAL_1556;
  reg [31:0] _RAND_93;
  reg  _EVAL_1563;
  reg [31:0] _RAND_94;
  reg  _EVAL_1567;
  reg [31:0] _RAND_95;
  reg  _EVAL_1585;
  reg [31:0] _RAND_96;
  reg [31:0] _EVAL_1589;
  reg [31:0] _RAND_97;
  reg  _EVAL_1593;
  reg [31:0] _RAND_98;
  reg  _EVAL_1608;
  reg [31:0] _RAND_99;
  reg  _EVAL_1620;
  reg [31:0] _RAND_100;
  reg [31:0] _EVAL_1632;
  reg [31:0] _RAND_101;
  reg [1:0] _EVAL_1666;
  reg [31:0] _RAND_102;
  reg [31:0] _EVAL_1688;
  reg [31:0] _RAND_103;
  reg [1:0] _EVAL_1700;
  reg [31:0] _RAND_104;
  reg [31:0] _EVAL_1725;
  reg [31:0] _RAND_105;
  reg  _EVAL_1733;
  reg [31:0] _RAND_106;
  reg  _EVAL_1743;
  reg [31:0] _RAND_107;
  reg  _EVAL_1763;
  reg [31:0] _RAND_108;
  reg  _EVAL_1769;
  reg [31:0] _RAND_109;
  reg  _EVAL_1770;
  reg [31:0] _RAND_110;
  reg  _EVAL_1792;
  reg [31:0] _RAND_111;
  reg  _EVAL_1808;
  reg [31:0] _RAND_112;
  reg  _EVAL_1869;
  reg [31:0] _RAND_113;
  reg  _EVAL_1877;
  reg [31:0] _RAND_114;
  reg  _EVAL_1895;
  reg [31:0] _RAND_115;
  reg  _EVAL_1899;
  reg [31:0] _RAND_116;
  reg  _EVAL_1929;
  reg [31:0] _RAND_117;
  reg [29:0] _EVAL_1942;
  reg [31:0] _RAND_118;
  reg [29:0] _EVAL_1952;
  reg [31:0] _RAND_119;
  reg  _EVAL_1956;
  reg [31:0] _RAND_120;
  reg [29:0] _EVAL_1978;
  reg [31:0] _RAND_121;
  reg  _EVAL_1982;
  reg [31:0] _RAND_122;
  reg  _EVAL_1986;
  reg [31:0] _RAND_123;
  reg  _EVAL_2002;
  reg [31:0] _RAND_124;
  reg  _EVAL_2033;
  reg [31:0] _RAND_125;
  reg  _EVAL_2047;
  reg [31:0] _RAND_126;
  reg  _EVAL_2063;
  reg [31:0] _RAND_127;
  reg  _EVAL_2074;
  reg [31:0] _RAND_128;
  reg  _EVAL_2084;
  reg [31:0] _RAND_129;
  reg [31:0] _EVAL_2090;
  reg [31:0] _RAND_130;
  reg [33:0] _EVAL_2106;
  reg [63:0] _RAND_131;
  reg  _EVAL_2131;
  reg [31:0] _RAND_132;
  reg  _EVAL_2152;
  reg [31:0] _RAND_133;
  reg  _EVAL_2158;
  reg [31:0] _RAND_134;
  reg  _EVAL_2159;
  reg [31:0] _RAND_135;
  reg [5:0] _EVAL_2177;
  reg [31:0] _RAND_136;
  reg  _EVAL_2180;
  reg [31:0] _RAND_137;
  reg [1:0] _EVAL_2181;
  reg [31:0] _RAND_138;
  reg  _EVAL_2190;
  reg [31:0] _RAND_139;
  reg [29:0] _EVAL_2210;
  reg [31:0] _RAND_140;
  reg  _EVAL_2220;
  reg [31:0] _RAND_141;
  reg [29:0] _EVAL_2224;
  reg [31:0] _RAND_142;
  reg [1:0] _EVAL_2226;
  reg [31:0] _RAND_143;
  reg [1:0] _EVAL_2227;
  reg [31:0] _RAND_144;
  reg  _EVAL_2230;
  reg [31:0] _RAND_145;
  reg  _EVAL_2232;
  reg [31:0] _RAND_146;
  reg  _EVAL_2238;
  reg [31:0] _RAND_147;
  wire  _EVAL_197;
  wire  _EVAL_500;
  wire [6:0] _EVAL_233;
  wire [31:0] _EVAL_2201;
  wire [31:0] _EVAL_580;
  wire [31:0] _EVAL_1969;
  wire [1:0] _EVAL_206;
  wire  _EVAL_652;
  wire [31:0] _EVAL_667;
  wire [31:0] _EVAL_2009;
  wire [31:0] _EVAL_1121;
  wire  _EVAL_1524;
  wire  _EVAL_278;
  wire  _EVAL_295;
  wire  _EVAL_980;
  wire  _EVAL_1444;
  wire  _EVAL_1338;
  wire  _EVAL_844;
  wire  _EVAL_259;
  wire  _EVAL_1336;
  wire  _EVAL_256;
  wire  _EVAL_529;
  wire  _EVAL_1989;
  wire  _EVAL_451;
  wire  _EVAL_1925;
  wire  _EVAL_982;
  wire  _EVAL_1704;
  wire  _EVAL_1076;
  wire  _EVAL_2209;
  wire  _EVAL_882;
  wire  _EVAL_732;
  wire  _EVAL_1587;
  wire  _EVAL_1735;
  wire  _EVAL_1388;
  wire  _EVAL_1824;
  wire  _EVAL_1848;
  wire  _EVAL_1441;
  wire  _EVAL_1144;
  wire  _EVAL_993;
  wire  _EVAL_2184;
  wire  _EVAL_1417;
  wire  _EVAL_1904;
  wire  _EVAL_1679;
  wire  _EVAL_1045;
  wire  _EVAL_1689;
  wire  _EVAL_835;
  wire  _EVAL_2010;
  wire  _EVAL_242;
  wire  _EVAL_511;
  wire  _EVAL_810;
  wire  _EVAL_1379;
  wire  _EVAL_1550;
  wire  _EVAL_1943;
  wire  _EVAL_1398;
  wire  _EVAL_662;
  wire  _EVAL_806;
  wire  _EVAL_1407;
  wire  _EVAL_1878;
  wire  _EVAL_1472;
  wire  _EVAL_248;
  wire  _EVAL_660;
  wire  _EVAL_415;
  wire  _EVAL_1400;
  wire  _EVAL_236;
  wire  _EVAL_1906;
  wire  _EVAL_247;
  wire  _EVAL_931;
  wire  _EVAL_2087;
  wire  _EVAL_962;
  wire  _EVAL_2025;
  wire  _EVAL_907;
  wire  _EVAL_892;
  wire  _EVAL_2019;
  wire  _EVAL_805;
  wire  _EVAL_1742;
  wire  _EVAL_1783;
  wire  _EVAL_1060;
  wire  _EVAL_1880;
  wire  _EVAL_595;
  wire  _EVAL_2237;
  wire  _EVAL_2135;
  wire  _EVAL_479;
  wire  _EVAL_1393;
  wire  _EVAL_1273;
  wire  _EVAL_874;
  wire  _EVAL_1579;
  wire  _EVAL_541;
  wire  _EVAL_1811;
  wire  _EVAL_1779;
  wire  _EVAL_1411;
  wire  _EVAL_638;
  wire  _EVAL_1874;
  wire  _EVAL_1490;
  wire  _EVAL_1253;
  wire  _EVAL_1951;
  wire  _EVAL_1142;
  wire  _EVAL_311;
  wire  _EVAL_223;
  wire  _EVAL_255;
  wire  _EVAL_1075;
  wire  _EVAL_1150;
  wire  _EVAL_304;
  wire  _EVAL_1745;
  wire  _EVAL_385;
  wire  _EVAL_969;
  wire  _EVAL_801;
  wire  _EVAL_276;
  wire  _EVAL_1569;
  wire  _EVAL_1056;
  wire  _EVAL_571;
  wire  _EVAL_2064;
  wire  _EVAL_1820;
  wire  _EVAL_1139;
  wire  _EVAL_942;
  wire  _EVAL_450;
  wire  _EVAL_409;
  wire  _EVAL_1708;
  wire  _EVAL_483;
  wire  _EVAL_1103;
  wire  _EVAL_266;
  wire  _EVAL_187;
  wire  _EVAL_1232;
  wire  _EVAL_1739;
  wire  _EVAL_1269;
  wire  _EVAL_632;
  wire  _EVAL_1633;
  wire  _EVAL_735;
  wire  _EVAL_230;
  wire  _EVAL_1164;
  wire  _EVAL_784;
  wire  _EVAL_1129;
  wire  _EVAL_683;
  wire  _EVAL_729;
  wire  _EVAL_1865;
  wire  _EVAL_2137;
  wire  _EVAL_232;
  wire  _EVAL_626;
  wire  _EVAL_1694;
  wire  _EVAL_796;
  wire  _EVAL_175;
  wire  _EVAL_1815;
  wire  _EVAL_1271;
  wire  _EVAL_1592;
  wire  _EVAL_2194;
  wire  _EVAL_693;
  wire  _EVAL_1805;
  wire  _EVAL_1420;
  wire  _EVAL_1830;
  wire  _EVAL_1582;
  wire  _EVAL_1183;
  wire  _EVAL_948;
  wire  _EVAL_2234;
  wire  _EVAL_591;
  wire  _EVAL_1220;
  wire  _EVAL_2225;
  wire  _EVAL_1881;
  wire  _EVAL_572;
  wire  _EVAL_1225;
  wire  _EVAL_217;
  wire  _EVAL_2175;
  wire  _EVAL_1626;
  wire  _EVAL_518;
  wire  _EVAL_1322;
  wire  _EVAL_1208;
  wire  _EVAL_1663;
  wire  _EVAL_1004;
  wire  _EVAL_1509;
  wire  _EVAL_403;
  wire  _EVAL_1019;
  wire  _EVAL_1449;
  wire  _EVAL_793;
  wire  _EVAL_1718;
  wire  _EVAL_1570;
  wire  _EVAL_615;
  wire  _EVAL_2188;
  wire  _EVAL_1602;
  wire  _EVAL_1349;
  wire  _EVAL_1983;
  wire  _EVAL_329;
  wire  _EVAL_1506;
  wire  _EVAL_1064;
  wire  _EVAL_1822;
  wire  _EVAL_908;
  wire  _EVAL_1671;
  wire  _EVAL_1796;
  wire  _EVAL_1730;
  wire  _EVAL_371;
  wire  _EVAL_313;
  wire  _EVAL_2115;
  wire  _EVAL_1298;
  wire  _EVAL_273;
  wire  _EVAL_369;
  wire  _EVAL_1780;
  wire  _EVAL_1938;
  wire  _EVAL_2172;
  wire  _EVAL_2193;
  wire  _EVAL_1558;
  wire  _EVAL_2007;
  wire  _EVAL_2005;
  wire  _EVAL_988;
  wire  _EVAL_2097;
  wire  _EVAL_1580;
  wire  _EVAL_1009;
  wire  _EVAL_193;
  wire  _EVAL_1052;
  wire  _EVAL_918;
  wire  _EVAL_937;
  wire  _EVAL_1658;
  wire  _EVAL_1467;
  wire  _EVAL_228;
  wire  _EVAL_1465;
  wire  _EVAL_360;
  wire  _EVAL_352;
  wire  _EVAL_2099;
  wire  _EVAL_1186;
  wire  _EVAL_1014;
  wire [31:0] _EVAL_953;
  wire [31:0] _EVAL_257;
  wire [31:0] _EVAL_428;
  wire [31:0] _EVAL_1038;
  wire  _EVAL_284;
  wire  _EVAL_1736;
  wire [15:0] _EVAL_2079;
  wire [15:0] _EVAL_1026;
  wire [31:0] _EVAL_2059;
  wire [31:0] _EVAL_1289;
  wire [31:0] _EVAL_1348;
  wire [31:0] _EVAL_1454;
  wire [31:0] _EVAL_497;
  wire  _EVAL_1997;
  wire [23:0] _EVAL_1888;
  wire [7:0] _EVAL_912;
  wire [1:0] _EVAL_1547;
  wire  _EVAL_1747;
  wire  _EVAL_461;
  wire [30:0] _EVAL_1092;
  wire [30:0] _EVAL_1577;
  wire [30:0] _EVAL_578;
  wire [30:0] _EVAL_246;
  wire [30:0] _EVAL_1433;
  wire [32:0] _EVAL_1141;
  wire  _EVAL_375;
  wire  _EVAL_1773;
  wire  _EVAL_2092;
  wire  _EVAL_309;
  wire  _EVAL_1722;
  wire  _EVAL_1310;
  wire [101:0] _EVAL_821;
  wire [1:0] _EVAL_1054;
  wire  _EVAL_753;
  wire  _EVAL_1765;
  wire [31:0] _EVAL_914;
  wire [31:0] _EVAL_1329;
  wire  _EVAL_1326;
  wire  _EVAL_898;
  wire  _EVAL_1112;
  wire [31:0] _EVAL_1859;
  wire  _EVAL_1043;
  wire  _EVAL_1902;
  wire [31:0] _EVAL_439;
  wire  _EVAL_1905;
  wire  _EVAL_739;
  wire  _EVAL_1849;
  wire  _EVAL_1937;
  wire [3:0] _EVAL_1621;
  wire [3:0] _EVAL_530;
  wire [31:0] _EVAL_1964;
  wire [31:0] _EVAL_579;
  wire  _EVAL_1334;
  wire [7:0] _EVAL_744;
  wire  _EVAL_750;
  wire  _EVAL_679;
  wire  _EVAL_2057;
  wire  _EVAL_1650;
  wire  _EVAL_1999;
  wire  _EVAL_1087;
  wire  _EVAL_1380;
  wire [3:0] _EVAL_1615;
  wire [3:0] _EVAL_778;
  wire  _EVAL_1046;
  wire  _EVAL_1855;
  wire  _EVAL_620;
  wire  _EVAL_939;
  wire  _EVAL_386;
  wire [1:0] _EVAL_845;
  wire  _EVAL_2017;
  wire  _EVAL_1520;
  wire [29:0] _EVAL_1919;
  wire  _EVAL_826;
  wire [1:0] _EVAL_913;
  wire [31:0] _EVAL_916;
  wire  _EVAL_283;
  wire  _EVAL_1188;
  wire  _EVAL_227;
  wire  _EVAL_343;
  wire  _EVAL_2116;
  wire  _EVAL_891;
  wire  _EVAL_2008;
  wire  _EVAL_2168;
  wire  _EVAL_1098;
  wire  _EVAL_1228;
  wire [1:0] _EVAL_1051;
  wire [1:0] _EVAL_1809;
  wire [1:0] _EVAL_1481;
  wire  _EVAL_697;
  wire  _EVAL_460;
  wire  _EVAL_462;
  wire  _EVAL_431;
  wire  _EVAL_1707;
  wire  _EVAL_2046;
  wire  _EVAL_1428;
  wire  _EVAL_719;
  wire  _EVAL_1115;
  wire  _EVAL_2085;
  wire  _EVAL_1539;
  wire  _EVAL_1609;
  wire  _EVAL_820;
  wire  _EVAL_495;
  wire  _EVAL_1842;
  wire [6:0] _EVAL_1669;
  wire [31:0] _EVAL_1517;
  wire [31:0] _EVAL_2174;
  wire [31:0] _EVAL_1816;
  wire [31:0] _EVAL_850;
  wire [31:0] _EVAL_1495;
  wire [31:0] _EVAL_222;
  wire [31:0] _EVAL_649;
  wire [31:0] _EVAL_1828;
  wire  _EVAL_1767;
  wire [30:0] _EVAL_1100;
  wire [31:0] _EVAL_1737;
  wire [31:0] _EVAL_180;
  wire [14:0] _EVAL_1496;
  wire [6:0] _EVAL_521;
  wire [18:0] _EVAL_689;
  wire [101:0] _EVAL_1003;
  wire [31:0] _EVAL_482;
  wire [31:0] _EVAL_1061;
  wire [31:0] _EVAL_2021;
  wire  _EVAL_755;
  wire  _EVAL_502;
  wire [6:0] _EVAL_549;
  wire [31:0] _EVAL_1970;
  wire [31:0] _EVAL_281;
  wire [31:0] _EVAL_1401;
  wire [31:0] _EVAL_1681;
  wire [31:0] _EVAL_2062;
  wire  _EVAL_569;
  wire [15:0] _EVAL_1656;
  wire [31:0] _EVAL_168;
  wire [31:0] _EVAL_2215;
  wire  _EVAL_1031;
  wire [31:0] _EVAL_630;
  wire [31:0] _EVAL_903;
  wire  _EVAL_1752;
  wire [31:0] _EVAL_503;
  wire [31:0] _EVAL_994;
  wire  _EVAL_1291;
  wire [31:0] _EVAL_2204;
  wire [31:0] _EVAL_771;
  wire [31:0] _EVAL_1315;
  wire [31:0] _EVAL_1893;
  wire [31:0] _EVAL_1946;
  wire [31:0] _EVAL_2182;
  wire [31:0] _EVAL_1463;
  wire  _EVAL_2208;
  wire [31:0] _EVAL_1635;
  wire [31:0] _EVAL_220;
  wire  _EVAL_262;
  wire  _EVAL_868;
  wire [31:0] _EVAL_342;
  wire [31:0] _EVAL_1664;
  wire  _EVAL_1833;
  wire [11:0] _EVAL_1190;
  wire [31:0] _EVAL_1256;
  wire [31:0] _EVAL_210;
  wire [31:0] _EVAL_188;
  wire  _EVAL_1297;
  wire [31:0] _EVAL_173;
  wire [31:0] _EVAL_711;
  wire [31:0] _EVAL_1032;
  wire [31:0] _EVAL_831;
  wire [31:0] _EVAL_1293;
  wire  _EVAL_2143;
  wire [31:0] _EVAL_1320;
  wire [31:0] _EVAL_885;
  wire  _EVAL_1713;
  wire [4:0] _EVAL_940;
  wire [31:0] _EVAL_487;
  wire [31:0] _EVAL_377;
  wire  _EVAL_772;
  wire [2:0] _EVAL_1288;
  wire [31:0] _EVAL_1127;
  wire [31:0] _EVAL_1347;
  wire [7:0] _EVAL_684;
  wire [7:0] _EVAL_2122;
  wire [31:0] _EVAL_1731;
  wire [31:0] _EVAL_2011;
  wire [63:0] _EVAL_817;
  wire  _EVAL_531;
  wire [63:0] _EVAL_2070;
  wire [63:0] _EVAL_656;
  wire [63:0] _EVAL_2112;
  wire  _EVAL_1559;
  wire [63:0] _EVAL_720;
  wire [63:0] _EVAL_1514;
  wire [63:0] _EVAL_2102;
  wire  _EVAL_1923;
  wire  _EVAL_1627;
  wire  _EVAL_1746;
  wire  _EVAL_1913;
  wire  _EVAL_749;
  wire [7:0] _EVAL_430;
  wire  _EVAL_2163;
  wire [7:0] _EVAL_857;
  wire [1:0] _EVAL_1143;
  wire  _EVAL_1515;
  wire [31:0] _EVAL_635;
  wire [31:0] _EVAL_1759;
  wire [6:0] _EVAL_1588;
  wire [31:0] _EVAL_688;
  wire [31:0] _EVAL_1359;
  wire [31:0] _EVAL_1096;
  wire [31:0] _EVAL_1236;
  wire  _EVAL_2162;
  wire  _EVAL_1408;
  wire [30:0] _EVAL_946;
  wire [6:0] _EVAL_318;
  wire [31:0] _EVAL_1945;
  wire [31:0] _EVAL_1889;
  wire  _EVAL_1445;
  wire  _EVAL_1702;
  wire  _EVAL_2073;
  wire  _EVAL_270;
  wire  _EVAL_1590;
  wire  _EVAL_1286;
  wire  _EVAL_412;
  wire  _EVAL_1050;
  wire  _EVAL_1151;
  wire  _EVAL_830;
  wire  _EVAL_1091;
  wire  _EVAL_1644;
  wire [15:0] _EVAL_1680;
  wire [7:0] _EVAL_1741;
  wire  _EVAL_243;
  wire  _EVAL_484;
  wire [31:0] _EVAL_1504;
  wire  _EVAL_1389;
  wire  _EVAL_396;
  wire  _EVAL_707;
  wire [39:0] _EVAL_2114;
  wire [31:0] _EVAL_1972;
  wire [39:0] _EVAL_658;
  wire  _EVAL_402;
  wire [29:0] _EVAL_474;
  wire [29:0] _EVAL_1074;
  wire [29:0] _EVAL_2032;
  wire [29:0] _EVAL_169;
  wire [29:0] _EVAL_1623;
  wire  _EVAL_1426;
  wire  _EVAL_666;
  wire [31:0] _EVAL_738;
  wire [63:0] _EVAL_769;
  wire [63:0] _EVAL_1640;
  wire  _EVAL_1358;
  wire [39:0] _EVAL_981;
  wire [39:0] _EVAL_445;
  wire [63:0] _EVAL_251;
  wire [63:0] _EVAL_1474;
  wire  _EVAL_2066;
  wire [39:0] _EVAL_449;
  wire [63:0] _EVAL_1535;
  wire [63:0] _EVAL_876;
  wire  _EVAL_1374;
  wire [7:0] _EVAL_389;
  wire [7:0] _EVAL_1174;
  wire [63:0] _EVAL_1988;
  wire [63:0] _EVAL_1021;
  wire  _EVAL_800;
  wire [7:0] _EVAL_977;
  wire [63:0] _EVAL_2236;
  wire [63:0] _EVAL_1631;
  wire  _EVAL_1617;
  wire [31:0] _EVAL_870;
  wire [63:0] _EVAL_459;
  wire [63:0] _EVAL_1748;
  wire  _EVAL_1437;
  wire [39:0] _EVAL_1122;
  wire [63:0] _EVAL_583;
  wire [63:0] _EVAL_1350;
  wire  _EVAL_316;
  wire [39:0] _EVAL_340;
  wire [63:0] _EVAL_1678;
  wire [63:0] _EVAL_1977;
  wire  _EVAL_1386;
  wire [7:0] _EVAL_2069;
  wire [7:0] _EVAL_1789;
  wire [63:0] _EVAL_680;
  wire [63:0] _EVAL_1578;
  wire  _EVAL_1560;
  wire [7:0] _EVAL_1448;
  wire [63:0] _EVAL_1571;
  wire [63:0] _EVAL_457;
  wire  _EVAL_677;
  wire [31:0] _EVAL_1873;
  wire [63:0] _EVAL_1311;
  wire [63:0] _EVAL_702;
  wire  _EVAL_425;
  wire [63:0] _EVAL_1784;
  wire [63:0] _EVAL_705;
  wire  _EVAL_323;
  wire [63:0] _EVAL_550;
  wire [63:0] _EVAL_322;
  wire  _EVAL_1657;
  wire [31:0] _EVAL_1724;
  wire [31:0] _EVAL_1471;
  wire [63:0] _EVAL_1077;
  wire [63:0] _EVAL_1568;
  wire  _EVAL_1872;
  wire [31:0] _EVAL_881;
  wire [31:0] _EVAL_1272;
  wire [63:0] _EVAL_1613;
  wire [63:0] _EVAL_1117;
  wire  _EVAL_596;
  wire [31:0] _EVAL_607;
  wire [63:0] _EVAL_258;
  wire [63:0] _EVAL_192;
  wire  _EVAL_212;
  wire [31:0] _EVAL_394;
  wire [63:0] _EVAL_1431;
  wire [63:0] _EVAL_1936;
  wire  _EVAL_1213;
  wire [7:0] _EVAL_2104;
  wire [7:0] _EVAL_1364;
  wire [15:0] _EVAL_2094;
  wire [31:0] _EVAL_525;
  wire [31:0] _EVAL_742;
  wire [63:0] _EVAL_321;
  wire [63:0] _EVAL_362;
  wire [7:0] _EVAL_1296;
  wire [7:0] _EVAL_888;
  wire [15:0] _EVAL_737;
  wire [31:0] _EVAL_548;
  wire [31:0] _EVAL_1548;
  wire [63:0] _EVAL_1887;
  wire [63:0] _EVAL_359;
  wire  _EVAL_1396;
  wire [29:0] _EVAL_1086;
  wire [63:0] _EVAL_478;
  wire [63:0] _EVAL_419;
  wire  _EVAL_237;
  wire  _EVAL_1307;
  wire [29:0] _EVAL_1321;
  wire [29:0] _EVAL_1645;
  wire [29:0] _EVAL_752;
  wire [29:0] _EVAL_1507;
  wire [29:0] _EVAL_339;
  wire [29:0] _EVAL_1890;
  wire [63:0] _EVAL_646;
  wire [63:0] _EVAL_1948;
  wire  _EVAL_780;
  wire  _EVAL_681;
  wire [29:0] _EVAL_1101;
  wire [29:0] _EVAL_198;
  wire [29:0] _EVAL_1907;
  wire [29:0] _EVAL_1118;
  wire [29:0] _EVAL_1278;
  wire [29:0] _EVAL_1171;
  wire [63:0] _EVAL_798;
  wire [63:0] _EVAL_1668;
  wire  _EVAL_539;
  wire  _EVAL_2151;
  wire [29:0] _EVAL_947;
  wire [29:0] _EVAL_1629;
  wire [29:0] _EVAL_411;
  wire [29:0] _EVAL_1961;
  wire [29:0] _EVAL_347;
  wire [29:0] _EVAL_1492;
  wire [63:0] _EVAL_1018;
  wire [63:0] _EVAL_854;
  wire  _EVAL_1647;
  wire  _EVAL_1306;
  wire [29:0] _EVAL_298;
  wire [29:0] _EVAL_1628;
  wire [29:0] _EVAL_2018;
  wire [29:0] _EVAL_896;
  wire [29:0] _EVAL_970;
  wire [29:0] _EVAL_517;
  wire [63:0] _EVAL_1202;
  wire [63:0] _EVAL_1238;
  wire  _EVAL_1418;
  wire [29:0] _EVAL_887;
  wire [29:0] _EVAL_1406;
  wire [29:0] _EVAL_2239;
  wire [29:0] _EVAL_1979;
  wire [29:0] _EVAL_2156;
  wire [29:0] _EVAL_509;
  wire [63:0] _EVAL_811;
  wire [63:0] _EVAL_546;
  wire  _EVAL_1285;
  wire  _EVAL_984;
  wire [29:0] _EVAL_775;
  wire [29:0] _EVAL_1832;
  wire [29:0] _EVAL_682;
  wire [29:0] _EVAL_2150;
  wire [29:0] _EVAL_641;
  wire [63:0] _EVAL_895;
  wire [63:0] _EVAL_1625;
  wire  _EVAL_279;
  wire [29:0] _EVAL_1891;
  wire [29:0] _EVAL_655;
  wire [29:0] _EVAL_224;
  wire [29:0] _EVAL_1015;
  wire [29:0] _EVAL_1508;
  wire [29:0] _EVAL_395;
  wire [63:0] _EVAL_1672;
  wire [63:0] _EVAL_2187;
  wire  _EVAL_1864;
  wire [31:0] _EVAL_280;
  wire [63:0] _EVAL_1372;
  wire [63:0] _EVAL_1404;
  wire  _EVAL_747;
  wire [31:0] _EVAL_1659;
  wire [63:0] _EVAL_293;
  wire [63:0] _EVAL_176;
  wire  _EVAL_2155;
  wire [31:0] _EVAL_1468;
  wire [63:0] _EVAL_387;
  wire [63:0] _EVAL_1442;
  wire  _EVAL_1500;
  wire [31:0] _EVAL_1361;
  wire [63:0] _EVAL_1475;
  wire [63:0] _EVAL_351;
  wire  _EVAL_1715;
  wire  _EVAL_2120;
  wire  _EVAL_1831;
  wire  _EVAL_733;
  wire  _EVAL_924;
  wire  _EVAL_797;
  wire  _EVAL_1120;
  wire  _EVAL_848;
  wire  _EVAL_832;
  wire  _EVAL_1260;
  wire  _EVAL_405;
  wire  _EVAL_1696;
  wire  _EVAL_538;
  wire  _EVAL_1540;
  wire  _EVAL_1387;
  wire  _EVAL_901;
  wire  _EVAL_2207;
  wire  _EVAL_1427;
  wire  _EVAL_1959;
  wire  _EVAL_1469;
  wire  _EVAL_2054;
  wire  _EVAL_418;
  wire  _EVAL_1482;
  wire  _EVAL_512;
  wire  _EVAL_1163;
  wire  _EVAL_392;
  wire  _EVAL_1330;
  wire  _EVAL_625;
  wire  _EVAL_260;
  wire  _EVAL_761;
  wire  _EVAL_1875;
  wire  _EVAL_1345;
  wire  _EVAL_2030;
  wire  _EVAL_1840;
  wire  _EVAL_1160;
  wire  _EVAL_957;
  wire  _EVAL_612;
  wire  _EVAL_337;
  wire  _EVAL_1565;
  wire  _EVAL_987;
  wire  _EVAL_324;
  wire  _EVAL_657;
  wire  _EVAL_274;
  wire  _EVAL_437;
  wire  _EVAL_1799;
  wire  _EVAL_2056;
  wire  _EVAL_884;
  wire  _EVAL_2071;
  wire  _EVAL_781;
  wire  _EVAL_254;
  wire  _EVAL_547;
  wire  _EVAL_315;
  wire  _EVAL_1430;
  wire  _EVAL_299;
  wire  _EVAL_1219;
  wire  _EVAL_327;
  wire  _EVAL_672;
  wire  _EVAL_2179;
  wire  _EVAL_527;
  wire  _EVAL_435;
  wire  _EVAL_1584;
  wire  _EVAL_961;
  wire  _EVAL_426;
  wire  _EVAL_622;
  wire [7:0] _EVAL_974;
  wire [39:0] _EVAL_899;
  wire [33:0] _EVAL_2154;
  wire [5:0] _EVAL_534;
  wire [6:0] _EVAL_1575;
  wire  _EVAL_1156;
  wire [33:0] _EVAL_1800;
  wire  _EVAL_1900;
  wire  _EVAL_1234;
  wire  _EVAL_1851;
  wire  _EVAL_676;
  wire  _EVAL_1137;
  wire  _EVAL_1764;
  wire  _EVAL_2229;
  wire  _EVAL_1035;
  wire  _EVAL_822;
  wire  _EVAL_1184;
  wire  _EVAL_1231;
  wire  _EVAL_1850;
  wire  _EVAL_1082;
  wire  _EVAL_356;
  wire  _EVAL_1966;
  wire  _EVAL_399;
  wire  _EVAL_889;
  wire  _EVAL_1598;
  wire  _EVAL_545;
  wire  _EVAL_400;
  wire  _EVAL_314;
  wire  _EVAL_380;
  wire  _EVAL_1155;
  wire  _EVAL_2125;
  wire  _EVAL_1931;
  wire  _EVAL_782;
  wire  _EVAL_1597;
  wire  _EVAL_1001;
  wire  _EVAL_1630;
  wire  _EVAL_905;
  wire  _EVAL_919;
  wire  _EVAL_1455;
  wire  _EVAL_1287;
  wire  _EVAL_893;
  wire  _EVAL_2136;
  wire  _EVAL_867;
  wire  _EVAL_2012;
  wire  _EVAL_1667;
  wire  _EVAL_2100;
  wire  _EVAL_823;
  wire  _EVAL_1157;
  wire  _EVAL_1554;
  wire  _EVAL_2080;
  wire  _EVAL_567;
  wire  _EVAL_963;
  wire  _EVAL_673;
  wire  _EVAL_345;
  wire  _EVAL_2127;
  wire  _EVAL_1189;
  wire  _EVAL_1453;
  wire  _EVAL_1246;
  wire  _EVAL_1818;
  wire  _EVAL_1594;
  wire  _EVAL_1512;
  wire  _EVAL_971;
  wire  _EVAL_190;
  wire  _EVAL_2050;
  wire  _EVAL_1502;
  wire  _EVAL_2138;
  wire  _EVAL_954;
  wire  _EVAL_902;
  wire  _EVAL_1491;
  wire  _EVAL_1994;
  wire  _EVAL_1879;
  wire  _EVAL_1526;
  wire  _EVAL_786;
  wire  _EVAL_1402;
  wire  _EVAL_1804;
  wire  _EVAL_448;
  wire  _EVAL_1538;
  wire  _EVAL_1362;
  wire  _EVAL_1016;
  wire  _EVAL_508;
  wire  _EVAL_1884;
  wire  _EVAL_1203;
  wire  _EVAL_185;
  wire  _EVAL_215;
  wire  _EVAL_1114;
  wire  _EVAL_979;
  wire  _EVAL_486;
  wire  _EVAL_1486;
  wire  _EVAL_1673;
  wire  _EVAL_1965;
  wire  _EVAL_1244;
  wire  _EVAL_470;
  wire  _EVAL_344;
  wire  _EVAL_1882;
  wire  _EVAL_2157;
  wire  _EVAL_967;
  wire  _EVAL_2118;
  wire  _EVAL_2013;
  wire  _EVAL_1709;
  wire  _EVAL_1553;
  wire  _EVAL_746;
  wire  _EVAL_496;
  wire  _EVAL_1384;
  wire  _EVAL_1369;
  wire  _EVAL_1483;
  wire  _EVAL_2211;
  wire  _EVAL_1939;
  wire  _EVAL_807;
  wire  _EVAL_384;
  wire  _EVAL_231;
  wire  _EVAL_1519;
  wire  _EVAL_566;
  wire  _EVAL_1912;
  wire  _EVAL_1023;
  wire  _EVAL_196;
  wire  _EVAL_2049;
  wire  _EVAL_968;
  wire  _EVAL_1968;
  wire  _EVAL_1920;
  wire  _EVAL_647;
  wire  _EVAL_932;
  wire  _EVAL_1774;
  wire  _EVAL_700;
  wire  _EVAL_1182;
  wire  _EVAL_1149;
  wire  _EVAL_1534;
  wire  _EVAL_1017;
  wire  _EVAL_776;
  wire  _EVAL_648;
  wire  _EVAL_374;
  wire  _EVAL_558;
  wire  _EVAL_1761;
  wire  _EVAL_1180;
  wire  _EVAL_1601;
  wire  _EVAL_205;
  wire  _EVAL_2218;
  wire  _EVAL_643;
  wire  _EVAL_492;
  wire  _EVAL_2200;
  wire  _EVAL_532;
  wire  _EVAL_287;
  wire  _EVAL_244;
  wire  _EVAL_1754;
  wire  _EVAL_731;
  wire  _EVAL_973;
  wire  _EVAL_208;
  wire  _EVAL_1211;
  wire  _EVAL_670;
  wire  _EVAL_1595;
  wire  _EVAL_1973;
  wire [1:0] _EVAL_602;
  wire  _EVAL_1785;
  wire  _EVAL_1125;
  wire  _EVAL_1266;
  wire  _EVAL_997;
  wire  _EVAL_843;
  wire  _EVAL_1217;
  wire  _EVAL_2235;
  wire [1:0] _EVAL_1693;
  wire [31:0] _EVAL_357;
  wire [31:0] _EVAL_1777;
  wire  _EVAL_1762;
  wire  _EVAL_2035;
  wire  _EVAL_1606;
  wire  _EVAL_1104;
  wire  _EVAL_787;
  wire  _EVAL_2003;
  wire  _EVAL_1085;
  wire [1:0] _EVAL_1871;
  wire  _EVAL_1562;
  wire  _EVAL_2124;
  wire  _EVAL_331;
  wire  _EVAL_1300;
  wire  _EVAL_1356;
  wire  _EVAL_328;
  wire [30:0] _EVAL_1235;
  wire [30:0] _EVAL_829;
  wire [30:0] _EVAL_1207;
  wire [6:0] _EVAL_1357;
  wire [31:0] _EVAL_1605;
  wire [31:0] _EVAL_1674;
  wire [31:0] _EVAL_1072;
  wire [31:0] _EVAL_1107;
  wire  _EVAL_1801;
  wire [14:0] _EVAL_1793;
  wire  _EVAL_1922;
  wire  _EVAL_1012;
  wire  _EVAL_2101;
  wire  _EVAL_1294;
  wire  _EVAL_2149;
  wire  _EVAL_674;
  wire  _EVAL_1305;
  wire  _EVAL_1279;
  wire  _EVAL_408;
  wire  _EVAL_866;
  wire  _EVAL_1566;
  wire  _EVAL_2228;
  wire  _EVAL_1478;
  wire  _EVAL_434;
  wire  _EVAL_1088;
  wire  _EVAL_1957;
  wire  _EVAL_1819;
  wire  _EVAL_1457;
  wire  _EVAL_199;
  wire  _EVAL_1254;
  wire  _EVAL_543;
  wire  _EVAL_2241;
  wire  _EVAL_1053;
  wire  _EVAL_1020;
  wire  _EVAL_1042;
  wire  _EVAL_1991;
  wire  _EVAL_1610;
  wire  _EVAL_455;
  wire  _EVAL_1838;
  wire  _EVAL_489;
  wire  _EVAL_1634;
  wire  _EVAL_1503;
  wire  _EVAL_1586;
  wire  _EVAL_1414;
  wire  _EVAL_1259;
  wire  _EVAL_1940;
  wire  _EVAL_1199;
  wire  _EVAL_2213;
  wire  _EVAL_211;
  wire  _EVAL_1797;
  wire  _EVAL_985;
  wire  _EVAL_792;
  wire  _EVAL_862;
  wire  _EVAL_1111;
  wire  _EVAL_1181;
  wire  _EVAL_370;
  wire  _EVAL_2240;
  wire  _EVAL_2006;
  wire  _EVAL_1084;
  wire  _EVAL_292;
  wire  _EVAL_2167;
  wire  _EVAL_1896;
  wire  _EVAL_184;
  wire  _EVAL_644;
  wire  _EVAL_708;
  wire  _EVAL_2095;
  wire  _EVAL_467;
  wire  _EVAL_1108;
  wire  _EVAL_354;
  wire  _EVAL_1751;
  wire [31:0] _EVAL_616;
  wire [31:0] _EVAL_219;
  wire  _EVAL_803;
  wire  _EVAL_650;
  wire [31:0] _EVAL_513;
  wire  _EVAL_209;
  wire [30:0] _EVAL_730;
  wire [30:0] _EVAL_424;
  wire [30:0] _EVAL_2108;
  wire [30:0] _EVAL_765;
  wire [30:0] _EVAL_1573;
  wire  _EVAL_654;
  wire  _EVAL_1910;
  wire [30:0] _EVAL_1886;
  wire [30:0] _EVAL_1652;
  wire  _EVAL_1825;
  wire  _EVAL_1123;
  wire  _EVAL_1541;
  wire  _EVAL_1292;
  wire [11:0] _EVAL_1355;
  wire [11:0] _EVAL_1395;
  wire  _EVAL_1200;
  wire  _EVAL_336;
  wire [2:0] _EVAL_691;
  wire  _EVAL_1028;
  wire  _EVAL_846;
  wire [24:0] _EVAL_1771;
  wire [4:0] _EVAL_573;
  wire [6:0] _EVAL_1130;
  wire [31:0] _EVAL_777;
  wire [29:0] _EVAL_2145;
  wire [31:0] _EVAL_526;
  wire [31:0] _EVAL_1639;
  wire [31:0] _EVAL_604;
  wire [31:0] _EVAL_561;
  wire [63:0] _EVAL_452;
  wire [57:0] _EVAL_1695;
  wire [5:0] _EVAL_440;
  wire [6:0] _EVAL_1049;
  wire  _EVAL_1914;
  wire [57:0] _EVAL_1845;
  wire  _EVAL_996;
  wire  _EVAL_250;
  wire [1:0] _EVAL_507;
  wire  _EVAL_1954;
  wire  _EVAL_1543;
  wire [1:0] _EVAL_659;
  wire  _EVAL_1523;
  wire  _EVAL_736;
  wire  _EVAL_310;
  wire  _EVAL_855;
  wire  _EVAL_174;
  wire  _EVAL_1533;
  wire [1:0] _EVAL_2161;
  wire [39:0] _EVAL_878;
  wire  _EVAL_201;
  wire  _EVAL_1146;
  wire  _EVAL_490;
  wire  _EVAL_1518;
  wire  _EVAL_364;
  wire  _EVAL_1720;
  wire [1:0] _EVAL_383;
  wire  _EVAL_2110;
  wire  _EVAL_1010;
  wire  _EVAL_404;
  wire  _EVAL_1251;
  wire  _EVAL_1960;
  wire  _EVAL_999;
  wire  _EVAL_2202;
  wire  _EVAL_858;
  wire [1:0] _EVAL_1136;
  wire  _EVAL_2027;
  wire [30:0] _EVAL_1373;
  wire  _EVAL_1781;
  wire  _EVAL_1210;
  wire  _EVAL_2221;
  wire  _EVAL_605;
  wire  _EVAL_1981;
  wire  _EVAL_1489;
  wire  _EVAL_909;
  wire [30:0] _EVAL_636;
  wire  _EVAL_2023;
  wire  _EVAL_2243;
  wire  _EVAL_2028;
  wire  _EVAL_1648;
  wire  _EVAL_935;
  wire  _EVAL_964;
  wire [31:0] _EVAL_2144;
  wire  _EVAL_1394;
  wire  _EVAL_998;
  wire  _EVAL_2192;
  wire  _EVAL_1921;
  wire [3:0] _EVAL_756;
  wire [3:0] _EVAL_1823;
  wire [3:0] _EVAL_510;
  wire [3:0] _EVAL_2223;
  wire [3:0] _EVAL_740;
  wire [3:0] _EVAL_2123;
  wire [3:0] _EVAL_1603;
  wire [3:0] _EVAL_2191;
  wire [3:0] _EVAL_1377;
  wire [3:0] _EVAL_1926;
  wire [3:0] _EVAL_358;
  wire [3:0] _EVAL_1464;
  wire [3:0] _EVAL_794;
  wire [3:0] _EVAL_923;
  wire [3:0] _EVAL_466;
  wire [3:0] _EVAL_1853;
  wire [3:0] _EVAL_1980;
  wire [3:0] _EVAL_709;
  wire [3:0] _EVAL_763;
  wire  _EVAL_1083;
  wire  _EVAL_271;
  wire  _EVAL_1461;
  wire [31:0] _EVAL_1302;
  wire  _EVAL_1079;
  wire  _EVAL_1058;
  wire  _EVAL_1551;
  wire  _EVAL_2024;
  wire  _EVAL_1416;
  wire  _EVAL_253;
  wire  _EVAL_2081;
  wire  _EVAL_1027;
  wire  _EVAL_1641;
  wire [31:0] _EVAL_577;
  wire [39:0] _EVAL_477;
  wire [5:0] _EVAL_504;
  wire [6:0] _EVAL_2089;
  wire  _EVAL_1317;
  wire  _EVAL_1264;
  wire  _EVAL_249;
  wire [30:0] _EVAL_2043;
  wire [30:0] _EVAL_1090;
  wire  _EVAL_883;
  wire  _EVAL_865;
  wire  _EVAL_2078;
  wire  _EVAL_1949;
  wire [7:0] _EVAL_1863;
  wire [39:0] _EVAL_773;
  wire [39:0] _EVAL_229;
  wire [39:0] _EVAL_443;
  wire  _EVAL_1941;
  wire [39:0] _EVAL_2082;
  wire  _EVAL_239;
  wire [5:0] _EVAL_995;
  wire [31:0] _EVAL_277;
  wire [31:0] _EVAL_213;
  wire  _EVAL_1908;
  wire  _EVAL_505;
  wire  _EVAL_1172;
  wire  _EVAL_307;
  wire [1:0] _EVAL_767;
  wire [1:0] _EVAL_1583;
  wire [1:0] _EVAL_2139;
  wire [1:0] _EVAL_302;
  wire [1:0] _EVAL_1498;
  wire  _EVAL_1194;
  wire  _EVAL_1536;
  wire [26:0] _EVAL_1721;
  wire [31:0] _EVAL_827;
  wire [31:0] _EVAL_718;
  wire [31:0] _EVAL_2173;
  wire [1:0] _EVAL_2183;
  wire [1:0] _EVAL_960;
  wire  _EVAL_1410;
  wire  _EVAL_959;
  wire  _EVAL_863;
  wire  _EVAL_1216;
  wire  _EVAL_1473;
  wire  _EVAL_1030;
  wire  _EVAL_1233;
  wire  _EVAL_390;
  wire  _EVAL_195;
  wire [5:0] _EVAL_522;
  wire [63:0] _EVAL_724;
  wire [63:0] _EVAL_2001;
  wire [31:0] _EVAL_282;
  wire  _EVAL_1451;
  wire  _EVAL_2130;
  wire [31:0] _EVAL_427;
  wire [31:0] _EVAL_2132;
  wire [1:0] _EVAL_2140;
  wire  _EVAL_1229;
  wire [30:0] _EVAL_1147;
  wire [1:0] _EVAL_275;
  wire  _EVAL_864;
  wire  _EVAL_1170;
  wire  _EVAL_678;
  wire  _EVAL_570;
  wire [31:0] _EVAL_920;
  wire [63:0] _EVAL_225;
  wire [57:0] _EVAL_1723;
  wire [33:0] _EVAL_1976;
  wire [4:0] _EVAL_1383;
  wire [31:0] _EVAL_713;
  wire  _EVAL_1856;
  wire  _EVAL_665;
  wire  _EVAL_1165;
  wire [31:0] _EVAL_1255;
  wire  _EVAL_722;
  wire  _EVAL_2219;
  wire  _EVAL_1131;
  wire  _EVAL_353;
  wire  _EVAL_1276;
  wire  _EVAL_1332;
  wire [30:0] _EVAL_1552;
  wire [30:0] _EVAL_2113;
  wire [30:0] _EVAL_1852;
  wire [1:0] _EVAL_816;
  wire  _EVAL_991;
  wire  _EVAL_1102;
  wire [31:0] _EVAL_1529;
  wire [63:0] _EVAL_619;
  wire [63:0] _EVAL_699;
  wire [6:0] _EVAL_717;
  wire [63:0] _EVAL_904;
  wire [63:0] _EVAL_886;
  wire [63:0] _EVAL_1328;
  wire  _EVAL_1827;
  wire  _EVAL_1275;
  wire [33:0] _EVAL_465;
  wire [33:0] _EVAL_533;
  wire  _EVAL_851;
  wire  _EVAL_1008;
  wire  _EVAL_2142;
  wire  _EVAL_653;
  wire [31:0] _EVAL_669;
  wire [31:0] _EVAL_1932;
  wire  _EVAL_349;
  wire [4:0] _EVAL_1343;
  wire [4:0] _EVAL_779;
  wire [31:0] _EVAL_1685;
  wire [31:0] _EVAL_1033;
  wire [31:0] _EVAL_2195;
  wire [3:0] _EVAL_1924;
  wire [3:0] _EVAL_441;
  wire [3:0] _EVAL_2129;
  wire [3:0] _EVAL_1067;
  wire  _EVAL_2222;
  wire [31:0] _EVAL_1443;
  wire [30:0] _EVAL_341;
  wire [32:0] _EVAL_1782;
  wire  _EVAL_828;
  wire [57:0] _EVAL_2077;
  wire  _EVAL_2029;
  wire  _EVAL_1145;
  wire  _EVAL_1025;
  wire [30:0] _EVAL_1044;
  wire [30:0] _EVAL_1813;
  wire [30:0] _EVAL_458;
  wire [31:0] _EVAL_506;
  wire [31:0] _EVAL_741;
  wire [32:0] _EVAL_1312;
  wire  _EVAL_1093;
  wire  _EVAL_1655;
  wire [31:0] _EVAL_1126;
  wire  _EVAL_928;
  wire [31:0] _EVAL_877;
  wire  _EVAL_808;
  wire  _EVAL_2160;
  wire [31:0] _EVAL_608;
  wire  _EVAL_2121;
  wire [30:0] _EVAL_303;
  wire [30:0] _EVAL_320;
  wire  _EVAL_559;
  wire [30:0] _EVAL_1459;
  wire [30:0] _EVAL_1876;
  wire [30:0] _EVAL_1649;
  wire [30:0] _EVAL_1691;
  wire  _EVAL_2015;
  wire [31:0] _EVAL_1791;
  wire [31:0] _EVAL_2068;
  wire [30:0] _EVAL_2165;
  wire [30:0] _EVAL_2185;
  wire [32:0] _EVAL_2169;
  wire  _EVAL_535;
  wire  _EVAL_1353;
  wire  _EVAL_1661;
  wire [31:0] _EVAL_639;
  wire  _EVAL_1772;
  wire  _EVAL_1953;
  wire [63:0] _EVAL_675;
  wire [63:0] _EVAL_330;
  wire  _EVAL_813;
  wire  _EVAL_1177;
  wire [31:0] _EVAL_2091;
  wire  _EVAL_2067;
  wire [30:0] _EVAL_790;
  wire [30:0] _EVAL_743;
  wire [30:0] _EVAL_716;
  wire [30:0] _EVAL_871;
  wire [57:0] _EVAL_1403;
  wire  _EVAL_565;
  wire [57:0] _EVAL_1947;
  wire [11:0] _EVAL_2147;
  wire  _EVAL_471;
  wire [31:0] _EVAL_476;
  wire [31:0] _EVAL_516;
  wire  _EVAL_1963;
  wire [31:0] _EVAL_1717;
  wire [31:0] _EVAL_326;
  wire [33:0] _EVAL_2153;
  wire [31:0] _EVAL_2205;
  wire [3:0] _EVAL_348;
  wire [31:0] _EVAL_809;
  wire  _EVAL_1158;
  wire  _EVAL_177;
  wire [32:0] _EVAL_728;
  wire  _EVAL_1843;
  wire  _EVAL_1642;
  wire [31:0] _EVAL_265;
  wire  _EVAL_1928;
  wire  _EVAL_624;
  wire [32:0] _EVAL_2133;
  wire [63:0] _EVAL_869;
  wire [32:0] _EVAL_1927;
  wire [39:0] _EVAL_186;
  wire [39:0] _EVAL_860;
  wire [1:0] _EVAL_1993;
  wire  _EVAL_1836;
  wire [1:0] _EVAL_1788;
  wire [31:0] _EVAL_2170;
  wire [31:0] _EVAL_906;
  wire  _EVAL_1159;
  wire  _EVAL_1371;
  wire  _EVAL_574;
  wire  _EVAL_1624;
  wire [32:0] _EVAL_2086;
  wire  _EVAL_204;
  wire [31:0] _EVAL_2065;
  wire [31:0] _EVAL_363;
  wire [1:0] _EVAL_651;
  assign _EVAL_197 = _EVAL_18 == 12'hc97;
  assign _EVAL_500 = _EVAL_23[1];
  assign _EVAL_233 = {_EVAL_2152,1'h0,1'h0,_EVAL_1743,_EVAL_2063,_EVAL_2002,_EVAL_1929};
  assign _EVAL_2201 = {4'h2,_EVAL_1769,14'h400,_EVAL_692,_EVAL_203,2'h0,_EVAL_1700,_EVAL_233};
  assign _EVAL_580 = _EVAL_500 ? _EVAL_2201 : 32'h0;
  assign _EVAL_1969 = _EVAL_580 | _EVAL_87;
  assign _EVAL_206 = _EVAL_23[1:0];
  assign _EVAL_652 = _EVAL_206 == 2'h3;
  assign _EVAL_667 = _EVAL_652 ? _EVAL_87 : 32'h0;
  assign _EVAL_2009 = ~ _EVAL_667;
  assign _EVAL_1121 = _EVAL_1969 & _EVAL_2009;
  assign _EVAL_1524 = _EVAL_18 == 12'h7a0;
  assign _EVAL_278 = _EVAL_18 == 12'h7a1;
  assign _EVAL_295 = _EVAL_1524 | _EVAL_278;
  assign _EVAL_980 = _EVAL_18 == 12'h7a2;
  assign _EVAL_1444 = _EVAL_295 | _EVAL_980;
  assign _EVAL_1338 = _EVAL_18 == 12'h301;
  assign _EVAL_844 = _EVAL_1444 | _EVAL_1338;
  assign _EVAL_259 = _EVAL_18 == 12'h300;
  assign _EVAL_1336 = _EVAL_844 | _EVAL_259;
  assign _EVAL_256 = _EVAL_18 == 12'h305;
  assign _EVAL_529 = _EVAL_1336 | _EVAL_256;
  assign _EVAL_1989 = _EVAL_18 == 12'h344;
  assign _EVAL_451 = _EVAL_529 | _EVAL_1989;
  assign _EVAL_1925 = _EVAL_18 == 12'h304;
  assign _EVAL_982 = _EVAL_451 | _EVAL_1925;
  assign _EVAL_1704 = _EVAL_18 == 12'h340;
  assign _EVAL_1076 = _EVAL_982 | _EVAL_1704;
  assign _EVAL_2209 = _EVAL_18 == 12'h341;
  assign _EVAL_882 = _EVAL_1076 | _EVAL_2209;
  assign _EVAL_732 = _EVAL_18 == 12'h343;
  assign _EVAL_1587 = _EVAL_882 | _EVAL_732;
  assign _EVAL_1735 = _EVAL_18 == 12'h342;
  assign _EVAL_1388 = _EVAL_1587 | _EVAL_1735;
  assign _EVAL_1824 = _EVAL_18 == 12'hf14;
  assign _EVAL_1848 = _EVAL_1388 | _EVAL_1824;
  assign _EVAL_1441 = _EVAL_18 == 12'h7b0;
  assign _EVAL_1144 = _EVAL_1848 | _EVAL_1441;
  assign _EVAL_993 = _EVAL_18 == 12'h7b1;
  assign _EVAL_2184 = _EVAL_1144 | _EVAL_993;
  assign _EVAL_1417 = _EVAL_18 == 12'h7b2;
  assign _EVAL_1904 = _EVAL_2184 | _EVAL_1417;
  assign _EVAL_1679 = _EVAL_18 == 12'h1;
  assign _EVAL_1045 = _EVAL_1904 | _EVAL_1679;
  assign _EVAL_1689 = _EVAL_18 == 12'h2;
  assign _EVAL_835 = _EVAL_1045 | _EVAL_1689;
  assign _EVAL_2010 = _EVAL_18 == 12'h3;
  assign _EVAL_242 = _EVAL_835 | _EVAL_2010;
  assign _EVAL_511 = _EVAL_18 == 12'hb00;
  assign _EVAL_810 = _EVAL_242 | _EVAL_511;
  assign _EVAL_1379 = _EVAL_18 == 12'hb02;
  assign _EVAL_1550 = _EVAL_810 | _EVAL_1379;
  assign _EVAL_1943 = _EVAL_18 == 12'h323;
  assign _EVAL_1398 = _EVAL_1550 | _EVAL_1943;
  assign _EVAL_662 = _EVAL_18 == 12'hb03;
  assign _EVAL_806 = _EVAL_1398 | _EVAL_662;
  assign _EVAL_1407 = _EVAL_18 == 12'hc03;
  assign _EVAL_1878 = _EVAL_806 | _EVAL_1407;
  assign _EVAL_1472 = _EVAL_18 == 12'hb83;
  assign _EVAL_248 = _EVAL_1878 | _EVAL_1472;
  assign _EVAL_660 = _EVAL_18 == 12'hc83;
  assign _EVAL_415 = _EVAL_248 | _EVAL_660;
  assign _EVAL_1400 = _EVAL_18 == 12'h324;
  assign _EVAL_236 = _EVAL_415 | _EVAL_1400;
  assign _EVAL_1906 = _EVAL_18 == 12'hb04;
  assign _EVAL_247 = _EVAL_236 | _EVAL_1906;
  assign _EVAL_931 = _EVAL_18 == 12'hc04;
  assign _EVAL_2087 = _EVAL_247 | _EVAL_931;
  assign _EVAL_962 = _EVAL_18 == 12'hb84;
  assign _EVAL_2025 = _EVAL_2087 | _EVAL_962;
  assign _EVAL_907 = _EVAL_18 == 12'hc84;
  assign _EVAL_892 = _EVAL_2025 | _EVAL_907;
  assign _EVAL_2019 = _EVAL_18 == 12'h325;
  assign _EVAL_805 = _EVAL_892 | _EVAL_2019;
  assign _EVAL_1742 = _EVAL_18 == 12'hb05;
  assign _EVAL_1783 = _EVAL_805 | _EVAL_1742;
  assign _EVAL_1060 = _EVAL_18 == 12'hc05;
  assign _EVAL_1880 = _EVAL_1783 | _EVAL_1060;
  assign _EVAL_595 = _EVAL_18 == 12'hb85;
  assign _EVAL_2237 = _EVAL_1880 | _EVAL_595;
  assign _EVAL_2135 = _EVAL_18 == 12'hc85;
  assign _EVAL_479 = _EVAL_2237 | _EVAL_2135;
  assign _EVAL_1393 = _EVAL_18 == 12'h326;
  assign _EVAL_1273 = _EVAL_479 | _EVAL_1393;
  assign _EVAL_874 = _EVAL_18 == 12'hb06;
  assign _EVAL_1579 = _EVAL_1273 | _EVAL_874;
  assign _EVAL_541 = _EVAL_18 == 12'hc06;
  assign _EVAL_1811 = _EVAL_1579 | _EVAL_541;
  assign _EVAL_1779 = _EVAL_18 == 12'hb86;
  assign _EVAL_1411 = _EVAL_1811 | _EVAL_1779;
  assign _EVAL_638 = _EVAL_18 == 12'hc86;
  assign _EVAL_1874 = _EVAL_1411 | _EVAL_638;
  assign _EVAL_1490 = _EVAL_18 == 12'h327;
  assign _EVAL_1253 = _EVAL_1874 | _EVAL_1490;
  assign _EVAL_1951 = _EVAL_18 == 12'hb07;
  assign _EVAL_1142 = _EVAL_1253 | _EVAL_1951;
  assign _EVAL_311 = _EVAL_18 == 12'hc07;
  assign _EVAL_223 = _EVAL_1142 | _EVAL_311;
  assign _EVAL_255 = _EVAL_18 == 12'hb87;
  assign _EVAL_1075 = _EVAL_223 | _EVAL_255;
  assign _EVAL_1150 = _EVAL_18 == 12'hc87;
  assign _EVAL_304 = _EVAL_1075 | _EVAL_1150;
  assign _EVAL_1745 = _EVAL_18 == 12'h328;
  assign _EVAL_385 = _EVAL_304 | _EVAL_1745;
  assign _EVAL_969 = _EVAL_18 == 12'hb08;
  assign _EVAL_801 = _EVAL_385 | _EVAL_969;
  assign _EVAL_276 = _EVAL_18 == 12'hc08;
  assign _EVAL_1569 = _EVAL_801 | _EVAL_276;
  assign _EVAL_1056 = _EVAL_18 == 12'hb88;
  assign _EVAL_571 = _EVAL_1569 | _EVAL_1056;
  assign _EVAL_2064 = _EVAL_18 == 12'hc88;
  assign _EVAL_1820 = _EVAL_571 | _EVAL_2064;
  assign _EVAL_1139 = _EVAL_18 == 12'h329;
  assign _EVAL_942 = _EVAL_1820 | _EVAL_1139;
  assign _EVAL_450 = _EVAL_18 == 12'hb09;
  assign _EVAL_409 = _EVAL_942 | _EVAL_450;
  assign _EVAL_1708 = _EVAL_18 == 12'hc09;
  assign _EVAL_483 = _EVAL_409 | _EVAL_1708;
  assign _EVAL_1103 = _EVAL_18 == 12'hb89;
  assign _EVAL_266 = _EVAL_483 | _EVAL_1103;
  assign _EVAL_187 = _EVAL_18 == 12'hc89;
  assign _EVAL_1232 = _EVAL_266 | _EVAL_187;
  assign _EVAL_1739 = _EVAL_18 == 12'h32a;
  assign _EVAL_1269 = _EVAL_1232 | _EVAL_1739;
  assign _EVAL_632 = _EVAL_18 == 12'hb0a;
  assign _EVAL_1633 = _EVAL_1269 | _EVAL_632;
  assign _EVAL_735 = _EVAL_18 == 12'hc0a;
  assign _EVAL_230 = _EVAL_1633 | _EVAL_735;
  assign _EVAL_1164 = _EVAL_18 == 12'hb8a;
  assign _EVAL_784 = _EVAL_230 | _EVAL_1164;
  assign _EVAL_1129 = _EVAL_18 == 12'hc8a;
  assign _EVAL_683 = _EVAL_784 | _EVAL_1129;
  assign _EVAL_729 = _EVAL_18 == 12'h32b;
  assign _EVAL_1865 = _EVAL_683 | _EVAL_729;
  assign _EVAL_2137 = _EVAL_18 == 12'hb0b;
  assign _EVAL_232 = _EVAL_1865 | _EVAL_2137;
  assign _EVAL_626 = _EVAL_18 == 12'hc0b;
  assign _EVAL_1694 = _EVAL_232 | _EVAL_626;
  assign _EVAL_796 = _EVAL_18 == 12'hb8b;
  assign _EVAL_175 = _EVAL_1694 | _EVAL_796;
  assign _EVAL_1815 = _EVAL_18 == 12'hc8b;
  assign _EVAL_1271 = _EVAL_175 | _EVAL_1815;
  assign _EVAL_1592 = _EVAL_18 == 12'h32c;
  assign _EVAL_2194 = _EVAL_1271 | _EVAL_1592;
  assign _EVAL_693 = _EVAL_18 == 12'hb0c;
  assign _EVAL_1805 = _EVAL_2194 | _EVAL_693;
  assign _EVAL_1420 = _EVAL_18 == 12'hc0c;
  assign _EVAL_1830 = _EVAL_1805 | _EVAL_1420;
  assign _EVAL_1582 = _EVAL_18 == 12'hb8c;
  assign _EVAL_1183 = _EVAL_1830 | _EVAL_1582;
  assign _EVAL_948 = _EVAL_18 == 12'hc8c;
  assign _EVAL_2234 = _EVAL_1183 | _EVAL_948;
  assign _EVAL_591 = _EVAL_18 == 12'h32d;
  assign _EVAL_1220 = _EVAL_2234 | _EVAL_591;
  assign _EVAL_2225 = _EVAL_18 == 12'hb0d;
  assign _EVAL_1881 = _EVAL_1220 | _EVAL_2225;
  assign _EVAL_572 = _EVAL_18 == 12'hc0d;
  assign _EVAL_1225 = _EVAL_1881 | _EVAL_572;
  assign _EVAL_217 = _EVAL_18 == 12'hb8d;
  assign _EVAL_2175 = _EVAL_1225 | _EVAL_217;
  assign _EVAL_1626 = _EVAL_18 == 12'hc8d;
  assign _EVAL_518 = _EVAL_2175 | _EVAL_1626;
  assign _EVAL_1322 = _EVAL_18 == 12'h32e;
  assign _EVAL_1208 = _EVAL_518 | _EVAL_1322;
  assign _EVAL_1663 = _EVAL_18 == 12'hb0e;
  assign _EVAL_1004 = _EVAL_1208 | _EVAL_1663;
  assign _EVAL_1509 = _EVAL_18 == 12'hc0e;
  assign _EVAL_403 = _EVAL_1004 | _EVAL_1509;
  assign _EVAL_1019 = _EVAL_18 == 12'hb8e;
  assign _EVAL_1449 = _EVAL_403 | _EVAL_1019;
  assign _EVAL_793 = _EVAL_18 == 12'hc8e;
  assign _EVAL_1718 = _EVAL_1449 | _EVAL_793;
  assign _EVAL_1570 = _EVAL_18 == 12'h32f;
  assign _EVAL_615 = _EVAL_1718 | _EVAL_1570;
  assign _EVAL_2188 = _EVAL_18 == 12'hb0f;
  assign _EVAL_1602 = _EVAL_615 | _EVAL_2188;
  assign _EVAL_1349 = _EVAL_18 == 12'hc0f;
  assign _EVAL_1983 = _EVAL_1602 | _EVAL_1349;
  assign _EVAL_329 = _EVAL_18 == 12'hb8f;
  assign _EVAL_1506 = _EVAL_1983 | _EVAL_329;
  assign _EVAL_1064 = _EVAL_18 == 12'hc8f;
  assign _EVAL_1822 = _EVAL_1506 | _EVAL_1064;
  assign _EVAL_908 = _EVAL_18 == 12'h330;
  assign _EVAL_1671 = _EVAL_1822 | _EVAL_908;
  assign _EVAL_1796 = _EVAL_18 == 12'hb10;
  assign _EVAL_1730 = _EVAL_1671 | _EVAL_1796;
  assign _EVAL_371 = _EVAL_18 == 12'hc10;
  assign _EVAL_313 = _EVAL_1730 | _EVAL_371;
  assign _EVAL_2115 = _EVAL_18 == 12'hb90;
  assign _EVAL_1298 = _EVAL_313 | _EVAL_2115;
  assign _EVAL_273 = _EVAL_18 == 12'hc90;
  assign _EVAL_369 = _EVAL_1298 | _EVAL_273;
  assign _EVAL_1780 = _EVAL_18 == 12'h331;
  assign _EVAL_1938 = _EVAL_369 | _EVAL_1780;
  assign _EVAL_2172 = _EVAL_18 == 12'hb11;
  assign _EVAL_2193 = _EVAL_1938 | _EVAL_2172;
  assign _EVAL_1558 = _EVAL_18 == 12'hc11;
  assign _EVAL_2007 = _EVAL_2193 | _EVAL_1558;
  assign _EVAL_2005 = _EVAL_18 == 12'hb91;
  assign _EVAL_988 = _EVAL_2007 | _EVAL_2005;
  assign _EVAL_2097 = _EVAL_18 == 12'hc91;
  assign _EVAL_1580 = _EVAL_988 | _EVAL_2097;
  assign _EVAL_1009 = _EVAL_18 == 12'h332;
  assign _EVAL_193 = _EVAL_1580 | _EVAL_1009;
  assign _EVAL_1052 = _EVAL_18 == 12'hb12;
  assign _EVAL_918 = _EVAL_193 | _EVAL_1052;
  assign _EVAL_937 = _EVAL_18 == 12'hc12;
  assign _EVAL_1658 = _EVAL_918 | _EVAL_937;
  assign _EVAL_1467 = _EVAL_18 == 12'hb92;
  assign _EVAL_228 = _EVAL_1658 | _EVAL_1467;
  assign _EVAL_1465 = _EVAL_18 == 12'hc92;
  assign _EVAL_360 = _EVAL_228 | _EVAL_1465;
  assign _EVAL_352 = _EVAL_23 == 3'h5;
  assign _EVAL_2099 = _EVAL_23 == 3'h6;
  assign _EVAL_1186 = _EVAL_23 == 3'h7;
  assign _EVAL_1014 = _EVAL_102 == 12'h3;
  assign _EVAL_953 = _EVAL_500 ? _EVAL_84 : 32'h0;
  assign _EVAL_257 = _EVAL_953 | _EVAL_87;
  assign _EVAL_428 = _EVAL_257 & _EVAL_2009;
  assign _EVAL_1038 = ~ _EVAL_428;
  assign _EVAL_284 = _EVAL_317 <= 2'h1;
  assign _EVAL_1736 = _EVAL_284 | _EVAL_442;
  assign _EVAL_2079 = {4'h0,_EVAL_77,1'h0,2'h0,_EVAL_6,1'h0,2'h0,_EVAL_165,1'h0,2'h0};
  assign _EVAL_1026 = _EVAL_2079 & 16'h888;
  assign _EVAL_2059 = {{16'd0}, _EVAL_1026};
  assign _EVAL_1289 = _EVAL_2059 & _EVAL_2090;
  assign _EVAL_1348 = ~ _EVAL_1289;
  assign _EVAL_1454 = ~ _EVAL_1348;
  assign _EVAL_497 = _EVAL_1736 ? _EVAL_1454 : 32'h0;
  assign _EVAL_1997 = _EVAL_497[15];
  assign _EVAL_1888 = _EVAL_428[31:8];
  assign _EVAL_912 = _EVAL_1888[7:0];
  assign _EVAL_1547 = _EVAL_912[4:3];
  assign _EVAL_1747 = _EVAL_1547[1];
  assign _EVAL_461 = _EVAL_1479[0];
  assign _EVAL_1092 = {_EVAL_182,_EVAL_461};
  assign _EVAL_1577 = _EVAL_1092 | 31'hf;
  assign _EVAL_578 = _EVAL_1577 + 31'h1;
  assign _EVAL_246 = ~ _EVAL_578;
  assign _EVAL_1433 = _EVAL_1577 & _EVAL_246;
  assign _EVAL_1141 = {_EVAL_1433,2'h3};
  assign _EVAL_375 = 2'h2 == _EVAL_631;
  assign _EVAL_1773 = _EVAL_1769 == 1'h0;
  assign _EVAL_2092 = _EVAL_1773 | _EVAL_2084;
  assign _EVAL_309 = _EVAL_375 & _EVAL_2092;
  assign _EVAL_1722 = _EVAL_102 == 12'h7a2;
  assign _EVAL_1310 = _EVAL_102 == 12'h300;
  assign _EVAL_821 = {{70'd0}, _EVAL_428};
  assign _EVAL_1054 = _EVAL_821[12:11];
  assign _EVAL_753 = _EVAL_1054[0];
  assign _EVAL_1765 = _EVAL_23 == 3'h4;
  assign _EVAL_914 = {_EVAL_102, 20'h0};
  assign _EVAL_1329 = _EVAL_914 & 32'ha0400000;
  assign _EVAL_1326 = _EVAL_1329 == 32'h20000000;
  assign _EVAL_898 = _EVAL_1765 & _EVAL_1326;
  assign _EVAL_1112 = _EVAL_102[10];
  assign _EVAL_1859 = _EVAL_914 & 32'h20100000;
  assign _EVAL_1043 = _EVAL_1859 == 32'h0;
  assign _EVAL_1902 = _EVAL_1765 & _EVAL_1043;
  assign _EVAL_439 = _EVAL_914 & 32'h10100000;
  assign _EVAL_1905 = _EVAL_439 == 32'h100000;
  assign _EVAL_739 = _EVAL_1765 & _EVAL_1905;
  assign _EVAL_1849 = _EVAL_1902 | _EVAL_739;
  assign _EVAL_1937 = _EVAL_1849 | _EVAL_155;
  assign _EVAL_1621 = {{2'd0}, _EVAL_317};
  assign _EVAL_530 = _EVAL_1621 + 4'h8;
  assign _EVAL_1964 = _EVAL_739 ? 32'h3 : _EVAL_78;
  assign _EVAL_579 = _EVAL_1902 ? {{28'd0}, _EVAL_530} : _EVAL_1964;
  assign _EVAL_1334 = _EVAL_579[31];
  assign _EVAL_744 = _EVAL_579[7:0];
  assign _EVAL_750 = _EVAL_744 == 8'he;
  assign _EVAL_679 = _EVAL_1334 & _EVAL_750;
  assign _EVAL_2057 = _EVAL_1073 | _EVAL_679;
  assign _EVAL_1650 = _EVAL_1334 == 1'h0;
  assign _EVAL_1999 = _EVAL_1650 & _EVAL_750;
  assign _EVAL_1087 = _EVAL_2057 | _EVAL_1999;
  assign _EVAL_1380 = _EVAL_1650 & _EVAL_739;
  assign _EVAL_1615 = {_EVAL_2033,1'h0,1'h0,_EVAL_594};
  assign _EVAL_778 = _EVAL_1615 >> _EVAL_317;
  assign _EVAL_1046 = _EVAL_778[0];
  assign _EVAL_1855 = _EVAL_1380 & _EVAL_1046;
  assign _EVAL_620 = _EVAL_1087 | _EVAL_1855;
  assign _EVAL_939 = _EVAL_620 | _EVAL_2084;
  assign _EVAL_386 = _EVAL_317[0];
  assign _EVAL_845 = _EVAL_386 ? 2'h3 : 2'h0;
  assign _EVAL_2017 = _EVAL_102 == 12'h343;
  assign _EVAL_1520 = _EVAL_1 > 2'h0;
  assign _EVAL_1919 = _EVAL_1978 | 30'h7;
  assign _EVAL_826 = _EVAL_102 == 12'h7a0;
  assign _EVAL_913 = _EVAL_826 ? _EVAL_631 : 2'h0;
  assign _EVAL_916 = {{30'd0}, _EVAL_913};
  assign _EVAL_283 = _EVAL_102 == 12'h7a1;
  assign _EVAL_1188 = 2'h1 == _EVAL_631 ? _EVAL_1899 : _EVAL_551;
  assign _EVAL_227 = 2'h2 == _EVAL_631 ? _EVAL_1769 : _EVAL_1188;
  assign _EVAL_343 = 2'h3 == _EVAL_631 ? _EVAL_1763 : _EVAL_227;
  assign _EVAL_2116 = 2'h1 == _EVAL_631 ? _EVAL_1956 : _EVAL_1366;
  assign _EVAL_891 = 2'h2 == _EVAL_631 ? _EVAL_692 : _EVAL_2116;
  assign _EVAL_2008 = 2'h3 == _EVAL_631 ? _EVAL_1877 : _EVAL_891;
  assign _EVAL_2168 = 2'h1 == _EVAL_631 ? _EVAL_1895 : _EVAL_2220;
  assign _EVAL_1098 = 2'h2 == _EVAL_631 ? _EVAL_203 : _EVAL_2168;
  assign _EVAL_1228 = 2'h3 == _EVAL_631 ? 1'h0 : _EVAL_1098;
  assign _EVAL_1051 = 2'h1 == _EVAL_631 ? _EVAL_194 : _EVAL_1425;
  assign _EVAL_1809 = 2'h2 == _EVAL_631 ? _EVAL_1700 : _EVAL_1051;
  assign _EVAL_1481 = 2'h3 == _EVAL_631 ? _EVAL_1494 : _EVAL_1809;
  assign _EVAL_697 = 2'h1 == _EVAL_631 ? _EVAL_1138 : _EVAL_1261;
  assign _EVAL_460 = 2'h2 == _EVAL_631 ? _EVAL_2152 : _EVAL_697;
  assign _EVAL_462 = 2'h3 == _EVAL_631 ? _EVAL_1376 : _EVAL_460;
  assign _EVAL_431 = 2'h1 == _EVAL_631 ? _EVAL_346 : _EVAL_361;
  assign _EVAL_1707 = 2'h2 == _EVAL_631 ? _EVAL_1743 : _EVAL_431;
  assign _EVAL_2046 = 2'h3 == _EVAL_631 ? _EVAL_1421 : _EVAL_1707;
  assign _EVAL_1428 = 2'h1 == _EVAL_631 ? _EVAL_2190 : _EVAL_1986;
  assign _EVAL_719 = 2'h2 == _EVAL_631 ? _EVAL_2063 : _EVAL_1428;
  assign _EVAL_1115 = 2'h3 == _EVAL_631 ? _EVAL_381 : _EVAL_719;
  assign _EVAL_2085 = 2'h1 == _EVAL_631 ? _EVAL_297 : _EVAL_178;
  assign _EVAL_1539 = 2'h2 == _EVAL_631 ? _EVAL_2002 : _EVAL_2085;
  assign _EVAL_1609 = 2'h3 == _EVAL_631 ? _EVAL_1808 : _EVAL_1539;
  assign _EVAL_820 = 2'h1 == _EVAL_631 ? _EVAL_436 : _EVAL_1556;
  assign _EVAL_495 = 2'h2 == _EVAL_631 ? _EVAL_1929 : _EVAL_820;
  assign _EVAL_1842 = 2'h3 == _EVAL_631 ? _EVAL_1241 : _EVAL_495;
  assign _EVAL_1669 = {_EVAL_462,1'h0,1'h0,_EVAL_2046,_EVAL_1115,_EVAL_1609,_EVAL_1842};
  assign _EVAL_1517 = {4'h2,_EVAL_343,14'h400,_EVAL_2008,_EVAL_1228,2'h0,_EVAL_1481,_EVAL_1669};
  assign _EVAL_2174 = _EVAL_283 ? _EVAL_1517 : 32'h0;
  assign _EVAL_1816 = _EVAL_916 | _EVAL_2174;
  assign _EVAL_850 = 2'h1 == _EVAL_631 ? _EVAL_1223 : _EVAL_1063;
  assign _EVAL_1495 = 2'h2 == _EVAL_631 ? _EVAL_900 : _EVAL_850;
  assign _EVAL_222 = 2'h3 == _EVAL_631 ? _EVAL_1725 : _EVAL_1495;
  assign _EVAL_649 = _EVAL_1722 ? _EVAL_222 : 32'h0;
  assign _EVAL_1828 = _EVAL_1816 | _EVAL_649;
  assign _EVAL_1767 = _EVAL_102 == 12'h301;
  assign _EVAL_1100 = _EVAL_1767 ? 31'h40901125 : 31'h0;
  assign _EVAL_1737 = {{1'd0}, _EVAL_1100};
  assign _EVAL_180 = _EVAL_1828 | _EVAL_1737;
  assign _EVAL_1496 = {_EVAL_120,_EVAL_71,_EVAL_8,_EVAL_91,_EVAL_61,_EVAL_36,_EVAL_95};
  assign _EVAL_521 = {_EVAL_52,_EVAL_122,_EVAL_27,_EVAL_111,_EVAL_63,_EVAL_139,_EVAL_94};
  assign _EVAL_689 = {_EVAL_48,_EVAL_124,_EVAL_135,_EVAL_22,_EVAL_73,_EVAL_68,_EVAL_143,_EVAL_130,_EVAL_521};
  assign _EVAL_1003 = {_EVAL_39,_EVAL_92,_EVAL_118,_EVAL_21,_EVAL_76,_EVAL_69,_EVAL_127,_EVAL_138,_EVAL_1496,_EVAL_689};
  assign _EVAL_482 = _EVAL_1003[31:0];
  assign _EVAL_1061 = _EVAL_1310 ? _EVAL_482 : 32'h0;
  assign _EVAL_2021 = _EVAL_180 | _EVAL_1061;
  assign _EVAL_755 = _EVAL_102 == 12'h305;
  assign _EVAL_502 = _EVAL_1239[0];
  assign _EVAL_549 = _EVAL_502 ? 7'h7e : 7'h2;
  assign _EVAL_1970 = {{25'd0}, _EVAL_549};
  assign _EVAL_281 = ~ _EVAL_1970;
  assign _EVAL_1401 = _EVAL_1239 & _EVAL_281;
  assign _EVAL_1681 = _EVAL_755 ? _EVAL_1401 : 32'h0;
  assign _EVAL_2062 = _EVAL_2021 | _EVAL_1681;
  assign _EVAL_569 = _EVAL_102 == 12'h344;
  assign _EVAL_1656 = _EVAL_569 ? _EVAL_1026 : 16'h0;
  assign _EVAL_168 = {{16'd0}, _EVAL_1656};
  assign _EVAL_2215 = _EVAL_2062 | _EVAL_168;
  assign _EVAL_1031 = _EVAL_102 == 12'h304;
  assign _EVAL_630 = _EVAL_1031 ? _EVAL_2090 : 32'h0;
  assign _EVAL_903 = _EVAL_2215 | _EVAL_630;
  assign _EVAL_1752 = _EVAL_102 == 12'h340;
  assign _EVAL_503 = _EVAL_1752 ? _EVAL_1688 : 32'h0;
  assign _EVAL_994 = _EVAL_903 | _EVAL_503;
  assign _EVAL_1291 = _EVAL_102 == 12'h341;
  assign _EVAL_2204 = ~ _EVAL_978;
  assign _EVAL_771 = _EVAL_2204 | 32'h1;
  assign _EVAL_1315 = ~ _EVAL_771;
  assign _EVAL_1893 = _EVAL_1291 ? _EVAL_1315 : 32'h0;
  assign _EVAL_1946 = _EVAL_994 | _EVAL_1893;
  assign _EVAL_2182 = _EVAL_2017 ? _EVAL_745 : 32'h0;
  assign _EVAL_1463 = _EVAL_1946 | _EVAL_2182;
  assign _EVAL_2208 = _EVAL_102 == 12'h342;
  assign _EVAL_1635 = _EVAL_2208 ? _EVAL_422 : 32'h0;
  assign _EVAL_220 = _EVAL_1463 | _EVAL_1635;
  assign _EVAL_262 = _EVAL_102 == 12'hf14;
  assign _EVAL_868 = _EVAL_262 ? _EVAL_86 : 1'h0;
  assign _EVAL_342 = {{31'd0}, _EVAL_868};
  assign _EVAL_1664 = _EVAL_220 | _EVAL_342;
  assign _EVAL_1833 = _EVAL_102 == 12'h7b0;
  assign _EVAL_1190 = {2'h0,1'h0,_EVAL_597,3'h0,_EVAL_762,_EVAL_1466};
  assign _EVAL_1256 = {4'h4,12'h0,_EVAL_2033,2'h0,_EVAL_594,_EVAL_1190};
  assign _EVAL_210 = _EVAL_1833 ? _EVAL_1256 : 32'h0;
  assign _EVAL_188 = _EVAL_1664 | _EVAL_210;
  assign _EVAL_1297 = _EVAL_102 == 12'h7b1;
  assign _EVAL_173 = ~ _EVAL_1589;
  assign _EVAL_711 = _EVAL_173 | 32'h1;
  assign _EVAL_1032 = ~ _EVAL_711;
  assign _EVAL_831 = _EVAL_1297 ? _EVAL_1032 : 32'h0;
  assign _EVAL_1293 = _EVAL_188 | _EVAL_831;
  assign _EVAL_2143 = _EVAL_102 == 12'h7b2;
  assign _EVAL_1320 = _EVAL_2143 ? _EVAL_1632 : 32'h0;
  assign _EVAL_885 = _EVAL_1293 | _EVAL_1320;
  assign _EVAL_1713 = _EVAL_102 == 12'h1;
  assign _EVAL_940 = _EVAL_1713 ? _EVAL_584 : 5'h0;
  assign _EVAL_487 = {{27'd0}, _EVAL_940};
  assign _EVAL_377 = _EVAL_885 | _EVAL_487;
  assign _EVAL_772 = _EVAL_102 == 12'h2;
  assign _EVAL_1288 = _EVAL_772 ? _EVAL_1458 : 3'h0;
  assign _EVAL_1127 = {{29'd0}, _EVAL_1288};
  assign _EVAL_1347 = _EVAL_377 | _EVAL_1127;
  assign _EVAL_684 = {_EVAL_1458,_EVAL_584};
  assign _EVAL_2122 = _EVAL_1014 ? _EVAL_684 : 8'h0;
  assign _EVAL_1731 = {{24'd0}, _EVAL_2122};
  assign _EVAL_2011 = _EVAL_1347 | _EVAL_1731;
  assign _EVAL_817 = {{32'd0}, _EVAL_2011};
  assign _EVAL_531 = _EVAL_102 == 12'hb00;
  assign _EVAL_2070 = {_EVAL_1212,_EVAL_1419};
  assign _EVAL_656 = _EVAL_531 ? _EVAL_2070 : 64'h0;
  assign _EVAL_2112 = _EVAL_817 | _EVAL_656;
  assign _EVAL_1559 = _EVAL_102 == 12'hb02;
  assign _EVAL_720 = {_EVAL_751,_EVAL_1249};
  assign _EVAL_1514 = _EVAL_1559 ? _EVAL_720 : 64'h0;
  assign _EVAL_2102 = _EVAL_2112 | _EVAL_1514;
  assign _EVAL_1923 = _EVAL_2099 | _EVAL_1186;
  assign _EVAL_1627 = _EVAL_1923 | _EVAL_352;
  assign _EVAL_1746 = _EVAL_102 == 12'h3a1;
  assign _EVAL_1913 = _EVAL_333 == 1'h0;
  assign _EVAL_749 = _EVAL_1746 & _EVAL_1913;
  assign _EVAL_430 = _EVAL_428[31:24];
  assign _EVAL_2163 = _EVAL_430[7];
  assign _EVAL_857 = _EVAL_428[7:0];
  assign _EVAL_1143 = _EVAL_857[4:3];
  assign _EVAL_1515 = _EVAL_1143[1];
  assign _EVAL_635 = ~ _EVAL;
  assign _EVAL_1759 = _EVAL_635 | 32'h1;
  assign _EVAL_1588 = {_EVAL_1261,1'h0,1'h0,_EVAL_361,_EVAL_1986,_EVAL_178,_EVAL_1556};
  assign _EVAL_688 = {4'h2,_EVAL_551,14'h400,_EVAL_1366,_EVAL_2220,2'h0,_EVAL_1425,_EVAL_1588};
  assign _EVAL_1359 = _EVAL_500 ? _EVAL_688 : 32'h0;
  assign _EVAL_1096 = _EVAL_1359 | _EVAL_87;
  assign _EVAL_1236 = _EVAL_1096 & _EVAL_2009;
  assign _EVAL_2162 = _EVAL_1236[12];
  assign _EVAL_1408 = _EVAL_1011[0];
  assign _EVAL_946 = {_EVAL_1942,_EVAL_1408};
  assign _EVAL_318 = {_EVAL_1138,1'h0,1'h0,_EVAL_346,_EVAL_2190,_EVAL_297,_EVAL_436};
  assign _EVAL_1945 = {4'h2,_EVAL_1899,14'h400,_EVAL_1956,_EVAL_1895,2'h0,_EVAL_194,_EVAL_318};
  assign _EVAL_1889 = _EVAL_500 ? _EVAL_1945 : 32'h0;
  assign _EVAL_1445 = 2'h0 == _EVAL_631;
  assign _EVAL_1702 = _EVAL_551 == 1'h0;
  assign _EVAL_2073 = _EVAL_1702 | _EVAL_2084;
  assign _EVAL_270 = _EVAL_1445 & _EVAL_2073;
  assign _EVAL_1590 = _EVAL_428[2];
  assign _EVAL_1286 = 2'h1 == _EVAL_631;
  assign _EVAL_412 = _EVAL_1899 == 1'h0;
  assign _EVAL_1050 = _EVAL_412 | _EVAL_2084;
  assign _EVAL_1151 = _EVAL_1286 & _EVAL_1050;
  assign _EVAL_830 = _EVAL_428[1];
  assign _EVAL_1091 = _EVAL_1555 == 1'h0;
  assign _EVAL_1644 = _EVAL_1746 & _EVAL_1091;
  assign _EVAL_1680 = _EVAL_428[31:16];
  assign _EVAL_1741 = _EVAL_1680[7:0];
  assign _EVAL_243 = _EVAL_1741[2];
  assign _EVAL_484 = _EVAL_102 == 12'h3b7;
  assign _EVAL_1504 = _EVAL_1282 & 32'h1f;
  assign _EVAL_1389 = _EVAL_1895 == 1'h0;
  assign _EVAL_396 = _EVAL_1899 | _EVAL_1389;
  assign _EVAL_707 = _EVAL_428[0];
  assign _EVAL_2114 = {_EVAL_2106,_EVAL_2177};
  assign _EVAL_1972 = _EVAL_2114[31:0];
  assign _EVAL_658 = {_EVAL_857,_EVAL_1972};
  assign _EVAL_402 = _EVAL_2181[1];
  assign _EVAL_474 = _EVAL_842 | 30'h7;
  assign _EVAL_1074 = ~ _EVAL_842;
  assign _EVAL_2032 = _EVAL_1074 | 30'hf;
  assign _EVAL_169 = ~ _EVAL_2032;
  assign _EVAL_1623 = _EVAL_402 ? _EVAL_474 : _EVAL_169;
  assign _EVAL_1426 = _EVAL_1440[1];
  assign _EVAL_666 = _EVAL_102 == 12'h323;
  assign _EVAL_738 = _EVAL_666 ? _EVAL_537 : 32'h0;
  assign _EVAL_769 = {{32'd0}, _EVAL_738};
  assign _EVAL_1640 = _EVAL_2102 | _EVAL_769;
  assign _EVAL_1358 = _EVAL_102 == 12'hb03;
  assign _EVAL_981 = {_EVAL_171,_EVAL_305};
  assign _EVAL_445 = _EVAL_1358 ? _EVAL_981 : 40'h0;
  assign _EVAL_251 = {{24'd0}, _EVAL_445};
  assign _EVAL_1474 = _EVAL_1640 | _EVAL_251;
  assign _EVAL_2066 = _EVAL_102 == 12'hc03;
  assign _EVAL_449 = _EVAL_2066 ? _EVAL_981 : 40'h0;
  assign _EVAL_1535 = {{24'd0}, _EVAL_449};
  assign _EVAL_876 = _EVAL_1474 | _EVAL_1535;
  assign _EVAL_1374 = _EVAL_102 == 12'hb83;
  assign _EVAL_389 = _EVAL_981[39:32];
  assign _EVAL_1174 = _EVAL_1374 ? _EVAL_389 : 8'h0;
  assign _EVAL_1988 = {{56'd0}, _EVAL_1174};
  assign _EVAL_1021 = _EVAL_876 | _EVAL_1988;
  assign _EVAL_800 = _EVAL_102 == 12'hc83;
  assign _EVAL_977 = _EVAL_800 ? _EVAL_389 : 8'h0;
  assign _EVAL_2236 = {{56'd0}, _EVAL_977};
  assign _EVAL_1631 = _EVAL_1021 | _EVAL_2236;
  assign _EVAL_1617 = _EVAL_102 == 12'h324;
  assign _EVAL_870 = _EVAL_1617 ? _EVAL_1048 : 32'h0;
  assign _EVAL_459 = {{32'd0}, _EVAL_870};
  assign _EVAL_1748 = _EVAL_1631 | _EVAL_459;
  assign _EVAL_1437 = _EVAL_102 == 12'hb04;
  assign _EVAL_1122 = _EVAL_1437 ? _EVAL_2114 : 40'h0;
  assign _EVAL_583 = {{24'd0}, _EVAL_1122};
  assign _EVAL_1350 = _EVAL_1748 | _EVAL_583;
  assign _EVAL_316 = _EVAL_102 == 12'hc04;
  assign _EVAL_340 = _EVAL_316 ? _EVAL_2114 : 40'h0;
  assign _EVAL_1678 = {{24'd0}, _EVAL_340};
  assign _EVAL_1977 = _EVAL_1350 | _EVAL_1678;
  assign _EVAL_1386 = _EVAL_102 == 12'hb84;
  assign _EVAL_2069 = _EVAL_2114[39:32];
  assign _EVAL_1789 = _EVAL_1386 ? _EVAL_2069 : 8'h0;
  assign _EVAL_680 = {{56'd0}, _EVAL_1789};
  assign _EVAL_1578 = _EVAL_1977 | _EVAL_680;
  assign _EVAL_1560 = _EVAL_102 == 12'hc84;
  assign _EVAL_1448 = _EVAL_1560 ? _EVAL_2069 : 8'h0;
  assign _EVAL_1571 = {{56'd0}, _EVAL_1448};
  assign _EVAL_457 = _EVAL_1578 | _EVAL_1571;
  assign _EVAL_677 = _EVAL_102 == 12'h306;
  assign _EVAL_1873 = _EVAL_677 ? _EVAL_1504 : 32'h0;
  assign _EVAL_1311 = {{32'd0}, _EVAL_1873};
  assign _EVAL_702 = _EVAL_457 | _EVAL_1311;
  assign _EVAL_425 = _EVAL_102 == 12'hc00;
  assign _EVAL_1784 = _EVAL_425 ? _EVAL_2070 : 64'h0;
  assign _EVAL_705 = _EVAL_702 | _EVAL_1784;
  assign _EVAL_323 = _EVAL_102 == 12'hc02;
  assign _EVAL_550 = _EVAL_323 ? _EVAL_720 : 64'h0;
  assign _EVAL_322 = _EVAL_705 | _EVAL_550;
  assign _EVAL_1657 = _EVAL_102 == 12'hb80;
  assign _EVAL_1724 = _EVAL_2070[63:32];
  assign _EVAL_1471 = _EVAL_1657 ? _EVAL_1724 : 32'h0;
  assign _EVAL_1077 = {{32'd0}, _EVAL_1471};
  assign _EVAL_1568 = _EVAL_322 | _EVAL_1077;
  assign _EVAL_1872 = _EVAL_102 == 12'hb82;
  assign _EVAL_881 = _EVAL_720[63:32];
  assign _EVAL_1272 = _EVAL_1872 ? _EVAL_881 : 32'h0;
  assign _EVAL_1613 = {{32'd0}, _EVAL_1272};
  assign _EVAL_1117 = _EVAL_1568 | _EVAL_1613;
  assign _EVAL_596 = _EVAL_102 == 12'hc80;
  assign _EVAL_607 = _EVAL_596 ? _EVAL_1724 : 32'h0;
  assign _EVAL_258 = {{32'd0}, _EVAL_607};
  assign _EVAL_192 = _EVAL_1117 | _EVAL_258;
  assign _EVAL_212 = _EVAL_102 == 12'hc82;
  assign _EVAL_394 = _EVAL_212 ? _EVAL_881 : 32'h0;
  assign _EVAL_1431 = {{32'd0}, _EVAL_394};
  assign _EVAL_1936 = _EVAL_192 | _EVAL_1431;
  assign _EVAL_1213 = _EVAL_102 == 12'h3a0;
  assign _EVAL_2104 = {_EVAL_181,2'h0,_EVAL_491,_EVAL_941,_EVAL_1193,_EVAL_2238};
  assign _EVAL_1364 = {_EVAL_2232,2'h0,_EVAL_2181,_EVAL_992,_EVAL_1022,_EVAL_1770};
  assign _EVAL_2094 = {_EVAL_1593,2'h0,_EVAL_2227,_EVAL_1608,_EVAL_1792,_EVAL_334,_EVAL_1364};
  assign _EVAL_525 = {_EVAL_611,2'h0,_EVAL_1479,_EVAL_710,_EVAL_1062,_EVAL_958,_EVAL_2104,_EVAL_2094};
  assign _EVAL_742 = _EVAL_1213 ? _EVAL_525 : 32'h0;
  assign _EVAL_321 = {{32'd0}, _EVAL_742};
  assign _EVAL_362 = _EVAL_1936 | _EVAL_321;
  assign _EVAL_1296 = {_EVAL_1555,2'h0,_EVAL_715,_EVAL_2131,_EVAL_2180,_EVAL_1733};
  assign _EVAL_888 = {_EVAL_1168,2'h0,_EVAL_2226,_EVAL_523,_EVAL_1499,_EVAL_1620};
  assign _EVAL_737 = {_EVAL_1585,2'h0,_EVAL_1440,_EVAL_1167,_EVAL_2047,_EVAL_1563,_EVAL_888};
  assign _EVAL_548 = {_EVAL_333,2'h0,_EVAL_1011,_EVAL_1869,_EVAL_207,_EVAL_1385,_EVAL_1296,_EVAL_737};
  assign _EVAL_1548 = _EVAL_1746 ? _EVAL_548 : 32'h0;
  assign _EVAL_1887 = {{32'd0}, _EVAL_1548};
  assign _EVAL_359 = _EVAL_362 | _EVAL_1887;
  assign _EVAL_1396 = _EVAL_102 == 12'h3b0;
  assign _EVAL_1086 = _EVAL_1396 ? _EVAL_1623 : 30'h0;
  assign _EVAL_478 = {{34'd0}, _EVAL_1086};
  assign _EVAL_419 = _EVAL_359 | _EVAL_478;
  assign _EVAL_237 = _EVAL_102 == 12'h3b1;
  assign _EVAL_1307 = _EVAL_2227[1];
  assign _EVAL_1321 = _EVAL_2224 | 30'h7;
  assign _EVAL_1645 = ~ _EVAL_2224;
  assign _EVAL_752 = _EVAL_1645 | 30'hf;
  assign _EVAL_1507 = ~ _EVAL_752;
  assign _EVAL_339 = _EVAL_1307 ? _EVAL_1321 : _EVAL_1507;
  assign _EVAL_1890 = _EVAL_237 ? _EVAL_339 : 30'h0;
  assign _EVAL_646 = {{34'd0}, _EVAL_1890};
  assign _EVAL_1948 = _EVAL_419 | _EVAL_646;
  assign _EVAL_780 = _EVAL_102 == 12'h3b2;
  assign _EVAL_681 = _EVAL_491[1];
  assign _EVAL_1101 = _EVAL_1952 | 30'h7;
  assign _EVAL_198 = ~ _EVAL_1952;
  assign _EVAL_1907 = _EVAL_198 | 30'hf;
  assign _EVAL_1118 = ~ _EVAL_1907;
  assign _EVAL_1278 = _EVAL_681 ? _EVAL_1101 : _EVAL_1118;
  assign _EVAL_1171 = _EVAL_780 ? _EVAL_1278 : 30'h0;
  assign _EVAL_798 = {{34'd0}, _EVAL_1171};
  assign _EVAL_1668 = _EVAL_1948 | _EVAL_798;
  assign _EVAL_539 = _EVAL_102 == 12'h3b3;
  assign _EVAL_2151 = _EVAL_1479[1];
  assign _EVAL_947 = _EVAL_182 | 30'h7;
  assign _EVAL_1629 = ~ _EVAL_182;
  assign _EVAL_411 = _EVAL_1629 | 30'hf;
  assign _EVAL_1961 = ~ _EVAL_411;
  assign _EVAL_347 = _EVAL_2151 ? _EVAL_947 : _EVAL_1961;
  assign _EVAL_1492 = _EVAL_539 ? _EVAL_347 : 30'h0;
  assign _EVAL_1018 = {{34'd0}, _EVAL_1492};
  assign _EVAL_854 = _EVAL_1668 | _EVAL_1018;
  assign _EVAL_1647 = _EVAL_102 == 12'h3b4;
  assign _EVAL_1306 = _EVAL_2226[1];
  assign _EVAL_298 = _EVAL_2210 | 30'h7;
  assign _EVAL_1628 = ~ _EVAL_2210;
  assign _EVAL_2018 = _EVAL_1628 | 30'hf;
  assign _EVAL_896 = ~ _EVAL_2018;
  assign _EVAL_970 = _EVAL_1306 ? _EVAL_298 : _EVAL_896;
  assign _EVAL_517 = _EVAL_1647 ? _EVAL_970 : 30'h0;
  assign _EVAL_1202 = {{34'd0}, _EVAL_517};
  assign _EVAL_1238 = _EVAL_854 | _EVAL_1202;
  assign _EVAL_1418 = _EVAL_102 == 12'h3b5;
  assign _EVAL_887 = _EVAL_286 | 30'h7;
  assign _EVAL_1406 = ~ _EVAL_286;
  assign _EVAL_2239 = _EVAL_1406 | 30'hf;
  assign _EVAL_1979 = ~ _EVAL_2239;
  assign _EVAL_2156 = _EVAL_1426 ? _EVAL_887 : _EVAL_1979;
  assign _EVAL_509 = _EVAL_1418 ? _EVAL_2156 : 30'h0;
  assign _EVAL_811 = {{34'd0}, _EVAL_509};
  assign _EVAL_546 = _EVAL_1238 | _EVAL_811;
  assign _EVAL_1285 = _EVAL_102 == 12'h3b6;
  assign _EVAL_984 = _EVAL_715[1];
  assign _EVAL_775 = ~ _EVAL_1978;
  assign _EVAL_1832 = _EVAL_775 | 30'hf;
  assign _EVAL_682 = ~ _EVAL_1832;
  assign _EVAL_2150 = _EVAL_984 ? _EVAL_1919 : _EVAL_682;
  assign _EVAL_641 = _EVAL_1285 ? _EVAL_2150 : 30'h0;
  assign _EVAL_895 = {{34'd0}, _EVAL_641};
  assign _EVAL_1625 = _EVAL_546 | _EVAL_895;
  assign _EVAL_279 = _EVAL_1011[1];
  assign _EVAL_1891 = _EVAL_1942 | 30'h7;
  assign _EVAL_655 = ~ _EVAL_1942;
  assign _EVAL_224 = _EVAL_655 | 30'hf;
  assign _EVAL_1015 = ~ _EVAL_224;
  assign _EVAL_1508 = _EVAL_279 ? _EVAL_1891 : _EVAL_1015;
  assign _EVAL_395 = _EVAL_484 ? _EVAL_1508 : 30'h0;
  assign _EVAL_1672 = {{34'd0}, _EVAL_395};
  assign _EVAL_2187 = _EVAL_1625 | _EVAL_1672;
  assign _EVAL_1864 = _EVAL_102 == 12'h7c1;
  assign _EVAL_280 = _EVAL_1864 ? _EVAL_1532 : 32'h0;
  assign _EVAL_1372 = {{32'd0}, _EVAL_280};
  assign _EVAL_1404 = _EVAL_2187 | _EVAL_1372;
  assign _EVAL_747 = _EVAL_102 == 12'hf11;
  assign _EVAL_1659 = _EVAL_747 ? 32'h489 : 32'h0;
  assign _EVAL_293 = {{32'd0}, _EVAL_1659};
  assign _EVAL_176 = _EVAL_1404 | _EVAL_293;
  assign _EVAL_2155 = _EVAL_102 == 12'hf12;
  assign _EVAL_1468 = _EVAL_2155 ? 32'h80000007 : 32'h0;
  assign _EVAL_387 = {{32'd0}, _EVAL_1468};
  assign _EVAL_1442 = _EVAL_176 | _EVAL_387;
  assign _EVAL_1500 = _EVAL_102 == 12'hf13;
  assign _EVAL_1361 = _EVAL_1500 ? 32'h20191204 : 32'h0;
  assign _EVAL_1475 = {{32'd0}, _EVAL_1361};
  assign _EVAL_351 = _EVAL_1442 | _EVAL_1475;
  assign _EVAL_1715 = _EVAL_1168 == 1'h0;
  assign _EVAL_2120 = _EVAL_1746 & _EVAL_1715;
  assign _EVAL_1831 = _EVAL_857[0];
  assign _EVAL_733 = _EVAL_984 == 1'h0;
  assign _EVAL_924 = _EVAL_715[0];
  assign _EVAL_797 = _EVAL_733 & _EVAL_924;
  assign _EVAL_1120 = _EVAL_1555 & _EVAL_797;
  assign _EVAL_848 = _EVAL_1585 | _EVAL_1120;
  assign _EVAL_832 = _EVAL_848 == 1'h0;
  assign _EVAL_1260 = _EVAL_1418 & _EVAL_832;
  assign _EVAL_405 = _EVAL_18 >= 12'hc80;
  assign _EVAL_1696 = _EVAL_18 == 12'h333;
  assign _EVAL_538 = _EVAL_360 | _EVAL_1696;
  assign _EVAL_1540 = _EVAL_18 == 12'hb13;
  assign _EVAL_1387 = _EVAL_538 | _EVAL_1540;
  assign _EVAL_901 = _EVAL_18 == 12'hc13;
  assign _EVAL_2207 = _EVAL_1387 | _EVAL_901;
  assign _EVAL_1427 = _EVAL_18 == 12'hb93;
  assign _EVAL_1959 = _EVAL_2207 | _EVAL_1427;
  assign _EVAL_1469 = _EVAL_18 == 12'hc93;
  assign _EVAL_2054 = _EVAL_1959 | _EVAL_1469;
  assign _EVAL_418 = _EVAL_18 == 12'h334;
  assign _EVAL_1482 = _EVAL_2054 | _EVAL_418;
  assign _EVAL_512 = _EVAL_18 == 12'hb14;
  assign _EVAL_1163 = _EVAL_1482 | _EVAL_512;
  assign _EVAL_392 = _EVAL_18 == 12'hc14;
  assign _EVAL_1330 = _EVAL_1163 | _EVAL_392;
  assign _EVAL_625 = _EVAL_18 == 12'hb94;
  assign _EVAL_260 = _EVAL_1330 | _EVAL_625;
  assign _EVAL_761 = _EVAL_18 == 12'hc94;
  assign _EVAL_1875 = _EVAL_260 | _EVAL_761;
  assign _EVAL_1345 = _EVAL_18 == 12'h335;
  assign _EVAL_2030 = _EVAL_1875 | _EVAL_1345;
  assign _EVAL_1840 = _EVAL_18 == 12'hb15;
  assign _EVAL_1160 = _EVAL_2030 | _EVAL_1840;
  assign _EVAL_957 = _EVAL_18 == 12'hc15;
  assign _EVAL_612 = _EVAL_1160 | _EVAL_957;
  assign _EVAL_337 = _EVAL_18 == 12'hb95;
  assign _EVAL_1565 = _EVAL_612 | _EVAL_337;
  assign _EVAL_987 = _EVAL_18 == 12'hc95;
  assign _EVAL_324 = _EVAL_1565 | _EVAL_987;
  assign _EVAL_657 = _EVAL_18 == 12'h336;
  assign _EVAL_274 = _EVAL_324 | _EVAL_657;
  assign _EVAL_437 = _EVAL_18 == 12'hb16;
  assign _EVAL_1799 = _EVAL_274 | _EVAL_437;
  assign _EVAL_2056 = _EVAL_18 == 12'hc16;
  assign _EVAL_884 = _EVAL_1799 | _EVAL_2056;
  assign _EVAL_2071 = _EVAL_18 == 12'hb96;
  assign _EVAL_781 = _EVAL_884 | _EVAL_2071;
  assign _EVAL_254 = _EVAL_18 == 12'hc96;
  assign _EVAL_547 = _EVAL_781 | _EVAL_254;
  assign _EVAL_315 = _EVAL_18 == 12'h337;
  assign _EVAL_1430 = _EVAL_547 | _EVAL_315;
  assign _EVAL_299 = _EVAL_18 == 12'hb17;
  assign _EVAL_1219 = _EVAL_1430 | _EVAL_299;
  assign _EVAL_327 = _EVAL_18 == 12'hc17;
  assign _EVAL_672 = _EVAL_1219 | _EVAL_327;
  assign _EVAL_2179 = _EVAL_18 == 12'hb97;
  assign _EVAL_527 = _EVAL_672 | _EVAL_2179;
  assign _EVAL_435 = _EVAL_527 | _EVAL_197;
  assign _EVAL_1584 = _EVAL_18 == 12'h338;
  assign _EVAL_961 = _EVAL_435 | _EVAL_1584;
  assign _EVAL_426 = _EVAL_18 == 12'hb18;
  assign _EVAL_622 = _EVAL_961 | _EVAL_426;
  assign _EVAL_974 = _EVAL_981[39:32];
  assign _EVAL_899 = {_EVAL_974,_EVAL_428};
  assign _EVAL_2154 = _EVAL_899[39:6];
  assign _EVAL_534 = {{4'd0}, _EVAL_41};
  assign _EVAL_1575 = _EVAL_305 + _EVAL_534;
  assign _EVAL_1156 = _EVAL_1575[6];
  assign _EVAL_1800 = _EVAL_171 + 34'h1;
  assign _EVAL_1900 = _EVAL_18[10];
  assign _EVAL_1234 = _EVAL_18 == 12'hc18;
  assign _EVAL_1851 = _EVAL_622 | _EVAL_1234;
  assign _EVAL_676 = _EVAL_18 == 12'hb98;
  assign _EVAL_1137 = _EVAL_1851 | _EVAL_676;
  assign _EVAL_1764 = _EVAL_18 == 12'hc98;
  assign _EVAL_2229 = _EVAL_1137 | _EVAL_1764;
  assign _EVAL_1035 = _EVAL_18 == 12'h339;
  assign _EVAL_822 = _EVAL_2229 | _EVAL_1035;
  assign _EVAL_1184 = _EVAL_18 == 12'hb19;
  assign _EVAL_1231 = _EVAL_822 | _EVAL_1184;
  assign _EVAL_1850 = _EVAL_18 == 12'hc19;
  assign _EVAL_1082 = _EVAL_1231 | _EVAL_1850;
  assign _EVAL_356 = _EVAL_18 == 12'hb99;
  assign _EVAL_1966 = _EVAL_1082 | _EVAL_356;
  assign _EVAL_399 = _EVAL_18 == 12'hc99;
  assign _EVAL_889 = _EVAL_1966 | _EVAL_399;
  assign _EVAL_1598 = _EVAL_18 == 12'h33a;
  assign _EVAL_545 = _EVAL_889 | _EVAL_1598;
  assign _EVAL_400 = _EVAL_18 == 12'hb1a;
  assign _EVAL_314 = _EVAL_545 | _EVAL_400;
  assign _EVAL_380 = _EVAL_18 == 12'hc1a;
  assign _EVAL_1155 = _EVAL_314 | _EVAL_380;
  assign _EVAL_2125 = _EVAL_18 == 12'hb9a;
  assign _EVAL_1931 = _EVAL_1155 | _EVAL_2125;
  assign _EVAL_782 = _EVAL_18 == 12'hc9a;
  assign _EVAL_1597 = _EVAL_1931 | _EVAL_782;
  assign _EVAL_1001 = _EVAL_18 == 12'h33b;
  assign _EVAL_1630 = _EVAL_1597 | _EVAL_1001;
  assign _EVAL_905 = _EVAL_18 == 12'hb1b;
  assign _EVAL_919 = _EVAL_1630 | _EVAL_905;
  assign _EVAL_1455 = _EVAL_18 == 12'hc1b;
  assign _EVAL_1287 = _EVAL_919 | _EVAL_1455;
  assign _EVAL_893 = _EVAL_18 == 12'hb9b;
  assign _EVAL_2136 = _EVAL_1287 | _EVAL_893;
  assign _EVAL_867 = _EVAL_18 == 12'hc9b;
  assign _EVAL_2012 = _EVAL_2136 | _EVAL_867;
  assign _EVAL_1667 = _EVAL_18 == 12'h33c;
  assign _EVAL_2100 = _EVAL_2012 | _EVAL_1667;
  assign _EVAL_823 = _EVAL_18 == 12'hb1c;
  assign _EVAL_1157 = _EVAL_2100 | _EVAL_823;
  assign _EVAL_1554 = _EVAL_18 == 12'hc1c;
  assign _EVAL_2080 = _EVAL_1157 | _EVAL_1554;
  assign _EVAL_567 = _EVAL_18 == 12'hb9c;
  assign _EVAL_963 = _EVAL_2080 | _EVAL_567;
  assign _EVAL_673 = _EVAL_18 == 12'hc9c;
  assign _EVAL_345 = _EVAL_963 | _EVAL_673;
  assign _EVAL_2127 = _EVAL_18 == 12'h33d;
  assign _EVAL_1189 = _EVAL_345 | _EVAL_2127;
  assign _EVAL_1453 = _EVAL_18 == 12'hb1d;
  assign _EVAL_1246 = _EVAL_1189 | _EVAL_1453;
  assign _EVAL_1818 = _EVAL_18 == 12'hc1d;
  assign _EVAL_1594 = _EVAL_1246 | _EVAL_1818;
  assign _EVAL_1512 = _EVAL_18 == 12'hb9d;
  assign _EVAL_971 = _EVAL_1594 | _EVAL_1512;
  assign _EVAL_190 = _EVAL_18 == 12'hc9d;
  assign _EVAL_2050 = _EVAL_971 | _EVAL_190;
  assign _EVAL_1502 = _EVAL_18 == 12'h33e;
  assign _EVAL_2138 = _EVAL_2050 | _EVAL_1502;
  assign _EVAL_954 = _EVAL_18 == 12'hb1e;
  assign _EVAL_902 = _EVAL_2138 | _EVAL_954;
  assign _EVAL_1491 = _EVAL_18 == 12'hc1e;
  assign _EVAL_1994 = _EVAL_902 | _EVAL_1491;
  assign _EVAL_1879 = _EVAL_18 == 12'hb9e;
  assign _EVAL_1526 = _EVAL_1994 | _EVAL_1879;
  assign _EVAL_786 = _EVAL_18 == 12'hc9e;
  assign _EVAL_1402 = _EVAL_1526 | _EVAL_786;
  assign _EVAL_1804 = _EVAL_18 == 12'h33f;
  assign _EVAL_448 = _EVAL_1402 | _EVAL_1804;
  assign _EVAL_1538 = _EVAL_18 == 12'hb1f;
  assign _EVAL_1362 = _EVAL_448 | _EVAL_1538;
  assign _EVAL_1016 = _EVAL_18 == 12'hc1f;
  assign _EVAL_508 = _EVAL_1362 | _EVAL_1016;
  assign _EVAL_1884 = _EVAL_18 == 12'hb9f;
  assign _EVAL_1203 = _EVAL_508 | _EVAL_1884;
  assign _EVAL_185 = _EVAL_18 == 12'hc9f;
  assign _EVAL_215 = _EVAL_1203 | _EVAL_185;
  assign _EVAL_1114 = _EVAL_18 == 12'h306;
  assign _EVAL_979 = _EVAL_215 | _EVAL_1114;
  assign _EVAL_486 = _EVAL_18 == 12'hc00;
  assign _EVAL_1486 = _EVAL_979 | _EVAL_486;
  assign _EVAL_1673 = _EVAL_18 == 12'hc02;
  assign _EVAL_1965 = _EVAL_1486 | _EVAL_1673;
  assign _EVAL_1244 = _EVAL_18 == 12'hb80;
  assign _EVAL_470 = _EVAL_1965 | _EVAL_1244;
  assign _EVAL_344 = _EVAL_18 == 12'hb82;
  assign _EVAL_1882 = _EVAL_470 | _EVAL_344;
  assign _EVAL_2157 = _EVAL_18 == 12'hc80;
  assign _EVAL_967 = _EVAL_1882 | _EVAL_2157;
  assign _EVAL_2118 = _EVAL_18 == 12'hc82;
  assign _EVAL_2013 = _EVAL_967 | _EVAL_2118;
  assign _EVAL_1709 = _EVAL_18 == 12'h3a0;
  assign _EVAL_1553 = _EVAL_2013 | _EVAL_1709;
  assign _EVAL_746 = _EVAL_18 == 12'h3a1;
  assign _EVAL_496 = _EVAL_1553 | _EVAL_746;
  assign _EVAL_1384 = _EVAL_18 == 12'h3a2;
  assign _EVAL_1369 = _EVAL_496 | _EVAL_1384;
  assign _EVAL_1483 = _EVAL_18 == 12'h3a3;
  assign _EVAL_2211 = _EVAL_1369 | _EVAL_1483;
  assign _EVAL_1939 = _EVAL_18 == 12'h3b0;
  assign _EVAL_807 = _EVAL_2211 | _EVAL_1939;
  assign _EVAL_384 = _EVAL_18 == 12'h3b1;
  assign _EVAL_231 = _EVAL_807 | _EVAL_384;
  assign _EVAL_1519 = _EVAL_18 == 12'h3b2;
  assign _EVAL_566 = _EVAL_231 | _EVAL_1519;
  assign _EVAL_1912 = _EVAL_18 == 12'h3b3;
  assign _EVAL_1023 = _EVAL_566 | _EVAL_1912;
  assign _EVAL_196 = _EVAL_18 == 12'h3b4;
  assign _EVAL_2049 = _EVAL_1023 | _EVAL_196;
  assign _EVAL_968 = _EVAL_18 == 12'h3b5;
  assign _EVAL_1968 = _EVAL_2049 | _EVAL_968;
  assign _EVAL_1920 = _EVAL_18 == 12'h3b6;
  assign _EVAL_647 = _EVAL_1968 | _EVAL_1920;
  assign _EVAL_932 = _EVAL_18 == 12'h3b7;
  assign _EVAL_1774 = _EVAL_647 | _EVAL_932;
  assign _EVAL_700 = _EVAL_18 == 12'h3b8;
  assign _EVAL_1182 = _EVAL_1774 | _EVAL_700;
  assign _EVAL_1149 = _EVAL_18 == 12'h3b9;
  assign _EVAL_1534 = _EVAL_1182 | _EVAL_1149;
  assign _EVAL_1017 = _EVAL_18 == 12'h3ba;
  assign _EVAL_776 = _EVAL_1534 | _EVAL_1017;
  assign _EVAL_648 = _EVAL_18 == 12'h3bb;
  assign _EVAL_374 = _EVAL_776 | _EVAL_648;
  assign _EVAL_558 = _EVAL_18 == 12'h3bc;
  assign _EVAL_1761 = _EVAL_374 | _EVAL_558;
  assign _EVAL_1180 = _EVAL_18 == 12'h3bd;
  assign _EVAL_1601 = _EVAL_1761 | _EVAL_1180;
  assign _EVAL_205 = _EVAL_18 == 12'h3be;
  assign _EVAL_2218 = _EVAL_1601 | _EVAL_205;
  assign _EVAL_643 = _EVAL_18 == 12'h3bf;
  assign _EVAL_492 = _EVAL_2218 | _EVAL_643;
  assign _EVAL_2200 = _EVAL_18 == 12'h7c1;
  assign _EVAL_532 = _EVAL_492 | _EVAL_2200;
  assign _EVAL_287 = _EVAL_18 == 12'hf11;
  assign _EVAL_244 = _EVAL_532 | _EVAL_287;
  assign _EVAL_1754 = _EVAL_18 == 12'hf12;
  assign _EVAL_731 = _EVAL_244 | _EVAL_1754;
  assign _EVAL_973 = _EVAL_1236[11];
  assign _EVAL_208 = _EVAL_973 & _EVAL_1389;
  assign _EVAL_1211 = _EVAL_1236[27];
  assign _EVAL_670 = _EVAL_1211 & _EVAL_2084;
  assign _EVAL_1595 = _EVAL_670 | _EVAL_412;
  assign _EVAL_1973 = _EVAL_208 & _EVAL_1595;
  assign _EVAL_602 = _EVAL_821[14:13];
  assign _EVAL_1785 = _EVAL_47 ? 1'h1 : _EVAL_74;
  assign _EVAL_1125 = _EVAL_1713 ? 1'h1 : _EVAL_1785;
  assign _EVAL_1266 = _EVAL_772 ? 1'h1 : _EVAL_1125;
  assign _EVAL_997 = _EVAL_1014 ? 1'h1 : _EVAL_1266;
  assign _EVAL_843 = _EVAL_1627 ? _EVAL_997 : _EVAL_1785;
  assign _EVAL_1217 = _EVAL_428[3];
  assign _EVAL_2235 = _EVAL_1741[1];
  assign _EVAL_1693 = _EVAL_428[8:7];
  assign _EVAL_357 = _EVAL_1889 | _EVAL_87;
  assign _EVAL_1777 = _EVAL_357 & _EVAL_2009;
  assign _EVAL_1762 = _EVAL_1777[27];
  assign _EVAL_2035 = _EVAL_1762 & _EVAL_2084;
  assign _EVAL_1606 = _EVAL_2220 == 1'h0;
  assign _EVAL_1104 = _EVAL_551 | _EVAL_1606;
  assign _EVAL_787 = _EVAL_2035 & _EVAL_1104;
  assign _EVAL_2003 = _EVAL_1777[12];
  assign _EVAL_1085 = _EVAL_857[2];
  assign _EVAL_1871 = _EVAL_1741[4:3];
  assign _EVAL_1562 = _EVAL_279 == 1'h0;
  assign _EVAL_2124 = _EVAL_1562 & _EVAL_1408;
  assign _EVAL_331 = _EVAL_333 & _EVAL_2124;
  assign _EVAL_1300 = _EVAL_1555 | _EVAL_331;
  assign _EVAL_1356 = _EVAL_1300 == 1'h0;
  assign _EVAL_328 = _EVAL_1285 & _EVAL_1356;
  assign _EVAL_1235 = {_EVAL_1978,_EVAL_924};
  assign _EVAL_829 = _EVAL_1235 | 31'hf;
  assign _EVAL_1207 = _EVAL_829 + 31'h1;
  assign _EVAL_1357 = {_EVAL_1376,1'h0,1'h0,_EVAL_1421,_EVAL_381,_EVAL_1808,_EVAL_1241};
  assign _EVAL_1605 = {4'h2,_EVAL_1763,14'h400,_EVAL_1877,1'h0,2'h0,_EVAL_1494,_EVAL_1357};
  assign _EVAL_1674 = _EVAL_500 ? _EVAL_1605 : 32'h0;
  assign _EVAL_1072 = _EVAL_1674 | _EVAL_87;
  assign _EVAL_1107 = _EVAL_1072 & _EVAL_2009;
  assign _EVAL_1801 = _EVAL_1107[27];
  assign _EVAL_1793 = {_EVAL_109, 14'h0};
  assign _EVAL_1922 = _EVAL_1793[14];
  assign _EVAL_1012 = _EVAL_1793[13];
  assign _EVAL_2101 = _EVAL_1922 | _EVAL_1012;
  assign _EVAL_1294 = _EVAL_1793[12];
  assign _EVAL_2149 = _EVAL_2101 | _EVAL_1294;
  assign _EVAL_674 = _EVAL_1793[11];
  assign _EVAL_1305 = _EVAL_2149 | _EVAL_674;
  assign _EVAL_1279 = _EVAL_1793[3];
  assign _EVAL_408 = _EVAL_1305 | _EVAL_1279;
  assign _EVAL_866 = _EVAL_1793[7];
  assign _EVAL_1566 = _EVAL_408 | _EVAL_866;
  assign _EVAL_2228 = _EVAL_1793[9];
  assign _EVAL_1478 = _EVAL_1566 | _EVAL_2228;
  assign _EVAL_434 = _EVAL_1793[1];
  assign _EVAL_1088 = _EVAL_1478 | _EVAL_434;
  assign _EVAL_1957 = _EVAL_1793[5];
  assign _EVAL_1819 = _EVAL_1088 | _EVAL_1957;
  assign _EVAL_1457 = _EVAL_1793[8];
  assign _EVAL_199 = _EVAL_1819 | _EVAL_1457;
  assign _EVAL_1254 = _EVAL_1793[0];
  assign _EVAL_543 = _EVAL_199 | _EVAL_1254;
  assign _EVAL_2241 = _EVAL_1793[4];
  assign _EVAL_1053 = _EVAL_543 | _EVAL_2241;
  assign _EVAL_1020 = _EVAL_1053 | _EVAL_1997;
  assign _EVAL_1042 = _EVAL_497[14];
  assign _EVAL_1991 = _EVAL_1020 | _EVAL_1042;
  assign _EVAL_1610 = _EVAL_497[13];
  assign _EVAL_455 = _EVAL_1991 | _EVAL_1610;
  assign _EVAL_1838 = _EVAL_497[12];
  assign _EVAL_489 = _EVAL_455 | _EVAL_1838;
  assign _EVAL_1634 = _EVAL_497[11];
  assign _EVAL_1503 = _EVAL_489 | _EVAL_1634;
  assign _EVAL_1586 = _EVAL_497[3];
  assign _EVAL_1414 = _EVAL_1503 | _EVAL_1586;
  assign _EVAL_1259 = _EVAL_497[7];
  assign _EVAL_1940 = _EVAL_1414 | _EVAL_1259;
  assign _EVAL_1199 = _EVAL_497[9];
  assign _EVAL_2213 = _EVAL_1940 | _EVAL_1199;
  assign _EVAL_211 = _EVAL_497[1];
  assign _EVAL_1797 = _EVAL_2213 | _EVAL_211;
  assign _EVAL_985 = _EVAL_497[5];
  assign _EVAL_792 = _EVAL_1797 | _EVAL_985;
  assign _EVAL_862 = _EVAL_497[8];
  assign _EVAL_1111 = _EVAL_792 | _EVAL_862;
  assign _EVAL_1181 = _EVAL_430[1];
  assign _EVAL_370 = _EVAL_1763 == 1'h0;
  assign _EVAL_2240 = _EVAL_370 | _EVAL_2084;
  assign _EVAL_2006 = _EVAL_333 | _EVAL_331;
  assign _EVAL_1084 = _EVAL_1441 | _EVAL_993;
  assign _EVAL_292 = _EVAL_1121[27];
  assign _EVAL_2167 = _EVAL_292 & _EVAL_2084;
  assign _EVAL_1896 = _EVAL_2167 & _EVAL_396;
  assign _EVAL_184 = _EVAL_1121[12];
  assign _EVAL_644 = _EVAL_1307 == 1'h0;
  assign _EVAL_708 = _EVAL_2227[0];
  assign _EVAL_2095 = _EVAL_644 & _EVAL_708;
  assign _EVAL_467 = _EVAL_1593 & _EVAL_2095;
  assign _EVAL_1108 = _EVAL_2232 | _EVAL_467;
  assign _EVAL_354 = _EVAL_1108 == 1'h0;
  assign _EVAL_1751 = _EVAL_1396 & _EVAL_354;
  assign _EVAL_616 = _EVAL_1751 ? _EVAL_428 : {{2'd0}, _EVAL_842};
  assign _EVAL_219 = _EVAL_1627 ? _EVAL_616 : {{2'd0}, _EVAL_842};
  assign _EVAL_803 = _EVAL_1741[0];
  assign _EVAL_650 = _EVAL_2235 & _EVAL_803;
  assign _EVAL_513 = _EVAL_914 & 32'h30000000;
  assign _EVAL_209 = _EVAL_491[0];
  assign _EVAL_730 = {_EVAL_1952,_EVAL_209};
  assign _EVAL_424 = _EVAL_730 | 31'hf;
  assign _EVAL_2108 = _EVAL_424 + 31'h1;
  assign _EVAL_765 = ~ _EVAL_2108;
  assign _EVAL_1573 = _EVAL_424 & _EVAL_765;
  assign _EVAL_654 = _EVAL_912[0];
  assign _EVAL_1910 = _EVAL_2226[0];
  assign _EVAL_1886 = {_EVAL_2210,_EVAL_1910};
  assign _EVAL_1652 = _EVAL_1886 | 31'hf;
  assign _EVAL_1825 = _EVAL_1896 | _EVAL_370;
  assign _EVAL_1123 = _EVAL_1585 == 1'h0;
  assign _EVAL_1541 = _EVAL_1746 & _EVAL_1123;
  assign _EVAL_1292 = _EVAL_912[7];
  assign _EVAL_1355 = _EVAL_739 ? 12'h800 : 12'h808;
  assign _EVAL_1395 = _EVAL_2084 ? _EVAL_1355 : 12'h800;
  assign _EVAL_1200 = _EVAL_1401[0];
  assign _EVAL_336 = _EVAL_1200 & _EVAL_1334;
  assign _EVAL_691 = _EVAL_744[7:5];
  assign _EVAL_1028 = _EVAL_691 == 3'h0;
  assign _EVAL_846 = _EVAL_336 & _EVAL_1028;
  assign _EVAL_1771 = _EVAL_1401[31:7];
  assign _EVAL_573 = _EVAL_579[4:0];
  assign _EVAL_1130 = {_EVAL_573, 2'h0};
  assign _EVAL_777 = {_EVAL_1771,_EVAL_1130};
  assign _EVAL_2145 = _EVAL_1401[31:2];
  assign _EVAL_526 = {_EVAL_2145, 2'h0};
  assign _EVAL_1639 = _EVAL_846 ? _EVAL_777 : _EVAL_526;
  assign _EVAL_604 = _EVAL_939 ? {{20'd0}, _EVAL_1395} : _EVAL_1639;
  assign _EVAL_561 = _EVAL_720[63:32];
  assign _EVAL_452 = {_EVAL_561,_EVAL_428};
  assign _EVAL_1695 = _EVAL_452[63:6];
  assign _EVAL_440 = {{4'd0}, _EVAL_1};
  assign _EVAL_1049 = _EVAL_1249 + _EVAL_440;
  assign _EVAL_1914 = _EVAL_1049[6];
  assign _EVAL_1845 = _EVAL_751 + 58'h1;
  assign _EVAL_996 = _EVAL_428[6];
  assign _EVAL_250 = _EVAL_1741[7];
  assign _EVAL_507 = _EVAL_430[4:3];
  assign _EVAL_1954 = _EVAL_507[1];
  assign _EVAL_1543 = _EVAL_507 != 2'h0;
  assign _EVAL_659 = {_EVAL_1954,_EVAL_1543};
  assign _EVAL_1523 = _EVAL_513 == 32'h10000000;
  assign _EVAL_736 = _EVAL_1765 & _EVAL_1523;
  assign _EVAL_310 = _EVAL_18 == 12'hf13;
  assign _EVAL_855 = _EVAL_731 | _EVAL_310;
  assign _EVAL_174 = _EVAL_1871[1];
  assign _EVAL_1533 = _EVAL_1871 != 2'h0;
  assign _EVAL_2161 = {_EVAL_174,_EVAL_1533};
  assign _EVAL_878 = _EVAL_1358 ? _EVAL_899 : {{33'd0}, _EVAL_1575};
  assign _EVAL_201 = _EVAL_611 == 1'h0;
  assign _EVAL_1146 = _EVAL_1213 & _EVAL_201;
  assign _EVAL_490 = _EVAL_2084 == 1'h0;
  assign _EVAL_1518 = _EVAL_2232 == 1'h0;
  assign _EVAL_364 = _EVAL_1213 & _EVAL_1518;
  assign _EVAL_1720 = _EVAL_1143 != 2'h0;
  assign _EVAL_383 = {_EVAL_1515,_EVAL_1720};
  assign _EVAL_2110 = _EVAL_2151 == 1'h0;
  assign _EVAL_1010 = _EVAL_2110 & _EVAL_461;
  assign _EVAL_404 = 2'h3 == _EVAL_631;
  assign _EVAL_1251 = _EVAL_404 & _EVAL_2240;
  assign _EVAL_1960 = _EVAL_611 & _EVAL_1010;
  assign _EVAL_999 = _EVAL_1593 == 1'h0;
  assign _EVAL_2202 = _EVAL_1213 & _EVAL_999;
  assign _EVAL_858 = _EVAL_1547 != 2'h0;
  assign _EVAL_1136 = {_EVAL_1747,_EVAL_858};
  assign _EVAL_2027 = _EVAL_2181[0];
  assign _EVAL_1373 = {_EVAL_842,_EVAL_2027};
  assign _EVAL_1781 = _EVAL_181 == 1'h0;
  assign _EVAL_1210 = _EVAL_1213 & _EVAL_1781;
  assign _EVAL_2221 = _EVAL_1801 & _EVAL_2084;
  assign _EVAL_605 = _EVAL_203 == 1'h0;
  assign _EVAL_1981 = _EVAL_1769 | _EVAL_605;
  assign _EVAL_1489 = _EVAL_2221 & _EVAL_1981;
  assign _EVAL_909 = _EVAL_1107[12];
  assign _EVAL_636 = {_EVAL_2224,_EVAL_708};
  assign _EVAL_2023 = _EVAL_1777[11];
  assign _EVAL_2243 = _EVAL_681 == 1'h0;
  assign _EVAL_2028 = _EVAL_2243 & _EVAL_209;
  assign _EVAL_1648 = _EVAL_181 & _EVAL_2028;
  assign _EVAL_935 = _EVAL_1593 | _EVAL_1648;
  assign _EVAL_964 = _EVAL_935 == 1'h0;
  assign _EVAL_2144 = _EVAL_2070[63:32];
  assign _EVAL_1394 = _EVAL_105 == 1'h0;
  assign _EVAL_998 = _EVAL_736 & _EVAL_1394;
  assign _EVAL_2192 = _EVAL_998 & _EVAL_490;
  assign _EVAL_1921 = _EVAL_497[0];
  assign _EVAL_756 = _EVAL_1921 ? 4'h0 : 4'h4;
  assign _EVAL_1823 = _EVAL_862 ? 4'h8 : _EVAL_756;
  assign _EVAL_510 = _EVAL_985 ? 4'h5 : _EVAL_1823;
  assign _EVAL_2223 = _EVAL_211 ? 4'h1 : _EVAL_510;
  assign _EVAL_740 = _EVAL_1199 ? 4'h9 : _EVAL_2223;
  assign _EVAL_2123 = _EVAL_1259 ? 4'h7 : _EVAL_740;
  assign _EVAL_1603 = _EVAL_1586 ? 4'h3 : _EVAL_2123;
  assign _EVAL_2191 = _EVAL_1634 ? 4'hb : _EVAL_1603;
  assign _EVAL_1377 = _EVAL_1838 ? 4'hc : _EVAL_2191;
  assign _EVAL_1926 = _EVAL_1610 ? 4'hd : _EVAL_1377;
  assign _EVAL_358 = _EVAL_1042 ? 4'he : _EVAL_1926;
  assign _EVAL_1464 = _EVAL_1997 ? 4'hf : _EVAL_358;
  assign _EVAL_794 = _EVAL_2241 ? 4'h4 : _EVAL_1464;
  assign _EVAL_923 = _EVAL_1254 ? 4'h0 : _EVAL_794;
  assign _EVAL_466 = _EVAL_1457 ? 4'h8 : _EVAL_923;
  assign _EVAL_1853 = _EVAL_1957 ? 4'h5 : _EVAL_466;
  assign _EVAL_1980 = _EVAL_434 ? 4'h1 : _EVAL_1853;
  assign _EVAL_709 = _EVAL_2228 ? 4'h9 : _EVAL_1980;
  assign _EVAL_763 = _EVAL_866 ? 4'h7 : _EVAL_709;
  assign _EVAL_1083 = _EVAL_912[1];
  assign _EVAL_271 = _EVAL_1083 & _EVAL_654;
  assign _EVAL_1461 = _EVAL_237 & _EVAL_964;
  assign _EVAL_1302 = _EVAL_1461 ? _EVAL_428 : {{2'd0}, _EVAL_2224};
  assign _EVAL_1079 = _EVAL_2220 | _EVAL_203;
  assign _EVAL_1058 = _EVAL_1079 == 1'h0;
  assign _EVAL_1551 = _EVAL_2023 & _EVAL_1058;
  assign _EVAL_2024 = _EVAL_857[1];
  assign _EVAL_1416 = _EVAL_2024 & _EVAL_1831;
  assign _EVAL_253 = _EVAL_1306 == 1'h0;
  assign _EVAL_2081 = _EVAL_253 & _EVAL_1910;
  assign _EVAL_1027 = _EVAL_1168 & _EVAL_2081;
  assign _EVAL_1641 = _EVAL_611 | _EVAL_1027;
  assign _EVAL_577 = _EVAL_981[31:0];
  assign _EVAL_477 = {_EVAL_857,_EVAL_577};
  assign _EVAL_504 = {{4'd0}, _EVAL_49};
  assign _EVAL_2089 = _EVAL_2177 + _EVAL_504;
  assign _EVAL_1317 = _EVAL_2089[6];
  assign _EVAL_1264 = _EVAL_430[0];
  assign _EVAL_249 = _EVAL_1181 & _EVAL_1264;
  assign _EVAL_2043 = _EVAL_946 | 31'hf;
  assign _EVAL_1090 = _EVAL_2043 + 31'h1;
  assign _EVAL_883 = _EVAL_1426 == 1'h0;
  assign _EVAL_865 = _EVAL_1440[0];
  assign _EVAL_2078 = _EVAL_883 & _EVAL_865;
  assign _EVAL_1949 = _EVAL_1585 & _EVAL_2078;
  assign _EVAL_1863 = _EVAL_2114[39:32];
  assign _EVAL_773 = {_EVAL_1863,_EVAL_428};
  assign _EVAL_229 = _EVAL_1437 ? _EVAL_773 : {{33'd0}, _EVAL_2089};
  assign _EVAL_443 = _EVAL_1386 ? _EVAL_658 : _EVAL_229;
  assign _EVAL_1941 = _EVAL_497[4];
  assign _EVAL_2082 = _EVAL_1627 ? _EVAL_443 : {{33'd0}, _EVAL_2089};
  assign _EVAL_239 = _EVAL_148 == 1'h0;
  assign _EVAL_995 = {{5'd0}, _EVAL_239};
  assign _EVAL_277 = _EVAL_1260 ? _EVAL_428 : {{2'd0}, _EVAL_286};
  assign _EVAL_213 = _EVAL_1627 ? _EVAL_277 : {{2'd0}, _EVAL_286};
  assign _EVAL_1908 = _EVAL_857[7];
  assign _EVAL_505 = _EVAL_1168 | _EVAL_1949;
  assign _EVAL_1172 = _EVAL_505 == 1'h0;
  assign _EVAL_307 = _EVAL_1647 & _EVAL_1172;
  assign _EVAL_767 = _EVAL_1112 ? _EVAL_1466 : _EVAL_267;
  assign _EVAL_1583 = _EVAL_490 ? 2'h3 : _EVAL_317;
  assign _EVAL_2139 = _EVAL_939 ? _EVAL_1583 : 2'h3;
  assign _EVAL_302 = _EVAL_1937 ? _EVAL_2139 : _EVAL_317;
  assign _EVAL_1498 = _EVAL_898 ? _EVAL_767 : _EVAL_302;
  assign _EVAL_1194 = _EVAL_1498[0];
  assign _EVAL_1536 = _EVAL_1084 | _EVAL_1417;
  assign _EVAL_1721 = _EVAL_428[31:5];
  assign _EVAL_827 = _EVAL_772 ? _EVAL_428 : {{29'd0}, _EVAL_1458};
  assign _EVAL_718 = _EVAL_1014 ? {{5'd0}, _EVAL_1721} : _EVAL_827;
  assign _EVAL_2173 = _EVAL_1627 ? _EVAL_718 : {{29'd0}, _EVAL_1458};
  assign _EVAL_2183 = _EVAL_1999 ? 2'h2 : 2'h1;
  assign _EVAL_960 = _EVAL_679 ? 2'h3 : _EVAL_2183;
  assign _EVAL_1410 = _EVAL_912[2];
  assign _EVAL_959 = _EVAL_102 >= 12'hb00;
  assign _EVAL_863 = _EVAL_102 < 12'hb20;
  assign _EVAL_1216 = _EVAL_959 & _EVAL_863;
  assign _EVAL_1473 = _EVAL_102 >= 12'hb80;
  assign _EVAL_1030 = _EVAL_102 < 12'hba0;
  assign _EVAL_1233 = _EVAL_1473 & _EVAL_1030;
  assign _EVAL_390 = _EVAL_1216 | _EVAL_1233;
  assign _EVAL_195 = _EVAL_1627 & _EVAL_390;
  assign _EVAL_522 = _EVAL_102[5:0];
  assign _EVAL_724 = 64'h1 << _EVAL_522;
  assign _EVAL_2001 = _EVAL_195 ? _EVAL_724 : 64'h0;
  assign _EVAL_282 = _EVAL_428 & 32'h888;
  assign _EVAL_1451 = _EVAL_18 < 12'hca0;
  assign _EVAL_2130 = _EVAL_405 & _EVAL_1451;
  assign _EVAL_427 = ~ _EVAL_1759;
  assign _EVAL_2132 = _EVAL_428 & 32'h8000000f;
  assign _EVAL_2140 = _EVAL_428[1:0];
  assign _EVAL_1229 = _EVAL_2140[0];
  assign _EVAL_1147 = ~ _EVAL_1207;
  assign _EVAL_275 = {{1'd0}, _EVAL_926};
  assign _EVAL_864 = _EVAL_787 | _EVAL_1773;
  assign _EVAL_1170 = _EVAL_1551 & _EVAL_864;
  assign _EVAL_678 = _EVAL_428[12];
  assign _EVAL_570 = _EVAL_821[7];
  assign _EVAL_920 = _EVAL_720[31:0];
  assign _EVAL_225 = {_EVAL_428,_EVAL_920};
  assign _EVAL_1723 = _EVAL_225[63:6];
  assign _EVAL_1976 = _EVAL_2106 + 34'h1;
  assign _EVAL_1383 = _EVAL_18[4:0];
  assign _EVAL_713 = _EVAL_1504 >> _EVAL_1383;
  assign _EVAL_1856 = _EVAL_713[0];
  assign _EVAL_665 = _EVAL_2006 == 1'h0;
  assign _EVAL_1165 = _EVAL_484 & _EVAL_665;
  assign _EVAL_1255 = _EVAL_428 & 32'h10007;
  assign _EVAL_722 = _EVAL_18 == 12'hffc;
  assign _EVAL_2219 = _EVAL_855 | _EVAL_722;
  assign _EVAL_1131 = _EVAL_1121[11];
  assign _EVAL_353 = _EVAL_18 >= 12'hc00;
  assign _EVAL_1276 = _EVAL_18 < 12'hc20;
  assign _EVAL_1332 = _EVAL_353 & _EVAL_1276;
  assign _EVAL_1552 = _EVAL_1652 + 31'h1;
  assign _EVAL_2113 = ~ _EVAL_1552;
  assign _EVAL_1852 = _EVAL_1652 & _EVAL_2113;
  assign _EVAL_816 = _EVAL_18[9:8];
  assign _EVAL_991 = _EVAL_317 < _EVAL_816;
  assign _EVAL_1102 = _EVAL_1 > 2'h1;
  assign _EVAL_1529 = _EVAL_2070[31:0];
  assign _EVAL_619 = {_EVAL_428,_EVAL_1529};
  assign _EVAL_699 = {_EVAL_2144,_EVAL_428};
  assign _EVAL_717 = _EVAL_1419 + _EVAL_995;
  assign _EVAL_904 = _EVAL_531 ? _EVAL_699 : {{57'd0}, _EVAL_717};
  assign _EVAL_886 = _EVAL_1657 ? _EVAL_619 : _EVAL_904;
  assign _EVAL_1328 = _EVAL_1627 ? _EVAL_886 : {{57'd0}, _EVAL_717};
  assign _EVAL_1827 = _EVAL_2219 == 1'h0;
  assign _EVAL_1275 = _EVAL_991 | _EVAL_1827;
  assign _EVAL_465 = _EVAL_658[39:6];
  assign _EVAL_533 = _EVAL_773[39:6];
  assign _EVAL_851 = _EVAL_1536 & _EVAL_490;
  assign _EVAL_1008 = _EVAL_317 > 2'h1;
  assign _EVAL_2142 = _EVAL_1008 | _EVAL_1856;
  assign _EVAL_653 = _EVAL_2142 == 1'h0;
  assign _EVAL_669 = {_EVAL_18, 20'h0};
  assign _EVAL_1932 = _EVAL_669 & 32'ha0400000;
  assign _EVAL_349 = _EVAL_1932 == 32'h20000000;
  assign _EVAL_1343 = _EVAL_584 | _EVAL_144;
  assign _EVAL_779 = _EVAL_47 ? _EVAL_1343 : _EVAL_584;
  assign _EVAL_1685 = _EVAL_1713 ? _EVAL_428 : {{27'd0}, _EVAL_779};
  assign _EVAL_1033 = _EVAL_1014 ? _EVAL_428 : _EVAL_1685;
  assign _EVAL_2195 = _EVAL_1627 ? _EVAL_1033 : {{27'd0}, _EVAL_779};
  assign _EVAL_1924 = _EVAL_1279 ? 4'h3 : _EVAL_763;
  assign _EVAL_441 = _EVAL_674 ? 4'hb : _EVAL_1924;
  assign _EVAL_2129 = _EVAL_1294 ? 4'hc : _EVAL_441;
  assign _EVAL_1067 = _EVAL_1012 ? 4'hd : _EVAL_2129;
  assign _EVAL_2222 = _EVAL_821[17];
  assign _EVAL_1443 = _EVAL_1165 ? _EVAL_428 : {{2'd0}, _EVAL_1942};
  assign _EVAL_341 = _EVAL_829 & _EVAL_1147;
  assign _EVAL_1782 = {_EVAL_341,2'h3};
  assign _EVAL_828 = _EVAL_821[3];
  assign _EVAL_2077 = _EVAL_619[63:6];
  assign _EVAL_2029 = _EVAL_1332 | _EVAL_2130;
  assign _EVAL_1145 = _EVAL_2029 & _EVAL_653;
  assign _EVAL_1025 = _EVAL_1275 | _EVAL_1145;
  assign _EVAL_1044 = {_EVAL_286,_EVAL_865};
  assign _EVAL_1813 = _EVAL_1044 | 31'hf;
  assign _EVAL_458 = _EVAL_1813 + 31'h1;
  assign _EVAL_506 = _EVAL_1038 | 32'h1;
  assign _EVAL_741 = ~ _EVAL_506;
  assign _EVAL_1312 = {_EVAL_1852,2'h3};
  assign _EVAL_1093 = _EVAL_430[2];
  assign _EVAL_1655 = _EVAL_1111 | _EVAL_1921;
  assign _EVAL_1126 = _EVAL_328 ? _EVAL_428 : {{2'd0}, _EVAL_1978};
  assign _EVAL_928 = _EVAL_428[15];
  assign _EVAL_877 = _EVAL_914 & 32'ha0200000;
  assign _EVAL_808 = _EVAL_877 == 32'h20000000;
  assign _EVAL_2160 = _EVAL_1765 & _EVAL_808;
  assign _EVAL_608 = _EVAL_307 ? _EVAL_428 : {{2'd0}, _EVAL_2210};
  assign _EVAL_2121 = _EVAL_1 >= 2'h1;
  assign _EVAL_303 = ~ _EVAL_458;
  assign _EVAL_320 = _EVAL_1813 & _EVAL_303;
  assign _EVAL_559 = _EVAL_1641 == 1'h0;
  assign _EVAL_1459 = _EVAL_1373 | 31'hf;
  assign _EVAL_1876 = _EVAL_1459 + 31'h1;
  assign _EVAL_1649 = ~ _EVAL_1876;
  assign _EVAL_1691 = _EVAL_1459 & _EVAL_1649;
  assign _EVAL_2015 = _EVAL_46 & _EVAL_134;
  assign _EVAL_1791 = _EVAL_826 ? _EVAL_428 : {{30'd0}, _EVAL_631};
  assign _EVAL_2068 = _EVAL_1627 ? _EVAL_1302 : {{2'd0}, _EVAL_2224};
  assign _EVAL_2165 = ~ _EVAL_1090;
  assign _EVAL_2185 = _EVAL_2043 & _EVAL_2165;
  assign _EVAL_2169 = {_EVAL_2185,2'h3};
  assign _EVAL_535 = _EVAL_181 | _EVAL_1960;
  assign _EVAL_1353 = _EVAL_535 == 1'h0;
  assign _EVAL_1661 = _EVAL_1[0];
  assign _EVAL_639 = _EVAL_428 & 32'h3ffff03;
  assign _EVAL_1772 = _EVAL_349 & _EVAL_1900;
  assign _EVAL_1953 = _EVAL_1772 & _EVAL_490;
  assign _EVAL_675 = _EVAL_1559 ? _EVAL_452 : {{57'd0}, _EVAL_1049};
  assign _EVAL_330 = _EVAL_1872 ? _EVAL_225 : _EVAL_675;
  assign _EVAL_813 = _EVAL_1131 & _EVAL_1389;
  assign _EVAL_1177 = _EVAL_813 & _EVAL_1825;
  assign _EVAL_2091 = _EVAL_1627 ? _EVAL_608 : {{2'd0}, _EVAL_2210};
  assign _EVAL_2067 = _EVAL_1381 & _EVAL_490;
  assign _EVAL_790 = _EVAL_636 | 31'hf;
  assign _EVAL_743 = _EVAL_790 + 31'h1;
  assign _EVAL_716 = ~ _EVAL_743;
  assign _EVAL_871 = _EVAL_790 & _EVAL_716;
  assign _EVAL_1403 = _EVAL_699[63:6];
  assign _EVAL_565 = _EVAL_717[6];
  assign _EVAL_1947 = _EVAL_1212 + 58'h1;
  assign _EVAL_2147 = _EVAL_18 & 12'ha00;
  assign _EVAL_471 = _EVAL_1661 | _EVAL_1937;
  assign _EVAL_476 = _EVAL_1532 & 32'hfffefff8;
  assign _EVAL_516 = _EVAL_1255 | _EVAL_476;
  assign _EVAL_1963 = _EVAL_780 & _EVAL_1353;
  assign _EVAL_1717 = _EVAL_1963 ? _EVAL_428 : {{2'd0}, _EVAL_1952};
  assign _EVAL_326 = _EVAL_1627 ? _EVAL_1717 : {{2'd0}, _EVAL_1952};
  assign _EVAL_2153 = _EVAL_477[39:6];
  assign _EVAL_2205 = _EVAL_1627 ? _EVAL_1791 : {{30'd0}, _EVAL_631};
  assign _EVAL_348 = _EVAL_1922 ? 4'he : _EVAL_1067;
  assign _EVAL_809 = {{28'd0}, _EVAL_348};
  assign _EVAL_1158 = _EVAL_1289 != 32'h0;
  assign _EVAL_177 = _EVAL_1158 | _EVAL_109;
  assign _EVAL_728 = {_EVAL_871,2'h3};
  assign _EVAL_1843 = _EVAL_177 | _EVAL_1937;
  assign _EVAL_1642 = _EVAL_135 == 2'h3;
  assign _EVAL_265 = _EVAL_1627 ? _EVAL_1126 : {{2'd0}, _EVAL_1978};
  assign _EVAL_1928 = _EVAL_1655 | _EVAL_1941;
  assign _EVAL_624 = _EVAL_1928 & _EVAL_1394;
  assign _EVAL_2133 = {_EVAL_1573,2'h3};
  assign _EVAL_869 = _EVAL_1627 ? _EVAL_330 : {{57'd0}, _EVAL_1049};
  assign _EVAL_1927 = {_EVAL_1691,2'h3};
  assign _EVAL_186 = _EVAL_1374 ? _EVAL_477 : _EVAL_878;
  assign _EVAL_860 = _EVAL_1627 ? _EVAL_186 : {{33'd0}, _EVAL_1575};
  assign _EVAL_1993 = _EVAL_939 ? {{1'd0}, _EVAL_926} : _EVAL_275;
  assign _EVAL_1836 = _EVAL_22 == 2'h3;
  assign _EVAL_1788 = _EVAL_1937 ? _EVAL_1993 : {{1'd0}, _EVAL_926};
  assign _EVAL_2170 = _EVAL_1112 ? _EVAL_1032 : _EVAL_1315;
  assign _EVAL_906 = _EVAL_1627 ? _EVAL_1443 : {{2'd0}, _EVAL_1942};
  assign _EVAL_1159 = _EVAL_2084 | _EVAL_92;
  assign _EVAL_1371 = _EVAL_1159 == 1'h0;
  assign _EVAL_574 = _EVAL_539 & _EVAL_559;
  assign _EVAL_1624 = _EVAL_624 | _EVAL_1073;
  assign _EVAL_2086 = {_EVAL_320,2'h3};
  assign _EVAL_204 = _EVAL_1025 | _EVAL_851;
  assign _EVAL_2065 = _EVAL_574 ? _EVAL_428 : {{2'd0}, _EVAL_182};
  assign _EVAL_363 = _EVAL_1627 ? _EVAL_2065 : {{2'd0}, _EVAL_182};
  assign _EVAL_651 = _EVAL_18[11:10];
  assign _EVAL_135 = _EVAL_1545;
  assign _EVAL_148 = _EVAL_645 | _EVAL_92;
  assign _EVAL_15 = _EVAL_1376;
  assign _EVAL_133 = _EVAL_297;
  assign _EVAL_54 = _EVAL_1942;
  assign _EVAL_92 = _EVAL_2159;
  assign _EVAL_40 = _EVAL_898 ? _EVAL_2170 : _EVAL_604;
  assign _EVAL_127 = _EVAL_1078;
  assign _EVAL_24 = _EVAL_1138;
  assign _EVAL_75 = _EVAL_2047;
  assign _EVAL_145 = _EVAL_1927[31:0];
  assign _EVAL_65 = _EVAL_692;
  assign _EVAL_147 = _EVAL_333;
  assign _EVAL_122 = _EVAL_2230;
  assign _EVAL_36 = _EVAL_1982;
  assign _EVAL_44 = 32'h80000000 + _EVAL_809;
  assign _EVAL_67 = _EVAL_1929;
  assign _EVAL_27 = _EVAL_2074;
  assign _EVAL_11 = _EVAL_1986;
  assign _EVAL_12 = _EVAL_1700;
  assign _EVAL_112 = _EVAL_2190;
  assign _EVAL_19 = _EVAL_1869;
  assign _EVAL_56 = _EVAL_1555;
  assign _EVAL_99 = _EVAL_1458;
  assign _EVAL_21 = _EVAL_760;
  assign _EVAL_76 = _EVAL_317;
  assign _EVAL_151 = _EVAL_1011;
  assign _EVAL_17 = _EVAL_941;
  assign _EVAL_156 = _EVAL_2210;
  assign _EVAL_104 = _EVAL_710;
  assign _EVAL_66 = _EVAL_182;
  assign _EVAL_68 = _EVAL_1666;
  assign _EVAL_120 = 2'h1;
  assign _EVAL_22 = _EVAL_252;
  assign _EVAL_42 = _EVAL_651 == 2'h3;
  assign _EVAL_57 = _EVAL_1241;
  assign _EVAL_136 = _EVAL_2169[31:0];
  assign _EVAL_159 = _EVAL_1479;
  assign _EVAL_73 = _EVAL_267;
  assign _EVAL_37 = _EVAL_842;
  assign _EVAL_7 = _EVAL_1062;
  assign _EVAL_38 = _EVAL_207;
  assign _EVAL_8 = _EVAL_463;
  assign _EVAL_2 = _EVAL_1782[31:0];
  assign _EVAL_26 = _EVAL_2220;
  assign _EVAL_31 = _EVAL_1425;
  assign _EVAL_14 = _EVAL_1048;
  assign _EVAL_132 = _EVAL_1223;
  assign _EVAL_157 = _EVAL_611;
  assign _EVAL_62 = _EVAL_436;
  assign _EVAL_142 = _EVAL_2224;
  assign _EVAL_10 = _EVAL_1193;
  assign _EVAL_28 = _EVAL_1770;
  assign _EVAL_100 = _EVAL_1440;
  assign _EVAL_161 = _EVAL_1743;
  assign _EVAL_82 = _EVAL_2227;
  assign _EVAL_9 = _EVAL_1593;
  assign _EVAL_98 = _EVAL_334;
  assign _EVAL_118 = 32'h40901125;
  assign _EVAL_108 = _EVAL_2063;
  assign _EVAL_20 = _EVAL_1877;
  assign _EVAL_166 = _EVAL_2086[31:0];
  assign _EVAL_158 = _EVAL_1312[31:0];
  assign _EVAL_103 = _EVAL_2131;
  assign _EVAL_3 = _EVAL_178;
  assign _EVAL_116 = _EVAL_346;
  assign _EVAL_83 = _EVAL_2001[31:0];
  assign _EVAL_4 = _EVAL_579[7:0];
  assign _EVAL_34 = _EVAL_1808;
  assign _EVAL_71 = _EVAL_69;
  assign _EVAL_96 = _EVAL_1141[31:0];
  assign _EVAL_88 = {_EVAL_2084,_EVAL_317};
  assign _EVAL_140 = _EVAL_1520 | _EVAL_25;
  assign _EVAL_46 = _EVAL_2147 == 12'h0;
  assign _EVAL_114 = _EVAL_1022;
  assign _EVAL_131 = _EVAL_1421;
  assign _EVAL_160 = _EVAL_1725;
  assign _EVAL_105 = _EVAL_762 & _EVAL_490;
  assign _EVAL_79 = _EVAL_1366;
  assign _EVAL_106 = _EVAL_1620;
  assign _EVAL_134 = _EVAL_22 == 2'h0;
  assign _EVAL_154 = _EVAL_2180;
  assign _EVAL_52 = _EVAL_1178;
  assign _EVAL_90 = _EVAL_204 | _EVAL_2015;
  assign _EVAL_91 = _EVAL_944;
  assign _EVAL_167 = _EVAL_900;
  assign _EVAL_130 = _EVAL_1162;
  assign _EVAL_70 = _EVAL_1624 & _EVAL_1371;
  assign _EVAL_97 = _EVAL_2232;
  assign _EVAL_63 = _EVAL_726;
  assign _EVAL_138 = 2'h0;
  assign _EVAL_84 = _EVAL_351[31:0];
  assign _EVAL_59 = _EVAL_361;
  assign _EVAL_30 = {_EVAL_2084,_EVAL_317};
  assign _EVAL_61 = _EVAL_2158;
  assign _EVAL_81 = _EVAL_2238;
  assign _EVAL_80 = _EVAL_537;
  assign _EVAL_13 = _EVAL_381;
  assign _EVAL_93 = _EVAL_2002;
  assign _EVAL_45 = _EVAL_715;
  assign _EVAL_33 = _EVAL_1168;
  assign _EVAL_128 = _EVAL_203;
  assign _EVAL_113 = _EVAL_728[31:0];
  assign _EVAL_107 = _EVAL_1556;
  assign _EVAL_137 = _EVAL_1792;
  assign _EVAL_72 = _EVAL_1102 | _EVAL_163;
  assign _EVAL_153 = _EVAL_992;
  assign _EVAL_85 = _EVAL_991 | _EVAL_1953;
  assign _EVAL_89 = _EVAL_1849 | _EVAL_898;
  assign _EVAL_95 = _EVAL_1354;
  assign _EVAL_124 = _EVAL_1381;
  assign _EVAL_48 = _EVAL_795;
  assign _EVAL_126 = _EVAL_2133[31:0];
  assign _EVAL_39 = _EVAL_2084;
  assign _EVAL_152 = _EVAL_1261;
  assign _EVAL_55 = _EVAL_2226;
  assign _EVAL_69 = _EVAL_1836 | _EVAL_1642;
  assign _EVAL_94 = _EVAL_1567;
  assign _EVAL_141 = _EVAL_1956;
  assign _EVAL_43 = _EVAL_491;
  assign _EVAL_25 = _EVAL_1849 | _EVAL_155;
  assign _EVAL_125 = _EVAL_1499;
  assign _EVAL_29 = _EVAL_1494;
  assign _EVAL_32 = _EVAL_181;
  assign _EVAL_139 = _EVAL_990;
  assign _EVAL_164 = _EVAL_958;
  assign _EVAL_119 = _EVAL_523;
  assign _EVAL_121 = _EVAL_2181;
  assign _EVAL_5 = _EVAL_1385;
  assign _EVAL_115 = _EVAL_579[7:0];
  assign _EVAL_163 = _EVAL_2121 & _EVAL_1937;
  assign _EVAL_35 = _EVAL_194;
  assign _EVAL_58 = _EVAL_1733;
  assign _EVAL_0 = _EVAL_1978;
  assign _EVAL_143 = _EVAL_926;
  assign _EVAL_162 = _EVAL_286;
  assign _EVAL_129 = _EVAL_1608;
  assign _EVAL_111 = _EVAL_442;
  assign _EVAL_16 = _EVAL_1585;
  assign _EVAL_51 = _EVAL_1532;
  assign _EVAL_64 = _EVAL_1063;
  assign _EVAL_149 = _EVAL_1167;
  assign _EVAL_150 = _EVAL_1895;
  assign _EVAL_101 = _EVAL_1952;
  assign _EVAL_123 = _EVAL_2070[31:0];
  assign _EVAL_110 = _EVAL_1563;
  assign _EVAL_60 = _EVAL_2152;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _EVAL_171 = _RAND_0[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_178 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_181 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_182 = _RAND_3[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_194 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_203 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_207 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_252 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_267 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_286 = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_297 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_305 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_317 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_333 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_334 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_346 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_361 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_381 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_422 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_436 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_442 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_463 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_491 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_523 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_528 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_537 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_551 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_584 = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_594 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_597 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_609 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_611 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_631 = _RAND_32[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_645 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_692 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_710 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_715 = _RAND_36[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_726 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_745 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _EVAL_751 = _RAND_39[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_759 = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_760 = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_762 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_795 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_842 = _RAND_44[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_900 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_926 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_941 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_944 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_958 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_978 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_990 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_992 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1011 = _RAND_53[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1022 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1048 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1062 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1063 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1073 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1078 = _RAND_59[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1138 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1162 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1167 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1168 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1178 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1193 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  _EVAL_1212 = _RAND_66[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1223 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1239 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1241 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1249 = _RAND_70[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1261 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1282 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1344 = _RAND_73[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1354 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1366 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1376 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1381 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1385 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1392 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1419 = _RAND_80[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1421 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1424 = _RAND_82[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1425 = _RAND_83[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1440 = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1458 = _RAND_85[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1466 = _RAND_86[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1479 = _RAND_87[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1494 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1499 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1532 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1545 = _RAND_91[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1555 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1556 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1563 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1567 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1585 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1589 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1593 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1608 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1620 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1632 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1666 = _RAND_102[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1688 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1700 = _RAND_104[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1725 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1733 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_1743 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1763 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_1769 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1770 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1792 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1808 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1869 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _EVAL_1877 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_1895 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1899 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1929 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1942 = _RAND_118[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_1952 = _RAND_119[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1956 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1978 = _RAND_121[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1982 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1986 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_2002 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_2033 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_2047 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_2063 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_2074 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_2084 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_2090 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {2{`RANDOM}};
  _EVAL_2106 = _RAND_131[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_2131 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_2152 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_2158 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_2159 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_2177 = _RAND_136[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_2180 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_2181 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_2190 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_2210 = _RAND_140[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_2220 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _EVAL_2224 = _RAND_142[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2226 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _EVAL_2227 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _EVAL_2230 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2232 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _EVAL_2238 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_53) begin
    if (_EVAL_1627) begin
      if (_EVAL_1374) begin
        _EVAL_171 <= _EVAL_2153;
      end else begin
        if (_EVAL_1358) begin
          _EVAL_171 <= _EVAL_2154;
        end else begin
          if (_EVAL_1156) begin
            _EVAL_171 <= _EVAL_1800;
          end
        end
      end
    end else begin
      if (_EVAL_1156) begin
        _EVAL_171 <= _EVAL_1800;
      end
    end
    if (_EVAL_146) begin
      _EVAL_178 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_270) begin
          if (_EVAL_283) begin
            _EVAL_178 <= _EVAL_830;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_181 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1210) begin
          _EVAL_181 <= _EVAL_250;
        end
      end
    end
    _EVAL_182 <= _EVAL_363[29:0];
    if (_EVAL_1627) begin
      if (_EVAL_1151) begin
        if (_EVAL_283) begin
          _EVAL_194 <= _EVAL_1693;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_203 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_309) begin
          if (_EVAL_283) begin
            _EVAL_203 <= _EVAL_1177;
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_749) begin
        _EVAL_207 <= _EVAL_249;
      end
    end
    if (_EVAL_146) begin
      _EVAL_252 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1310) begin
          _EVAL_252 <= _EVAL_602;
        end else begin
          if (_EVAL_843) begin
            _EVAL_252 <= 2'h3;
          end
        end
      end else begin
        if (_EVAL_843) begin
          _EVAL_252 <= 2'h3;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_267 <= 2'h3;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1310) begin
          if (_EVAL_753) begin
            _EVAL_267 <= 2'h3;
          end else begin
            _EVAL_267 <= 2'h0;
          end
        end else begin
          if (_EVAL_898) begin
            if (_EVAL_1112) begin
              if (_EVAL_1937) begin
                if (!(_EVAL_939)) begin
                  if (_EVAL_386) begin
                    _EVAL_267 <= 2'h3;
                  end else begin
                    _EVAL_267 <= 2'h0;
                  end
                end
              end
            end else begin
              _EVAL_267 <= 2'h0;
            end
          end else begin
            if (_EVAL_1937) begin
              if (!(_EVAL_939)) begin
                if (_EVAL_386) begin
                  _EVAL_267 <= 2'h3;
                end else begin
                  _EVAL_267 <= 2'h0;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_898) begin
          if (_EVAL_1112) begin
            if (_EVAL_1937) begin
              if (!(_EVAL_939)) begin
                if (_EVAL_386) begin
                  _EVAL_267 <= 2'h3;
                end else begin
                  _EVAL_267 <= 2'h0;
                end
              end
            end
          end else begin
            _EVAL_267 <= 2'h0;
          end
        end else begin
          if (_EVAL_1937) begin
            if (!(_EVAL_939)) begin
              if (_EVAL_386) begin
                _EVAL_267 <= 2'h3;
              end else begin
                _EVAL_267 <= 2'h0;
              end
            end
          end
        end
      end
    end
    _EVAL_286 <= _EVAL_213[29:0];
    if (_EVAL_146) begin
      _EVAL_297 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1151) begin
          if (_EVAL_283) begin
            _EVAL_297 <= _EVAL_830;
          end
        end
      end
    end
    _EVAL_305 <= _EVAL_860[5:0];
    if (_EVAL_146) begin
      _EVAL_317 <= 2'h3;
    end else begin
      if (_EVAL_1194) begin
        _EVAL_317 <= 2'h3;
      end else begin
        _EVAL_317 <= 2'h0;
      end
    end
    if (_EVAL_146) begin
      _EVAL_333 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_749) begin
          _EVAL_333 <= _EVAL_2163;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2202) begin
        _EVAL_334 <= _EVAL_654;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1151) begin
        if (_EVAL_283) begin
          _EVAL_346 <= _EVAL_1217;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_270) begin
        if (_EVAL_283) begin
          _EVAL_361 <= _EVAL_1217;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_381 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1251) begin
          if (_EVAL_283) begin
            _EVAL_381 <= _EVAL_1590;
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2208) begin
        _EVAL_422 <= _EVAL_2132;
      end else begin
        if (_EVAL_1937) begin
          if (!(_EVAL_939)) begin
            if (_EVAL_1902) begin
              _EVAL_422 <= {{28'd0}, _EVAL_530};
            end else begin
              if (_EVAL_739) begin
                _EVAL_422 <= 32'h3;
              end else begin
                _EVAL_422 <= _EVAL_78;
              end
            end
          end
        end
      end
    end else begin
      if (_EVAL_1937) begin
        if (!(_EVAL_939)) begin
          if (_EVAL_1902) begin
            _EVAL_422 <= {{28'd0}, _EVAL_530};
          end else begin
            if (_EVAL_739) begin
              _EVAL_422 <= 32'h3;
            end else begin
              _EVAL_422 <= _EVAL_78;
            end
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_436 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1151) begin
          if (_EVAL_283) begin
            _EVAL_436 <= _EVAL_707;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_442 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1310) begin
          _EVAL_442 <= _EVAL_828;
        end else begin
          if (_EVAL_898) begin
            if (_EVAL_1112) begin
              if (_EVAL_1937) begin
                if (!(_EVAL_939)) begin
                  _EVAL_442 <= 1'h0;
                end
              end
            end else begin
              _EVAL_442 <= _EVAL_1162;
            end
          end else begin
            if (_EVAL_1937) begin
              if (!(_EVAL_939)) begin
                _EVAL_442 <= 1'h0;
              end
            end
          end
        end
      end else begin
        if (_EVAL_898) begin
          if (_EVAL_1112) begin
            if (_EVAL_1937) begin
              if (!(_EVAL_939)) begin
                _EVAL_442 <= 1'h0;
              end
            end
          end else begin
            _EVAL_442 <= _EVAL_1162;
          end
        end else begin
          if (_EVAL_1937) begin
            if (!(_EVAL_939)) begin
              _EVAL_442 <= 1'h0;
            end
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_463 <= 8'h0;
    end
    if (_EVAL_146) begin
      _EVAL_491 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1210) begin
          _EVAL_491 <= _EVAL_2161;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2120) begin
        _EVAL_523 <= _EVAL_1085;
      end
    end
    if (_EVAL_146) begin
      _EVAL_528 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_537 <= 32'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_666) begin
          _EVAL_537 <= _EVAL_639;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_551 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_270) begin
          if (_EVAL_283) begin
            _EVAL_551 <= _EVAL_670;
          end
        end
      end
    end
    _EVAL_584 <= _EVAL_2195[4:0];
    if (_EVAL_146) begin
      _EVAL_594 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1833) begin
          _EVAL_594 <= _EVAL_678;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_597 <= 3'h0;
    end else begin
      if (_EVAL_1937) begin
        if (_EVAL_939) begin
          if (_EVAL_490) begin
            if (_EVAL_1073) begin
              _EVAL_597 <= 3'h4;
            end else begin
              _EVAL_597 <= {{1'd0}, _EVAL_960};
            end
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_609 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_611 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1146) begin
          _EVAL_611 <= _EVAL_2163;
        end
      end
    end
    _EVAL_631 <= _EVAL_2205[1:0];
    if (_EVAL_146) begin
      _EVAL_692 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_309) begin
          if (_EVAL_283) begin
            if (_EVAL_1896) begin
              _EVAL_692 <= _EVAL_184;
            end else begin
              _EVAL_692 <= 1'h0;
            end
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1146) begin
        _EVAL_710 <= _EVAL_1093;
      end
    end
    if (_EVAL_146) begin
      _EVAL_715 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1644) begin
          _EVAL_715 <= _EVAL_2161;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_726 <= 1'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_2017) begin
        _EVAL_745 <= _EVAL_428;
      end else begin
        if (_EVAL_1937) begin
          if (!(_EVAL_939)) begin
            _EVAL_745 <= _EVAL_117;
          end
        end
      end
    end else begin
      if (_EVAL_1937) begin
        if (!(_EVAL_939)) begin
          _EVAL_745 <= _EVAL_117;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_751 <= 58'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1872) begin
          _EVAL_751 <= _EVAL_1723;
        end else begin
          if (_EVAL_1559) begin
            _EVAL_751 <= _EVAL_1695;
          end else begin
            if (_EVAL_1914) begin
              _EVAL_751 <= _EVAL_1845;
            end
          end
        end
      end else begin
        if (_EVAL_1914) begin
          _EVAL_751 <= _EVAL_1845;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_759 <= 2'h0;
    end
    if (_EVAL_2067) begin
      _EVAL_760 <= _EVAL_267;
    end else begin
      _EVAL_760 <= _EVAL_317;
    end
    if (_EVAL_146) begin
      _EVAL_762 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1833) begin
          _EVAL_762 <= _EVAL_1590;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_795 <= 1'h0;
    end
    _EVAL_842 <= _EVAL_219[29:0];
    if (_EVAL_1627) begin
      if (_EVAL_309) begin
        if (_EVAL_1722) begin
          _EVAL_900 <= _EVAL_428;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_926 <= 1'h0;
    end else begin
      _EVAL_926 <= _EVAL_1788[0];
    end
    if (_EVAL_1627) begin
      if (_EVAL_1210) begin
        _EVAL_941 <= _EVAL_243;
      end
    end
    if (_EVAL_146) begin
      _EVAL_944 <= 1'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_1146) begin
        _EVAL_958 <= _EVAL_1264;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1291) begin
        _EVAL_978 <= _EVAL_741;
      end else begin
        if (_EVAL_1937) begin
          if (!(_EVAL_939)) begin
            _EVAL_978 <= _EVAL_427;
          end
        end
      end
    end else begin
      if (_EVAL_1937) begin
        if (!(_EVAL_939)) begin
          _EVAL_978 <= _EVAL_427;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_990 <= 1'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_364) begin
        _EVAL_992 <= _EVAL_1085;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1011 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_749) begin
          _EVAL_1011 <= _EVAL_659;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_364) begin
        _EVAL_1022 <= _EVAL_1416;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1048 <= 32'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1617) begin
          _EVAL_1048 <= _EVAL_639;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1146) begin
        _EVAL_1062 <= _EVAL_249;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_270) begin
        if (_EVAL_1722) begin
          _EVAL_1063 <= _EVAL_428;
        end
      end
    end
    if (_EVAL_1394) begin
      _EVAL_1073 <= 1'h0;
    end else begin
      if (_EVAL_471) begin
        _EVAL_1073 <= 1'h1;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1078 <= 27'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_1151) begin
        if (_EVAL_283) begin
          _EVAL_1138 <= _EVAL_996;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1162 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1310) begin
          _EVAL_1162 <= _EVAL_570;
        end else begin
          if (_EVAL_898) begin
            if (_EVAL_1112) begin
              if (_EVAL_1937) begin
                if (!(_EVAL_939)) begin
                  _EVAL_1162 <= _EVAL_442;
                end
              end
            end else begin
              _EVAL_1162 <= 1'h1;
            end
          end else begin
            if (_EVAL_1937) begin
              if (!(_EVAL_939)) begin
                _EVAL_1162 <= _EVAL_442;
              end
            end
          end
        end
      end else begin
        if (_EVAL_898) begin
          if (_EVAL_1112) begin
            if (_EVAL_1937) begin
              if (!(_EVAL_939)) begin
                _EVAL_1162 <= _EVAL_442;
              end
            end
          end else begin
            _EVAL_1162 <= 1'h1;
          end
        end else begin
          if (_EVAL_1937) begin
            if (!(_EVAL_939)) begin
              _EVAL_1162 <= _EVAL_442;
            end
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1541) begin
        _EVAL_1167 <= _EVAL_1410;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1168 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_2120) begin
          _EVAL_1168 <= _EVAL_1908;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1178 <= 1'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_1210) begin
        _EVAL_1193 <= _EVAL_650;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1151) begin
        if (_EVAL_1722) begin
          _EVAL_1223 <= _EVAL_428;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1239 <= 32'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_755) begin
          _EVAL_1239 <= _EVAL_428;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1241 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1251) begin
          if (_EVAL_283) begin
            _EVAL_1241 <= _EVAL_707;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1249 <= 6'h0;
    end else begin
      _EVAL_1249 <= _EVAL_869[5:0];
    end
    if (_EVAL_1627) begin
      if (_EVAL_270) begin
        if (_EVAL_283) begin
          _EVAL_1261 <= _EVAL_996;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_677) begin
        _EVAL_1282 <= _EVAL_428;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1344 <= 2'h0;
    end
    if (_EVAL_146) begin
      _EVAL_1354 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_1366 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_270) begin
          if (_EVAL_283) begin
            if (_EVAL_670) begin
              _EVAL_1366 <= _EVAL_2162;
            end else begin
              _EVAL_1366 <= 1'h0;
            end
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1251) begin
        if (_EVAL_283) begin
          _EVAL_1376 <= _EVAL_996;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1381 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1310) begin
          _EVAL_1381 <= _EVAL_2222;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_749) begin
        _EVAL_1385 <= _EVAL_1264;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1392 <= 32'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_1251) begin
        if (_EVAL_283) begin
          _EVAL_1421 <= _EVAL_1217;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1424 <= 2'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_270) begin
        if (_EVAL_283) begin
          _EVAL_1425 <= _EVAL_1693;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1440 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1541) begin
          _EVAL_1440 <= _EVAL_1136;
        end
      end
    end
    _EVAL_1458 <= _EVAL_2173[2:0];
    if (_EVAL_146) begin
      _EVAL_1466 <= 2'h3;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1833) begin
          if (_EVAL_1229) begin
            _EVAL_1466 <= 2'h3;
          end else begin
            _EVAL_1466 <= 2'h0;
          end
        end else begin
          if (_EVAL_1937) begin
            if (_EVAL_939) begin
              if (_EVAL_490) begin
                _EVAL_1466 <= _EVAL_845;
              end
            end
          end
        end
      end else begin
        if (_EVAL_1937) begin
          if (_EVAL_939) begin
            if (_EVAL_490) begin
              _EVAL_1466 <= _EVAL_845;
            end
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1479 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1146) begin
          _EVAL_1479 <= _EVAL_659;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1251) begin
        if (_EVAL_283) begin
          _EVAL_1494 <= _EVAL_1693;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2120) begin
        _EVAL_1499 <= _EVAL_1416;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1532 <= 32'h10007;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1864) begin
          _EVAL_1532 <= _EVAL_516;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1545 <= 2'h0;
    end
    if (_EVAL_146) begin
      _EVAL_1555 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1644) begin
          _EVAL_1555 <= _EVAL_250;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1556 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_270) begin
          if (_EVAL_283) begin
            _EVAL_1556 <= _EVAL_707;
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1541) begin
        _EVAL_1563 <= _EVAL_654;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1567 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_1585 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1541) begin
          _EVAL_1585 <= _EVAL_1292;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1297) begin
        _EVAL_1589 <= _EVAL_741;
      end else begin
        if (_EVAL_1937) begin
          if (_EVAL_939) begin
            if (_EVAL_490) begin
              _EVAL_1589 <= _EVAL_427;
            end
          end
        end
      end
    end else begin
      if (_EVAL_1937) begin
        if (_EVAL_939) begin
          if (_EVAL_490) begin
            _EVAL_1589 <= _EVAL_427;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1593 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_2202) begin
          _EVAL_1593 <= _EVAL_1292;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2202) begin
        _EVAL_1608 <= _EVAL_1410;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2120) begin
        _EVAL_1620 <= _EVAL_1831;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2143) begin
        _EVAL_1632 <= _EVAL_428;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1666 <= 2'h0;
    end
    if (_EVAL_1627) begin
      if (_EVAL_1752) begin
        _EVAL_1688 <= _EVAL_428;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_309) begin
        if (_EVAL_283) begin
          _EVAL_1700 <= _EVAL_1693;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1251) begin
        if (_EVAL_1722) begin
          _EVAL_1725 <= _EVAL_428;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1644) begin
        _EVAL_1733 <= _EVAL_803;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_309) begin
        if (_EVAL_283) begin
          _EVAL_1743 <= _EVAL_1217;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1763 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1251) begin
          if (_EVAL_283) begin
            _EVAL_1763 <= _EVAL_1489;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1769 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_309) begin
          if (_EVAL_283) begin
            _EVAL_1769 <= _EVAL_1896;
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_364) begin
        _EVAL_1770 <= _EVAL_1831;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_2202) begin
        _EVAL_1792 <= _EVAL_271;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1808 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1251) begin
          if (_EVAL_283) begin
            _EVAL_1808 <= _EVAL_830;
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_749) begin
        _EVAL_1869 <= _EVAL_1093;
      end
    end
    if (_EVAL_146) begin
      _EVAL_1877 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1251) begin
          if (_EVAL_283) begin
            if (_EVAL_1489) begin
              _EVAL_1877 <= _EVAL_909;
            end else begin
              _EVAL_1877 <= 1'h0;
            end
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1895 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1151) begin
          if (_EVAL_283) begin
            _EVAL_1895 <= _EVAL_1170;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1899 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1151) begin
          if (_EVAL_283) begin
            _EVAL_1899 <= _EVAL_787;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1929 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_309) begin
          if (_EVAL_283) begin
            _EVAL_1929 <= _EVAL_707;
          end
        end
      end
    end
    _EVAL_1942 <= _EVAL_906[29:0];
    _EVAL_1952 <= _EVAL_326[29:0];
    if (_EVAL_146) begin
      _EVAL_1956 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1151) begin
          if (_EVAL_283) begin
            if (_EVAL_787) begin
              _EVAL_1956 <= _EVAL_2003;
            end else begin
              _EVAL_1956 <= 1'h0;
            end
          end
        end
      end
    end
    _EVAL_1978 <= _EVAL_265[29:0];
    if (_EVAL_146) begin
      _EVAL_1982 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_1986 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_270) begin
          if (_EVAL_283) begin
            _EVAL_1986 <= _EVAL_1590;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2002 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_309) begin
          if (_EVAL_283) begin
            _EVAL_2002 <= _EVAL_830;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2033 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1833) begin
          _EVAL_2033 <= _EVAL_928;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1541) begin
        _EVAL_2047 <= _EVAL_271;
      end
    end
    if (_EVAL_146) begin
      _EVAL_2063 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_309) begin
          if (_EVAL_283) begin
            _EVAL_2063 <= _EVAL_1590;
          end
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2074 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_2084 <= 1'h0;
    end else begin
      if (_EVAL_898) begin
        if (_EVAL_1112) begin
          _EVAL_2084 <= 1'h0;
        end else begin
          if (_EVAL_1937) begin
            if (_EVAL_939) begin
              if (_EVAL_490) begin
                _EVAL_2084 <= 1'h1;
              end
            end
          end
        end
      end else begin
        if (_EVAL_1937) begin
          if (_EVAL_939) begin
            if (_EVAL_490) begin
              _EVAL_2084 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1031) begin
        _EVAL_2090 <= _EVAL_282;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1386) begin
        _EVAL_2106 <= _EVAL_465;
      end else begin
        if (_EVAL_1437) begin
          _EVAL_2106 <= _EVAL_533;
        end else begin
          if (_EVAL_1317) begin
            _EVAL_2106 <= _EVAL_1976;
          end
        end
      end
    end else begin
      if (_EVAL_1317) begin
        _EVAL_2106 <= _EVAL_1976;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1644) begin
        _EVAL_2131 <= _EVAL_243;
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_309) begin
        if (_EVAL_283) begin
          _EVAL_2152 <= _EVAL_996;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2158 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_2159 <= 1'h0;
    end else begin
      if (_EVAL_2160) begin
        _EVAL_2159 <= 1'h1;
      end
    end
    _EVAL_2177 <= _EVAL_2082[5:0];
    if (_EVAL_1627) begin
      if (_EVAL_1644) begin
        _EVAL_2180 <= _EVAL_650;
      end
    end
    if (_EVAL_146) begin
      _EVAL_2181 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_364) begin
          _EVAL_2181 <= _EVAL_383;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2190 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1151) begin
          if (_EVAL_283) begin
            _EVAL_2190 <= _EVAL_1590;
          end
        end
      end
    end
    _EVAL_2210 <= _EVAL_2091[29:0];
    if (_EVAL_146) begin
      _EVAL_2220 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_270) begin
          if (_EVAL_283) begin
            _EVAL_2220 <= _EVAL_1973;
          end
        end
      end
    end
    _EVAL_2224 <= _EVAL_2068[29:0];
    if (_EVAL_146) begin
      _EVAL_2226 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_2120) begin
          _EVAL_2226 <= _EVAL_383;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2227 <= 2'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_2202) begin
          _EVAL_2227 <= _EVAL_1136;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_2230 <= 1'h0;
    end
    if (_EVAL_146) begin
      _EVAL_2232 <= 1'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_364) begin
          _EVAL_2232 <= _EVAL_1908;
        end
      end
    end
    if (_EVAL_1627) begin
      if (_EVAL_1210) begin
        _EVAL_2238 <= _EVAL_803;
      end
    end
  end
  always @(posedge _EVAL_50) begin
    if (_EVAL_146) begin
      _EVAL_645 <= 1'h0;
    end else begin
      if (_EVAL_1843) begin
        _EVAL_645 <= 1'h0;
      end else begin
        if (_EVAL_2192) begin
          _EVAL_645 <= 1'h1;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1212 <= 58'h0;
    end else begin
      if (_EVAL_1627) begin
        if (_EVAL_1657) begin
          _EVAL_1212 <= _EVAL_2077;
        end else begin
          if (_EVAL_531) begin
            _EVAL_1212 <= _EVAL_1403;
          end else begin
            if (_EVAL_565) begin
              _EVAL_1212 <= _EVAL_1947;
            end
          end
        end
      end else begin
        if (_EVAL_565) begin
          _EVAL_1212 <= _EVAL_1947;
        end
      end
    end
    if (_EVAL_146) begin
      _EVAL_1419 <= 6'h0;
    end else begin
      _EVAL_1419 <= _EVAL_1328[5:0];
    end
  end
endmodule
