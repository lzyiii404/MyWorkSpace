//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_299(
  input  [31:0] _EVAL,
  input  [2:0]  _EVAL_0,
  output [4:0]  _EVAL_1,
  output [32:0] _EVAL_2,
  input         _EVAL_3
);
  wire  round__EVAL;
  wire [6:0] round__EVAL_0;
  wire [2:0] round__EVAL_1;
  wire  round__EVAL_2;
  wire [32:0] round__EVAL_3;
  wire [32:0] round__EVAL_4;
  wire [4:0] round__EVAL_5;
  wire [15:0] _EVAL_21;
  wire [7:0] _EVAL_108;
  wire [3:0] _EVAL_90;
  wire  _EVAL_45;
  wire [31:0] _EVAL_139;
  wire [15:0] _EVAL_152;
  wire [15:0] _EVAL_140;
  wire [7:0] _EVAL_61;
  wire [3:0] _EVAL_66;
  wire  _EVAL_129;
  wire [7:0] _EVAL_39;
  wire [3:0] _EVAL_53;
  wire  _EVAL_22;
  wire [15:0] _EVAL_11;
  wire [7:0] _EVAL_159;
  wire [3:0] _EVAL_24;
  wire  _EVAL_112;
  wire [3:0] _EVAL_10;
  wire  _EVAL_57;
  wire [7:0] _EVAL_80;
  wire [3:0] _EVAL_15;
  wire  _EVAL_18;
  wire [3:0] _EVAL_47;
  wire  _EVAL_134;
  wire  _EVAL_149;
  wire  _EVAL_49;
  wire [1:0] _EVAL_27;
  wire [3:0] _EVAL_42;
  wire  _EVAL_177;
  wire  _EVAL_36;
  wire  _EVAL_98;
  wire [1:0] _EVAL_86;
  wire [1:0] _EVAL_101;
  wire [3:0] _EVAL_50;
  wire  _EVAL_158;
  wire  _EVAL_170;
  wire  _EVAL_92;
  wire [1:0] _EVAL_164;
  wire [1:0] _EVAL_131;
  wire [7:0] _EVAL_54;
  wire [3:0] _EVAL_71;
  wire  _EVAL_127;
  wire  _EVAL_114;
  wire  _EVAL_14;
  wire  _EVAL_166;
  wire [1:0] _EVAL_23;
  wire [1:0] _EVAL_16;
  wire [3:0] _EVAL_106;
  wire  _EVAL_4;
  wire  _EVAL_151;
  wire  _EVAL_143;
  wire [1:0] _EVAL_78;
  wire [1:0] _EVAL_8;
  wire [1:0] _EVAL_91;
  wire [2:0] _EVAL_100;
  wire [7:0] _EVAL_173;
  wire [3:0] _EVAL_63;
  wire  _EVAL_124;
  wire  _EVAL_146;
  wire  _EVAL_31;
  wire  _EVAL_155;
  wire  _EVAL_160;
  wire [1:0] _EVAL_9;
  wire [1:0] _EVAL_33;
  wire [1:0] _EVAL_169;
  wire [2:0] _EVAL_123;
  wire  _EVAL_133;
  wire  _EVAL_30;
  wire [31:0] _EVAL_153;
  wire [31:0] _EVAL_137;
  wire  _EVAL_32;
  wire [7:0] _EVAL_34;
  wire  _EVAL_156;
  wire [3:0] _EVAL_162;
  wire  _EVAL_118;
  wire  _EVAL_161;
  wire  _EVAL_7;
  wire  _EVAL_176;
  wire [1:0] _EVAL_82;
  wire [1:0] _EVAL_58;
  wire [3:0] _EVAL_38;
  wire  _EVAL_97;
  wire  _EVAL_144;
  wire  _EVAL_163;
  wire [1:0] _EVAL_67;
  wire [1:0] _EVAL_171;
  wire [1:0] _EVAL_6;
  wire [2:0] _EVAL_5;
  wire  _EVAL_132;
  wire  _EVAL_73;
  wire [1:0] _EVAL_109;
  wire [1:0] _EVAL_56;
  wire  _EVAL_60;
  wire  _EVAL_148;
  wire [1:0] _EVAL_83;
  wire [1:0] _EVAL_96;
  wire [1:0] _EVAL_55;
  wire [2:0] _EVAL_95;
  wire [2:0] _EVAL_68;
  wire [3:0] _EVAL_117;
  wire  _EVAL_147;
  wire  _EVAL_81;
  wire [1:0] _EVAL_88;
  wire  _EVAL_13;
  wire  _EVAL_138;
  wire [1:0] _EVAL_93;
  wire [1:0] _EVAL_44;
  wire [1:0] _EVAL_77;
  wire [2:0] _EVAL_130;
  wire [3:0] _EVAL_105;
  wire  _EVAL_75;
  wire  _EVAL_107;
  wire  _EVAL_113;
  wire  _EVAL_125;
  wire [1:0] _EVAL_70;
  wire [1:0] _EVAL_19;
  wire  _EVAL_104;
  wire  _EVAL_12;
  wire [1:0] _EVAL_37;
  wire [1:0] _EVAL_76;
  wire [1:0] _EVAL_103;
  wire [2:0] _EVAL_43;
  wire [2:0] _EVAL_115;
  wire [3:0] _EVAL_141;
  wire [3:0] _EVAL_41;
  wire [4:0] _EVAL_25;
  wire  _EVAL_136;
  wire  _EVAL_79;
  wire  _EVAL_17;
  wire [1:0] _EVAL_154;
  wire [1:0] _EVAL_167;
  wire [1:0] _EVAL_126;
  wire [2:0] _EVAL_150;
  wire  _EVAL_172;
  wire  _EVAL_64;
  wire [2:0] _EVAL_111;
  wire [3:0] _EVAL_120;
  wire  _EVAL_51;
  wire  _EVAL_145;
  wire  _EVAL_89;
  wire  _EVAL_65;
  wire [1:0] _EVAL_59;
  wire [1:0] _EVAL_135;
  wire [3:0] _EVAL_52;
  wire  _EVAL_74;
  wire  _EVAL_28;
  wire  _EVAL_157;
  wire [1:0] _EVAL_128;
  wire [1:0] _EVAL_85;
  wire [1:0] _EVAL_20;
  wire [2:0] _EVAL_119;
  wire [2:0] _EVAL_26;
  wire [3:0] _EVAL_121;
  wire [3:0] _EVAL_46;
  wire [4:0] _EVAL_102;
  wire [4:0] _EVAL_48;
  wire  _EVAL_99;
  wire  _EVAL_29;
  wire  _EVAL_40;
  wire [31:0] _EVAL_87;
  wire  _EVAL_116;
  wire  _EVAL_110;
  wire [4:0] _EVAL_94;
  wire [4:0] _EVAL_62;
  wire [4:0] _EVAL_69;
  wire [4:0] _EVAL_72;
  wire [5:0] _EVAL_175;
  wire [62:0] _EVAL_122;
  wire [62:0] _EVAL_35;
  wire [62:0] _EVAL_174;
  wire [31:0] _EVAL_142;
  wire  _EVAL_84;
  SiFive__EVAL_298 round (
    ._EVAL(round__EVAL),
    ._EVAL_0(round__EVAL_0),
    ._EVAL_1(round__EVAL_1),
    ._EVAL_2(round__EVAL_2),
    ._EVAL_3(round__EVAL_3),
    ._EVAL_4(round__EVAL_4),
    ._EVAL_5(round__EVAL_5)
  );
  assign _EVAL_21 = _EVAL[31:16];
  assign _EVAL_108 = _EVAL_21[7:0];
  assign _EVAL_90 = _EVAL_108[3:0];
  assign _EVAL_45 = _EVAL_90[3];
  assign _EVAL_139 = ~ _EVAL;
  assign _EVAL_152 = _EVAL_139[15:0];
  assign _EVAL_140 = _EVAL[15:0];
  assign _EVAL_61 = _EVAL_140[15:8];
  assign _EVAL_66 = _EVAL_61[7:4];
  assign _EVAL_129 = _EVAL_66 != 4'h0;
  assign _EVAL_39 = _EVAL_152[15:8];
  assign _EVAL_53 = _EVAL_39[3:0];
  assign _EVAL_22 = _EVAL_53[1];
  assign _EVAL_11 = _EVAL_139[31:16];
  assign _EVAL_159 = _EVAL_11[7:0];
  assign _EVAL_24 = _EVAL_159[3:0];
  assign _EVAL_112 = _EVAL_24[1];
  assign _EVAL_10 = _EVAL_39[7:4];
  assign _EVAL_57 = _EVAL_10 != 4'h0;
  assign _EVAL_80 = _EVAL_140[7:0];
  assign _EVAL_15 = _EVAL_80[7:4];
  assign _EVAL_18 = _EVAL_15 != 4'h0;
  assign _EVAL_47 = _EVAL_159[7:4];
  assign _EVAL_134 = _EVAL_47[3];
  assign _EVAL_149 = _EVAL_10[2];
  assign _EVAL_49 = _EVAL_10[1];
  assign _EVAL_27 = _EVAL_149 ? 2'h2 : {{1'd0}, _EVAL_49};
  assign _EVAL_42 = _EVAL_108[7:4];
  assign _EVAL_177 = _EVAL_42[3];
  assign _EVAL_36 = _EVAL_42[2];
  assign _EVAL_98 = _EVAL_42[1];
  assign _EVAL_86 = _EVAL_36 ? 2'h2 : {{1'd0}, _EVAL_98};
  assign _EVAL_101 = _EVAL_177 ? 2'h3 : _EVAL_86;
  assign _EVAL_50 = _EVAL_80[3:0];
  assign _EVAL_158 = _EVAL_50[3];
  assign _EVAL_170 = _EVAL_50[2];
  assign _EVAL_92 = _EVAL_50[1];
  assign _EVAL_164 = _EVAL_170 ? 2'h2 : {{1'd0}, _EVAL_92};
  assign _EVAL_131 = _EVAL_158 ? 2'h3 : _EVAL_164;
  assign _EVAL_54 = _EVAL_21[15:8];
  assign _EVAL_71 = _EVAL_54[7:4];
  assign _EVAL_127 = _EVAL_71 != 4'h0;
  assign _EVAL_114 = _EVAL_71[3];
  assign _EVAL_14 = _EVAL_71[2];
  assign _EVAL_166 = _EVAL_71[1];
  assign _EVAL_23 = _EVAL_14 ? 2'h2 : {{1'd0}, _EVAL_166};
  assign _EVAL_16 = _EVAL_114 ? 2'h3 : _EVAL_23;
  assign _EVAL_106 = _EVAL_54[3:0];
  assign _EVAL_4 = _EVAL_106[3];
  assign _EVAL_151 = _EVAL_106[2];
  assign _EVAL_143 = _EVAL_106[1];
  assign _EVAL_78 = _EVAL_151 ? 2'h2 : {{1'd0}, _EVAL_143};
  assign _EVAL_8 = _EVAL_4 ? 2'h3 : _EVAL_78;
  assign _EVAL_91 = _EVAL_127 ? _EVAL_16 : _EVAL_8;
  assign _EVAL_100 = {_EVAL_127,_EVAL_91};
  assign _EVAL_173 = _EVAL_152[7:0];
  assign _EVAL_63 = _EVAL_173[3:0];
  assign _EVAL_124 = _EVAL_63[2];
  assign _EVAL_146 = _EVAL_47[1];
  assign _EVAL_31 = _EVAL_15[3];
  assign _EVAL_155 = _EVAL_15[2];
  assign _EVAL_160 = _EVAL_15[1];
  assign _EVAL_9 = _EVAL_155 ? 2'h2 : {{1'd0}, _EVAL_160};
  assign _EVAL_33 = _EVAL_31 ? 2'h3 : _EVAL_9;
  assign _EVAL_169 = _EVAL_18 ? _EVAL_33 : _EVAL_131;
  assign _EVAL_123 = {_EVAL_18,_EVAL_169};
  assign _EVAL_133 = _EVAL[31];
  assign _EVAL_30 = _EVAL_3 & _EVAL_133;
  assign _EVAL_153 = 32'h0 - _EVAL;
  assign _EVAL_137 = _EVAL_30 ? _EVAL_153 : _EVAL;
  assign _EVAL_32 = _EVAL_11 != 16'h0;
  assign _EVAL_34 = _EVAL_11[15:8];
  assign _EVAL_156 = _EVAL_34 != 8'h0;
  assign _EVAL_162 = _EVAL_34[7:4];
  assign _EVAL_118 = _EVAL_162 != 4'h0;
  assign _EVAL_161 = _EVAL_162[3];
  assign _EVAL_7 = _EVAL_162[2];
  assign _EVAL_176 = _EVAL_162[1];
  assign _EVAL_82 = _EVAL_7 ? 2'h2 : {{1'd0}, _EVAL_176};
  assign _EVAL_58 = _EVAL_161 ? 2'h3 : _EVAL_82;
  assign _EVAL_38 = _EVAL_34[3:0];
  assign _EVAL_97 = _EVAL_38[3];
  assign _EVAL_144 = _EVAL_38[2];
  assign _EVAL_163 = _EVAL_38[1];
  assign _EVAL_67 = _EVAL_144 ? 2'h2 : {{1'd0}, _EVAL_163};
  assign _EVAL_171 = _EVAL_97 ? 2'h3 : _EVAL_67;
  assign _EVAL_6 = _EVAL_118 ? _EVAL_58 : _EVAL_171;
  assign _EVAL_5 = {_EVAL_118,_EVAL_6};
  assign _EVAL_132 = _EVAL_47 != 4'h0;
  assign _EVAL_73 = _EVAL_47[2];
  assign _EVAL_109 = _EVAL_73 ? 2'h2 : {{1'd0}, _EVAL_146};
  assign _EVAL_56 = _EVAL_134 ? 2'h3 : _EVAL_109;
  assign _EVAL_60 = _EVAL_24[3];
  assign _EVAL_148 = _EVAL_24[2];
  assign _EVAL_83 = _EVAL_148 ? 2'h2 : {{1'd0}, _EVAL_112};
  assign _EVAL_96 = _EVAL_60 ? 2'h3 : _EVAL_83;
  assign _EVAL_55 = _EVAL_132 ? _EVAL_56 : _EVAL_96;
  assign _EVAL_95 = {_EVAL_132,_EVAL_55};
  assign _EVAL_68 = _EVAL_156 ? _EVAL_5 : _EVAL_95;
  assign _EVAL_117 = {_EVAL_156,_EVAL_68};
  assign _EVAL_147 = _EVAL_39 != 8'h0;
  assign _EVAL_81 = _EVAL_10[3];
  assign _EVAL_88 = _EVAL_81 ? 2'h3 : _EVAL_27;
  assign _EVAL_13 = _EVAL_53[3];
  assign _EVAL_138 = _EVAL_53[2];
  assign _EVAL_93 = _EVAL_138 ? 2'h2 : {{1'd0}, _EVAL_22};
  assign _EVAL_44 = _EVAL_13 ? 2'h3 : _EVAL_93;
  assign _EVAL_77 = _EVAL_57 ? _EVAL_88 : _EVAL_44;
  assign _EVAL_130 = {_EVAL_57,_EVAL_77};
  assign _EVAL_105 = _EVAL_173[7:4];
  assign _EVAL_75 = _EVAL_105 != 4'h0;
  assign _EVAL_107 = _EVAL_105[3];
  assign _EVAL_113 = _EVAL_105[2];
  assign _EVAL_125 = _EVAL_105[1];
  assign _EVAL_70 = _EVAL_113 ? 2'h2 : {{1'd0}, _EVAL_125};
  assign _EVAL_19 = _EVAL_107 ? 2'h3 : _EVAL_70;
  assign _EVAL_104 = _EVAL_63[3];
  assign _EVAL_12 = _EVAL_63[1];
  assign _EVAL_37 = _EVAL_124 ? 2'h2 : {{1'd0}, _EVAL_12};
  assign _EVAL_76 = _EVAL_104 ? 2'h3 : _EVAL_37;
  assign _EVAL_103 = _EVAL_75 ? _EVAL_19 : _EVAL_76;
  assign _EVAL_43 = {_EVAL_75,_EVAL_103};
  assign _EVAL_115 = _EVAL_147 ? _EVAL_130 : _EVAL_43;
  assign _EVAL_141 = {_EVAL_147,_EVAL_115};
  assign _EVAL_41 = _EVAL_32 ? _EVAL_117 : _EVAL_141;
  assign _EVAL_25 = {_EVAL_32,_EVAL_41};
  assign _EVAL_136 = _EVAL_42 != 4'h0;
  assign _EVAL_79 = _EVAL_90[2];
  assign _EVAL_17 = _EVAL_90[1];
  assign _EVAL_154 = _EVAL_79 ? 2'h2 : {{1'd0}, _EVAL_17};
  assign _EVAL_167 = _EVAL_45 ? 2'h3 : _EVAL_154;
  assign _EVAL_126 = _EVAL_136 ? _EVAL_101 : _EVAL_167;
  assign _EVAL_150 = {_EVAL_136,_EVAL_126};
  assign _EVAL_172 = _EVAL_21 != 16'h0;
  assign _EVAL_64 = _EVAL_54 != 8'h0;
  assign _EVAL_111 = _EVAL_64 ? _EVAL_100 : _EVAL_150;
  assign _EVAL_120 = {_EVAL_64,_EVAL_111};
  assign _EVAL_51 = _EVAL_61 != 8'h0;
  assign _EVAL_145 = _EVAL_66[3];
  assign _EVAL_89 = _EVAL_66[2];
  assign _EVAL_65 = _EVAL_66[1];
  assign _EVAL_59 = _EVAL_89 ? 2'h2 : {{1'd0}, _EVAL_65};
  assign _EVAL_135 = _EVAL_145 ? 2'h3 : _EVAL_59;
  assign _EVAL_52 = _EVAL_61[3:0];
  assign _EVAL_74 = _EVAL_52[3];
  assign _EVAL_28 = _EVAL_52[2];
  assign _EVAL_157 = _EVAL_52[1];
  assign _EVAL_128 = _EVAL_28 ? 2'h2 : {{1'd0}, _EVAL_157};
  assign _EVAL_85 = _EVAL_74 ? 2'h3 : _EVAL_128;
  assign _EVAL_20 = _EVAL_129 ? _EVAL_135 : _EVAL_85;
  assign _EVAL_119 = {_EVAL_129,_EVAL_20};
  assign _EVAL_26 = _EVAL_51 ? _EVAL_119 : _EVAL_123;
  assign _EVAL_121 = {_EVAL_51,_EVAL_26};
  assign _EVAL_46 = _EVAL_172 ? _EVAL_120 : _EVAL_121;
  assign _EVAL_102 = {_EVAL_172,_EVAL_46};
  assign _EVAL_48 = _EVAL_30 ? _EVAL_25 : _EVAL_102;
  assign _EVAL_99 = _EVAL[0];
  assign _EVAL_29 = _EVAL_99 == 1'h0;
  assign _EVAL_40 = _EVAL_30 & _EVAL_29;
  assign _EVAL_87 = _EVAL_139 & _EVAL_153;
  assign _EVAL_116 = _EVAL_87 == 32'h0;
  assign _EVAL_110 = _EVAL_40 & _EVAL_116;
  assign _EVAL_94 = ~ _EVAL_48;
  assign _EVAL_62 = _EVAL_94 - 5'h1;
  assign _EVAL_69 = _EVAL_110 ? _EVAL_62 : _EVAL_94;
  assign _EVAL_72 = ~ _EVAL_69;
  assign _EVAL_175 = {1'h1,_EVAL_72};
  assign _EVAL_122 = {{31'd0}, _EVAL_137};
  assign _EVAL_35 = _EVAL_122 << _EVAL_94;
  assign _EVAL_174 = _EVAL_35 >> _EVAL_110;
  assign _EVAL_142 = _EVAL_174[31:0];
  assign _EVAL_84 = _EVAL_142[31];
  assign round__EVAL_1 = _EVAL_0;
  assign round__EVAL_0 = {1'b0,$signed(_EVAL_175)};
  assign _EVAL_2 = round__EVAL_4;
  assign round__EVAL_2 = _EVAL_84 == 1'h0;
  assign round__EVAL_3 = {{1'd0}, _EVAL_142};
  assign round__EVAL = _EVAL_3 & _EVAL_133;
  assign _EVAL_1 = round__EVAL_5;
endmodule
