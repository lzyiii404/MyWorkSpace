//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_224_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [7:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [3:0]  _EVAL_20,
  input  [31:0] _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input  [31:0] _EVAL_24,
  input  [31:0] _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [3:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input  [2:0]  _EVAL_33
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_44;
  reg [31:0] _RAND_0;
  reg  _EVAL_56;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_116;
  reg [31:0] _RAND_2;
  reg  _EVAL_118;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_150;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_168;
  reg [31:0] _RAND_5;
  reg [31:0] _EVAL_180;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_214;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_220;
  reg [31:0] _RAND_8;
  reg [1:0] _EVAL_270;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_300;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_320;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_348;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_374;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_384;
  reg [31:0] _RAND_14;
  reg [31:0] _EVAL_431;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_433;
  reg [31:0] _RAND_16;
  reg [4:0] _EVAL_449;
  reg [31:0] _RAND_17;
  reg [1:0] _EVAL_483;
  reg [31:0] _RAND_18;
  reg [2:0] _EVAL_502;
  reg [31:0] _RAND_19;
  reg [4:0] _EVAL_535;
  reg [31:0] _RAND_20;
  reg [3:0] _EVAL_562;
  reg [31:0] _RAND_21;
  reg [4:0] _EVAL_592;
  reg [31:0] _RAND_22;
  reg [2:0] _EVAL_598;
  reg [31:0] _RAND_23;
  reg [7:0] _EVAL_623;
  reg [31:0] _RAND_24;
  reg [2:0] _EVAL_628;
  reg [31:0] _RAND_25;
  reg [4:0] _EVAL_630;
  reg [31:0] _RAND_26;
  reg [3:0] _EVAL_639;
  reg [31:0] _RAND_27;
  wire  _EVAL_43;
  wire  _EVAL_566;
  wire  _EVAL_450;
  wire  _EVAL_610;
  wire [31:0] _EVAL_47;
  wire [31:0] _EVAL_380;
  wire [32:0] _EVAL_262;
  wire [31:0] _EVAL_63;
  wire [32:0] _EVAL_552;
  wire [32:0] _EVAL_627;
  wire [32:0] _EVAL_364;
  wire  _EVAL_606;
  wire [31:0] _EVAL_519;
  wire [32:0] _EVAL_391;
  wire [32:0] _EVAL_420;
  wire [32:0] _EVAL_361;
  wire  _EVAL_454;
  wire  _EVAL_599;
  wire [31:0] _EVAL_589;
  wire [32:0] _EVAL_467;
  wire [32:0] _EVAL_138;
  wire [32:0] _EVAL_289;
  wire  _EVAL_165;
  wire  _EVAL_513;
  wire [31:0] _EVAL_94;
  wire [32:0] _EVAL_547;
  wire [32:0] _EVAL_74;
  wire [32:0] _EVAL_573;
  wire  _EVAL_617;
  wire  _EVAL_225;
  wire [31:0] _EVAL_488;
  wire [32:0] _EVAL_83;
  wire [32:0] _EVAL_344;
  wire [32:0] _EVAL_45;
  wire  _EVAL_564;
  wire  _EVAL_652;
  wire [32:0] _EVAL_624;
  wire [32:0] _EVAL_193;
  wire [32:0] _EVAL_245;
  wire  _EVAL_311;
  wire  _EVAL_337;
  wire [31:0] _EVAL_269;
  wire [32:0] _EVAL_473;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_50;
  wire  _EVAL_279;
  wire  _EVAL_81;
  wire [31:0] _EVAL_607;
  wire [32:0] _EVAL_609;
  wire [32:0] _EVAL_343;
  wire [32:0] _EVAL_286;
  wire  _EVAL_46;
  wire  _EVAL_435;
  wire [31:0] _EVAL_99;
  wire [32:0] _EVAL_649;
  wire [32:0] _EVAL_338;
  wire [32:0] _EVAL_405;
  wire  _EVAL_586;
  wire  _EVAL_243;
  wire  _EVAL_582;
  wire  _EVAL_176;
  wire  _EVAL_230;
  wire  _EVAL_315;
  wire  _EVAL_531;
  wire  _EVAL_618;
  wire [22:0] _EVAL_126;
  wire [7:0] _EVAL_256;
  wire [7:0] _EVAL_61;
  wire [4:0] _EVAL_472;
  wire [4:0] _EVAL_137;
  wire  _EVAL_264;
  wire  _EVAL_539;
  wire [22:0] _EVAL_55;
  wire [7:0] _EVAL_553;
  wire [7:0] _EVAL_232;
  wire [4:0] _EVAL_451;
  wire [4:0] _EVAL_86;
  wire  _EVAL_164;
  wire [1:0] _EVAL_572;
  wire [3:0] _EVAL_386;
  wire [2:0] _EVAL_87;
  wire [2:0] _EVAL_219;
  wire  _EVAL_182;
  wire  _EVAL_37;
  wire  _EVAL_128;
  wire  _EVAL_144;
  wire  _EVAL_325;
  wire  _EVAL_69;
  wire  _EVAL_400;
  wire [22:0] _EVAL_387;
  wire [7:0] _EVAL_226;
  wire [7:0] _EVAL_643;
  wire [31:0] _EVAL_490;
  wire [31:0] _EVAL_353;
  wire [31:0] _EVAL_203;
  wire [32:0] _EVAL_274;
  wire [32:0] _EVAL_428;
  wire [32:0] _EVAL_479;
  wire [31:0] _EVAL_597;
  wire  _EVAL_481;
  wire  _EVAL_197;
  wire  _EVAL_258;
  wire [31:0] _EVAL_530;
  wire [32:0] _EVAL_629;
  wire [32:0] _EVAL_356;
  wire [32:0] _EVAL_192;
  wire  _EVAL_35;
  wire  _EVAL_500;
  wire  _EVAL_359;
  wire  _EVAL_275;
  wire  _EVAL_278;
  wire  _EVAL_51;
  wire  _EVAL_382;
  wire  _EVAL_542;
  wire  _EVAL_580;
  wire  _EVAL_48;
  wire  _EVAL_561;
  wire  _EVAL_72;
  wire  _EVAL_257;
  wire  _EVAL_70;
  wire  _EVAL_312;
  wire  _EVAL_108;
  wire [1:0] _EVAL_213;
  wire [1:0] _EVAL_581;
  wire [1:0] _EVAL_308;
  wire  _EVAL_75;
  wire  _EVAL_558;
  wire  _EVAL_68;
  wire  _EVAL_299;
  wire  _EVAL_267;
  wire  _EVAL_565;
  wire  _EVAL_587;
  wire [7:0] _EVAL_367;
  wire  _EVAL_465;
  wire  _EVAL_127;
  wire  _EVAL_134;
  wire [7:0] _EVAL_196;
  wire  _EVAL_570;
  wire  _EVAL_332;
  wire  _EVAL_155;
  wire  _EVAL_555;
  wire  _EVAL_79;
  wire  _EVAL_89;
  wire  _EVAL_326;
  wire  _EVAL_252;
  wire [31:0] _EVAL_236;
  wire [32:0] _EVAL_266;
  wire [31:0] _EVAL_457;
  wire  _EVAL_368;
  wire  _EVAL_616;
  wire  _EVAL_498;
  wire  _EVAL_462;
  wire  _EVAL_579;
  wire  _EVAL_307;
  wire  _EVAL_430;
  wire  _EVAL_503;
  wire  _EVAL_438;
  wire  _EVAL_216;
  wire  _EVAL_591;
  wire  _EVAL_244;
  wire  _EVAL_76;
  wire  _EVAL_418;
  wire  _EVAL_115;
  wire  _EVAL_396;
  wire  _EVAL_588;
  wire  _EVAL_363;
  wire  _EVAL_480;
  wire  _EVAL_294;
  wire  _EVAL_296;
  wire  _EVAL_303;
  wire  _EVAL_634;
  wire  _EVAL_575;
  wire  _EVAL_324;
  wire  _EVAL_611;
  wire  _EVAL_268;
  wire  _EVAL_522;
  wire  _EVAL_527;
  wire  _EVAL_183;
  wire  _EVAL_548;
  wire  _EVAL_120;
  wire  _EVAL_439;
  wire  _EVAL_442;
  wire  _EVAL_246;
  wire  _EVAL_210;
  wire  _EVAL_97;
  wire  _EVAL_306;
  wire  _EVAL_166;
  wire  _EVAL_365;
  wire  _EVAL_233;
  wire  _EVAL_549;
  wire  _EVAL_77;
  wire  _EVAL_596;
  wire  _EVAL_254;
  wire  _EVAL_189;
  wire  _EVAL_301;
  wire  _EVAL_122;
  wire [7:0] _EVAL_119;
  wire  _EVAL_205;
  wire  _EVAL_401;
  wire [31:0] _EVAL_234;
  wire [32:0] _EVAL_407;
  wire [32:0] _EVAL_64;
  wire [32:0] _EVAL_349;
  wire  _EVAL_569;
  wire [31:0] _EVAL_619;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_355;
  wire [32:0] _EVAL_376;
  wire  _EVAL_71;
  wire  _EVAL_421;
  wire [31:0] _EVAL_82;
  wire [32:0] _EVAL_277;
  wire [32:0] _EVAL_358;
  wire [32:0] _EVAL_466;
  wire  _EVAL_577;
  wire  _EVAL_574;
  wire  _EVAL_259;
  wire  _EVAL_492;
  wire  _EVAL_313;
  wire  _EVAL_170;
  wire  _EVAL_477;
  wire [7:0] _EVAL_283;
  wire [31:0] _EVAL_327;
  wire [32:0] _EVAL_536;
  wire [32:0] _EVAL_153;
  wire [32:0] _EVAL_362;
  wire  _EVAL_373;
  wire  _EVAL_132;
  wire  _EVAL_600;
  wire  _EVAL_217;
  wire  _EVAL_455;
  wire  _EVAL_96;
  wire  _EVAL_145;
  wire  _EVAL_517;
  wire [31:0] _EVAL_404;
  wire [32:0] _EVAL_637;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_80;
  wire [32:0] _EVAL_228;
  wire [32:0] _EVAL_395;
  wire  _EVAL_221;
  wire  _EVAL_408;
  wire  _EVAL_162;
  wire  _EVAL_478;
  wire [32:0] _EVAL_141;
  wire  _EVAL_124;
  wire  _EVAL_114;
  wire  _EVAL_642;
  wire  _EVAL_285;
  wire  _EVAL_49;
  wire  _EVAL_463;
  wire  _EVAL_171;
  wire  _EVAL_567;
  wire  _EVAL_528;
  wire  _EVAL_626;
  wire  _EVAL_135;
  wire  _EVAL_281;
  wire  _EVAL_330;
  wire [4:0] _EVAL_88;
  wire  _EVAL_621;
  wire  _EVAL_511;
  wire  _EVAL_508;
  wire  _EVAL_341;
  wire  _EVAL_131;
  wire  _EVAL_650;
  wire  _EVAL_631;
  wire  _EVAL_406;
  wire [4:0] _EVAL_340;
  wire [4:0] _EVAL_354;
  wire  _EVAL_571;
  wire  _EVAL_328;
  wire  _EVAL_100;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire [7:0] _EVAL_347;
  wire  _EVAL_392;
  wire  _EVAL_215;
  wire  _EVAL_298;
  wire  _EVAL_510;
  wire  _EVAL_211;
  wire [1:0] _EVAL_471;
  wire  _EVAL_550;
  wire  _EVAL_422;
  wire  _EVAL_370;
  wire  _EVAL_154;
  wire [32:0] _EVAL_414;
  wire [32:0] _EVAL_429;
  wire [32:0] _EVAL_302;
  wire  _EVAL_556;
  wire  _EVAL_181;
  wire [32:0] _EVAL_417;
  wire [32:0] _EVAL_93;
  wire  _EVAL_411;
  wire  _EVAL_85;
  wire [31:0] _EVAL_351;
  wire [32:0] _EVAL_184;
  wire [32:0] _EVAL_419;
  wire [32:0] _EVAL_653;
  wire  _EVAL_436;
  wire  _EVAL_398;
  wire  _EVAL_292;
  wire  _EVAL_635;
  wire  _EVAL_540;
  wire  _EVAL_515;
  wire [32:0] _EVAL_161;
  wire [32:0] _EVAL_187;
  wire [32:0] _EVAL_65;
  wire  _EVAL_106;
  wire  _EVAL_57;
  wire [32:0] _EVAL_142;
  wire [32:0] _EVAL_537;
  wire  _EVAL_272;
  wire  _EVAL_255;
  wire  _EVAL_375;
  wire  _EVAL_484;
  wire [32:0] _EVAL_113;
  wire [32:0] _EVAL_524;
  wire  _EVAL_223;
  wire  _EVAL_448;
  wire  _EVAL_546;
  wire  _EVAL_319;
  wire  _EVAL_445;
  wire  _EVAL_101;
  wire  _EVAL_251;
  wire  _EVAL_282;
  wire  _EVAL_147;
  wire  _EVAL_622;
  wire [1:0] _EVAL_146;
  wire [1:0] _EVAL_437;
  wire [1:0] _EVAL_424;
  wire  _EVAL_159;
  wire  _EVAL_453;
  wire  _EVAL_209;
  wire  _EVAL_276;
  wire  _EVAL_167;
  wire [7:0] _EVAL_434;
  wire  _EVAL_645;
  wire  _EVAL_190;
  wire  _EVAL_333;
  wire [31:0] _EVAL_194;
  wire  _EVAL_521;
  wire  _EVAL_321;
  wire  _EVAL_111;
  wire [7:0] _EVAL_107;
  wire  _EVAL_416;
  wire  _EVAL_73;
  wire  _EVAL_432;
  wire  _EVAL_632;
  wire  _EVAL_494;
  wire  _EVAL_242;
  wire  _EVAL_310;
  wire  _EVAL_177;
  wire [31:0] _EVAL_284;
  wire  _EVAL_633;
  wire [31:0] _EVAL_227;
  wire [32:0] _EVAL_560;
  wire [32:0] _EVAL_316;
  wire [32:0] _EVAL_496;
  wire  _EVAL_648;
  wire  _EVAL_174;
  wire  _EVAL_602;
  wire  _EVAL_148;
  wire [31:0] _EVAL_638;
  wire [32:0] _EVAL_309;
  wire [32:0] _EVAL_644;
  wire [32:0] _EVAL_497;
  wire  _EVAL_188;
  wire  _EVAL_157;
  wire [31:0] _EVAL_533;
  wire [32:0] _EVAL_468;
  wire [32:0] _EVAL_92;
  wire [32:0] _EVAL_204;
  wire  _EVAL_393;
  wire  _EVAL_91;
  wire [31:0] _EVAL_288;
  wire [32:0] _EVAL_425;
  wire [32:0] _EVAL_41;
  wire [32:0] _EVAL_379;
  wire  _EVAL_231;
  wire  _EVAL_200;
  wire  _EVAL_493;
  wire [32:0] _EVAL_293;
  wire  _EVAL_377;
  wire  _EVAL_186;
  wire  _EVAL_608;
  wire  _EVAL_604;
  wire [31:0] _EVAL_636;
  wire [32:0] _EVAL_280;
  wire [32:0] _EVAL_504;
  wire [32:0] _EVAL_95;
  wire  _EVAL_175;
  wire  _EVAL_265;
  wire [31:0] _EVAL_149;
  wire [32:0] _EVAL_249;
  wire [32:0] _EVAL_640;
  wire [32:0] _EVAL_495;
  wire  _EVAL_485;
  wire  _EVAL_207;
  wire  _EVAL_104;
  wire  _EVAL_646;
  wire  _EVAL_461;
  wire  _EVAL_287;
  wire  _EVAL_331;
  wire  _EVAL_603;
  wire  _EVAL_84;
  wire  _EVAL_169;
  wire  _EVAL_427;
  wire  _EVAL_525;
  wire  _EVAL_291;
  wire  _EVAL_509;
  wire  _EVAL_40;
  wire  _EVAL_66;
  wire  _EVAL_62;
  wire  _EVAL_601;
  wire  _EVAL_423;
  wire  _EVAL_42;
  wire  _EVAL_518;
  wire [4:0] _EVAL_641;
  wire  _EVAL_551;
  wire  _EVAL_512;
  wire  _EVAL_173;
  wire  _EVAL_334;
  wire  _EVAL_520;
  wire  _EVAL_505;
  wire  _EVAL_459;
  wire  _EVAL_526;
  wire  _EVAL_317;
  wire  _EVAL_378;
  wire  _EVAL_229;
  wire  _EVAL_516;
  wire  _EVAL_152;
  wire  _EVAL_538;
  wire  _EVAL_314;
  wire  _EVAL_198;
  wire  _EVAL_476;
  wire [7:0] _EVAL_290;
  wire [7:0] _EVAL_615;
  wire [7:0] _EVAL_237;
  wire [7:0] _EVAL_143;
  wire  _EVAL_410;
  wire  _EVAL_222;
  wire  _EVAL_199;
  wire  _EVAL_501;
  wire  _EVAL_241;
  wire  _EVAL_160;
  wire  _EVAL_532;
  wire  _EVAL_585;
  wire [7:0] _EVAL_506;
  wire [7:0] _EVAL_60;
  wire  _EVAL_139;
  wire  _EVAL_67;
  wire  _EVAL_178;
  wire  _EVAL_253;
  wire  _EVAL_620;
  wire  _EVAL_151;
  wire  _EVAL_595;
  wire  _EVAL_412;
  wire  _EVAL_38;
  wire  _EVAL_58;
  wire  _EVAL_594;
  wire  _EVAL_305;
  wire  _EVAL_369;
  wire  _EVAL_415;
  wire  _EVAL_413;
  wire  _EVAL_447;
  wire  _EVAL_475;
  wire  _EVAL_563;
  wire [4:0] _EVAL_179;
  wire  _EVAL_191;
  wire  _EVAL_590;
  wire  _EVAL_469;
  wire  _EVAL_271;
  wire  _EVAL_339;
  wire  _EVAL_125;
  wire  _EVAL_409;
  wire  _EVAL_105;
  wire  _EVAL_240;
  wire  _EVAL_456;
  wire  _EVAL_583;
  wire  _EVAL_371;
  wire  _EVAL_36;
  wire  _EVAL_593;
  wire  _EVAL_52;
  wire  _EVAL_129;
  wire  _EVAL_458;
  wire  _EVAL_614;
  wire  _EVAL_444;
  wire [31:0] _EVAL_460;
  wire  _EVAL_499;
  wire  _EVAL_578;
  wire  _EVAL_238;
  wire  _EVAL_295;
  wire  _EVAL_136;
  wire  _EVAL_112;
  wire  _EVAL_185;
  wire  _EVAL_397;
  wire  _EVAL_441;
  wire [7:0] _EVAL_557;
  wire  _EVAL_346;
  wire  _EVAL_208;
  wire  _EVAL_117;
  wire  _EVAL_133;
  wire  _EVAL_78;
  wire  _EVAL_366;
  wire  _EVAL_98;
  wire  _EVAL_474;
  wire  _EVAL_541;
  wire  _EVAL_464;
  wire  _EVAL_486;
  wire  _EVAL_59;
  wire  _EVAL_206;
  wire  _EVAL_651;
  wire  _EVAL_394;
  wire  _EVAL_357;
  wire  _EVAL_559;
  wire  _EVAL_263;
  wire  _EVAL_224;
  wire  _EVAL_545;
  wire  _EVAL_201;
  wire  _EVAL_426;
  wire  _EVAL_568;
  wire  _EVAL_514;
  wire  _EVAL_543;
  wire  _EVAL_491;
  wire  _EVAL_470;
  wire  _EVAL_123;
  wire [1:0] _EVAL_323;
  wire  _EVAL_297;
  wire  _EVAL_372;
  wire  _EVAL_235;
  wire  _EVAL_388;
  wire  _EVAL_446;
  wire  _EVAL_212;
  wire  _EVAL_335;
  wire [4:0] _EVAL_261;
  wire  _EVAL_329;
  wire  _EVAL_273;
  wire  _EVAL_195;
  wire  _EVAL_452;
  wire  _EVAL_239;
  wire  _EVAL_342;
  wire  _EVAL_39;
  wire  _EVAL_440;
  wire  _EVAL_383;
  wire  _EVAL_360;
  wire  _EVAL_247;
  wire  _EVAL_523;
  wire  _EVAL_647;
  wire  _EVAL_443;
  wire  _EVAL_389;
  wire [1:0] _EVAL_304;
  wire [1:0] _EVAL_34;
  wire  _EVAL_385;
  wire  _EVAL_554;
  wire  _EVAL_487;
  wire  _EVAL_121;
  wire  _EVAL_218;
  wire  _EVAL_352;
  wire  _EVAL_534;
  wire  _EVAL_489;
  wire  _EVAL_336;
  wire  _EVAL_318;
  wire  _EVAL_53;
  wire  _EVAL_322;
  wire  _EVAL_613;
  wire  _EVAL_625;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_43 = _EVAL_6 <= 3'h2;
  assign _EVAL_566 = _EVAL_26 & _EVAL_30;
  assign _EVAL_450 = _EVAL_32 & _EVAL_22;
  assign _EVAL_610 = _EVAL_566 | _EVAL_450;
  assign _EVAL_47 = _EVAL_180 + 32'h1;
  assign _EVAL_380 = _EVAL_24 ^ 32'h1800000;
  assign _EVAL_262 = {1'b0,$signed(_EVAL_380)};
  assign _EVAL_63 = _EVAL_21 ^ 32'h40000000;
  assign _EVAL_552 = {1'b0,$signed(_EVAL_63)};
  assign _EVAL_627 = $signed(_EVAL_552) & $signed(-33'sh2000);
  assign _EVAL_364 = $signed(_EVAL_627);
  assign _EVAL_606 = $signed(_EVAL_364) == $signed(33'sh0);
  assign _EVAL_519 = _EVAL_21 ^ 32'h80000000;
  assign _EVAL_391 = {1'b0,$signed(_EVAL_519)};
  assign _EVAL_420 = $signed(_EVAL_391) & $signed(-33'sh20000);
  assign _EVAL_361 = $signed(_EVAL_420);
  assign _EVAL_454 = $signed(_EVAL_361) == $signed(33'sh0);
  assign _EVAL_599 = _EVAL_606 | _EVAL_454;
  assign _EVAL_589 = _EVAL_21 ^ 32'h3000;
  assign _EVAL_467 = {1'b0,$signed(_EVAL_589)};
  assign _EVAL_138 = $signed(_EVAL_467) & $signed(-33'sh1000);
  assign _EVAL_289 = $signed(_EVAL_138);
  assign _EVAL_165 = $signed(_EVAL_289) == $signed(33'sh0);
  assign _EVAL_513 = _EVAL_599 | _EVAL_165;
  assign _EVAL_94 = _EVAL_21 ^ 32'hc000000;
  assign _EVAL_547 = {1'b0,$signed(_EVAL_94)};
  assign _EVAL_74 = $signed(_EVAL_547) & $signed(-33'sh4000000);
  assign _EVAL_573 = $signed(_EVAL_74);
  assign _EVAL_617 = $signed(_EVAL_573) == $signed(33'sh0);
  assign _EVAL_225 = _EVAL_513 | _EVAL_617;
  assign _EVAL_488 = _EVAL_21 ^ 32'h2000000;
  assign _EVAL_83 = {1'b0,$signed(_EVAL_488)};
  assign _EVAL_344 = $signed(_EVAL_83) & $signed(-33'sh10000);
  assign _EVAL_45 = $signed(_EVAL_344);
  assign _EVAL_564 = $signed(_EVAL_45) == $signed(33'sh0);
  assign _EVAL_652 = _EVAL_225 | _EVAL_564;
  assign _EVAL_624 = {1'b0,$signed(_EVAL_21)};
  assign _EVAL_193 = $signed(_EVAL_624) & $signed(-33'sh1000);
  assign _EVAL_245 = $signed(_EVAL_193);
  assign _EVAL_311 = $signed(_EVAL_245) == $signed(33'sh0);
  assign _EVAL_337 = _EVAL_652 | _EVAL_311;
  assign _EVAL_269 = _EVAL_21 ^ 32'h1800000;
  assign _EVAL_473 = {1'b0,$signed(_EVAL_269)};
  assign _EVAL_163 = $signed(_EVAL_473) & $signed(-33'sh8000);
  assign _EVAL_50 = $signed(_EVAL_163);
  assign _EVAL_279 = $signed(_EVAL_50) == $signed(33'sh0);
  assign _EVAL_81 = _EVAL_337 | _EVAL_279;
  assign _EVAL_607 = _EVAL_21 ^ 32'h1900000;
  assign _EVAL_609 = {1'b0,$signed(_EVAL_607)};
  assign _EVAL_343 = $signed(_EVAL_609) & $signed(-33'sh2000);
  assign _EVAL_286 = $signed(_EVAL_343);
  assign _EVAL_46 = $signed(_EVAL_286) == $signed(33'sh0);
  assign _EVAL_435 = _EVAL_81 | _EVAL_46;
  assign _EVAL_99 = _EVAL_21 ^ 32'h4000;
  assign _EVAL_649 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_338 = $signed(_EVAL_649) & $signed(-33'sh1000);
  assign _EVAL_405 = $signed(_EVAL_338);
  assign _EVAL_586 = $signed(_EVAL_405) == $signed(33'sh0);
  assign _EVAL_243 = _EVAL_435 | _EVAL_586;
  assign _EVAL_582 = _EVAL_29 == 3'h0;
  assign _EVAL_176 = 4'h6 == _EVAL_28;
  assign _EVAL_230 = _EVAL_582 ? _EVAL_176 : 1'h0;
  assign _EVAL_315 = _EVAL_374 == 5'h0;
  assign _EVAL_531 = _EVAL_15[2];
  assign _EVAL_618 = _EVAL_531 == 1'h0;
  assign _EVAL_126 = 23'hff << _EVAL_28;
  assign _EVAL_256 = _EVAL_126[7:0];
  assign _EVAL_61 = ~ _EVAL_256;
  assign _EVAL_472 = _EVAL_61[7:3];
  assign _EVAL_137 = _EVAL_374 - 5'h1;
  assign _EVAL_264 = _EVAL_630 == 5'h0;
  assign _EVAL_539 = _EVAL_7[0];
  assign _EVAL_55 = 23'hff << _EVAL_20;
  assign _EVAL_553 = _EVAL_55[7:0];
  assign _EVAL_232 = ~ _EVAL_553;
  assign _EVAL_451 = _EVAL_232[7:3];
  assign _EVAL_86 = _EVAL_630 - 5'h1;
  assign _EVAL_164 = _EVAL_33 == 3'h4;
  assign _EVAL_572 = _EVAL_28[1:0];
  assign _EVAL_386 = 4'h1 << _EVAL_572;
  assign _EVAL_87 = _EVAL_386[2:0];
  assign _EVAL_219 = _EVAL_87 | 3'h1;
  assign _EVAL_182 = _EVAL_219[1];
  assign _EVAL_37 = _EVAL_9 == 1'h0;
  assign _EVAL_128 = _EVAL_37 | _EVAL_5;
  assign _EVAL_144 = _EVAL_128 == 1'h0;
  assign _EVAL_325 = _EVAL_14 != 2'h2;
  assign _EVAL_69 = _EVAL_325 | _EVAL_5;
  assign _EVAL_400 = _EVAL_69 == 1'h0;
  assign _EVAL_387 = 23'hff << _EVAL_4;
  assign _EVAL_226 = _EVAL_387[7:0];
  assign _EVAL_643 = ~ _EVAL_226;
  assign _EVAL_490 = {{24'd0}, _EVAL_643};
  assign _EVAL_353 = _EVAL_21 & _EVAL_490;
  assign _EVAL_203 = _EVAL_25 ^ 32'h20000000;
  assign _EVAL_274 = {1'b0,$signed(_EVAL_203)};
  assign _EVAL_428 = $signed(_EVAL_274) & $signed(-33'sh2000);
  assign _EVAL_479 = $signed(_EVAL_428);
  assign _EVAL_597 = _EVAL_24 ^ 32'h1900000;
  assign _EVAL_481 = _EVAL_28 == _EVAL_116;
  assign _EVAL_197 = _EVAL_481 | _EVAL_5;
  assign _EVAL_258 = _EVAL_28 <= 4'h6;
  assign _EVAL_530 = _EVAL_24 ^ 32'h80000000;
  assign _EVAL_629 = {1'b0,$signed(_EVAL_530)};
  assign _EVAL_356 = $signed(_EVAL_629) & $signed(-33'sh20000);
  assign _EVAL_192 = $signed(_EVAL_356);
  assign _EVAL_35 = $signed(_EVAL_192) == $signed(33'sh0);
  assign _EVAL_500 = _EVAL_258 & _EVAL_35;
  assign _EVAL_359 = _EVAL_500 | _EVAL_5;
  assign _EVAL_275 = _EVAL_6 <= 3'h4;
  assign _EVAL_278 = _EVAL_275 | _EVAL_5;
  assign _EVAL_51 = _EVAL_384 == 5'h0;
  assign _EVAL_382 = _EVAL_51 == 1'h0;
  assign _EVAL_542 = _EVAL_30 & _EVAL_382;
  assign _EVAL_580 = _EVAL_219[2];
  assign _EVAL_48 = _EVAL_449 == 5'h0;
  assign _EVAL_561 = _EVAL_450 & _EVAL_48;
  assign _EVAL_72 = _EVAL_7[2];
  assign _EVAL_257 = _EVAL_7[1];
  assign _EVAL_70 = _EVAL_257 == 1'h0;
  assign _EVAL_312 = _EVAL_72 & _EVAL_70;
  assign _EVAL_108 = _EVAL_561 & _EVAL_312;
  assign _EVAL_213 = 2'h1 << _EVAL_19;
  assign _EVAL_581 = _EVAL_108 ? _EVAL_213 : 2'h0;
  assign _EVAL_308 = _EVAL_270 >> _EVAL_19;
  assign _EVAL_75 = _EVAL_4 <= 4'h6;
  assign _EVAL_558 = _EVAL_75 & _EVAL_454;
  assign _EVAL_68 = _EVAL_12 == 3'h0;
  assign _EVAL_299 = 3'h1 <= _EVAL_12;
  assign _EVAL_267 = _EVAL_68 | _EVAL_299;
  assign _EVAL_565 = _EVAL_33 == 3'h5;
  assign _EVAL_587 = _EVAL_18 & _EVAL_565;
  assign _EVAL_367 = 8'h1 << _EVAL_0;
  assign _EVAL_465 = _EVAL_15 == 3'h1;
  assign _EVAL_127 = _EVAL_7 == 3'h0;
  assign _EVAL_134 = _EVAL_22 & _EVAL_127;
  assign _EVAL_196 = ~ _EVAL_3;
  assign _EVAL_570 = _EVAL_196 == 8'h0;
  assign _EVAL_332 = _EVAL_570 | _EVAL_5;
  assign _EVAL_155 = _EVAL_332 == 1'h0;
  assign _EVAL_555 = _EVAL_6 != 3'h0;
  assign _EVAL_79 = _EVAL_555 | _EVAL_5;
  assign _EVAL_89 = _EVAL_79 == 1'h0;
  assign _EVAL_326 = _EVAL_33 == 3'h6;
  assign _EVAL_252 = _EVAL_18 & _EVAL_326;
  assign _EVAL_236 = _EVAL_24 ^ 32'h20000000;
  assign _EVAL_266 = {1'b0,$signed(_EVAL_236)};
  assign _EVAL_457 = _EVAL_25 ^ 32'h1800000;
  assign _EVAL_368 = _EVAL_28 >= 4'h3;
  assign _EVAL_616 = _EVAL_24[2];
  assign _EVAL_498 = _EVAL_580 & _EVAL_616;
  assign _EVAL_462 = _EVAL_368 | _EVAL_498;
  assign _EVAL_579 = _EVAL_24[1];
  assign _EVAL_307 = _EVAL_616 & _EVAL_579;
  assign _EVAL_430 = _EVAL_182 & _EVAL_307;
  assign _EVAL_503 = _EVAL_462 | _EVAL_430;
  assign _EVAL_438 = _EVAL_219[0];
  assign _EVAL_216 = _EVAL_24[0];
  assign _EVAL_591 = _EVAL_307 & _EVAL_216;
  assign _EVAL_244 = _EVAL_438 & _EVAL_591;
  assign _EVAL_76 = _EVAL_503 | _EVAL_244;
  assign _EVAL_418 = _EVAL_216 == 1'h0;
  assign _EVAL_115 = _EVAL_307 & _EVAL_418;
  assign _EVAL_396 = _EVAL_438 & _EVAL_115;
  assign _EVAL_588 = _EVAL_503 | _EVAL_396;
  assign _EVAL_363 = _EVAL_579 == 1'h0;
  assign _EVAL_480 = _EVAL_616 & _EVAL_363;
  assign _EVAL_294 = _EVAL_182 & _EVAL_480;
  assign _EVAL_296 = _EVAL_462 | _EVAL_294;
  assign _EVAL_303 = _EVAL_480 & _EVAL_216;
  assign _EVAL_634 = _EVAL_438 & _EVAL_303;
  assign _EVAL_575 = _EVAL_296 | _EVAL_634;
  assign _EVAL_324 = _EVAL_480 & _EVAL_418;
  assign _EVAL_611 = _EVAL_438 & _EVAL_324;
  assign _EVAL_268 = _EVAL_296 | _EVAL_611;
  assign _EVAL_522 = _EVAL_616 == 1'h0;
  assign _EVAL_527 = _EVAL_580 & _EVAL_522;
  assign _EVAL_183 = _EVAL_368 | _EVAL_527;
  assign _EVAL_548 = _EVAL_522 & _EVAL_579;
  assign _EVAL_120 = _EVAL_182 & _EVAL_548;
  assign _EVAL_439 = _EVAL_183 | _EVAL_120;
  assign _EVAL_442 = _EVAL_548 & _EVAL_216;
  assign _EVAL_246 = _EVAL_438 & _EVAL_442;
  assign _EVAL_210 = _EVAL_439 | _EVAL_246;
  assign _EVAL_97 = _EVAL_548 & _EVAL_418;
  assign _EVAL_306 = _EVAL_438 & _EVAL_97;
  assign _EVAL_166 = _EVAL_439 | _EVAL_306;
  assign _EVAL_365 = _EVAL_522 & _EVAL_363;
  assign _EVAL_233 = _EVAL_182 & _EVAL_365;
  assign _EVAL_549 = _EVAL_183 | _EVAL_233;
  assign _EVAL_77 = _EVAL_365 & _EVAL_216;
  assign _EVAL_596 = _EVAL_438 & _EVAL_77;
  assign _EVAL_254 = _EVAL_549 | _EVAL_596;
  assign _EVAL_189 = _EVAL_365 & _EVAL_418;
  assign _EVAL_301 = _EVAL_438 & _EVAL_189;
  assign _EVAL_122 = _EVAL_549 | _EVAL_301;
  assign _EVAL_119 = {_EVAL_76,_EVAL_588,_EVAL_575,_EVAL_268,_EVAL_210,_EVAL_166,_EVAL_254,_EVAL_122};
  assign _EVAL_205 = _EVAL_3 == _EVAL_119;
  assign _EVAL_401 = _EVAL_205 | _EVAL_5;
  assign _EVAL_234 = _EVAL_24 ^ 32'h3000;
  assign _EVAL_407 = {1'b0,$signed(_EVAL_234)};
  assign _EVAL_64 = $signed(_EVAL_407) & $signed(-33'sh1000);
  assign _EVAL_349 = $signed(_EVAL_64);
  assign _EVAL_569 = $signed(_EVAL_349) == $signed(33'sh0);
  assign _EVAL_619 = _EVAL_24 ^ 32'hc000000;
  assign _EVAL_172 = {1'b0,$signed(_EVAL_619)};
  assign _EVAL_355 = $signed(_EVAL_172) & $signed(-33'sh4000000);
  assign _EVAL_376 = $signed(_EVAL_355);
  assign _EVAL_71 = $signed(_EVAL_376) == $signed(33'sh0);
  assign _EVAL_421 = _EVAL_569 | _EVAL_71;
  assign _EVAL_82 = _EVAL_24 ^ 32'h2000000;
  assign _EVAL_277 = {1'b0,$signed(_EVAL_82)};
  assign _EVAL_358 = $signed(_EVAL_277) & $signed(-33'sh10000);
  assign _EVAL_466 = $signed(_EVAL_358);
  assign _EVAL_577 = $signed(_EVAL_466) == $signed(33'sh0);
  assign _EVAL_574 = _EVAL_421 | _EVAL_577;
  assign _EVAL_259 = _EVAL_300 == 5'h0;
  assign _EVAL_492 = _EVAL_450 & _EVAL_259;
  assign _EVAL_313 = _EVAL_7 == 3'h6;
  assign _EVAL_170 = _EVAL_313 == 1'h0;
  assign _EVAL_477 = _EVAL_492 & _EVAL_170;
  assign _EVAL_283 = _EVAL_477 ? _EVAL_367 : 8'h0;
  assign _EVAL_327 = _EVAL_21 ^ 32'h20000000;
  assign _EVAL_536 = {1'b0,$signed(_EVAL_327)};
  assign _EVAL_153 = $signed(_EVAL_536) & $signed(-33'sh2000);
  assign _EVAL_362 = $signed(_EVAL_153);
  assign _EVAL_373 = $signed(_EVAL_362) == $signed(33'sh0);
  assign _EVAL_132 = _EVAL_243 | _EVAL_373;
  assign _EVAL_600 = 3'h1 <= _EVAL_29;
  assign _EVAL_217 = _EVAL_582 | _EVAL_600;
  assign _EVAL_455 = _EVAL_20 >= 4'h3;
  assign _EVAL_96 = _EVAL_2 <= 2'h2;
  assign _EVAL_145 = _EVAL_96 | _EVAL_5;
  assign _EVAL_517 = _EVAL_566 & _EVAL_51;
  assign _EVAL_404 = _EVAL_25 ^ 32'h2000000;
  assign _EVAL_637 = {1'b0,$signed(_EVAL_404)};
  assign _EVAL_130 = $signed(_EVAL_637) & $signed(-33'sh10000);
  assign _EVAL_80 = $signed(_EVAL_130);
  assign _EVAL_228 = {1'b0,$signed(_EVAL_457)};
  assign _EVAL_395 = $signed(_EVAL_228) & $signed(-33'sh8000);
  assign _EVAL_221 = plusarg_reader_out == 32'h0;
  assign _EVAL_408 = _EVAL_8 <= 3'h5;
  assign _EVAL_162 = _EVAL_408 | _EVAL_5;
  assign _EVAL_478 = _EVAL_162 == 1'h0;
  assign _EVAL_141 = $signed(_EVAL_395);
  assign _EVAL_124 = _EVAL_28 <= 4'h8;
  assign _EVAL_114 = _EVAL_353 == 32'h0;
  assign _EVAL_642 = _EVAL_114 | _EVAL_5;
  assign _EVAL_285 = _EVAL_642 == 1'h0;
  assign _EVAL_49 = _EVAL_15 == _EVAL_348;
  assign _EVAL_463 = _EVAL_49 | _EVAL_5;
  assign _EVAL_171 = _EVAL_463 == 1'h0;
  assign _EVAL_567 = _EVAL_278 == 1'h0;
  assign _EVAL_528 = _EVAL_14 <= 2'h2;
  assign _EVAL_626 = _EVAL_528 | _EVAL_5;
  assign _EVAL_135 = _EVAL_626 == 1'h0;
  assign _EVAL_281 = $signed(_EVAL_80) == $signed(33'sh0);
  assign _EVAL_330 = _EVAL_14 == 2'h0;
  assign _EVAL_88 = _EVAL_384 - 5'h1;
  assign _EVAL_621 = _EVAL_24 == _EVAL_214;
  assign _EVAL_511 = _EVAL_621 | _EVAL_5;
  assign _EVAL_508 = _EVAL_511 == 1'h0;
  assign _EVAL_341 = _EVAL_7 == 3'h5;
  assign _EVAL_131 = _EVAL_22 & _EVAL_341;
  assign _EVAL_650 = _EVAL_1 & _EVAL_18;
  assign _EVAL_631 = _EVAL_535 == 5'h0;
  assign _EVAL_406 = _EVAL_33[0];
  assign _EVAL_340 = _EVAL_643[7:3];
  assign _EVAL_354 = _EVAL_535 - 5'h1;
  assign _EVAL_571 = _EVAL_25 == _EVAL_431;
  assign _EVAL_328 = _EVAL_23 == 1'h0;
  assign _EVAL_100 = _EVAL_328 | _EVAL_5;
  assign _EVAL_102 = _EVAL_100 == 1'h0;
  assign _EVAL_103 = _EVAL_132 | _EVAL_5;
  assign _EVAL_347 = ~ _EVAL_119;
  assign _EVAL_392 = _EVAL_6 <= 3'h3;
  assign _EVAL_215 = _EVAL_392 | _EVAL_5;
  assign _EVAL_298 = _EVAL_215 == 1'h0;
  assign _EVAL_510 = _EVAL_33 == 3'h7;
  assign _EVAL_211 = _EVAL_18 & _EVAL_510;
  assign _EVAL_471 = _EVAL_581 | _EVAL_270;
  assign _EVAL_550 = _EVAL_0 == 3'h0;
  assign _EVAL_422 = 3'h1 <= _EVAL_0;
  assign _EVAL_370 = _EVAL_550 | _EVAL_422;
  assign _EVAL_154 = _EVAL_370 | _EVAL_5;
  assign _EVAL_414 = {1'b0,$signed(_EVAL_24)};
  assign _EVAL_429 = $signed(_EVAL_414) & $signed(-33'sh5000);
  assign _EVAL_302 = $signed(_EVAL_429);
  assign _EVAL_556 = $signed(_EVAL_302) == $signed(33'sh0);
  assign _EVAL_181 = _EVAL_574 | _EVAL_556;
  assign _EVAL_417 = $signed(_EVAL_262) & $signed(-33'sh8000);
  assign _EVAL_93 = $signed(_EVAL_417);
  assign _EVAL_411 = $signed(_EVAL_93) == $signed(33'sh0);
  assign _EVAL_85 = _EVAL_181 | _EVAL_411;
  assign _EVAL_351 = _EVAL_24 ^ 32'h40000000;
  assign _EVAL_184 = {1'b0,$signed(_EVAL_351)};
  assign _EVAL_419 = $signed(_EVAL_184) & $signed(-33'sh2000);
  assign _EVAL_653 = $signed(_EVAL_419);
  assign _EVAL_436 = $signed(_EVAL_653) == $signed(33'sh0);
  assign _EVAL_398 = _EVAL_436 | _EVAL_35;
  assign _EVAL_292 = _EVAL_398 | _EVAL_71;
  assign _EVAL_635 = _EVAL_292 | _EVAL_577;
  assign _EVAL_540 = _EVAL_635 | _EVAL_556;
  assign _EVAL_515 = _EVAL_540 | _EVAL_411;
  assign _EVAL_161 = {1'b0,$signed(_EVAL_597)};
  assign _EVAL_187 = $signed(_EVAL_161) & $signed(-33'sh2000);
  assign _EVAL_65 = $signed(_EVAL_187);
  assign _EVAL_106 = $signed(_EVAL_65) == $signed(33'sh0);
  assign _EVAL_57 = _EVAL_515 | _EVAL_106;
  assign _EVAL_142 = $signed(_EVAL_266) & $signed(-33'sh2000);
  assign _EVAL_537 = $signed(_EVAL_142);
  assign _EVAL_272 = $signed(_EVAL_537) == $signed(33'sh0);
  assign _EVAL_255 = _EVAL_57 | _EVAL_272;
  assign _EVAL_375 = _EVAL_12 == _EVAL_320;
  assign _EVAL_484 = _EVAL_145 == 1'h0;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_25)};
  assign _EVAL_524 = $signed(_EVAL_113) & $signed(-33'sh1000);
  assign _EVAL_223 = _EVAL_23 == _EVAL_56;
  assign _EVAL_448 = _EVAL_223 | _EVAL_5;
  assign _EVAL_546 = _EVAL_448 == 1'h0;
  assign _EVAL_319 = _EVAL_15 == 3'h3;
  assign _EVAL_445 = _EVAL_623 != 8'h0;
  assign _EVAL_101 = _EVAL_592 == 5'h0;
  assign _EVAL_251 = _EVAL_101 == 1'h0;
  assign _EVAL_282 = _EVAL_15 == 3'h0;
  assign _EVAL_147 = _EVAL_30 & _EVAL_282;
  assign _EVAL_622 = _EVAL_10 & _EVAL_11;
  assign _EVAL_146 = 2'h1 << _EVAL_13;
  assign _EVAL_437 = _EVAL_622 ? _EVAL_146 : 2'h0;
  assign _EVAL_424 = ~ _EVAL_437;
  assign _EVAL_159 = _EVAL_30 & _EVAL_465;
  assign _EVAL_453 = _EVAL_258 & _EVAL_255;
  assign _EVAL_209 = _EVAL_124 & _EVAL_569;
  assign _EVAL_276 = _EVAL_453 | _EVAL_209;
  assign _EVAL_167 = _EVAL_276 | _EVAL_5;
  assign _EVAL_434 = ~ _EVAL_283;
  assign _EVAL_645 = _EVAL_631 == 1'h0;
  assign _EVAL_190 = _EVAL_375 | _EVAL_5;
  assign _EVAL_333 = _EVAL_190 == 1'h0;
  assign _EVAL_194 = _EVAL_25 & 32'h3f;
  assign _EVAL_521 = _EVAL_194 == 32'h0;
  assign _EVAL_321 = _EVAL_521 | _EVAL_5;
  assign _EVAL_111 = _EVAL_8 == 3'h0;
  assign _EVAL_107 = _EVAL_623 >> _EVAL_29;
  assign _EVAL_416 = _EVAL_107[0];
  assign _EVAL_73 = _EVAL_416 == 1'h0;
  assign _EVAL_432 = _EVAL_73 | _EVAL_5;
  assign _EVAL_632 = _EVAL_432 == 1'h0;
  assign _EVAL_494 = _EVAL_4 == _EVAL_562;
  assign _EVAL_242 = _EVAL_16 == 1'h0;
  assign _EVAL_310 = _EVAL_242 | _EVAL_5;
  assign _EVAL_177 = _EVAL_310 == 1'h0;
  assign _EVAL_284 = {{24'd0}, _EVAL_61};
  assign _EVAL_633 = _EVAL_180 < plusarg_reader_out;
  assign _EVAL_227 = _EVAL_25 ^ 32'h40000000;
  assign _EVAL_560 = {1'b0,$signed(_EVAL_227)};
  assign _EVAL_316 = $signed(_EVAL_560) & $signed(-33'sh2000);
  assign _EVAL_496 = $signed(_EVAL_316);
  assign _EVAL_648 = _EVAL_2 == _EVAL_483;
  assign _EVAL_174 = _EVAL_648 | _EVAL_5;
  assign _EVAL_602 = _EVAL_174 == 1'h0;
  assign _EVAL_148 = $signed(_EVAL_496) == $signed(33'sh0);
  assign _EVAL_638 = _EVAL_25 ^ 32'h80000000;
  assign _EVAL_309 = {1'b0,$signed(_EVAL_638)};
  assign _EVAL_644 = $signed(_EVAL_309) & $signed(-33'sh20000);
  assign _EVAL_497 = $signed(_EVAL_644);
  assign _EVAL_188 = $signed(_EVAL_497) == $signed(33'sh0);
  assign _EVAL_157 = _EVAL_148 | _EVAL_188;
  assign _EVAL_533 = _EVAL_25 ^ 32'h3000;
  assign _EVAL_468 = {1'b0,$signed(_EVAL_533)};
  assign _EVAL_92 = $signed(_EVAL_468) & $signed(-33'sh1000);
  assign _EVAL_204 = $signed(_EVAL_92);
  assign _EVAL_393 = $signed(_EVAL_204) == $signed(33'sh0);
  assign _EVAL_91 = _EVAL_157 | _EVAL_393;
  assign _EVAL_288 = _EVAL_25 ^ 32'hc000000;
  assign _EVAL_425 = {1'b0,$signed(_EVAL_288)};
  assign _EVAL_41 = $signed(_EVAL_425) & $signed(-33'sh4000000);
  assign _EVAL_379 = $signed(_EVAL_41);
  assign _EVAL_231 = $signed(_EVAL_379) == $signed(33'sh0);
  assign _EVAL_200 = _EVAL_91 | _EVAL_231;
  assign _EVAL_493 = _EVAL_200 | _EVAL_281;
  assign _EVAL_293 = $signed(_EVAL_524);
  assign _EVAL_377 = $signed(_EVAL_293) == $signed(33'sh0);
  assign _EVAL_186 = _EVAL_493 | _EVAL_377;
  assign _EVAL_608 = $signed(_EVAL_141) == $signed(33'sh0);
  assign _EVAL_604 = _EVAL_186 | _EVAL_608;
  assign _EVAL_636 = _EVAL_25 ^ 32'h1900000;
  assign _EVAL_280 = {1'b0,$signed(_EVAL_636)};
  assign _EVAL_504 = $signed(_EVAL_280) & $signed(-33'sh2000);
  assign _EVAL_95 = $signed(_EVAL_504);
  assign _EVAL_175 = $signed(_EVAL_95) == $signed(33'sh0);
  assign _EVAL_265 = _EVAL_604 | _EVAL_175;
  assign _EVAL_149 = _EVAL_25 ^ 32'h4000;
  assign _EVAL_249 = {1'b0,$signed(_EVAL_149)};
  assign _EVAL_640 = $signed(_EVAL_249) & $signed(-33'sh1000);
  assign _EVAL_495 = $signed(_EVAL_640);
  assign _EVAL_485 = $signed(_EVAL_495) == $signed(33'sh0);
  assign _EVAL_207 = _EVAL_265 | _EVAL_485;
  assign _EVAL_104 = $signed(_EVAL_479) == $signed(33'sh0);
  assign _EVAL_646 = _EVAL_207 | _EVAL_104;
  assign _EVAL_461 = _EVAL_646 | _EVAL_5;
  assign _EVAL_287 = _EVAL_21 == _EVAL_44;
  assign _EVAL_331 = _EVAL_8 <= 3'h2;
  assign _EVAL_603 = _EVAL_331 | _EVAL_5;
  assign _EVAL_84 = _EVAL_603 == 1'h0;
  assign _EVAL_169 = _EVAL_33 == _EVAL_598;
  assign _EVAL_427 = _EVAL_308[0];
  assign _EVAL_525 = _EVAL_427 == 1'h0;
  assign _EVAL_291 = _EVAL_525 | _EVAL_5;
  assign _EVAL_509 = _EVAL_291 == 1'h0;
  assign _EVAL_40 = _EVAL_29 == _EVAL_433;
  assign _EVAL_66 = _EVAL_40 | _EVAL_5;
  assign _EVAL_62 = _EVAL_15 == 3'h7;
  assign _EVAL_601 = _EVAL_30 & _EVAL_62;
  assign _EVAL_423 = _EVAL_4 >= 4'h3;
  assign _EVAL_42 = _EVAL_15 == 3'h6;
  assign _EVAL_518 = _EVAL_33 == 3'h2;
  assign _EVAL_641 = _EVAL_300 - 5'h1;
  assign _EVAL_551 = _EVAL_423 | _EVAL_5;
  assign _EVAL_512 = _EVAL_551 == 1'h0;
  assign _EVAL_173 = _EVAL_267 | _EVAL_5;
  assign _EVAL_334 = _EVAL_445 == 1'h0;
  assign _EVAL_520 = _EVAL_334 | _EVAL_221;
  assign _EVAL_505 = _EVAL_520 | _EVAL_633;
  assign _EVAL_459 = _EVAL_505 | _EVAL_5;
  assign _EVAL_526 = _EVAL_459 == 1'h0;
  assign _EVAL_317 = _EVAL_0 == _EVAL_168;
  assign _EVAL_378 = _EVAL_317 | _EVAL_5;
  assign _EVAL_229 = _EVAL_359 == 1'h0;
  assign _EVAL_516 = _EVAL_287 | _EVAL_5;
  assign _EVAL_152 = _EVAL_17 == 1'h0;
  assign _EVAL_538 = _EVAL_15 == 3'h4;
  assign _EVAL_314 = _EVAL_30 & _EVAL_538;
  assign _EVAL_198 = _EVAL_330 | _EVAL_5;
  assign _EVAL_476 = _EVAL_566 & _EVAL_315;
  assign _EVAL_290 = 8'h1 << _EVAL_29;
  assign _EVAL_615 = _EVAL_476 ? _EVAL_290 : 8'h0;
  assign _EVAL_237 = _EVAL_623 | _EVAL_615;
  assign _EVAL_143 = _EVAL_237 & _EVAL_434;
  assign _EVAL_410 = _EVAL_321 == 1'h0;
  assign _EVAL_222 = _EVAL_15 == 3'h2;
  assign _EVAL_199 = _EVAL_615 != _EVAL_283;
  assign _EVAL_501 = _EVAL_615 != 8'h0;
  assign _EVAL_241 = _EVAL_501 == 1'h0;
  assign _EVAL_160 = _EVAL_199 | _EVAL_241;
  assign _EVAL_532 = _EVAL_160 | _EVAL_5;
  assign _EVAL_585 = _EVAL_532 == 1'h0;
  assign _EVAL_506 = _EVAL_615 | _EVAL_623;
  assign _EVAL_60 = _EVAL_506 >> _EVAL_0;
  assign _EVAL_139 = _EVAL_60[0];
  assign _EVAL_67 = _EVAL_139 | _EVAL_5;
  assign _EVAL_178 = _EVAL_67 == 1'h0;
  assign _EVAL_253 = _EVAL_217 | _EVAL_5;
  assign _EVAL_620 = _EVAL_197 == 1'h0;
  assign _EVAL_151 = _EVAL_7 == _EVAL_628;
  assign _EVAL_595 = _EVAL_151 | _EVAL_5;
  assign _EVAL_412 = _EVAL_595 == 1'h0;
  assign _EVAL_38 = _EVAL_230 | _EVAL_5;
  assign _EVAL_58 = _EVAL_38 == 1'h0;
  assign _EVAL_594 = _EVAL_20 == _EVAL_639;
  assign _EVAL_305 = _EVAL_594 | _EVAL_5;
  assign _EVAL_369 = _EVAL_305 == 1'h0;
  assign _EVAL_415 = _EVAL_378 == 1'h0;
  assign _EVAL_413 = _EVAL_15 == 3'h5;
  assign _EVAL_447 = _EVAL_30 & _EVAL_413;
  assign _EVAL_475 = _EVAL_7 == 3'h2;
  assign _EVAL_563 = _EVAL_22 & _EVAL_475;
  assign _EVAL_179 = _EVAL_449 - 5'h1;
  assign _EVAL_191 = _EVAL_7 <= 3'h6;
  assign _EVAL_590 = _EVAL_191 | _EVAL_5;
  assign _EVAL_469 = _EVAL_590 == 1'h0;
  assign _EVAL_271 = _EVAL_30 & _EVAL_222;
  assign _EVAL_339 = _EVAL_18 & _EVAL_164;
  assign _EVAL_125 = _EVAL_328 | _EVAL_16;
  assign _EVAL_409 = _EVAL_125 | _EVAL_5;
  assign _EVAL_105 = _EVAL_409 == 1'h0;
  assign _EVAL_240 = _EVAL_8 == _EVAL_150;
  assign _EVAL_456 = _EVAL_240 | _EVAL_5;
  assign _EVAL_583 = _EVAL_456 == 1'h0;
  assign _EVAL_371 = _EVAL_14 == _EVAL_220;
  assign _EVAL_36 = _EVAL_371 | _EVAL_5;
  assign _EVAL_593 = _EVAL_36 == 1'h0;
  assign _EVAL_52 = _EVAL_558 | _EVAL_5;
  assign _EVAL_129 = _EVAL_52 == 1'h0;
  assign _EVAL_458 = _EVAL_22 & _EVAL_313;
  assign _EVAL_614 = _EVAL_650 & _EVAL_631;
  assign _EVAL_444 = _EVAL_167 == 1'h0;
  assign _EVAL_460 = _EVAL_24 & _EVAL_284;
  assign _EVAL_499 = _EVAL_460 == 32'h0;
  assign _EVAL_578 = _EVAL_499 | _EVAL_5;
  assign _EVAL_238 = _EVAL_33 == 3'h1;
  assign _EVAL_295 = _EVAL_18 & _EVAL_238;
  assign _EVAL_136 = _EVAL_6 == 3'h0;
  assign _EVAL_112 = _EVAL_136 | _EVAL_5;
  assign _EVAL_185 = _EVAL_112 == 1'h0;
  assign _EVAL_397 = _EVAL_33 == 3'h0;
  assign _EVAL_441 = _EVAL_18 & _EVAL_397;
  assign _EVAL_557 = _EVAL_3 & _EVAL_347;
  assign _EVAL_346 = _EVAL_557 == 8'h0;
  assign _EVAL_208 = _EVAL_346 | _EVAL_5;
  assign _EVAL_117 = _EVAL_43 | _EVAL_5;
  assign _EVAL_133 = _EVAL_28 <= 4'h2;
  assign _EVAL_78 = _EVAL_85 | _EVAL_106;
  assign _EVAL_366 = _EVAL_78 | _EVAL_272;
  assign _EVAL_98 = _EVAL_133 & _EVAL_366;
  assign _EVAL_474 = _EVAL_98 | _EVAL_5;
  assign _EVAL_541 = _EVAL_450 & _EVAL_264;
  assign _EVAL_464 = _EVAL_19 == _EVAL_118;
  assign _EVAL_486 = _EVAL_516 == 1'h0;
  assign _EVAL_59 = _EVAL_18 & _EVAL_645;
  assign _EVAL_206 = _EVAL_464 | _EVAL_5;
  assign _EVAL_651 = _EVAL_455 | _EVAL_5;
  assign _EVAL_394 = _EVAL_6 == _EVAL_502;
  assign _EVAL_357 = _EVAL_394 | _EVAL_5;
  assign _EVAL_559 = _EVAL_357 == 1'h0;
  assign _EVAL_263 = _EVAL_206 == 1'h0;
  assign _EVAL_224 = _EVAL_154 == 1'h0;
  assign _EVAL_545 = _EVAL_173 == 1'h0;
  assign _EVAL_201 = _EVAL_571 | _EVAL_5;
  assign _EVAL_426 = _EVAL_201 == 1'h0;
  assign _EVAL_568 = 4'h6 == _EVAL_4;
  assign _EVAL_514 = _EVAL_68 ? _EVAL_568 : 1'h0;
  assign _EVAL_543 = _EVAL_514 | _EVAL_5;
  assign _EVAL_491 = _EVAL_543 == 1'h0;
  assign _EVAL_470 = _EVAL_198 == 1'h0;
  assign _EVAL_123 = _EVAL_474 == 1'h0;
  assign _EVAL_323 = _EVAL_471 >> _EVAL_13;
  assign _EVAL_297 = _EVAL_651 == 1'h0;
  assign _EVAL_372 = _EVAL_152 | _EVAL_5;
  assign _EVAL_235 = _EVAL_323[0];
  assign _EVAL_388 = _EVAL_494 | _EVAL_5;
  assign _EVAL_446 = _EVAL_388 == 1'h0;
  assign _EVAL_212 = _EVAL_117 == 1'h0;
  assign _EVAL_335 = _EVAL_31 & _EVAL_251;
  assign _EVAL_261 = _EVAL_592 - 5'h1;
  assign _EVAL_329 = _EVAL_209 | _EVAL_5;
  assign _EVAL_273 = _EVAL_111 | _EVAL_5;
  assign _EVAL_195 = _EVAL_273 == 1'h0;
  assign _EVAL_452 = _EVAL_401 == 1'h0;
  assign _EVAL_239 = _EVAL_103 == 1'h0;
  assign _EVAL_342 = _EVAL_368 | _EVAL_5;
  assign _EVAL_39 = _EVAL_342 == 1'h0;
  assign _EVAL_440 = _EVAL_169 | _EVAL_5;
  assign _EVAL_383 = _EVAL_440 == 1'h0;
  assign _EVAL_360 = _EVAL_578 == 1'h0;
  assign _EVAL_247 = _EVAL_372 == 1'h0;
  assign _EVAL_523 = _EVAL_208 == 1'h0;
  assign _EVAL_647 = _EVAL_7 == 3'h4;
  assign _EVAL_443 = _EVAL_22 & _EVAL_647;
  assign _EVAL_389 = _EVAL_7 == 3'h1;
  assign _EVAL_304 = _EVAL_270 | _EVAL_581;
  assign _EVAL_34 = _EVAL_304 & _EVAL_424;
  assign _EVAL_385 = _EVAL_22 & _EVAL_389;
  assign _EVAL_554 = _EVAL_264 == 1'h0;
  assign _EVAL_487 = _EVAL_329 == 1'h0;
  assign _EVAL_121 = _EVAL_235 | _EVAL_5;
  assign _EVAL_218 = _EVAL_121 == 1'h0;
  assign _EVAL_352 = _EVAL_66 == 1'h0;
  assign _EVAL_534 = _EVAL_30 & _EVAL_319;
  assign _EVAL_489 = _EVAL_30 & _EVAL_42;
  assign _EVAL_336 = _EVAL_27 & _EVAL_31;
  assign _EVAL_318 = _EVAL_461 == 1'h0;
  assign _EVAL_53 = _EVAL_18 & _EVAL_518;
  assign _EVAL_322 = _EVAL_22 & _EVAL_554;
  assign _EVAL_613 = _EVAL_336 & _EVAL_101;
  assign _EVAL_625 = _EVAL_253 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_44 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_56 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_116 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_118 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_150 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_168 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_180 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_214 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_220 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_270 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_300 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_320 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_348 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_374 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_384 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_431 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_433 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_449 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_483 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_502 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_535 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_562 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_592 = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_598 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_623 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_628 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_630 = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_639 = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_614) begin
      _EVAL_44 <= _EVAL_21;
    end
    if (_EVAL_541) begin
      _EVAL_56 <= _EVAL_23;
    end
    if (_EVAL_517) begin
      _EVAL_116 <= _EVAL_28;
    end
    if (_EVAL_541) begin
      _EVAL_118 <= _EVAL_19;
    end
    if (_EVAL_614) begin
      _EVAL_150 <= _EVAL_8;
    end
    if (_EVAL_541) begin
      _EVAL_168 <= _EVAL_0;
    end
    if (_EVAL_5) begin
      _EVAL_180 <= 32'h0;
    end else begin
      if (_EVAL_610) begin
        _EVAL_180 <= 32'h0;
      end else begin
        _EVAL_180 <= _EVAL_47;
      end
    end
    if (_EVAL_517) begin
      _EVAL_214 <= _EVAL_24;
    end
    if (_EVAL_541) begin
      _EVAL_220 <= _EVAL_14;
    end
    if (_EVAL_5) begin
      _EVAL_270 <= 2'h0;
    end else begin
      _EVAL_270 <= _EVAL_34;
    end
    if (_EVAL_5) begin
      _EVAL_300 <= 5'h0;
    end else begin
      if (_EVAL_450) begin
        if (_EVAL_259) begin
          if (_EVAL_539) begin
            _EVAL_300 <= _EVAL_451;
          end else begin
            _EVAL_300 <= 5'h0;
          end
        end else begin
          _EVAL_300 <= _EVAL_641;
        end
      end
    end
    if (_EVAL_614) begin
      _EVAL_320 <= _EVAL_12;
    end
    if (_EVAL_517) begin
      _EVAL_348 <= _EVAL_15;
    end
    if (_EVAL_5) begin
      _EVAL_374 <= 5'h0;
    end else begin
      if (_EVAL_566) begin
        if (_EVAL_315) begin
          if (_EVAL_618) begin
            _EVAL_374 <= _EVAL_472;
          end else begin
            _EVAL_374 <= 5'h0;
          end
        end else begin
          _EVAL_374 <= _EVAL_137;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_384 <= 5'h0;
    end else begin
      if (_EVAL_566) begin
        if (_EVAL_51) begin
          if (_EVAL_618) begin
            _EVAL_384 <= _EVAL_472;
          end else begin
            _EVAL_384 <= 5'h0;
          end
        end else begin
          _EVAL_384 <= _EVAL_88;
        end
      end
    end
    if (_EVAL_613) begin
      _EVAL_431 <= _EVAL_25;
    end
    if (_EVAL_517) begin
      _EVAL_433 <= _EVAL_29;
    end
    if (_EVAL_5) begin
      _EVAL_449 <= 5'h0;
    end else begin
      if (_EVAL_450) begin
        if (_EVAL_48) begin
          if (_EVAL_539) begin
            _EVAL_449 <= _EVAL_451;
          end else begin
            _EVAL_449 <= 5'h0;
          end
        end else begin
          _EVAL_449 <= _EVAL_179;
        end
      end
    end
    if (_EVAL_613) begin
      _EVAL_483 <= _EVAL_2;
    end
    if (_EVAL_517) begin
      _EVAL_502 <= _EVAL_6;
    end
    if (_EVAL_5) begin
      _EVAL_535 <= 5'h0;
    end else begin
      if (_EVAL_650) begin
        if (_EVAL_631) begin
          if (_EVAL_406) begin
            _EVAL_535 <= _EVAL_340;
          end else begin
            _EVAL_535 <= 5'h0;
          end
        end else begin
          _EVAL_535 <= _EVAL_354;
        end
      end
    end
    if (_EVAL_614) begin
      _EVAL_562 <= _EVAL_4;
    end
    if (_EVAL_5) begin
      _EVAL_592 <= 5'h0;
    end else begin
      if (_EVAL_336) begin
        if (_EVAL_101) begin
          _EVAL_592 <= 5'h0;
        end else begin
          _EVAL_592 <= _EVAL_261;
        end
      end
    end
    if (_EVAL_614) begin
      _EVAL_598 <= _EVAL_33;
    end
    if (_EVAL_5) begin
      _EVAL_623 <= 8'h0;
    end else begin
      _EVAL_623 <= _EVAL_143;
    end
    if (_EVAL_541) begin
      _EVAL_628 <= _EVAL_7;
    end
    if (_EVAL_5) begin
      _EVAL_630 <= 5'h0;
    end else begin
      if (_EVAL_450) begin
        if (_EVAL_264) begin
          if (_EVAL_539) begin
            _EVAL_630 <= _EVAL_451;
          end else begin
            _EVAL_630 <= 5'h0;
          end
        end else begin
          _EVAL_630 <= _EVAL_86;
        end
      end
    end
    if (_EVAL_541) begin
      _EVAL_639 <= _EVAL_20;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f7d2c76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccd725b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_383) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4179d4a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_567) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(507622a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_476 & _EVAL_632) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db8e8082)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94aa23ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(156b75a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ade4bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d651ae56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_523) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2875e6f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_400) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6431c6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(627a24e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_593) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb365ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f496c62c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_509) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f30e073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c5e032f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b9bc326)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6494ae03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83eb60a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2617b1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71c36f0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(647df33a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91728e2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_512) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8ffe85f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d388d4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30ba0ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38c791a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_410) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c228535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_622 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88839c49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_415) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91d2169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88556d5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(439d09fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9cc1ff5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8422d0fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd43360a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(877288e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9278f1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5d2e4d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_410) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdd9a8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_426) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_491) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(268f81ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_491) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_369) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4081ed60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f73908b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6108dc56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_567) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b0542c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ec1106)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_415) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e31a1e38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_585) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20d57402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e674439)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f36aa69b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db950160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_400) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2ec6c0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_593) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_512) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0b99621)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_487) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6e857f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e97dcb14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_622 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_333) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a46f68a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_512) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47d176d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8360dd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(356f40c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_333) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_484) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b949edda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_478) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c332ab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b0c0066)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bab97bbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(626324ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa49717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_508) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2d0645f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef00079c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc9d529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e5dc7e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64023f80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_469) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ed8ef28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_486) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70154fff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_512) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_620) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e9c2e54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cce5eb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8bc8953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f41173)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c160252)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_478) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59e3e26d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6dc2d89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_620) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9aa4eb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_583) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_523) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d1e376)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6bd9ed1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfc6ae59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d80c12e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cda701b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b13e0c49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_559) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_512) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94217273)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f852646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_478) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(850ad109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6477472)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_369) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39510f2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_491) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_546) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_486) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_469) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_400) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca6f9327)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_476 & _EVAL_632) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20a4e0e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_559) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aec4d13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_602) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18eb0076)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ecdf402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c499b618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5667e3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9384867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9e4e52b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_484) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_512) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e891973c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_512) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31089b17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_602) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73409ffb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7c14535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_583) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b25d2289)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7aef22a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95ee76a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_400) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13869c3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52afe86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb765d7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea95b829)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea41c1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3306a35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_491) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42b17a1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_478) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c937f74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40dc0f24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebb0724d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81fc407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7932b44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12ecd141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cae6a4f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5eb4686c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d966e05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dfb6d79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_546) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(599ead0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_509) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(955cd323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_383) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(578fcc5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_585) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b06f8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fc67ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd32af64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226fcfcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3ea3794)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ef5ebd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b965d57a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(261176de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_426) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c2cc3c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_508) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_545) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c913e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_512) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ba3271a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84c57422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
