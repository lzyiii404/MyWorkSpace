//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_172_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [6:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [6:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [29:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [2:0]  _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_27;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_28;
  reg [31:0] _RAND_1;
  reg [72:0] _EVAL_56;
  reg [95:0] _RAND_2;
  reg [3:0] _EVAL_67;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_81;
  reg [31:0] _RAND_4;
  reg [29:0] _EVAL_119;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_121;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_142;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_171;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_190;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_208;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_222;
  reg [31:0] _RAND_11;
  reg  _EVAL_247;
  reg [31:0] _RAND_12;
  reg [6:0] _EVAL_248;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_289;
  reg [31:0] _RAND_14;
  wire  _EVAL_126;
  wire  _EVAL_69;
  wire  _EVAL_75;
  wire [12:0] _EVAL_205;
  wire [5:0] _EVAL_183;
  wire  _EVAL_207;
  wire  _EVAL_236;
  wire  _EVAL_242;
  wire [29:0] _EVAL_158;
  wire  _EVAL_18;
  wire  _EVAL_215;
  wire  _EVAL_23;
  wire  _EVAL_83;
  wire  _EVAL_203;
  wire  _EVAL_160;
  wire  _EVAL_273;
  wire [1:0] _EVAL_155;
  wire [1:0] _EVAL_140;
  wire  _EVAL_147;
  wire  _EVAL_177;
  wire  _EVAL_141;
  wire  _EVAL_165;
  wire  _EVAL_76;
  wire  _EVAL_135;
  wire  _EVAL_108;
  wire  _EVAL_263;
  wire  _EVAL_102;
  wire  _EVAL_116;
  wire  _EVAL_148;
  wire  _EVAL_209;
  wire  _EVAL_249;
  wire  _EVAL_99;
  wire  _EVAL_104;
  wire  _EVAL_175;
  wire  _EVAL_30;
  wire [3:0] _EVAL_138;
  wire [3:0] _EVAL_255;
  wire [127:0] _EVAL_269;
  wire  _EVAL_62;
  wire  _EVAL_43;
  wire  _EVAL_90;
  wire  _EVAL_57;
  wire  _EVAL_294;
  wire  _EVAL_281;
  wire  _EVAL_241;
  wire  _EVAL_206;
  wire  _EVAL_297;
  wire [3:0] _EVAL_33;
  wire  _EVAL_68;
  wire  _EVAL_214;
  wire  _EVAL_41;
  wire  _EVAL_38;
  wire [12:0] _EVAL_239;
  wire [5:0] _EVAL_268;
  wire [5:0] _EVAL_109;
  wire [3:0] _EVAL_245;
  wire [5:0] _EVAL_35;
  wire  _EVAL_202;
  wire  _EVAL_167;
  wire  _EVAL_92;
  wire  _EVAL_260;
  wire  _EVAL_145;
  wire  _EVAL_221;
  wire  _EVAL_110;
  wire  _EVAL_106;
  wire  _EVAL_173;
  wire  _EVAL_277;
  wire  _EVAL_296;
  wire  _EVAL_265;
  wire  _EVAL_120;
  wire [3:0] _EVAL_233;
  wire  _EVAL_115;
  wire [2:0] _EVAL_179;
  wire  _EVAL_162;
  wire  _EVAL_285;
  wire  _EVAL_295;
  wire  _EVAL_298;
  wire  _EVAL_95;
  wire  _EVAL_86;
  wire  _EVAL_280;
  wire  _EVAL_40;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_85;
  wire  _EVAL_185;
  wire  _EVAL_78;
  wire  _EVAL_112;
  wire  _EVAL_146;
  wire  _EVAL_168;
  wire  _EVAL_216;
  wire  _EVAL_118;
  wire  _EVAL_25;
  wire  _EVAL_161;
  wire [3:0] _EVAL_163;
  wire  _EVAL_253;
  wire  _EVAL_53;
  wire [72:0] _EVAL_204;
  wire  _EVAL_258;
  wire  _EVAL_82;
  wire [3:0] _EVAL_176;
  wire  _EVAL_199;
  wire  _EVAL_164;
  wire  _EVAL_132;
  wire  _EVAL_191;
  wire  _EVAL_127;
  wire  _EVAL_29;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_144;
  wire  _EVAL_72;
  wire  _EVAL_97;
  wire  _EVAL_94;
  wire  _EVAL_299;
  wire  _EVAL_271;
  wire  _EVAL_47;
  wire  _EVAL_211;
  wire  _EVAL_303;
  wire  _EVAL_250;
  wire  _EVAL_243;
  wire  _EVAL_122;
  wire  _EVAL_259;
  wire  _EVAL_46;
  wire  _EVAL_105;
  wire [127:0] _EVAL_107;
  wire [127:0] _EVAL_87;
  wire [72:0] _EVAL_244;
  wire  _EVAL_180;
  wire  _EVAL_219;
  wire  _EVAL_212;
  wire  _EVAL_292;
  wire [3:0] _EVAL_61;
  wire  _EVAL_238;
  wire [2:0] _EVAL_151;
  wire  _EVAL_88;
  wire  _EVAL_210;
  wire  _EVAL_186;
  wire  _EVAL_237;
  wire  _EVAL_74;
  wire  _EVAL_80;
  wire  _EVAL_184;
  wire  _EVAL_284;
  wire  _EVAL_246;
  wire  _EVAL_231;
  wire  _EVAL_174;
  wire  _EVAL_129;
  wire  _EVAL_300;
  wire  _EVAL_178;
  wire  _EVAL_291;
  wire [127:0] _EVAL_124;
  wire [72:0] _EVAL_34;
  wire  _EVAL_282;
  wire [3:0] _EVAL_266;
  wire [3:0] _EVAL_20;
  wire  _EVAL_44;
  wire  _EVAL_187;
  wire  _EVAL_136;
  wire  _EVAL_26;
  wire  _EVAL_234;
  wire  _EVAL_274;
  wire  _EVAL_267;
  wire  _EVAL_152;
  wire  _EVAL_264;
  wire  _EVAL_189;
  wire  _EVAL_261;
  wire  _EVAL_278;
  wire [3:0] _EVAL_256;
  wire  _EVAL_194;
  wire  _EVAL_125;
  wire  _EVAL_45;
  wire  _EVAL_71;
  wire [30:0] _EVAL_293;
  wire [30:0] _EVAL_65;
  wire [72:0] _EVAL_130;
  wire  _EVAL_262;
  wire  _EVAL_50;
  wire  _EVAL_101;
  wire  _EVAL_52;
  wire  _EVAL_166;
  wire [3:0] _EVAL_98;
  wire  _EVAL_31;
  wire  _EVAL_232;
  wire [30:0] _EVAL_224;
  wire [72:0] _EVAL_139;
  wire  _EVAL_113;
  wire  _EVAL_77;
  wire  _EVAL_195;
  wire  _EVAL_37;
  wire  _EVAL_55;
  wire  _EVAL_100;
  wire  _EVAL_96;
  wire  _EVAL_22;
  wire  _EVAL_157;
  wire  _EVAL_301;
  wire  _EVAL_251;
  wire  _EVAL_276;
  wire  _EVAL_91;
  wire  _EVAL_111;
  wire  _EVAL_36;
  wire  _EVAL_48;
  wire  _EVAL_32;
  wire  _EVAL_39;
  wire  _EVAL_159;
  wire  _EVAL_170;
  wire  _EVAL_134;
  wire  _EVAL_188;
  wire  _EVAL_143;
  wire  _EVAL_225;
  wire  _EVAL_181;
  wire  _EVAL_64;
  wire  _EVAL_60;
  wire [29:0] _EVAL_154;
  wire [29:0] _EVAL_131;
  wire  _EVAL_272;
  wire  _EVAL_226;
  wire  _EVAL_283;
  wire  _EVAL_182;
  wire [72:0] _EVAL_128;
  wire  _EVAL_218;
  wire  _EVAL_287;
  wire  _EVAL_133;
  wire  _EVAL_252;
  wire  _EVAL_54;
  wire  _EVAL_223;
  wire  _EVAL_21;
  wire  _EVAL_93;
  wire  _EVAL_198;
  wire [31:0] _EVAL_51;
  wire  _EVAL_254;
  wire  _EVAL_217;
  wire  _EVAL_172;
  wire  _EVAL_235;
  wire  _EVAL_169;
  wire  _EVAL_84;
  wire  _EVAL_257;
  wire  _EVAL_63;
  wire  _EVAL_193;
  wire  _EVAL_49;
  wire  _EVAL_200;
  wire  _EVAL_156;
  wire  _EVAL_197;
  wire  _EVAL_17;
  wire  _EVAL_290;
  wire  _EVAL_279;
  wire  _EVAL_19;
  wire  _EVAL_153;
  wire [72:0] _EVAL_288;
  wire  _EVAL_201;
  wire  _EVAL_270;
  wire  _EVAL_302;
  wire  _EVAL_123;
  wire  _EVAL_286;
  wire  _EVAL_66;
  wire  _EVAL_229;
  wire  _EVAL_114;
  wire [72:0] _EVAL_73;
  wire  _EVAL_230;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_126 = _EVAL_13 == _EVAL_119;
  assign _EVAL_69 = _EVAL_126 | _EVAL;
  assign _EVAL_75 = _EVAL_69 == 1'h0;
  assign _EVAL_205 = 13'h3f << _EVAL_11;
  assign _EVAL_183 = _EVAL_205[5:0];
  assign _EVAL_207 = _EVAL_15 & _EVAL_2;
  assign _EVAL_236 = _EVAL_289 == 4'h0;
  assign _EVAL_242 = _EVAL_207 & _EVAL_236;
  assign _EVAL_158 = _EVAL_13 ^ 30'h20000000;
  assign _EVAL_18 = _EVAL_13[1];
  assign _EVAL_215 = _EVAL_18 == 1'h0;
  assign _EVAL_23 = _EVAL_13[0];
  assign _EVAL_83 = _EVAL_23 == 1'h0;
  assign _EVAL_203 = _EVAL_215 & _EVAL_83;
  assign _EVAL_160 = _EVAL_16 >= 3'h2;
  assign _EVAL_273 = _EVAL_16[0];
  assign _EVAL_155 = 2'h1 << _EVAL_273;
  assign _EVAL_140 = _EVAL_155 | 2'h1;
  assign _EVAL_147 = _EVAL_140[1];
  assign _EVAL_177 = _EVAL_147 & _EVAL_18;
  assign _EVAL_141 = _EVAL_160 | _EVAL_177;
  assign _EVAL_165 = _EVAL_140[0];
  assign _EVAL_76 = _EVAL_18 & _EVAL_23;
  assign _EVAL_135 = _EVAL_165 & _EVAL_76;
  assign _EVAL_108 = _EVAL_141 | _EVAL_135;
  assign _EVAL_263 = _EVAL_18 & _EVAL_83;
  assign _EVAL_102 = _EVAL_165 & _EVAL_263;
  assign _EVAL_116 = _EVAL_141 | _EVAL_102;
  assign _EVAL_148 = _EVAL_147 & _EVAL_215;
  assign _EVAL_209 = _EVAL_160 | _EVAL_148;
  assign _EVAL_249 = _EVAL_215 & _EVAL_23;
  assign _EVAL_99 = _EVAL_165 & _EVAL_249;
  assign _EVAL_104 = _EVAL_209 | _EVAL_99;
  assign _EVAL_175 = _EVAL_165 & _EVAL_203;
  assign _EVAL_30 = _EVAL_209 | _EVAL_175;
  assign _EVAL_138 = {_EVAL_108,_EVAL_116,_EVAL_104,_EVAL_30};
  assign _EVAL_255 = ~ _EVAL_138;
  assign _EVAL_269 = 128'h1 << _EVAL_10;
  assign _EVAL_62 = _EVAL_4 == 3'h4;
  assign _EVAL_43 = _EVAL_8 == _EVAL_81;
  assign _EVAL_90 = _EVAL_1 == 7'h48;
  assign _EVAL_57 = _EVAL_1 == 7'h40;
  assign _EVAL_294 = _EVAL_90 | _EVAL_57;
  assign _EVAL_281 = _EVAL_12 == _EVAL_138;
  assign _EVAL_241 = _EVAL_281 | _EVAL;
  assign _EVAL_206 = _EVAL_241 == 1'h0;
  assign _EVAL_297 = plusarg_reader_out == 32'h0;
  assign _EVAL_33 = _EVAL_289 - 4'h1;
  assign _EVAL_68 = _EVAL_8 == 3'h7;
  assign _EVAL_214 = _EVAL_2 & _EVAL_68;
  assign _EVAL_41 = _EVAL_8[2];
  assign _EVAL_38 = _EVAL_41 == 1'h0;
  assign _EVAL_239 = 13'h3f << _EVAL_16;
  assign _EVAL_268 = _EVAL_239[5:0];
  assign _EVAL_109 = ~ _EVAL_268;
  assign _EVAL_245 = _EVAL_109[5:2];
  assign _EVAL_35 = ~ _EVAL_183;
  assign _EVAL_202 = _EVAL_27 < plusarg_reader_out;
  assign _EVAL_167 = _EVAL_4 == 3'h6;
  assign _EVAL_92 = _EVAL_9 & _EVAL_167;
  assign _EVAL_260 = _EVAL_1 == 7'h20;
  assign _EVAL_145 = _EVAL_8 == 3'h2;
  assign _EVAL_221 = _EVAL_1 == _EVAL_28;
  assign _EVAL_110 = _EVAL_160 | _EVAL;
  assign _EVAL_106 = _EVAL_6 <= 3'h4;
  assign _EVAL_173 = _EVAL_106 | _EVAL;
  assign _EVAL_277 = _EVAL_173 == 1'h0;
  assign _EVAL_296 = _EVAL_10 == 7'h48;
  assign _EVAL_265 = _EVAL_10 == 7'h40;
  assign _EVAL_120 = _EVAL_296 | _EVAL_265;
  assign _EVAL_233 = _EVAL_10[6:3];
  assign _EVAL_115 = _EVAL_233 == 4'h8;
  assign _EVAL_179 = _EVAL_10[2:0];
  assign _EVAL_162 = 3'h1 <= _EVAL_179;
  assign _EVAL_285 = _EVAL_115 & _EVAL_162;
  assign _EVAL_295 = _EVAL_120 | _EVAL_285;
  assign _EVAL_298 = _EVAL_10 == 7'h20;
  assign _EVAL_95 = _EVAL_295 | _EVAL_298;
  assign _EVAL_86 = _EVAL_233 == 4'h0;
  assign _EVAL_280 = _EVAL_95 | _EVAL_86;
  assign _EVAL_40 = _EVAL_233 == 4'h1;
  assign _EVAL_149 = _EVAL_280 | _EVAL_40;
  assign _EVAL_150 = _EVAL_233 == 4'h2;
  assign _EVAL_85 = _EVAL_149 | _EVAL_150;
  assign _EVAL_185 = _EVAL_233 == 4'h3;
  assign _EVAL_78 = _EVAL_85 | _EVAL_185;
  assign _EVAL_112 = _EVAL_78 | _EVAL;
  assign _EVAL_146 = _EVAL_3 == 1'h0;
  assign _EVAL_168 = _EVAL_146 | _EVAL_7;
  assign _EVAL_216 = _EVAL_168 | _EVAL;
  assign _EVAL_118 = _EVAL_216 == 1'h0;
  assign _EVAL_25 = _EVAL_11 >= 3'h2;
  assign _EVAL_161 = _EVAL_25 | _EVAL;
  assign _EVAL_163 = ~ _EVAL_12;
  assign _EVAL_253 = _EVAL_163 == 4'h0;
  assign _EVAL_53 = _EVAL_253 | _EVAL;
  assign _EVAL_204 = _EVAL_56 >> _EVAL_1;
  assign _EVAL_258 = _EVAL_204[0];
  assign _EVAL_82 = _EVAL_43 | _EVAL;
  assign _EVAL_176 = _EVAL_12 & _EVAL_255;
  assign _EVAL_199 = _EVAL_176 == 4'h0;
  assign _EVAL_164 = _EVAL_199 | _EVAL;
  assign _EVAL_132 = _EVAL_164 == 1'h0;
  assign _EVAL_191 = _EVAL_6 <= 3'h3;
  assign _EVAL_127 = _EVAL_191 | _EVAL;
  assign _EVAL_29 = _EVAL_16 == _EVAL_171;
  assign _EVAL_58 = _EVAL_29 | _EVAL;
  assign _EVAL_59 = _EVAL_58 == 1'h0;
  assign _EVAL_144 = _EVAL_5 & _EVAL_9;
  assign _EVAL_72 = _EVAL_67 == 4'h0;
  assign _EVAL_97 = _EVAL_144 & _EVAL_72;
  assign _EVAL_94 = _EVAL_167 == 1'h0;
  assign _EVAL_299 = _EVAL_97 & _EVAL_94;
  assign _EVAL_271 = _EVAL_8 == 3'h3;
  assign _EVAL_47 = _EVAL_2 & _EVAL_271;
  assign _EVAL_211 = _EVAL_258 == 1'h0;
  assign _EVAL_303 = _EVAL_211 | _EVAL;
  assign _EVAL_250 = _EVAL_303 == 1'h0;
  assign _EVAL_243 = _EVAL_3 == _EVAL_247;
  assign _EVAL_122 = _EVAL_243 | _EVAL;
  assign _EVAL_259 = _EVAL_6 != 3'h0;
  assign _EVAL_46 = _EVAL_142 == 4'h0;
  assign _EVAL_105 = _EVAL_207 & _EVAL_46;
  assign _EVAL_107 = 128'h1 << _EVAL_1;
  assign _EVAL_87 = _EVAL_105 ? _EVAL_107 : 128'h0;
  assign _EVAL_244 = _EVAL_87[72:0];
  assign _EVAL_180 = _EVAL_244 != 73'h0;
  assign _EVAL_219 = _EVAL_222 == 4'h0;
  assign _EVAL_212 = _EVAL_219 == 1'h0;
  assign _EVAL_292 = _EVAL_221 | _EVAL;
  assign _EVAL_61 = _EVAL_1[6:3];
  assign _EVAL_238 = _EVAL_61 == 4'h8;
  assign _EVAL_151 = _EVAL_1[2:0];
  assign _EVAL_88 = 3'h1 <= _EVAL_151;
  assign _EVAL_210 = _EVAL_238 & _EVAL_88;
  assign _EVAL_186 = _EVAL_294 | _EVAL_210;
  assign _EVAL_237 = _EVAL_186 | _EVAL_260;
  assign _EVAL_74 = _EVAL_61 == 4'h0;
  assign _EVAL_80 = _EVAL_237 | _EVAL_74;
  assign _EVAL_184 = _EVAL_61 == 4'h1;
  assign _EVAL_284 = _EVAL_80 | _EVAL_184;
  assign _EVAL_246 = _EVAL_61 == 4'h2;
  assign _EVAL_231 = _EVAL_284 | _EVAL_246;
  assign _EVAL_174 = _EVAL_61 == 4'h3;
  assign _EVAL_129 = _EVAL_231 | _EVAL_174;
  assign _EVAL_300 = _EVAL_129 | _EVAL;
  assign _EVAL_178 = _EVAL_4[0];
  assign _EVAL_291 = _EVAL_9 & _EVAL_62;
  assign _EVAL_124 = _EVAL_299 ? _EVAL_269 : 128'h0;
  assign _EVAL_34 = _EVAL_124[72:0];
  assign _EVAL_282 = _EVAL_244 != _EVAL_34;
  assign _EVAL_266 = _EVAL_35[5:2];
  assign _EVAL_20 = _EVAL_67 - 4'h1;
  assign _EVAL_44 = _EVAL_4 == _EVAL_121;
  assign _EVAL_187 = _EVAL_44 | _EVAL;
  assign _EVAL_136 = _EVAL_187 == 1'h0;
  assign _EVAL_26 = _EVAL_56 != 73'h0;
  assign _EVAL_234 = _EVAL_26 == 1'h0;
  assign _EVAL_274 = _EVAL_234 | _EVAL_297;
  assign _EVAL_267 = _EVAL_274 | _EVAL_202;
  assign _EVAL_152 = _EVAL_267 | _EVAL;
  assign _EVAL_264 = _EVAL_146 | _EVAL;
  assign _EVAL_189 = _EVAL_264 == 1'h0;
  assign _EVAL_261 = _EVAL_0 == 1'h0;
  assign _EVAL_278 = _EVAL_261 | _EVAL;
  assign _EVAL_256 = _EVAL_222 - 4'h1;
  assign _EVAL_194 = _EVAL_6 == _EVAL_190;
  assign _EVAL_125 = 3'h6 == _EVAL_16;
  assign _EVAL_45 = _EVAL_57 ? _EVAL_125 : 1'h0;
  assign _EVAL_71 = _EVAL_45 | _EVAL;
  assign _EVAL_293 = {1'b0,$signed(_EVAL_158)};
  assign _EVAL_65 = $signed(_EVAL_293) & $signed(-31'sh2000);
  assign _EVAL_130 = ~ _EVAL_34;
  assign _EVAL_262 = _EVAL_11 == _EVAL_208;
  assign _EVAL_50 = _EVAL_262 | _EVAL;
  assign _EVAL_101 = _EVAL_50 == 1'h0;
  assign _EVAL_52 = _EVAL_8 == 3'h0;
  assign _EVAL_166 = _EVAL_2 & _EVAL_52;
  assign _EVAL_98 = _EVAL_142 - 4'h1;
  assign _EVAL_31 = _EVAL_4 == 3'h2;
  assign _EVAL_232 = _EVAL_9 & _EVAL_31;
  assign _EVAL_224 = $signed(_EVAL_65);
  assign _EVAL_139 = _EVAL_244 | _EVAL_56;
  assign _EVAL_113 = _EVAL_2 & _EVAL_145;
  assign _EVAL_77 = _EVAL_8 == 3'h4;
  assign _EVAL_195 = _EVAL_16 <= 3'h6;
  assign _EVAL_37 = $signed(_EVAL_224) == $signed(31'sh0);
  assign _EVAL_55 = _EVAL_195 & _EVAL_37;
  assign _EVAL_100 = _EVAL_55 | _EVAL;
  assign _EVAL_96 = _EVAL_100 == 1'h0;
  assign _EVAL_22 = _EVAL_4 <= 3'h6;
  assign _EVAL_157 = _EVAL_22 | _EVAL;
  assign _EVAL_301 = _EVAL_157 == 1'h0;
  assign _EVAL_251 = _EVAL_4 == 3'h0;
  assign _EVAL_276 = _EVAL_8 == 3'h1;
  assign _EVAL_91 = _EVAL_8 == 3'h5;
  assign _EVAL_111 = _EVAL_2 & _EVAL_91;
  assign _EVAL_36 = _EVAL_180 == 1'h0;
  assign _EVAL_48 = _EVAL_282 | _EVAL_36;
  assign _EVAL_32 = _EVAL_48 | _EVAL;
  assign _EVAL_39 = _EVAL_32 == 1'h0;
  assign _EVAL_159 = _EVAL_9 & _EVAL_251;
  assign _EVAL_170 = _EVAL_7 == 1'h0;
  assign _EVAL_134 = _EVAL_9 & _EVAL_212;
  assign _EVAL_188 = _EVAL_4 == 3'h5;
  assign _EVAL_143 = _EVAL_9 & _EVAL_188;
  assign _EVAL_225 = _EVAL_170 | _EVAL;
  assign _EVAL_181 = _EVAL_236 == 1'h0;
  assign _EVAL_64 = _EVAL_2 & _EVAL_181;
  assign _EVAL_60 = _EVAL_300 == 1'h0;
  assign _EVAL_154 = {{24'd0}, _EVAL_109};
  assign _EVAL_131 = _EVAL_13 & _EVAL_154;
  assign _EVAL_272 = _EVAL_131 == 30'h0;
  assign _EVAL_226 = _EVAL_272 | _EVAL;
  assign _EVAL_283 = _EVAL_226 == 1'h0;
  assign _EVAL_182 = _EVAL_259 | _EVAL;
  assign _EVAL_128 = _EVAL_139 >> _EVAL_10;
  assign _EVAL_218 = _EVAL_128[0];
  assign _EVAL_287 = _EVAL_225 == 1'h0;
  assign _EVAL_133 = _EVAL_207 | _EVAL_144;
  assign _EVAL_252 = _EVAL_8 == 3'h6;
  assign _EVAL_54 = _EVAL_2 & _EVAL_252;
  assign _EVAL_223 = _EVAL_4 == 3'h1;
  assign _EVAL_21 = _EVAL_218 | _EVAL;
  assign _EVAL_93 = _EVAL_21 == 1'h0;
  assign _EVAL_198 = _EVAL_122 == 1'h0;
  assign _EVAL_51 = _EVAL_27 + 32'h1;
  assign _EVAL_254 = _EVAL_2 & _EVAL_276;
  assign _EVAL_217 = _EVAL_278 == 1'h0;
  assign _EVAL_172 = _EVAL_292 == 1'h0;
  assign _EVAL_235 = _EVAL_6 <= 3'h2;
  assign _EVAL_169 = _EVAL_2 & _EVAL_77;
  assign _EVAL_84 = _EVAL_144 & _EVAL_219;
  assign _EVAL_257 = _EVAL_194 | _EVAL;
  assign _EVAL_63 = _EVAL_257 == 1'h0;
  assign _EVAL_193 = _EVAL_112 == 1'h0;
  assign _EVAL_49 = _EVAL_235 | _EVAL;
  assign _EVAL_200 = _EVAL_49 == 1'h0;
  assign _EVAL_156 = _EVAL_182 == 1'h0;
  assign _EVAL_197 = _EVAL_10 == _EVAL_248;
  assign _EVAL_17 = _EVAL_197 | _EVAL;
  assign _EVAL_290 = _EVAL == 1'h0;
  assign _EVAL_279 = _EVAL_6 == 3'h0;
  assign _EVAL_19 = _EVAL_152 == 1'h0;
  assign _EVAL_153 = _EVAL_82 == 1'h0;
  assign _EVAL_288 = _EVAL_56 | _EVAL_244;
  assign _EVAL_201 = _EVAL_110 == 1'h0;
  assign _EVAL_270 = _EVAL_17 == 1'h0;
  assign _EVAL_302 = _EVAL_279 | _EVAL;
  assign _EVAL_123 = _EVAL_71 == 1'h0;
  assign _EVAL_286 = _EVAL_127 == 1'h0;
  assign _EVAL_66 = _EVAL_161 == 1'h0;
  assign _EVAL_229 = _EVAL_9 & _EVAL_223;
  assign _EVAL_114 = _EVAL_302 == 1'h0;
  assign _EVAL_73 = _EVAL_288 & _EVAL_130;
  assign _EVAL_230 = _EVAL_53 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_27 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_28 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {3{`RANDOM}};
  _EVAL_56 = _RAND_2[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_67 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_81 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_119 = _RAND_5[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_121 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_142 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_171 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_190 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_208 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_222 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_247 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_248 = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_289 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL) begin
      _EVAL_27 <= 32'h0;
    end else begin
      if (_EVAL_133) begin
        _EVAL_27 <= 32'h0;
      end else begin
        _EVAL_27 <= _EVAL_51;
      end
    end
    if (_EVAL_242) begin
      _EVAL_28 <= _EVAL_1;
    end
    if (_EVAL) begin
      _EVAL_56 <= 73'h0;
    end else begin
      _EVAL_56 <= _EVAL_73;
    end
    if (_EVAL) begin
      _EVAL_67 <= 4'h0;
    end else begin
      if (_EVAL_144) begin
        if (_EVAL_72) begin
          if (_EVAL_178) begin
            _EVAL_67 <= _EVAL_266;
          end else begin
            _EVAL_67 <= 4'h0;
          end
        end else begin
          _EVAL_67 <= _EVAL_20;
        end
      end
    end
    if (_EVAL_242) begin
      _EVAL_81 <= _EVAL_8;
    end
    if (_EVAL_242) begin
      _EVAL_119 <= _EVAL_13;
    end
    if (_EVAL_84) begin
      _EVAL_121 <= _EVAL_4;
    end
    if (_EVAL) begin
      _EVAL_142 <= 4'h0;
    end else begin
      if (_EVAL_207) begin
        if (_EVAL_46) begin
          if (_EVAL_38) begin
            _EVAL_142 <= _EVAL_245;
          end else begin
            _EVAL_142 <= 4'h0;
          end
        end else begin
          _EVAL_142 <= _EVAL_98;
        end
      end
    end
    if (_EVAL_242) begin
      _EVAL_171 <= _EVAL_16;
    end
    if (_EVAL_242) begin
      _EVAL_190 <= _EVAL_6;
    end
    if (_EVAL_84) begin
      _EVAL_208 <= _EVAL_11;
    end
    if (_EVAL) begin
      _EVAL_222 <= 4'h0;
    end else begin
      if (_EVAL_144) begin
        if (_EVAL_219) begin
          if (_EVAL_178) begin
            _EVAL_222 <= _EVAL_266;
          end else begin
            _EVAL_222 <= 4'h0;
          end
        end else begin
          _EVAL_222 <= _EVAL_256;
        end
      end
    end
    if (_EVAL_84) begin
      _EVAL_247 <= _EVAL_3;
    end
    if (_EVAL_84) begin
      _EVAL_248 <= _EVAL_10;
    end
    if (_EVAL) begin
      _EVAL_289 <= 4'h0;
    end else begin
      if (_EVAL_207) begin
        if (_EVAL_236) begin
          if (_EVAL_38) begin
            _EVAL_289 <= _EVAL_245;
          end else begin
            _EVAL_289 <= 4'h0;
          end
        end else begin
          _EVAL_289 <= _EVAL_33;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(808af58c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d317a93b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0aeaf90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a4391e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(210d240b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4a75bd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(899a0b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf5bf044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30a3441c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25e8d8da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b780fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb8c432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(822cbee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4c3f0cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e6d1acc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ce43c39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a58cce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eb770b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83c68e65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb51a35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f66e62e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35736f01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b2703a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8835be42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a425f59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30da9593)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb64fa40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e746b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4a55021)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9ba313a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5af380a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(905e7e3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61a0bd46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ef356c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c4445ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7f4d543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b484f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc32fb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaba50a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(168ca410)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c1c8aa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78dc8ed3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be987ff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b84ce40c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(802f1cc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc0c798)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23370815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(394bcd60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c39d62f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6002024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57b385c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54063205)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5e56b62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(814c0bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad724b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61e0214f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a5de2af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feaa085e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f71a3ab6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c290e3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d317b874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0fcedf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71939e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(271be4c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0fb2f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4c241fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97738ff0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3216d65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c00bc045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2815b3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6632e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3815352f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16a7cada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb1501c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0950ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15f1993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5fc133d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f51584b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c16c105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a4d080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
