//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_168(
  output [2:0]  _EVAL,
  output [7:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output [31:0] _EVAL_5,
  input  [29:0] _EVAL_6,
  input  [31:0] _EVAL_7,
  output [3:0]  _EVAL_8,
  input  [3:0]  _EVAL_9,
  output [1:0]  _EVAL_10,
  output [1:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output [29:0] _EVAL_16,
  output        _EVAL_17,
  output [15:0] _EVAL_18,
  input  [3:0]  _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [15:0] _EVAL_21,
  input         _EVAL_22,
  output [29:0] _EVAL_23,
  output [3:0]  _EVAL_24,
  output        _EVAL_25,
  output [3:0]  _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  output [1:0]  _EVAL_31,
  output        _EVAL_32,
  output [3:0]  _EVAL_33,
  output        _EVAL_34,
  output [7:0]  _EVAL_35,
  input  [2:0]  _EVAL_36,
  output        _EVAL_37,
  input  [7:0]  _EVAL_38,
  input         _EVAL_39,
  output [31:0] _EVAL_40,
  input  [1:0]  _EVAL_41,
  input  [15:0] _EVAL_42,
  output [15:0] _EVAL_43,
  output [2:0]  _EVAL_44,
  input  [2:0]  _EVAL_45,
  output        _EVAL_46,
  input  [7:0]  _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49,
  output [15:0] _EVAL_50,
  input  [31:0] _EVAL_51,
  output        _EVAL_52,
  input  [15:0] _EVAL_53,
  input  [1:0]  _EVAL_54,
  output        _EVAL_55,
  output [1:0]  _EVAL_56,
  output [2:0]  _EVAL_57,
  input         _EVAL_58,
  input  [15:0] _EVAL_59,
  input  [3:0]  _EVAL_60,
  output        _EVAL_61,
  output [15:0] _EVAL_62,
  input  [29:0] _EVAL_63,
  input         _EVAL_64,
  output [2:0]  _EVAL_65,
  output [3:0]  _EVAL_66,
  input  [1:0]  _EVAL_67,
  input  [3:0]  _EVAL_68,
  input         _EVAL_69,
  output        _EVAL_70,
  output        _EVAL_71,
  output        _EVAL_72,
  output        _EVAL_73,
  input  [3:0]  _EVAL_74,
  output        _EVAL_75,
  input  [1:0]  _EVAL_76
);
  assign _EVAL_46 = _EVAL_58;
  assign _EVAL_0 = _EVAL_47;
  assign _EVAL_31 = _EVAL_54;
  assign _EVAL_73 = _EVAL_1;
  assign _EVAL_17 = _EVAL_14;
  assign _EVAL_32 = _EVAL_2;
  assign _EVAL_61 = _EVAL_69;
  assign _EVAL_16 = _EVAL_6;
  assign _EVAL_15 = _EVAL_3;
  assign _EVAL_37 = _EVAL_30;
  assign _EVAL_10 = _EVAL_76;
  assign _EVAL_44 = _EVAL_45;
  assign _EVAL_8 = _EVAL_60;
  assign _EVAL_70 = _EVAL_29;
  assign _EVAL_24 = _EVAL_19;
  assign _EVAL_35 = _EVAL_38;
  assign _EVAL_18 = _EVAL_53;
  assign _EVAL_25 = _EVAL_39;
  assign _EVAL_11 = _EVAL_41;
  assign _EVAL_65 = _EVAL_20;
  assign _EVAL_34 = _EVAL_13;
  assign _EVAL_26 = _EVAL_9;
  assign _EVAL_55 = _EVAL_48;
  assign _EVAL_50 = _EVAL_21;
  assign _EVAL_40 = _EVAL_51;
  assign _EVAL_52 = _EVAL_64;
  assign _EVAL_23 = _EVAL_63;
  assign _EVAL_75 = _EVAL_4;
  assign _EVAL_33 = _EVAL_68;
  assign _EVAL_49 = _EVAL_27;
  assign _EVAL_71 = _EVAL_22;
  assign _EVAL_62 = _EVAL_42;
  assign _EVAL = _EVAL_36;
  assign _EVAL_72 = _EVAL_28;
  assign _EVAL_5 = _EVAL_7;
  assign _EVAL_66 = _EVAL_74;
  assign _EVAL_43 = _EVAL_59;
  assign _EVAL_57 = _EVAL_12;
  assign _EVAL_56 = _EVAL_67;
endmodule
