//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_289(
  input         _EVAL,
  input  [4:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  input  [9:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input  [48:0] _EVAL_10,
  output [9:0]  _EVAL_11,
  output        _EVAL_12,
  input  [25:0] _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input  [2:0]  _EVAL_16,
  input         _EVAL_17,
  output [26:0] _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23
);
  wire [1:0] _EVAL_26;
  wire  _EVAL_209;
  wire [25:0] _EVAL_324;
  wire [25:0] _EVAL_271;
  wire [47:0] _EVAL_290;
  wire [74:0] _EVAL_24;
  wire [46:0] _EVAL_76;
  wire [49:0] _EVAL_261;
  wire [23:0] _EVAL_218;
  wire [23:0] _EVAL_317;
  wire  _EVAL_43;
  wire [50:0] _EVAL_238;
  wire [50:0] _EVAL_307;
  wire [50:0] _EVAL_173;
  wire [50:0] _EVAL_226;
  wire [50:0] _EVAL_160;
  wire  _EVAL_322;
  wire [1:0] _EVAL_132;
  wire  _EVAL_213;
  wire [1:0] _EVAL_217;
  wire  _EVAL_77;
  wire [1:0] _EVAL_116;
  wire  _EVAL_127;
  wire [1:0] _EVAL_32;
  wire  _EVAL_228;
  wire [1:0] _EVAL_254;
  wire  _EVAL_252;
  wire [1:0] _EVAL_267;
  wire  _EVAL_135;
  wire [1:0] _EVAL_178;
  wire  _EVAL_319;
  wire [1:0] _EVAL_253;
  wire  _EVAL_193;
  wire [1:0] _EVAL_129;
  wire  _EVAL_45;
  wire [1:0] _EVAL_256;
  wire  _EVAL_335;
  wire [1:0] _EVAL_49;
  wire  _EVAL_177;
  wire [1:0] _EVAL_104;
  wire  _EVAL_195;
  wire [5:0] _EVAL_118;
  wire [1:0] _EVAL_72;
  wire  _EVAL_263;
  wire [1:0] _EVAL_55;
  wire  _EVAL_326;
  wire [1:0] _EVAL_251;
  wire  _EVAL_65;
  wire [1:0] _EVAL_187;
  wire  _EVAL_310;
  wire [1:0] _EVAL_299;
  wire  _EVAL_265;
  wire [1:0] _EVAL_171;
  wire  _EVAL_30;
  wire [1:0] _EVAL_149;
  wire  _EVAL_152;
  wire [1:0] _EVAL_266;
  wire  _EVAL_120;
  wire [1:0] _EVAL_278;
  wire  _EVAL_147;
  wire [1:0] _EVAL_142;
  wire  _EVAL_258;
  wire [1:0] _EVAL_189;
  wire  _EVAL_172;
  wire [1:0] _EVAL_225;
  wire  _EVAL_293;
  wire [1:0] _EVAL_196;
  wire  _EVAL_316;
  wire [5:0] _EVAL_141;
  wire [12:0] _EVAL_229;
  wire [25:0] _EVAL_291;
  wire [15:0] _EVAL_243;
  wire [7:0] _EVAL_131;
  wire [15:0] _EVAL_309;
  wire [7:0] _EVAL_133;
  wire [15:0] _EVAL_111;
  wire [15:0] _EVAL_150;
  wire [15:0] _EVAL_184;
  wire [11:0] _EVAL_125;
  wire [15:0] _EVAL_134;
  wire [15:0] _EVAL_86;
  wire [11:0] _EVAL_47;
  wire [15:0] _EVAL_36;
  wire [15:0] _EVAL_288;
  wire [15:0] _EVAL_224;
  wire [13:0] _EVAL_227;
  wire [15:0] _EVAL_73;
  wire [15:0] _EVAL_210;
  wire [13:0] _EVAL_88;
  wire [15:0] _EVAL_219;
  wire [15:0] _EVAL_207;
  wire [15:0] _EVAL_119;
  wire [14:0] _EVAL_41;
  wire [15:0] _EVAL_198;
  wire [15:0] _EVAL_139;
  wire [14:0] _EVAL_107;
  wire [15:0] _EVAL_100;
  wire [15:0] _EVAL_186;
  wire [15:0] _EVAL_205;
  wire [9:0] _EVAL_235;
  wire [7:0] _EVAL_281;
  wire [3:0] _EVAL_113;
  wire [7:0] _EVAL_318;
  wire [3:0] _EVAL_190;
  wire [7:0] _EVAL_110;
  wire [7:0] _EVAL_234;
  wire [7:0] _EVAL_304;
  wire [5:0] _EVAL_48;
  wire [7:0] _EVAL_103;
  wire [7:0] _EVAL_327;
  wire [5:0] _EVAL_179;
  wire [7:0] _EVAL_334;
  wire [7:0] _EVAL_123;
  wire [7:0] _EVAL_90;
  wire [6:0] _EVAL_33;
  wire [7:0] _EVAL_53;
  wire [7:0] _EVAL_280;
  wire [6:0] _EVAL_211;
  wire [7:0] _EVAL_122;
  wire [7:0] _EVAL_64;
  wire [7:0] _EVAL_287;
  wire [1:0] _EVAL_212;
  wire  _EVAL_340;
  wire  _EVAL_126;
  wire [25:0] _EVAL_300;
  wire  _EVAL_168;
  wire  _EVAL_94;
  wire  _EVAL_44;
  wire  _EVAL_67;
  wire  _EVAL_283;
  wire  _EVAL_155;
  wire  _EVAL_237;
  wire  _EVAL_220;
  wire  _EVAL_329;
  wire  _EVAL_29;
  wire  _EVAL_244;
  wire  _EVAL_325;
  wire  _EVAL_39;
  wire  _EVAL_85;
  wire  _EVAL_54;
  wire  _EVAL_121;
  wire  _EVAL_233;
  wire  _EVAL_180;
  wire  _EVAL_276;
  wire [4:0] _EVAL_61;
  wire [4:0] _EVAL_42;
  wire [4:0] _EVAL_285;
  wire [4:0] _EVAL_146;
  wire [4:0] _EVAL_89;
  wire [4:0] _EVAL_50;
  wire [4:0] _EVAL_200;
  wire [4:0] _EVAL_246;
  wire [4:0] _EVAL_328;
  wire [4:0] _EVAL_197;
  wire [4:0] _EVAL_191;
  wire [4:0] _EVAL_130;
  wire [4:0] _EVAL_62;
  wire [4:0] _EVAL_40;
  wire [4:0] _EVAL_188;
  wire [4:0] _EVAL_320;
  wire [4:0] _EVAL_260;
  wire [4:0] _EVAL_151;
  wire  _EVAL_305;
  wire  _EVAL_78;
  wire  _EVAL_71;
  wire  _EVAL_303;
  wire  _EVAL_332;
  wire  _EVAL_286;
  wire  _EVAL_166;
  wire  _EVAL_313;
  wire  _EVAL_167;
  wire [4:0] _EVAL_214;
  wire [4:0] _EVAL_157;
  wire [4:0] _EVAL_272;
  wire [4:0] _EVAL_99;
  wire [4:0] _EVAL_25;
  wire [4:0] _EVAL_202;
  wire [4:0] _EVAL_63;
  wire [3:0] _EVAL_112;
  wire [3:0] _EVAL_159;
  wire [16:0] _EVAL_59;
  wire [5:0] _EVAL_289;
  wire [1:0] _EVAL_38;
  wire [49:0] _EVAL_174;
  wire [49:0] _EVAL_323;
  wire [49:0] _EVAL_162;
  wire [23:0] _EVAL_181;
  wire [26:0] _EVAL_156;
  wire [3:0] _EVAL_221;
  wire  _EVAL_270;
  wire [1:0] _EVAL_274;
  wire [9:0] _EVAL_204;
  wire  _EVAL_222;
  wire  _EVAL_315;
  wire  _EVAL_31;
  wire  _EVAL_257;
  wire  _EVAL_165;
  wire [3:0] _EVAL_108;
  wire [1:0] _EVAL_294;
  wire  _EVAL_240;
  wire  _EVAL_153;
  wire  _EVAL_75;
  wire  _EVAL_81;
  wire [80:0] _EVAL_302;
  wire [1:0] _EVAL_87;
  wire  _EVAL_284;
  wire  _EVAL_194;
  wire [24:0] _EVAL_138;
  wire  _EVAL_295;
  wire  _EVAL_301;
  wire [2:0] _EVAL_203;
  wire [2:0] _EVAL_201;
  wire [8:0] _EVAL_95;
  wire [5:0] _EVAL_338;
  wire [1:0] _EVAL_231;
  wire  _EVAL_161;
  wire [12:0] _EVAL_331;
  wire [1:0] _EVAL_199;
  wire  _EVAL_268;
  wire  _EVAL_175;
  wire  _EVAL_37;
  wire  _EVAL_57;
  wire [2:0] _EVAL_312;
  wire  _EVAL_70;
  wire  _EVAL_339;
  wire  _EVAL_216;
  wire  _EVAL_176;
  wire  _EVAL_51;
  wire  _EVAL_245;
  wire  _EVAL_143;
  wire  _EVAL_247;
  wire  _EVAL_140;
  wire [9:0] _EVAL_206;
  wire [3:0] _EVAL_169;
  wire  _EVAL_109;
  wire [3:0] _EVAL_83;
  wire [1:0] _EVAL_105;
  wire [3:0] _EVAL_35;
  wire  _EVAL_170;
  wire [113:0] _EVAL_232;
  wire [5:0] _EVAL_185;
  wire [113:0] _EVAL_223;
  wire [28:0] _EVAL_321;
  wire [2:0] _EVAL_154;
  wire  _EVAL_249;
  wire  _EVAL_311;
  wire [1:0] _EVAL_66;
  wire  _EVAL_262;
  wire [1:0] _EVAL_28;
  wire  _EVAL_136;
  wire [1:0] _EVAL_102;
  wire  _EVAL_163;
  wire [1:0] _EVAL_279;
  wire  _EVAL_264;
  wire [1:0] _EVAL_336;
  wire  _EVAL_92;
  wire [6:0] _EVAL_91;
  wire  _EVAL_308;
  wire  _EVAL_117;
  wire  _EVAL_337;
  wire  _EVAL_208;
  wire [5:0] _EVAL_80;
  wire [6:0] _EVAL_82;
  wire [6:0] _EVAL_250;
  wire  _EVAL_236;
  wire  _EVAL_192;
  wire  _EVAL_158;
  wire  _EVAL_69;
  wire [25:0] _EVAL_58;
  wire [26:0] _EVAL_34;
  wire [1:0] _EVAL_97;
  wire  _EVAL_27;
  wire [80:0] _EVAL_330;
  wire [28:0] _EVAL_215;
  wire [2:0] _EVAL_46;
  wire  _EVAL_230;
  wire [9:0] _EVAL_255;
  wire [1:0] _EVAL_56;
  wire  _EVAL_297;
  wire  _EVAL_333;
  wire [25:0] _EVAL_298;
  wire  _EVAL_84;
  wire [3:0] _EVAL_145;
  wire  _EVAL_314;
  wire [3:0] _EVAL_144;
  wire  _EVAL_93;
  wire [3:0] _EVAL_137;
  wire  _EVAL_275;
  wire [6:0] _EVAL_273;
  wire  _EVAL_101;
  wire  _EVAL_292;
  wire  _EVAL_182;
  wire  _EVAL_241;
  wire [5:0] _EVAL_148;
  wire [6:0] _EVAL_277;
  wire [6:0] _EVAL_164;
  wire  _EVAL_115;
  wire  _EVAL_106;
  wire  _EVAL_52;
  wire [26:0] _EVAL_242;
  wire  _EVAL_68;
  wire  _EVAL_306;
  wire  _EVAL_79;
  wire [6:0] _EVAL_248;
  wire [9:0] _EVAL_60;
  wire  _EVAL_96;
  wire  _EVAL_74;
  wire  _EVAL_296;
  wire [9:0] _EVAL_128;
  wire [9:0] _EVAL_239;
  wire  _EVAL_259;
  wire  _EVAL_124;
  wire  _EVAL_98;
  assign _EVAL_26 = _EVAL_13[25:24];
  assign _EVAL_209 = _EVAL_10[48];
  assign _EVAL_324 = _EVAL_13 + 26'h1;
  assign _EVAL_271 = _EVAL_209 ? _EVAL_324 : _EVAL_13;
  assign _EVAL_290 = _EVAL_10[47:0];
  assign _EVAL_24 = {_EVAL_271,_EVAL_290,_EVAL_17};
  assign _EVAL_76 = _EVAL_24[72:26];
  assign _EVAL_261 = {1'h0,_EVAL_26,_EVAL_76};
  assign _EVAL_218 = _EVAL_24[24:1];
  assign _EVAL_317 = ~ _EVAL_218;
  assign _EVAL_43 = _EVAL_24[51];
  assign _EVAL_238 = _EVAL_24[50:0];
  assign _EVAL_307 = ~ _EVAL_238;
  assign _EVAL_173 = {{50'd0}, _EVAL_23};
  assign _EVAL_226 = _EVAL_238 + _EVAL_173;
  assign _EVAL_160 = _EVAL_43 ? _EVAL_307 : _EVAL_226;
  assign _EVAL_322 = _EVAL_160[50];
  assign _EVAL_132 = _EVAL_160[49:48];
  assign _EVAL_213 = _EVAL_132 != 2'h0;
  assign _EVAL_217 = _EVAL_160[47:46];
  assign _EVAL_77 = _EVAL_217 != 2'h0;
  assign _EVAL_116 = _EVAL_160[45:44];
  assign _EVAL_127 = _EVAL_116 != 2'h0;
  assign _EVAL_32 = _EVAL_160[43:42];
  assign _EVAL_228 = _EVAL_32 != 2'h0;
  assign _EVAL_254 = _EVAL_160[41:40];
  assign _EVAL_252 = _EVAL_254 != 2'h0;
  assign _EVAL_267 = _EVAL_160[39:38];
  assign _EVAL_135 = _EVAL_267 != 2'h0;
  assign _EVAL_178 = _EVAL_160[37:36];
  assign _EVAL_319 = _EVAL_178 != 2'h0;
  assign _EVAL_253 = _EVAL_160[35:34];
  assign _EVAL_193 = _EVAL_253 != 2'h0;
  assign _EVAL_129 = _EVAL_160[33:32];
  assign _EVAL_45 = _EVAL_129 != 2'h0;
  assign _EVAL_256 = _EVAL_160[31:30];
  assign _EVAL_335 = _EVAL_256 != 2'h0;
  assign _EVAL_49 = _EVAL_160[29:28];
  assign _EVAL_177 = _EVAL_49 != 2'h0;
  assign _EVAL_104 = _EVAL_160[27:26];
  assign _EVAL_195 = _EVAL_104 != 2'h0;
  assign _EVAL_118 = {_EVAL_319,_EVAL_193,_EVAL_45,_EVAL_335,_EVAL_177,_EVAL_195};
  assign _EVAL_72 = _EVAL_160[25:24];
  assign _EVAL_263 = _EVAL_72 != 2'h0;
  assign _EVAL_55 = _EVAL_160[23:22];
  assign _EVAL_326 = _EVAL_55 != 2'h0;
  assign _EVAL_251 = _EVAL_160[21:20];
  assign _EVAL_65 = _EVAL_251 != 2'h0;
  assign _EVAL_187 = _EVAL_160[19:18];
  assign _EVAL_310 = _EVAL_187 != 2'h0;
  assign _EVAL_299 = _EVAL_160[17:16];
  assign _EVAL_265 = _EVAL_299 != 2'h0;
  assign _EVAL_171 = _EVAL_160[15:14];
  assign _EVAL_30 = _EVAL_171 != 2'h0;
  assign _EVAL_149 = _EVAL_160[13:12];
  assign _EVAL_152 = _EVAL_149 != 2'h0;
  assign _EVAL_266 = _EVAL_160[11:10];
  assign _EVAL_120 = _EVAL_266 != 2'h0;
  assign _EVAL_278 = _EVAL_160[9:8];
  assign _EVAL_147 = _EVAL_278 != 2'h0;
  assign _EVAL_142 = _EVAL_160[7:6];
  assign _EVAL_258 = _EVAL_142 != 2'h0;
  assign _EVAL_189 = _EVAL_160[5:4];
  assign _EVAL_172 = _EVAL_189 != 2'h0;
  assign _EVAL_225 = _EVAL_160[3:2];
  assign _EVAL_293 = _EVAL_225 != 2'h0;
  assign _EVAL_196 = _EVAL_160[1:0];
  assign _EVAL_316 = _EVAL_196 != 2'h0;
  assign _EVAL_141 = {_EVAL_120,_EVAL_147,_EVAL_258,_EVAL_172,_EVAL_293,_EVAL_316};
  assign _EVAL_229 = {_EVAL_263,_EVAL_326,_EVAL_65,_EVAL_310,_EVAL_265,_EVAL_30,_EVAL_152,_EVAL_141};
  assign _EVAL_291 = {_EVAL_322,_EVAL_213,_EVAL_77,_EVAL_127,_EVAL_228,_EVAL_252,_EVAL_135,_EVAL_118,_EVAL_229};
  assign _EVAL_243 = _EVAL_291[15:0];
  assign _EVAL_131 = _EVAL_243[15:8];
  assign _EVAL_309 = {{8'd0}, _EVAL_131};
  assign _EVAL_133 = _EVAL_243[7:0];
  assign _EVAL_111 = {_EVAL_133, 8'h0};
  assign _EVAL_150 = _EVAL_111 & 16'hff00;
  assign _EVAL_184 = _EVAL_309 | _EVAL_150;
  assign _EVAL_125 = _EVAL_184[15:4];
  assign _EVAL_134 = {{4'd0}, _EVAL_125};
  assign _EVAL_86 = _EVAL_134 & 16'hf0f;
  assign _EVAL_47 = _EVAL_184[11:0];
  assign _EVAL_36 = {_EVAL_47, 4'h0};
  assign _EVAL_288 = _EVAL_36 & 16'hf0f0;
  assign _EVAL_224 = _EVAL_86 | _EVAL_288;
  assign _EVAL_227 = _EVAL_224[15:2];
  assign _EVAL_73 = {{2'd0}, _EVAL_227};
  assign _EVAL_210 = _EVAL_73 & 16'h3333;
  assign _EVAL_88 = _EVAL_224[13:0];
  assign _EVAL_219 = {_EVAL_88, 2'h0};
  assign _EVAL_207 = _EVAL_219 & 16'hcccc;
  assign _EVAL_119 = _EVAL_210 | _EVAL_207;
  assign _EVAL_41 = _EVAL_119[15:1];
  assign _EVAL_198 = {{1'd0}, _EVAL_41};
  assign _EVAL_139 = _EVAL_198 & 16'h5555;
  assign _EVAL_107 = _EVAL_119[14:0];
  assign _EVAL_100 = {_EVAL_107, 1'h0};
  assign _EVAL_186 = _EVAL_100 & 16'haaaa;
  assign _EVAL_205 = _EVAL_139 | _EVAL_186;
  assign _EVAL_235 = _EVAL_291[25:16];
  assign _EVAL_281 = _EVAL_235[7:0];
  assign _EVAL_113 = _EVAL_281[7:4];
  assign _EVAL_318 = {{4'd0}, _EVAL_113};
  assign _EVAL_190 = _EVAL_281[3:0];
  assign _EVAL_110 = {_EVAL_190, 4'h0};
  assign _EVAL_234 = _EVAL_110 & 8'hf0;
  assign _EVAL_304 = _EVAL_318 | _EVAL_234;
  assign _EVAL_48 = _EVAL_304[7:2];
  assign _EVAL_103 = {{2'd0}, _EVAL_48};
  assign _EVAL_327 = _EVAL_103 & 8'h33;
  assign _EVAL_179 = _EVAL_304[5:0];
  assign _EVAL_334 = {_EVAL_179, 2'h0};
  assign _EVAL_123 = _EVAL_334 & 8'hcc;
  assign _EVAL_90 = _EVAL_327 | _EVAL_123;
  assign _EVAL_33 = _EVAL_90[7:1];
  assign _EVAL_53 = {{1'd0}, _EVAL_33};
  assign _EVAL_280 = _EVAL_53 & 8'h55;
  assign _EVAL_211 = _EVAL_90[6:0];
  assign _EVAL_122 = {_EVAL_211, 1'h0};
  assign _EVAL_64 = _EVAL_122 & 8'haa;
  assign _EVAL_287 = _EVAL_280 | _EVAL_64;
  assign _EVAL_212 = _EVAL_235[9:8];
  assign _EVAL_340 = _EVAL_212[0];
  assign _EVAL_126 = _EVAL_212[1];
  assign _EVAL_300 = {_EVAL_205,_EVAL_287,_EVAL_340,_EVAL_126};
  assign _EVAL_168 = _EVAL_300[0];
  assign _EVAL_94 = _EVAL_300[7];
  assign _EVAL_44 = _EVAL_300[8];
  assign _EVAL_67 = _EVAL_300[9];
  assign _EVAL_283 = _EVAL_300[10];
  assign _EVAL_155 = _EVAL_300[11];
  assign _EVAL_237 = _EVAL_300[12];
  assign _EVAL_220 = _EVAL_300[13];
  assign _EVAL_329 = _EVAL_300[14];
  assign _EVAL_29 = _EVAL_300[15];
  assign _EVAL_244 = _EVAL_300[16];
  assign _EVAL_325 = _EVAL_300[17];
  assign _EVAL_39 = _EVAL_300[18];
  assign _EVAL_85 = _EVAL_300[19];
  assign _EVAL_54 = _EVAL_300[20];
  assign _EVAL_121 = _EVAL_300[21];
  assign _EVAL_233 = _EVAL_300[22];
  assign _EVAL_180 = _EVAL_300[23];
  assign _EVAL_276 = _EVAL_300[24];
  assign _EVAL_61 = _EVAL_276 ? 5'h18 : 5'h19;
  assign _EVAL_42 = _EVAL_180 ? 5'h17 : _EVAL_61;
  assign _EVAL_285 = _EVAL_233 ? 5'h16 : _EVAL_42;
  assign _EVAL_146 = _EVAL_121 ? 5'h15 : _EVAL_285;
  assign _EVAL_89 = _EVAL_54 ? 5'h14 : _EVAL_146;
  assign _EVAL_50 = _EVAL_85 ? 5'h13 : _EVAL_89;
  assign _EVAL_200 = _EVAL_39 ? 5'h12 : _EVAL_50;
  assign _EVAL_246 = _EVAL_325 ? 5'h11 : _EVAL_200;
  assign _EVAL_328 = _EVAL_244 ? 5'h10 : _EVAL_246;
  assign _EVAL_197 = _EVAL_29 ? 5'hf : _EVAL_328;
  assign _EVAL_191 = _EVAL_329 ? 5'he : _EVAL_197;
  assign _EVAL_130 = _EVAL_220 ? 5'hd : _EVAL_191;
  assign _EVAL_62 = _EVAL_237 ? 5'hc : _EVAL_130;
  assign _EVAL_40 = _EVAL_155 ? 5'hb : _EVAL_62;
  assign _EVAL_188 = _EVAL_283 ? 5'ha : _EVAL_40;
  assign _EVAL_320 = _EVAL_67 ? 5'h9 : _EVAL_188;
  assign _EVAL_260 = _EVAL_44 ? 5'h8 : _EVAL_320;
  assign _EVAL_151 = _EVAL_94 ? 5'h7 : _EVAL_260;
  assign _EVAL_305 = _EVAL_20 | _EVAL;
  assign _EVAL_78 = _EVAL_305 & _EVAL_21;
  assign _EVAL_71 = _EVAL_78 == 1'h0;
  assign _EVAL_303 = _EVAL_300[1];
  assign _EVAL_332 = _EVAL_300[2];
  assign _EVAL_286 = _EVAL_300[3];
  assign _EVAL_166 = _EVAL_300[4];
  assign _EVAL_313 = _EVAL_300[5];
  assign _EVAL_167 = _EVAL_300[6];
  assign _EVAL_214 = _EVAL_167 ? 5'h6 : _EVAL_151;
  assign _EVAL_157 = _EVAL_313 ? 5'h5 : _EVAL_214;
  assign _EVAL_272 = _EVAL_166 ? 5'h4 : _EVAL_157;
  assign _EVAL_99 = _EVAL_286 ? 5'h3 : _EVAL_272;
  assign _EVAL_25 = _EVAL_332 ? 5'h2 : _EVAL_99;
  assign _EVAL_202 = _EVAL_303 ? 5'h1 : _EVAL_25;
  assign _EVAL_63 = _EVAL_168 ? 5'h0 : _EVAL_202;
  assign _EVAL_112 = _EVAL_63[4:1];
  assign _EVAL_159 = ~ _EVAL_112;
  assign _EVAL_59 = $signed(-17'sh10000) >>> _EVAL_159;
  assign _EVAL_289 = _EVAL_59[6:1];
  assign _EVAL_38 = _EVAL_289[5:4];
  assign _EVAL_174 = _EVAL_24[74:25];
  assign _EVAL_323 = ~ _EVAL_174;
  assign _EVAL_162 = _EVAL_23 ? _EVAL_323 : _EVAL_261;
  assign _EVAL_181 = _EVAL_162[23:0];
  assign _EVAL_156 = {_EVAL_181, 3'h0};
  assign _EVAL_221 = _EVAL_156[3:0];
  assign _EVAL_270 = _EVAL_221 != 4'h0;
  assign _EVAL_274 = {1'b0,$signed(_EVAL_23)};
  assign _EVAL_204 = {{8{_EVAL_274[1]}},_EVAL_274};
  assign _EVAL_222 = _EVAL_19 | _EVAL_14;
  assign _EVAL_315 = _EVAL_222 | _EVAL_5;
  assign _EVAL_31 = _EVAL_315 == 1'h0;
  assign _EVAL_257 = _EVAL_31 & _EVAL_71;
  assign _EVAL_165 = _EVAL_16 == 3'h2;
  assign _EVAL_108 = _EVAL_289[3:0];
  assign _EVAL_294 = _EVAL_108[3:2];
  assign _EVAL_240 = _EVAL_78 & _EVAL_165;
  assign _EVAL_153 = _EVAL_22 ^ _EVAL_23;
  assign _EVAL_75 = _EVAL_22 | _EVAL_153;
  assign _EVAL_81 = _EVAL_240 & _EVAL_75;
  assign _EVAL_302 = {{31'd0}, _EVAL_162};
  assign _EVAL_87 = _EVAL_108[1:0];
  assign _EVAL_284 = _EVAL_87[0];
  assign _EVAL_194 = _EVAL_317 != 24'h0;
  assign _EVAL_138 = _EVAL_24[25:1];
  assign _EVAL_295 = _EVAL_138 != 25'h0;
  assign _EVAL_301 = _EVAL_23 ? _EVAL_194 : _EVAL_295;
  assign _EVAL_203 = _EVAL_0[4:2];
  assign _EVAL_201 = ~ _EVAL_203;
  assign _EVAL_95 = $signed(-9'sh100) >>> _EVAL_201;
  assign _EVAL_338 = _EVAL_95[6:1];
  assign _EVAL_231 = _EVAL_338[5:4];
  assign _EVAL_161 = _EVAL_231[0];
  assign _EVAL_331 = _EVAL_291[12:0];
  assign _EVAL_199 = _EVAL_331[1:0];
  assign _EVAL_268 = _EVAL_199 != 2'h0;
  assign _EVAL_175 = _EVAL_1 == 1'h0;
  assign _EVAL_37 = _EVAL_175 & _EVAL_222;
  assign _EVAL_57 = _EVAL_37 & _EVAL_5;
  assign _EVAL_312 = _EVAL_156[26:24];
  assign _EVAL_70 = _EVAL_294[1];
  assign _EVAL_339 = _EVAL_222 & _EVAL_22;
  assign _EVAL_216 = _EVAL_5 & _EVAL_153;
  assign _EVAL_176 = _EVAL_339 | _EVAL_216;
  assign _EVAL_51 = _EVAL_165 == 1'h0;
  assign _EVAL_245 = _EVAL_78 & _EVAL_51;
  assign _EVAL_143 = _EVAL_245 & _EVAL_22;
  assign _EVAL_247 = _EVAL_143 & _EVAL_153;
  assign _EVAL_140 = _EVAL_176 | _EVAL_247;
  assign _EVAL_206 = $signed(_EVAL_7) - $signed(_EVAL_204);
  assign _EVAL_169 = _EVAL_156[7:4];
  assign _EVAL_109 = _EVAL_169 != 4'h0;
  assign _EVAL_83 = _EVAL_338[3:0];
  assign _EVAL_105 = _EVAL_83[3:2];
  assign _EVAL_35 = _EVAL_156[23:20];
  assign _EVAL_170 = _EVAL_35 != 4'h0;
  assign _EVAL_232 = {{63'd0}, _EVAL_160};
  assign _EVAL_185 = {_EVAL_63, 1'h0};
  assign _EVAL_223 = _EVAL_232 << _EVAL_185;
  assign _EVAL_321 = _EVAL_223[51:23];
  assign _EVAL_154 = _EVAL_321[2:0];
  assign _EVAL_249 = _EVAL_154 != 3'h0;
  assign _EVAL_311 = _EVAL_331[12];
  assign _EVAL_66 = _EVAL_331[11:10];
  assign _EVAL_262 = _EVAL_66 != 2'h0;
  assign _EVAL_28 = _EVAL_331[9:8];
  assign _EVAL_136 = _EVAL_28 != 2'h0;
  assign _EVAL_102 = _EVAL_331[7:6];
  assign _EVAL_163 = _EVAL_102 != 2'h0;
  assign _EVAL_279 = _EVAL_331[5:4];
  assign _EVAL_264 = _EVAL_279 != 2'h0;
  assign _EVAL_336 = _EVAL_331[3:2];
  assign _EVAL_92 = _EVAL_336 != 2'h0;
  assign _EVAL_91 = {_EVAL_311,_EVAL_262,_EVAL_136,_EVAL_163,_EVAL_264,_EVAL_92,_EVAL_268};
  assign _EVAL_308 = _EVAL_87[1];
  assign _EVAL_117 = _EVAL_294[0];
  assign _EVAL_337 = _EVAL_38[0];
  assign _EVAL_208 = _EVAL_38[1];
  assign _EVAL_80 = {_EVAL_284,_EVAL_308,_EVAL_117,_EVAL_70,_EVAL_337,_EVAL_208};
  assign _EVAL_82 = {{1'd0}, _EVAL_80};
  assign _EVAL_250 = _EVAL_91 & _EVAL_82;
  assign _EVAL_236 = _EVAL_250 != 7'h0;
  assign _EVAL_192 = _EVAL_249 | _EVAL_236;
  assign _EVAL_158 = _EVAL_19 & _EVAL;
  assign _EVAL_69 = _EVAL_2 | _EVAL_158;
  assign _EVAL_58 = _EVAL_321[28:3];
  assign _EVAL_34 = {_EVAL_58,_EVAL_192};
  assign _EVAL_97 = _EVAL_34[26:25];
  assign _EVAL_27 = _EVAL_20 & _EVAL_14;
  assign _EVAL_330 = _EVAL_302 << _EVAL_0;
  assign _EVAL_215 = _EVAL_330[49:21];
  assign _EVAL_46 = _EVAL_215[2:0];
  assign _EVAL_230 = _EVAL_46 != 3'h0;
  assign _EVAL_255 = $signed(_EVAL_206);
  assign _EVAL_56 = _EVAL_83[1:0];
  assign _EVAL_297 = _EVAL_56[1];
  assign _EVAL_333 = _EVAL_69 | _EVAL_27;
  assign _EVAL_298 = _EVAL_215[28:3];
  assign _EVAL_84 = _EVAL_312 != 3'h0;
  assign _EVAL_145 = _EVAL_156[19:16];
  assign _EVAL_314 = _EVAL_145 != 4'h0;
  assign _EVAL_144 = _EVAL_156[15:12];
  assign _EVAL_93 = _EVAL_144 != 4'h0;
  assign _EVAL_137 = _EVAL_156[11:8];
  assign _EVAL_275 = _EVAL_137 != 4'h0;
  assign _EVAL_273 = {_EVAL_84,_EVAL_170,_EVAL_314,_EVAL_93,_EVAL_275,_EVAL_109,_EVAL_270};
  assign _EVAL_101 = _EVAL_56[0];
  assign _EVAL_292 = _EVAL_105[0];
  assign _EVAL_182 = _EVAL_105[1];
  assign _EVAL_241 = _EVAL_231[1];
  assign _EVAL_148 = {_EVAL_101,_EVAL_297,_EVAL_292,_EVAL_182,_EVAL_161,_EVAL_241};
  assign _EVAL_277 = {{1'd0}, _EVAL_148};
  assign _EVAL_164 = _EVAL_273 & _EVAL_277;
  assign _EVAL_115 = _EVAL_164 != 7'h0;
  assign _EVAL_106 = _EVAL_230 | _EVAL_115;
  assign _EVAL_52 = _EVAL_106 | _EVAL_301;
  assign _EVAL_242 = {_EVAL_298,_EVAL_52};
  assign _EVAL_68 = _EVAL_97 == 2'h0;
  assign _EVAL_306 = _EVAL_22 ^ _EVAL_43;
  assign _EVAL_79 = _EVAL_68 ? _EVAL_165 : _EVAL_306;
  assign _EVAL_248 = {1'b0,$signed(_EVAL_185)};
  assign _EVAL_60 = {{3{_EVAL_248[6]}},_EVAL_248};
  assign _EVAL_96 = _EVAL_57 & _EVAL_23;
  assign _EVAL_74 = _EVAL_4 ? _EVAL_153 : _EVAL_79;
  assign _EVAL_296 = _EVAL_257 & _EVAL_74;
  assign _EVAL_128 = $signed(_EVAL_7) - $signed(_EVAL_60);
  assign _EVAL_239 = $signed(_EVAL_128);
  assign _EVAL_259 = _EVAL_4 == 1'h0;
  assign _EVAL_124 = _EVAL_259 & _EVAL_68;
  assign _EVAL_98 = _EVAL_140 | _EVAL_81;
  assign _EVAL_18 = _EVAL_4 ? _EVAL_242 : _EVAL_34;
  assign _EVAL_12 = _EVAL_78 | _EVAL_124;
  assign _EVAL_8 = _EVAL_98 | _EVAL_296;
  assign _EVAL_11 = _EVAL_4 ? $signed(_EVAL_255) : $signed(_EVAL_239);
  assign _EVAL_15 = _EVAL_333 | _EVAL_96;
  assign _EVAL_9 = _EVAL_222 | _EVAL_5;
  assign _EVAL_6 = _EVAL_1 | _EVAL_3;
endmodule
