//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_69(
  output        _EVAL,
  input         _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  input  [31:0] _EVAL_3,
  input  [31:0] _EVAL_4,
  input  [1:0]  _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  output [3:0]  _EVAL_8,
  output [4:0]  _EVAL_9,
  output        _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [4:0]  _EVAL_13,
  output [31:0] _EVAL_14,
  input         _EVAL_15,
  input  [7:0]  _EVAL_16,
  output        _EVAL_17,
  output [2:0]  _EVAL_18,
  output        _EVAL_19,
  output [3:0]  _EVAL_20,
  output        _EVAL_21,
  input  [7:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [31:0] _EVAL_25,
  input         _EVAL_26,
  output [2:0]  _EVAL_27,
  input         _EVAL_28,
  output [31:0] _EVAL_29,
  input  [2:0]  _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  input  [2:0]  _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  output [1:0]  _EVAL_37,
  input  [3:0]  _EVAL_38,
  output [31:0] _EVAL_39,
  output        _EVAL_40,
  output [1:0]  _EVAL_41,
  input  [3:0]  _EVAL_42,
  output [1:0]  _EVAL_43,
  input         _EVAL_44,
  output [1:0]  _EVAL_45
);
  wire  Queue__EVAL;
  wire  Queue__EVAL_0;
  wire [1:0] Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire [1:0] Queue__EVAL_4;
  wire [31:0] Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire [1:0] Queue__EVAL_9;
  wire [1:0] Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire [31:0] Queue__EVAL_12;
  wire  Queue_1__EVAL;
  wire [1:0] Queue_1__EVAL_0;
  wire [1:0] Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire [1:0] Queue_1__EVAL_4;
  wire [1:0] Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire  Queue_1__EVAL_8;
  reg  _EVAL_110;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_142;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_156;
  reg [31:0] _RAND_2;
  reg [7:0] _EVAL_179;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_200;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_223;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_232;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_245;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_254;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_256;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_298;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_319;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_325;
  reg [31:0] _RAND_12;
  reg  _EVAL_394;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_403;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_432;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_440;
  reg [31:0] _RAND_16;
  wire [15:0] _EVAL_341;
  wire [22:0] _EVAL_149;
  wire [22:0] _EVAL_170;
  wire [14:0] _EVAL_265;
  wire [15:0] _EVAL_235;
  wire [15:0] _EVAL_446;
  wire [15:0] _EVAL_333;
  wire [15:0] _EVAL_117;
  wire [15:0] _EVAL_424;
  wire [7:0] _EVAL_73;
  wire  _EVAL_242;
  wire [7:0] _EVAL_85;
  wire [7:0] _EVAL_216;
  wire [3:0] _EVAL_322;
  wire  _EVAL_402;
  wire [3:0] _EVAL_133;
  wire [3:0] _EVAL_46;
  wire [1:0] _EVAL_351;
  wire  _EVAL_313;
  wire [1:0] _EVAL_344;
  wire [1:0] _EVAL_53;
  wire  _EVAL_222;
  wire [3:0] _EVAL_354;
  wire  _EVAL_148;
  wire  _EVAL_88;
  wire [1:0] _EVAL_138;
  wire [1:0] _EVAL_260;
  wire  _EVAL_426;
  wire  _EVAL_127;
  wire [31:0] _EVAL_241;
  wire [32:0] _EVAL_379;
  wire [32:0] _EVAL_202;
  wire [32:0] _EVAL_229;
  wire  _EVAL_56;
  wire [31:0] _EVAL_201;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_188;
  wire [32:0] _EVAL_401;
  wire  _EVAL_391;
  wire  _EVAL_79;
  wire [31:0] _EVAL_324;
  wire [32:0] _EVAL_270;
  wire [32:0] _EVAL_122;
  wire [32:0] _EVAL_253;
  wire  _EVAL_350;
  wire  _EVAL_430;
  wire [31:0] _EVAL_349;
  wire [32:0] _EVAL_137;
  wire [32:0] _EVAL_378;
  wire [32:0] _EVAL_282;
  wire  _EVAL_52;
  wire  _EVAL_128;
  wire [32:0] _EVAL_436;
  wire [32:0] _EVAL_189;
  wire [32:0] _EVAL_250;
  wire  _EVAL_348;
  wire  _EVAL_310;
  wire [31:0] _EVAL_74;
  wire [32:0] _EVAL_102;
  wire [32:0] _EVAL_366;
  wire [32:0] _EVAL_103;
  wire  _EVAL_293;
  wire  _EVAL_197;
  wire [31:0] _EVAL_301;
  wire [32:0] _EVAL_288;
  wire [32:0] _EVAL_421;
  wire [32:0] _EVAL_269;
  wire  _EVAL_84;
  wire  _EVAL_66;
  wire [31:0] _EVAL_435;
  wire [32:0] _EVAL_417;
  wire [32:0] _EVAL_247;
  wire [32:0] _EVAL_316;
  wire  _EVAL_126;
  wire  _EVAL_150;
  wire  _EVAL_309;
  wire  _EVAL_60;
  wire [31:0] _EVAL_248;
  wire [32:0] _EVAL_80;
  wire [32:0] _EVAL_392;
  wire [32:0] _EVAL_387;
  wire  _EVAL_238;
  wire  _EVAL_75;
  wire  _EVAL_166;
  wire [1:0] _EVAL_427;
  wire [13:0] _EVAL_144;
  wire [13:0] _EVAL_220;
  wire [31:0] _EVAL_164;
  wire  _EVAL_277;
  wire  _EVAL_342;
  wire  _EVAL_139;
  wire  _EVAL_101;
  wire  _EVAL_225;
  wire  _EVAL_99;
  wire  _EVAL_327;
  wire  _EVAL_153;
  wire  _EVAL_190;
  wire  _EVAL_300;
  wire  _EVAL_251;
  wire [1:0] _EVAL_90;
  wire [1:0] _EVAL_174;
  wire [1:0] _EVAL_183;
  wire [3:0] _EVAL_161;
  wire [2:0] _EVAL_286;
  wire [3:0] _EVAL_358;
  wire [3:0] _EVAL_210;
  wire [2:0] _EVAL_259;
  wire [3:0] _EVAL_281;
  wire [3:0] _EVAL_203;
  wire [3:0] _EVAL_67;
  wire [1:0] _EVAL_346;
  wire [1:0] _EVAL_275;
  wire [1:0] _EVAL_154;
  wire [1:0] _EVAL_345;
  wire  _EVAL_311;
  wire  _EVAL_347;
  wire  _EVAL_240;
  wire  _EVAL_278;
  wire [15:0] _EVAL_112;
  wire [22:0] _EVAL_82;
  wire [22:0] _EVAL_303;
  wire [14:0] _EVAL_244;
  wire [15:0] _EVAL_420;
  wire [15:0] _EVAL_199;
  wire [15:0] _EVAL_398;
  wire [15:0] _EVAL_271;
  wire [15:0] _EVAL_119;
  wire [7:0] _EVAL_425;
  wire  _EVAL_121;
  wire [7:0] _EVAL_268;
  wire [7:0] _EVAL_314;
  wire [3:0] _EVAL_233;
  wire  _EVAL_176;
  wire [3:0] _EVAL_55;
  wire [3:0] _EVAL_339;
  wire [1:0] _EVAL_155;
  wire  _EVAL_437;
  wire [1:0] _EVAL_444;
  wire [1:0] _EVAL_239;
  wire  _EVAL_370;
  wire [3:0] _EVAL_135;
  wire  _EVAL_143;
  wire [1:0] _EVAL_147;
  wire [2:0] _EVAL_81;
  wire [2:0] _EVAL_302;
  wire [2:0] _EVAL_163;
  wire [2:0] _EVAL_167;
  wire [2:0] _EVAL_335;
  wire [2:0] _EVAL_360;
  wire  _EVAL_249;
  wire  _EVAL_266;
  wire  _EVAL_395;
  wire [3:0] _EVAL_390;
  wire  _EVAL_372;
  wire  _EVAL_317;
  wire  _EVAL_283;
  wire  _EVAL_380;
  wire  _EVAL_98;
  wire  _EVAL_192;
  wire  _EVAL_297;
  wire  _EVAL_272;
  wire [31:0] _EVAL_331;
  wire [32:0] _EVAL_304;
  wire [32:0] _EVAL_337;
  wire [32:0] _EVAL_400;
  wire  _EVAL_285;
  wire [31:0] _EVAL_375;
  wire [32:0] _EVAL_140;
  wire [32:0] _EVAL_58;
  wire [32:0] _EVAL_340;
  wire  _EVAL_175;
  wire [31:0] _EVAL_423;
  wire [32:0] _EVAL_118;
  wire [32:0] _EVAL_289;
  wire [32:0] _EVAL_442;
  wire  _EVAL_113;
  wire  _EVAL_194;
  wire [31:0] _EVAL_336;
  wire [32:0] _EVAL_204;
  wire [32:0] _EVAL_362;
  wire [32:0] _EVAL_371;
  wire  _EVAL_217;
  wire  _EVAL_261;
  wire  _EVAL_211;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_295;
  wire [32:0] _EVAL_94;
  wire  _EVAL_114;
  wire  _EVAL_385;
  wire [31:0] _EVAL_165;
  wire [32:0] _EVAL_359;
  wire [32:0] _EVAL_64;
  wire [32:0] _EVAL_274;
  wire  _EVAL_59;
  wire  _EVAL_125;
  wire [31:0] _EVAL_123;
  wire [32:0] _EVAL_330;
  wire [32:0] _EVAL_318;
  wire [32:0] _EVAL_407;
  wire  _EVAL_182;
  wire  _EVAL_416;
  wire  _EVAL_93;
  wire  _EVAL_445;
  wire  _EVAL_334;
  wire  _EVAL_169;
  wire [3:0] _EVAL_258;
  wire  _EVAL_105;
  wire  _EVAL_92;
  wire [2:0] _EVAL_246;
  wire [2:0] _EVAL_196;
  wire [2:0] _EVAL_257;
  wire [2:0] _EVAL_255;
  wire [1:0] _EVAL_77;
  wire  _EVAL_226;
  wire  _EVAL_363;
  wire [2:0] _EVAL_78;
  wire [2:0] _EVAL_262;
  wire [2:0] _EVAL_49;
  wire [2:0] _EVAL_280;
  wire [1:0] _EVAL_355;
  wire  _EVAL_195;
  wire  _EVAL_72;
  wire [1:0] _EVAL_219;
  wire [13:0] _EVAL_384;
  wire [13:0] _EVAL_132;
  wire  _EVAL_315;
  wire  _EVAL_83;
  wire  _EVAL_441;
  wire [22:0] _EVAL_48;
  wire [7:0] _EVAL_422;
  wire [7:0] _EVAL_54;
  wire  _EVAL_443;
  wire  _EVAL_208;
  wire  _EVAL_152;
  wire [31:0] _EVAL_187;
  wire [32:0] _EVAL_215;
  wire [32:0] _EVAL_198;
  wire [32:0] _EVAL_279;
  wire  _EVAL_120;
  wire  _EVAL_367;
  wire [3:0] _EVAL_61;
  wire  _EVAL_320;
  wire  _EVAL_411;
  wire  _EVAL_214;
  wire  _EVAL_414;
  wire  _EVAL_171;
  wire  _EVAL_68;
  wire [5:0] _EVAL_146;
  wire  _EVAL_65;
  wire  _EVAL_386;
  wire [7:0] _EVAL_184;
  wire  _EVAL_399;
  wire [2:0] _EVAL_206;
  wire  _EVAL_191;
  wire [2:0] _EVAL_160;
  wire  _EVAL_368;
  wire  _EVAL_299;
  wire  _EVAL_95;
  wire  _EVAL_180;
  wire [2:0] _EVAL_47;
  wire  _EVAL_51;
  wire  _EVAL_276;
  wire [31:0] _EVAL_89;
  wire [32:0] _EVAL_352;
  wire [32:0] _EVAL_338;
  wire [32:0] _EVAL_205;
  wire  _EVAL_447;
  wire  _EVAL_267;
  wire  _EVAL_70;
  wire [31:0] _EVAL_97;
  wire  _EVAL_212;
  wire  _EVAL_129;
  wire  _EVAL_159;
  wire  _EVAL_145;
  wire  _EVAL_224;
  wire  _EVAL_393;
  wire  _EVAL_236;
  wire  _EVAL_227;
  wire  _EVAL_185;
  wire  _EVAL_312;
  wire  _EVAL_100;
  wire [68:0] _EVAL_356;
  wire [83:0] _EVAL_369;
  wire [83:0] _EVAL_431;
  wire  _EVAL_69;
  wire  _EVAL_63;
  wire [2:0] _EVAL_116;
  wire  _EVAL_243;
  wire [5:0] _EVAL_263;
  wire [5:0] _EVAL_106;
  wire [2:0] _EVAL_264;
  wire [2:0] _EVAL_305;
  wire  _EVAL_86;
  wire [68:0] _EVAL_328;
  wire [83:0] _EVAL_71;
  wire [83:0] _EVAL_357;
  wire  _EVAL_439;
  wire  _EVAL_136;
  wire  _EVAL_221;
  wire [1:0] _EVAL_172;
  wire [2:0] _EVAL_228;
  wire [7:0] _EVAL_62;
  wire  _EVAL_230;
  wire [2:0] _EVAL_124;
  wire  _EVAL_291;
  wire [1:0] _EVAL_410;
  wire  _EVAL_406;
  wire [2:0] _EVAL_433;
  wire  _EVAL_412;
  wire  _EVAL_376;
  wire [2:0] _EVAL_353;
  wire  _EVAL_178;
  wire  _EVAL_173;
  wire  _EVAL_115;
  wire [2:0] _EVAL_292;
  wire  _EVAL_323;
  wire [1:0] _EVAL_287;
  wire  _EVAL_429;
  wire [83:0] _EVAL_134;
  SiFive__EVAL_67 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12)
  );
  SiFive__EVAL_68 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8)
  );
  assign _EVAL_341 = {_EVAL_22,8'hff};
  assign _EVAL_149 = {{7'd0}, _EVAL_341};
  assign _EVAL_170 = _EVAL_149 << _EVAL_12;
  assign _EVAL_265 = _EVAL_170[22:8];
  assign _EVAL_235 = {_EVAL_265, 1'h0};
  assign _EVAL_446 = _EVAL_235 | 16'h1;
  assign _EVAL_333 = {1'h0,_EVAL_265};
  assign _EVAL_117 = ~ _EVAL_333;
  assign _EVAL_424 = _EVAL_446 & _EVAL_117;
  assign _EVAL_73 = _EVAL_424[15:8];
  assign _EVAL_242 = _EVAL_73 != 8'h0;
  assign _EVAL_85 = _EVAL_424[7:0];
  assign _EVAL_216 = _EVAL_73 | _EVAL_85;
  assign _EVAL_322 = _EVAL_216[7:4];
  assign _EVAL_402 = _EVAL_322 != 4'h0;
  assign _EVAL_133 = _EVAL_216[3:0];
  assign _EVAL_46 = _EVAL_322 | _EVAL_133;
  assign _EVAL_351 = _EVAL_46[3:2];
  assign _EVAL_313 = _EVAL_351 != 2'h0;
  assign _EVAL_344 = _EVAL_46[1:0];
  assign _EVAL_53 = _EVAL_351 | _EVAL_344;
  assign _EVAL_222 = _EVAL_53[1];
  assign _EVAL_354 = {_EVAL_242,_EVAL_402,_EVAL_313,_EVAL_222};
  assign _EVAL_148 = _EVAL_354 >= 4'h2;
  assign _EVAL_88 = _EVAL_354[0];
  assign _EVAL_138 = 2'h1 << _EVAL_88;
  assign _EVAL_260 = _EVAL_138 | 2'h1;
  assign _EVAL_426 = _EVAL_260[1];
  assign _EVAL_127 = _EVAL_354 <= 4'h6;
  assign _EVAL_241 = _EVAL_25 ^ 32'h40000000;
  assign _EVAL_379 = {1'b0,$signed(_EVAL_241)};
  assign _EVAL_202 = $signed(_EVAL_379) & $signed(-33'sh2000);
  assign _EVAL_229 = $signed(_EVAL_202);
  assign _EVAL_56 = $signed(_EVAL_229) == $signed(33'sh0);
  assign _EVAL_201 = _EVAL_25 ^ 32'h80000000;
  assign _EVAL_104 = {1'b0,$signed(_EVAL_201)};
  assign _EVAL_188 = $signed(_EVAL_104) & $signed(-33'sh20000);
  assign _EVAL_401 = $signed(_EVAL_188);
  assign _EVAL_391 = $signed(_EVAL_401) == $signed(33'sh0);
  assign _EVAL_79 = _EVAL_56 | _EVAL_391;
  assign _EVAL_324 = _EVAL_25 ^ 32'hc000000;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_324)};
  assign _EVAL_122 = $signed(_EVAL_270) & $signed(-33'sh4000000);
  assign _EVAL_253 = $signed(_EVAL_122);
  assign _EVAL_350 = $signed(_EVAL_253) == $signed(33'sh0);
  assign _EVAL_430 = _EVAL_79 | _EVAL_350;
  assign _EVAL_349 = _EVAL_25 ^ 32'h2000000;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_349)};
  assign _EVAL_378 = $signed(_EVAL_137) & $signed(-33'sh10000);
  assign _EVAL_282 = $signed(_EVAL_378);
  assign _EVAL_52 = $signed(_EVAL_282) == $signed(33'sh0);
  assign _EVAL_128 = _EVAL_430 | _EVAL_52;
  assign _EVAL_436 = {1'b0,$signed(_EVAL_25)};
  assign _EVAL_189 = $signed(_EVAL_436) & $signed(-33'sh5000);
  assign _EVAL_250 = $signed(_EVAL_189);
  assign _EVAL_348 = $signed(_EVAL_250) == $signed(33'sh0);
  assign _EVAL_310 = _EVAL_128 | _EVAL_348;
  assign _EVAL_74 = _EVAL_25 ^ 32'h1800000;
  assign _EVAL_102 = {1'b0,$signed(_EVAL_74)};
  assign _EVAL_366 = $signed(_EVAL_102) & $signed(-33'sh8000);
  assign _EVAL_103 = $signed(_EVAL_366);
  assign _EVAL_293 = $signed(_EVAL_103) == $signed(33'sh0);
  assign _EVAL_197 = _EVAL_310 | _EVAL_293;
  assign _EVAL_301 = _EVAL_25 ^ 32'h1900000;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_301)};
  assign _EVAL_421 = $signed(_EVAL_288) & $signed(-33'sh2000);
  assign _EVAL_269 = $signed(_EVAL_421);
  assign _EVAL_84 = $signed(_EVAL_269) == $signed(33'sh0);
  assign _EVAL_66 = _EVAL_197 | _EVAL_84;
  assign _EVAL_435 = _EVAL_25 ^ 32'h20000000;
  assign _EVAL_417 = {1'b0,$signed(_EVAL_435)};
  assign _EVAL_247 = $signed(_EVAL_417) & $signed(-33'sh2000);
  assign _EVAL_316 = $signed(_EVAL_247);
  assign _EVAL_126 = $signed(_EVAL_316) == $signed(33'sh0);
  assign _EVAL_150 = _EVAL_66 | _EVAL_126;
  assign _EVAL_309 = _EVAL_127 & _EVAL_150;
  assign _EVAL_60 = _EVAL_354 <= 4'h8;
  assign _EVAL_248 = _EVAL_25 ^ 32'h3000;
  assign _EVAL_80 = {1'b0,$signed(_EVAL_248)};
  assign _EVAL_392 = $signed(_EVAL_80) & $signed(-33'sh1000);
  assign _EVAL_387 = $signed(_EVAL_392);
  assign _EVAL_238 = $signed(_EVAL_387) == $signed(33'sh0);
  assign _EVAL_75 = _EVAL_60 & _EVAL_238;
  assign _EVAL_166 = _EVAL_309 | _EVAL_75;
  assign _EVAL_427 = _EVAL_25[1:0];
  assign _EVAL_144 = {{12'd0}, _EVAL_427};
  assign _EVAL_220 = 14'h3000 | _EVAL_144;
  assign _EVAL_164 = _EVAL_166 ? _EVAL_25 : {{18'd0}, _EVAL_220};
  assign _EVAL_277 = _EVAL_164[1];
  assign _EVAL_342 = _EVAL_277 == 1'h0;
  assign _EVAL_139 = _EVAL_426 & _EVAL_342;
  assign _EVAL_101 = _EVAL_148 | _EVAL_139;
  assign _EVAL_225 = _EVAL_260[0];
  assign _EVAL_99 = _EVAL_164[0];
  assign _EVAL_327 = _EVAL_99 == 1'h0;
  assign _EVAL_153 = _EVAL_342 & _EVAL_327;
  assign _EVAL_190 = _EVAL_225 & _EVAL_153;
  assign _EVAL_300 = _EVAL_101 | _EVAL_190;
  assign _EVAL_251 = _EVAL_26 & _EVAL_15;
  assign _EVAL_90 = {_EVAL_251,_EVAL_23};
  assign _EVAL_174 = ~ _EVAL_319;
  assign _EVAL_183 = _EVAL_90 & _EVAL_174;
  assign _EVAL_161 = {_EVAL_183,_EVAL_251,_EVAL_23};
  assign _EVAL_286 = _EVAL_161[3:1];
  assign _EVAL_358 = {{1'd0}, _EVAL_286};
  assign _EVAL_210 = _EVAL_161 | _EVAL_358;
  assign _EVAL_259 = _EVAL_210[3:1];
  assign _EVAL_281 = {{1'd0}, _EVAL_259};
  assign _EVAL_203 = {_EVAL_319, 2'h0};
  assign _EVAL_67 = _EVAL_281 | _EVAL_203;
  assign _EVAL_346 = _EVAL_67[3:2];
  assign _EVAL_275 = _EVAL_67[1:0];
  assign _EVAL_154 = _EVAL_346 & _EVAL_275;
  assign _EVAL_345 = ~ _EVAL_154;
  assign _EVAL_311 = _EVAL_345[0];
  assign _EVAL_347 = _EVAL_311 & _EVAL_23;
  assign _EVAL_240 = _EVAL_345[1];
  assign _EVAL_278 = _EVAL_240 & _EVAL_251;
  assign _EVAL_112 = {_EVAL_16,8'hff};
  assign _EVAL_82 = {{7'd0}, _EVAL_112};
  assign _EVAL_303 = _EVAL_82 << _EVAL_33;
  assign _EVAL_244 = _EVAL_303[22:8];
  assign _EVAL_420 = {_EVAL_244, 1'h0};
  assign _EVAL_199 = _EVAL_420 | 16'h1;
  assign _EVAL_398 = {1'h0,_EVAL_244};
  assign _EVAL_271 = ~ _EVAL_398;
  assign _EVAL_119 = _EVAL_199 & _EVAL_271;
  assign _EVAL_425 = _EVAL_119[15:8];
  assign _EVAL_121 = _EVAL_425 != 8'h0;
  assign _EVAL_268 = _EVAL_119[7:0];
  assign _EVAL_314 = _EVAL_425 | _EVAL_268;
  assign _EVAL_233 = _EVAL_314[7:4];
  assign _EVAL_176 = _EVAL_233 != 4'h0;
  assign _EVAL_55 = _EVAL_314[3:0];
  assign _EVAL_339 = _EVAL_233 | _EVAL_55;
  assign _EVAL_155 = _EVAL_339[3:2];
  assign _EVAL_437 = _EVAL_155 != 2'h0;
  assign _EVAL_444 = _EVAL_339[1:0];
  assign _EVAL_239 = _EVAL_155 | _EVAL_444;
  assign _EVAL_370 = _EVAL_239[1];
  assign _EVAL_135 = {_EVAL_121,_EVAL_176,_EVAL_437,_EVAL_370};
  assign _EVAL_143 = Queue_1__EVAL_2;
  assign _EVAL_147 = Queue_1__EVAL_1;
  assign _EVAL_81 = 2'h1 == _EVAL_147 ? _EVAL_232 : _EVAL_200;
  assign _EVAL_302 = 2'h2 == _EVAL_147 ? _EVAL_256 : _EVAL_81;
  assign _EVAL_163 = 2'h3 == _EVAL_147 ? _EVAL_432 : _EVAL_302;
  assign _EVAL_167 = 2'h1 == _EVAL_147 ? _EVAL_223 : _EVAL_142;
  assign _EVAL_335 = 2'h2 == _EVAL_147 ? _EVAL_156 : _EVAL_167;
  assign _EVAL_360 = 2'h3 == _EVAL_147 ? _EVAL_245 : _EVAL_335;
  assign _EVAL_249 = _EVAL_163 != _EVAL_360;
  assign _EVAL_266 = _EVAL_143 & _EVAL_249;
  assign _EVAL_395 = _EVAL_44 & _EVAL_266;
  assign _EVAL_390 = 4'h1 << _EVAL_147;
  assign _EVAL_372 = _EVAL_390[1];
  assign _EVAL_317 = _EVAL_395 & _EVAL_372;
  assign _EVAL_283 = _EVAL_30[0];
  assign _EVAL_380 = Queue__EVAL_7;
  assign _EVAL_98 = Queue_1__EVAL_8;
  assign _EVAL_192 = _EVAL_283 ? _EVAL_380 : _EVAL_98;
  assign _EVAL_297 = _EVAL_192 & _EVAL_36;
  assign _EVAL_272 = _EVAL_394 ? _EVAL_23 : 1'h0;
  assign _EVAL_331 = _EVAL_3 ^ 32'h2000000;
  assign _EVAL_304 = {1'b0,$signed(_EVAL_331)};
  assign _EVAL_337 = $signed(_EVAL_304) & $signed(-33'sh10000);
  assign _EVAL_400 = $signed(_EVAL_337);
  assign _EVAL_285 = $signed(_EVAL_400) == $signed(33'sh0);
  assign _EVAL_375 = _EVAL_3 ^ 32'h40000000;
  assign _EVAL_140 = {1'b0,$signed(_EVAL_375)};
  assign _EVAL_58 = $signed(_EVAL_140) & $signed(-33'sh2000);
  assign _EVAL_340 = $signed(_EVAL_58);
  assign _EVAL_175 = $signed(_EVAL_340) == $signed(33'sh0);
  assign _EVAL_423 = _EVAL_3 ^ 32'h80000000;
  assign _EVAL_118 = {1'b0,$signed(_EVAL_423)};
  assign _EVAL_289 = $signed(_EVAL_118) & $signed(-33'sh20000);
  assign _EVAL_442 = $signed(_EVAL_289);
  assign _EVAL_113 = $signed(_EVAL_442) == $signed(33'sh0);
  assign _EVAL_194 = _EVAL_175 | _EVAL_113;
  assign _EVAL_336 = _EVAL_3 ^ 32'hc000000;
  assign _EVAL_204 = {1'b0,$signed(_EVAL_336)};
  assign _EVAL_362 = $signed(_EVAL_204) & $signed(-33'sh4000000);
  assign _EVAL_371 = $signed(_EVAL_362);
  assign _EVAL_217 = $signed(_EVAL_371) == $signed(33'sh0);
  assign _EVAL_261 = _EVAL_194 | _EVAL_217;
  assign _EVAL_211 = _EVAL_261 | _EVAL_285;
  assign _EVAL_130 = {1'b0,$signed(_EVAL_3)};
  assign _EVAL_295 = $signed(_EVAL_130) & $signed(-33'sh5000);
  assign _EVAL_94 = $signed(_EVAL_295);
  assign _EVAL_114 = $signed(_EVAL_94) == $signed(33'sh0);
  assign _EVAL_385 = _EVAL_211 | _EVAL_114;
  assign _EVAL_165 = _EVAL_3 ^ 32'h1800000;
  assign _EVAL_359 = {1'b0,$signed(_EVAL_165)};
  assign _EVAL_64 = $signed(_EVAL_359) & $signed(-33'sh8000);
  assign _EVAL_274 = $signed(_EVAL_64);
  assign _EVAL_59 = $signed(_EVAL_274) == $signed(33'sh0);
  assign _EVAL_125 = _EVAL_385 | _EVAL_59;
  assign _EVAL_123 = _EVAL_3 ^ 32'h1900000;
  assign _EVAL_330 = {1'b0,$signed(_EVAL_123)};
  assign _EVAL_318 = $signed(_EVAL_330) & $signed(-33'sh2000);
  assign _EVAL_407 = $signed(_EVAL_318);
  assign _EVAL_182 = $signed(_EVAL_407) == $signed(33'sh0);
  assign _EVAL_416 = _EVAL_125 | _EVAL_182;
  assign _EVAL_93 = _EVAL_179 == 8'h0;
  assign _EVAL_445 = _EVAL_93 ? _EVAL_311 : _EVAL_394;
  assign _EVAL_334 = _EVAL_0 & _EVAL_445;
  assign _EVAL_169 = _EVAL_334 & _EVAL_23;
  assign _EVAL_258 = 4'h1 << _EVAL_5;
  assign _EVAL_105 = _EVAL_258[1];
  assign _EVAL_92 = _EVAL_169 & _EVAL_105;
  assign _EVAL_246 = _EVAL_254 + 3'h1;
  assign _EVAL_196 = 2'h1 == _EVAL_5 ? _EVAL_254 : _EVAL_440;
  assign _EVAL_257 = 2'h2 == _EVAL_5 ? _EVAL_325 : _EVAL_196;
  assign _EVAL_255 = 2'h3 == _EVAL_5 ? _EVAL_403 : _EVAL_257;
  assign _EVAL_77 = _EVAL_255[1:0];
  assign _EVAL_226 = _EVAL_390[0];
  assign _EVAL_363 = _EVAL_395 & _EVAL_226;
  assign _EVAL_78 = _EVAL_200 + 3'h1;
  assign _EVAL_262 = 2'h1 == _EVAL_11 ? _EVAL_223 : _EVAL_142;
  assign _EVAL_49 = 2'h2 == _EVAL_11 ? _EVAL_156 : _EVAL_262;
  assign _EVAL_280 = 2'h3 == _EVAL_11 ? _EVAL_245 : _EVAL_49;
  assign _EVAL_355 = _EVAL_280[1:0];
  assign _EVAL_195 = _EVAL_110 ? _EVAL_251 : 1'h0;
  assign _EVAL_72 = _EVAL_272 | _EVAL_195;
  assign _EVAL_219 = _EVAL_3[1:0];
  assign _EVAL_384 = {{12'd0}, _EVAL_219};
  assign _EVAL_132 = 14'h3000 | _EVAL_384;
  assign _EVAL_315 = _EVAL_390[3];
  assign _EVAL_83 = _EVAL_395 & _EVAL_315;
  assign _EVAL_441 = _EVAL_23 | _EVAL_251;
  assign _EVAL_48 = 23'hff << _EVAL_38;
  assign _EVAL_422 = _EVAL_48[7:0];
  assign _EVAL_54 = ~ _EVAL_422;
  assign _EVAL_443 = _EVAL_32 | _EVAL_6;
  assign _EVAL_208 = _EVAL_93 ? _EVAL_240 : _EVAL_110;
  assign _EVAL_152 = _EVAL_0 & _EVAL_208;
  assign _EVAL_187 = _EVAL_3 ^ 32'h20000000;
  assign _EVAL_215 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_198 = $signed(_EVAL_215) & $signed(-33'sh2000);
  assign _EVAL_279 = $signed(_EVAL_198);
  assign _EVAL_120 = $signed(_EVAL_279) == $signed(33'sh0);
  assign _EVAL_367 = _EVAL_416 | _EVAL_120;
  assign _EVAL_61 = 4'h1 << _EVAL_11;
  assign _EVAL_320 = _EVAL_152 & _EVAL_15;
  assign _EVAL_411 = _EVAL_320 & _EVAL_35;
  assign _EVAL_214 = _EVAL_411 & _EVAL_26;
  assign _EVAL_414 = _EVAL_61[2];
  assign _EVAL_171 = _EVAL_214 & _EVAL_414;
  assign _EVAL_68 = _EVAL_258[3];
  assign _EVAL_146 = _EVAL_54[7:2];
  assign _EVAL_65 = _EVAL_93 ? _EVAL_441 : _EVAL_72;
  assign _EVAL_386 = _EVAL_0 & _EVAL_65;
  assign _EVAL_184 = {{7'd0}, _EVAL_386};
  assign _EVAL_399 = _EVAL_169 & _EVAL_68;
  assign _EVAL_206 = _EVAL_403 + 3'h1;
  assign _EVAL_191 = _EVAL_93 ? _EVAL_347 : _EVAL_394;
  assign _EVAL_160 = _EVAL_232 + 3'h1;
  assign _EVAL_368 = _EVAL_135 <= 4'h6;
  assign _EVAL_299 = _EVAL_368 & _EVAL_367;
  assign _EVAL_95 = _EVAL_61[0];
  assign _EVAL_180 = _EVAL_214 & _EVAL_95;
  assign _EVAL_47 = _EVAL_142 + 3'h1;
  assign _EVAL_51 = _EVAL_90 != 2'h0;
  assign _EVAL_276 = _EVAL_135 <= 4'h8;
  assign _EVAL_89 = _EVAL_3 ^ 32'h3000;
  assign _EVAL_352 = {1'b0,$signed(_EVAL_89)};
  assign _EVAL_338 = $signed(_EVAL_352) & $signed(-33'sh1000);
  assign _EVAL_205 = $signed(_EVAL_338);
  assign _EVAL_447 = $signed(_EVAL_205) == $signed(33'sh0);
  assign _EVAL_267 = _EVAL_276 & _EVAL_447;
  assign _EVAL_70 = _EVAL_299 | _EVAL_267;
  assign _EVAL_97 = _EVAL_70 ? _EVAL_3 : {{18'd0}, _EVAL_132};
  assign _EVAL_212 = _EVAL_426 & _EVAL_277;
  assign _EVAL_129 = _EVAL_148 | _EVAL_212;
  assign _EVAL_159 = _EVAL_277 & _EVAL_99;
  assign _EVAL_145 = _EVAL_225 & _EVAL_159;
  assign _EVAL_224 = _EVAL_129 | _EVAL_145;
  assign _EVAL_393 = _EVAL_277 & _EVAL_327;
  assign _EVAL_236 = _EVAL_225 & _EVAL_393;
  assign _EVAL_227 = _EVAL_129 | _EVAL_236;
  assign _EVAL_185 = _EVAL_342 & _EVAL_99;
  assign _EVAL_312 = _EVAL_225 & _EVAL_185;
  assign _EVAL_100 = _EVAL_101 | _EVAL_312;
  assign _EVAL_356 = {_EVAL_164,_EVAL_224,_EVAL_227,_EVAL_100,_EVAL_300,33'h0};
  assign _EVAL_369 = {6'h20,_EVAL_242,_EVAL_402,_EVAL_313,_EVAL_222,_EVAL_5,_EVAL_77,1'h0,_EVAL_356};
  assign _EVAL_431 = _EVAL_191 ? _EVAL_369 : 84'h0;
  assign _EVAL_69 = _EVAL_390[2];
  assign _EVAL_63 = _EVAL_395 & _EVAL_69;
  assign _EVAL_116 = _EVAL_256 + 3'h1;
  assign _EVAL_243 = _EVAL_298 == 6'h0;
  assign _EVAL_263 = _EVAL_283 ? _EVAL_146 : 6'h0;
  assign _EVAL_106 = _EVAL_298 - 6'h1;
  assign _EVAL_264 = _EVAL_432 + 3'h1;
  assign _EVAL_305 = _EVAL_223 + 3'h1;
  assign _EVAL_86 = _EVAL_93 ? _EVAL_278 : _EVAL_110;
  assign _EVAL_328 = {_EVAL_97,_EVAL_42,_EVAL_4,1'h0};
  assign _EVAL_71 = {6'h8,_EVAL_121,_EVAL_176,_EVAL_437,_EVAL_370,_EVAL_11,_EVAL_355,1'h1,_EVAL_328};
  assign _EVAL_357 = _EVAL_86 ? _EVAL_71 : 84'h0;
  assign _EVAL_439 = _EVAL_258[0];
  assign _EVAL_136 = _EVAL_258[2];
  assign _EVAL_221 = _EVAL_169 & _EVAL_136;
  assign _EVAL_172 = _EVAL_345 & _EVAL_90;
  assign _EVAL_228 = {_EVAL_172, 1'h0};
  assign _EVAL_62 = _EVAL_179 - _EVAL_184;
  assign _EVAL_230 = _EVAL_169 & _EVAL_439;
  assign _EVAL_124 = _EVAL_440 + 3'h1;
  assign _EVAL_291 = _EVAL_298 == 6'h1;
  assign _EVAL_410 = _EVAL_228[1:0];
  assign _EVAL_406 = _EVAL_61[3];
  assign _EVAL_433 = _EVAL_325 + 3'h1;
  assign _EVAL_412 = _EVAL_263 == 6'h0;
  assign _EVAL_376 = _EVAL_214 & _EVAL_406;
  assign _EVAL_353 = _EVAL_245 + 3'h1;
  assign _EVAL_178 = _EVAL_61[1];
  assign _EVAL_173 = _EVAL_214 & _EVAL_178;
  assign _EVAL_115 = _EVAL_93 & _EVAL_0;
  assign _EVAL_292 = _EVAL_156 + 3'h1;
  assign _EVAL_323 = _EVAL_115 & _EVAL_51;
  assign _EVAL_287 = _EVAL_172 | _EVAL_410;
  assign _EVAL_429 = _EVAL_283 == 1'h0;
  assign _EVAL_134 = _EVAL_431 | _EVAL_357;
  assign Queue_1__EVAL_6 = _EVAL_24;
  assign Queue__EVAL_3 = _EVAL_291 | _EVAL_412;
  assign _EVAL = Queue__EVAL_6;
  assign _EVAL_29 = _EVAL_134[68:37];
  assign Queue_1__EVAL_3 = _EVAL_28;
  assign _EVAL_19 = _EVAL_320 & _EVAL_35;
  assign _EVAL_45 = Queue_1__EVAL_1;
  assign _EVAL_18 = _EVAL_134[83:81];
  assign _EVAL_14 = _EVAL_134[32:1];
  assign Queue__EVAL_8 = _EVAL_24;
  assign _EVAL_7 = _EVAL_134[0];
  assign _EVAL_37 = Queue_1__EVAL_0;
  assign _EVAL_40 = _EVAL_283 ? _EVAL_380 : _EVAL_98;
  assign _EVAL_21 = _EVAL_143 & _EVAL_249;
  assign _EVAL_9 = _EVAL_134[73:69];
  assign Queue_1__EVAL_5 = _EVAL_13[4:3];
  assign Queue_1__EVAL = _EVAL_44 & _EVAL_249;
  assign _EVAL_20 = _EVAL_134[77:74];
  assign Queue__EVAL_11 = _EVAL_2;
  assign _EVAL_34 = Queue__EVAL_2;
  assign _EVAL_10 = _EVAL_152 & _EVAL_26;
  assign _EVAL_43 = Queue__EVAL_4;
  assign Queue__EVAL = _EVAL_28;
  assign Queue_1__EVAL_7 = _EVAL_36 & _EVAL_429;
  assign Queue__EVAL_9 = _EVAL_443 ? 2'h2 : 2'h0;
  assign _EVAL_31 = _EVAL_93 ? _EVAL_441 : _EVAL_72;
  assign _EVAL_39 = Queue__EVAL_5;
  assign Queue__EVAL_0 = _EVAL_36 & _EVAL_283;
  assign _EVAL_27 = _EVAL_134[80:78];
  assign Queue_1__EVAL_4 = _EVAL_443 ? 2'h2 : 2'h0;
  assign _EVAL_17 = _EVAL_0 & _EVAL_445;
  assign Queue__EVAL_10 = _EVAL_13[4:3];
  assign _EVAL_8 = _EVAL_134[36:33];
  assign Queue__EVAL_12 = _EVAL_1;
  assign _EVAL_41 = Queue__EVAL_1;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_110 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_142 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_156 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_179 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_200 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_223 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_232 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_245 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_254 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_256 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_298 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_319 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_325 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_394 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_403 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_432 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_440 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_24) begin
    if (_EVAL_28) begin
      _EVAL_110 <= 1'h0;
    end else begin
      if (_EVAL_93) begin
        _EVAL_110 <= _EVAL_278;
      end
    end
    if (_EVAL_28) begin
      _EVAL_142 <= 3'h0;
    end else begin
      if (_EVAL_180) begin
        _EVAL_142 <= _EVAL_47;
      end
    end
    if (_EVAL_28) begin
      _EVAL_156 <= 3'h0;
    end else begin
      if (_EVAL_171) begin
        _EVAL_156 <= _EVAL_292;
      end
    end
    if (_EVAL_28) begin
      _EVAL_179 <= 8'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_278) begin
          _EVAL_179 <= _EVAL_16;
        end else begin
          _EVAL_179 <= 8'h0;
        end
      end else begin
        _EVAL_179 <= _EVAL_62;
      end
    end
    if (_EVAL_28) begin
      _EVAL_200 <= 3'h0;
    end else begin
      if (_EVAL_363) begin
        _EVAL_200 <= _EVAL_78;
      end
    end
    if (_EVAL_28) begin
      _EVAL_223 <= 3'h0;
    end else begin
      if (_EVAL_173) begin
        _EVAL_223 <= _EVAL_305;
      end
    end
    if (_EVAL_28) begin
      _EVAL_232 <= 3'h0;
    end else begin
      if (_EVAL_317) begin
        _EVAL_232 <= _EVAL_160;
      end
    end
    if (_EVAL_28) begin
      _EVAL_245 <= 3'h0;
    end else begin
      if (_EVAL_376) begin
        _EVAL_245 <= _EVAL_353;
      end
    end
    if (_EVAL_28) begin
      _EVAL_254 <= 3'h0;
    end else begin
      if (_EVAL_92) begin
        _EVAL_254 <= _EVAL_246;
      end
    end
    if (_EVAL_28) begin
      _EVAL_256 <= 3'h0;
    end else begin
      if (_EVAL_63) begin
        _EVAL_256 <= _EVAL_116;
      end
    end
    if (_EVAL_28) begin
      _EVAL_298 <= 6'h0;
    end else begin
      if (_EVAL_297) begin
        if (_EVAL_243) begin
          if (_EVAL_283) begin
            _EVAL_298 <= _EVAL_146;
          end else begin
            _EVAL_298 <= 6'h0;
          end
        end else begin
          _EVAL_298 <= _EVAL_106;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_319 <= 2'h3;
    end else begin
      if (_EVAL_323) begin
        _EVAL_319 <= _EVAL_287;
      end
    end
    if (_EVAL_28) begin
      _EVAL_325 <= 3'h0;
    end else begin
      if (_EVAL_221) begin
        _EVAL_325 <= _EVAL_433;
      end
    end
    if (_EVAL_28) begin
      _EVAL_394 <= 1'h0;
    end else begin
      if (_EVAL_93) begin
        _EVAL_394 <= _EVAL_347;
      end
    end
    if (_EVAL_28) begin
      _EVAL_403 <= 3'h0;
    end else begin
      if (_EVAL_399) begin
        _EVAL_403 <= _EVAL_206;
      end
    end
    if (_EVAL_28) begin
      _EVAL_432 <= 3'h0;
    end else begin
      if (_EVAL_83) begin
        _EVAL_432 <= _EVAL_264;
      end
    end
    if (_EVAL_28) begin
      _EVAL_440 <= 3'h0;
    end else begin
      if (_EVAL_230) begin
        _EVAL_440 <= _EVAL_124;
      end
    end
  end
endmodule
