//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_309(
  input          _EVAL,
  output         _EVAL_0,
  input  [1:0]   _EVAL_1,
  output         _EVAL_2,
  output [2:0]   _EVAL_3,
  output         _EVAL_4,
  input          _EVAL_5,
  output         _EVAL_6,
  input          _EVAL_7,
  output         _EVAL_8,
  output [4:0]   _EVAL_9,
  input          _EVAL_10,
  input          _EVAL_11,
  input          _EVAL_12,
  output [4:0]   _EVAL_13,
  input          _EVAL_14,
  input          _EVAL_15,
  input          _EVAL_16,
  output         _EVAL_17,
  output [2:0]   _EVAL_18,
  input          _EVAL_19,
  output         _EVAL_20,
  output         _EVAL_21,
  output         _EVAL_22,
  input  [127:0] _EVAL_23,
  output [14:0]  _EVAL_24,
  input          _EVAL_25,
  output         _EVAL_26,
  output [4:0]   _EVAL_27,
  input          _EVAL_28,
  input  [127:0] _EVAL_29,
  output [2:0]   _EVAL_30,
  input  [4:0]   _EVAL_31,
  input          _EVAL_32,
  input          _EVAL_33,
  output         _EVAL_34,
  input          _EVAL_35,
  input          _EVAL_36,
  input          _EVAL_37,
  output         _EVAL_38,
  input  [14:0]  _EVAL_39,
  output         _EVAL_40,
  input  [14:0]  _EVAL_41,
  input          _EVAL_42,
  output         _EVAL_43,
  input          _EVAL_44,
  output         _EVAL_45,
  input          _EVAL_46,
  input  [2:0]   _EVAL_47,
  input  [4:0]   _EVAL_48,
  output         _EVAL_49,
  input          _EVAL_50,
  input          _EVAL_51,
  output         _EVAL_52,
  output         _EVAL_53,
  input          _EVAL_54,
  input          _EVAL_55,
  output         _EVAL_56,
  output         _EVAL_57,
  input  [4:0]   _EVAL_58,
  output         _EVAL_59,
  input          _EVAL_60,
  output         _EVAL_61,
  input  [4:0]   _EVAL_62,
  input  [6:0]   _EVAL_63,
  input          _EVAL_64,
  output         _EVAL_65,
  output         _EVAL_66,
  output         _EVAL_67,
  input          _EVAL_68,
  output [1:0]   _EVAL_69,
  output         _EVAL_70,
  input          _EVAL_71,
  input  [8:0]   _EVAL_72,
  output         _EVAL_73,
  output [4:0]   _EVAL_74,
  input          _EVAL_75,
  input          _EVAL_76,
  output [31:0]  _EVAL_77,
  output         _EVAL_78,
  output         _EVAL_79,
  input          _EVAL_80,
  output         _EVAL_81,
  input  [2:0]   _EVAL_82,
  output         _EVAL_83,
  output         _EVAL_84,
  output         _EVAL_85,
  input          _EVAL_86,
  input          _EVAL_87,
  input  [4:0]   _EVAL_88,
  input          _EVAL_89,
  output         _EVAL_90,
  output [4:0]   _EVAL_91,
  input  [2:0]   _EVAL_92,
  output         _EVAL_93,
  output         _EVAL_94,
  input          _EVAL_95,
  output         _EVAL_96,
  input          _EVAL_97,
  output [127:0] _EVAL_98,
  input          _EVAL_99,
  input          _EVAL_100,
  input  [2:0]   _EVAL_101,
  input  [31:0]  _EVAL_102,
  input  [1:0]   _EVAL_103,
  input          _EVAL_104,
  input          _EVAL_105,
  output         _EVAL_106,
  input  [8:0]   _EVAL_107,
  input          _EVAL_108,
  output [4:0]   _EVAL_109,
  input          _EVAL_110,
  output         _EVAL_111,
  output         _EVAL_112,
  output         _EVAL_113,
  input          _EVAL_114,
  input          _EVAL_115,
  input          _EVAL_116,
  input  [4:0]   _EVAL_117,
  output         _EVAL_118,
  input          _EVAL_119,
  input          _EVAL_120,
  output         _EVAL_121,
  input          _EVAL_122,
  output         _EVAL_123,
  output         _EVAL_124,
  output [14:0]  _EVAL_125,
  input  [2:0]   _EVAL_126,
  input  [31:0]  _EVAL_127,
  output [2:0]   _EVAL_128,
  output [6:0]   _EVAL_129,
  input          _EVAL_130,
  input          _EVAL_131,
  output         _EVAL_132,
  output [4:0]   _EVAL_133,
  output         _EVAL_134,
  input          _EVAL_135,
  output         _EVAL_136,
  input          _EVAL_137,
  output         _EVAL_138,
  input          _EVAL_139,
  output         _EVAL_140,
  output [4:0]   _EVAL_141,
  input          _EVAL_142,
  input          _EVAL_143,
  output         _EVAL_144,
  output [1:0]   _EVAL_145,
  output [31:0]  _EVAL_146,
  input          _EVAL_147,
  input  [6:0]   _EVAL_148,
  input  [2:0]   _EVAL_149,
  input          _EVAL_150,
  input          _EVAL_151,
  output [127:0] _EVAL_152,
  input          _EVAL_153,
  input  [4:0]   _EVAL_154,
  output         _EVAL_155,
  input          _EVAL_156,
  input          _EVAL_157,
  input          _EVAL_158,
  output         _EVAL_159,
  output         _EVAL_160,
  input          _EVAL_161,
  output         _EVAL_162,
  output [2:0]   _EVAL_163,
  input          _EVAL_164,
  output         _EVAL_165,
  output         _EVAL_166,
  input          _EVAL_167,
  input          _EVAL_168,
  input  [4:0]   _EVAL_169,
  output         _EVAL_170,
  output [6:0]   _EVAL_171,
  input          _EVAL_172,
  output         _EVAL_173,
  input          _EVAL_174,
  input          _EVAL_175,
  output         _EVAL_176,
  input          _EVAL_177,
  input          _EVAL_178,
  output         _EVAL_179,
  output         _EVAL_180,
  input          _EVAL_181,
  output         _EVAL_182,
  output [2:0]   _EVAL_183,
  input          _EVAL_184,
  output         _EVAL_185
);
  reg  _EVAL_186;
  reg [31:0] _RAND_0;
  reg [4:0] _EVAL_187;
  reg [31:0] _RAND_1;
  reg  _EVAL_188;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_192;
  reg [31:0] _RAND_3;
  reg  _EVAL_194;
  reg [31:0] _RAND_4;
  reg [31:0] _EVAL_196;
  reg [31:0] _RAND_5;
  reg [6:0] _EVAL_197;
  reg [31:0] _RAND_6;
  reg  _EVAL_199;
  reg [31:0] _RAND_7;
  reg  _EVAL_200;
  reg [31:0] _RAND_8;
  reg  _EVAL_201;
  reg [31:0] _RAND_9;
  reg  _EVAL_202;
  reg [31:0] _RAND_10;
  reg  _EVAL_203;
  reg [31:0] _RAND_11;
  reg  _EVAL_209;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_210;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_211;
  reg [31:0] _RAND_14;
  reg  _EVAL_215;
  reg [31:0] _RAND_15;
  reg [4:0] _EVAL_217;
  reg [31:0] _RAND_16;
  reg  _EVAL_218;
  reg [31:0] _RAND_17;
  reg  _EVAL_219;
  reg [31:0] _RAND_18;
  reg  _EVAL_221;
  reg [31:0] _RAND_19;
  reg  _EVAL_222;
  reg [31:0] _RAND_20;
  reg  _EVAL_223;
  reg [31:0] _RAND_21;
  reg [14:0] _EVAL_225;
  reg [31:0] _RAND_22;
  reg  _EVAL_229;
  reg [31:0] _RAND_23;
  reg [4:0] _EVAL_233;
  reg [31:0] _RAND_24;
  reg  _EVAL_234;
  reg [31:0] _RAND_25;
  reg  _EVAL_235;
  reg [31:0] _RAND_26;
  reg  _EVAL_237;
  reg [31:0] _RAND_27;
  reg  _EVAL_239;
  reg [31:0] _RAND_28;
  reg [31:0] _EVAL_240;
  reg [31:0] _RAND_29;
  reg  _EVAL_241;
  reg [31:0] _RAND_30;
  reg  _EVAL_242;
  reg [31:0] _RAND_31;
  reg  _EVAL_243;
  reg [31:0] _RAND_32;
  reg  _EVAL_244;
  reg [31:0] _RAND_33;
  reg  _EVAL_246;
  reg [31:0] _RAND_34;
  reg  _EVAL_247;
  reg [31:0] _RAND_35;
  reg  _EVAL_248;
  reg [31:0] _RAND_36;
  reg [4:0] _EVAL_251;
  reg [31:0] _RAND_37;
  reg [4:0] _EVAL_252;
  reg [31:0] _RAND_38;
  reg  _EVAL_254;
  reg [31:0] _RAND_39;
  reg  _EVAL_255;
  reg [31:0] _RAND_40;
  reg  _EVAL_256;
  reg [31:0] _RAND_41;
  reg [2:0] _EVAL_257;
  reg [31:0] _RAND_42;
  reg [4:0] _EVAL_259;
  reg [31:0] _RAND_43;
  reg [2:0] _EVAL_260;
  reg [31:0] _RAND_44;
  reg  _EVAL_263;
  reg [31:0] _RAND_45;
  reg  _EVAL_264;
  reg [31:0] _RAND_46;
  reg [31:0] _EVAL_267;
  reg [31:0] _RAND_47;
  reg  _EVAL_268;
  reg [31:0] _RAND_48;
  reg  _EVAL_269;
  reg [31:0] _RAND_49;
  reg  _EVAL_270;
  reg [31:0] _RAND_50;
  reg  _EVAL_271;
  reg [31:0] _RAND_51;
  reg  _EVAL_272;
  reg [31:0] _RAND_52;
  reg [31:0] _EVAL_274;
  reg [31:0] _RAND_53;
  reg  _EVAL_277;
  reg [31:0] _RAND_54;
  reg  _EVAL_278;
  reg [31:0] _RAND_55;
  reg [1:0] _EVAL_279;
  reg [31:0] _RAND_56;
  reg  _EVAL_280;
  reg [31:0] _RAND_57;
  reg  _EVAL_282;
  reg [31:0] _RAND_58;
  reg [2:0] _EVAL_284;
  reg [31:0] _RAND_59;
  reg  _EVAL_285;
  reg [31:0] _RAND_60;
  reg  _EVAL_286;
  reg [31:0] _RAND_61;
  reg  _EVAL_288;
  reg [31:0] _RAND_62;
  reg  _EVAL_289;
  reg [31:0] _RAND_63;
  reg  _EVAL_291;
  reg [31:0] _RAND_64;
  reg  _EVAL_294;
  reg [31:0] _RAND_65;
  reg  _EVAL_296;
  reg [31:0] _RAND_66;
  reg [6:0] _EVAL_297;
  reg [31:0] _RAND_67;
  reg  _EVAL_301;
  reg [31:0] _RAND_68;
  reg  _EVAL_302;
  reg [31:0] _RAND_69;
  reg  _EVAL_303;
  reg [31:0] _RAND_70;
  reg  _EVAL_304;
  reg [31:0] _RAND_71;
  reg  _EVAL_306;
  reg [31:0] _RAND_72;
  reg  _EVAL_307;
  reg [31:0] _RAND_73;
  reg  _EVAL_308;
  reg [31:0] _RAND_74;
  reg  _EVAL_309;
  reg [31:0] _RAND_75;
  reg  _EVAL_311;
  reg [31:0] _RAND_76;
  reg  _EVAL_312;
  reg [31:0] _RAND_77;
  reg  _EVAL_313;
  reg [31:0] _RAND_78;
  reg  _EVAL_315;
  reg [31:0] _RAND_79;
  reg [2:0] _EVAL_316;
  reg [31:0] _RAND_80;
  reg [8:0] _EVAL_317;
  reg [31:0] _RAND_81;
  reg  _EVAL_318;
  reg [31:0] _RAND_82;
  reg  _EVAL_322;
  reg [31:0] _RAND_83;
  reg  _EVAL_323;
  reg [31:0] _RAND_84;
  reg [31:0] _EVAL_328;
  reg [31:0] _RAND_85;
  reg  _EVAL_330;
  reg [31:0] _RAND_86;
  reg  _EVAL_331;
  reg [31:0] _RAND_87;
  reg  _EVAL_332;
  reg [31:0] _RAND_88;
  reg  _EVAL_333;
  reg [31:0] _RAND_89;
  reg  _EVAL_335;
  reg [31:0] _RAND_90;
  reg [2:0] _EVAL_336;
  reg [31:0] _RAND_91;
  reg [2:0] _EVAL_337;
  reg [31:0] _RAND_92;
  reg [4:0] _EVAL_338;
  reg [31:0] _RAND_93;
  reg  _EVAL_339;
  reg [31:0] _RAND_94;
  reg [127:0] _EVAL_340;
  reg [127:0] _RAND_95;
  reg [2:0] _EVAL_342;
  reg [31:0] _RAND_96;
  reg [2:0] _EVAL_343;
  reg [31:0] _RAND_97;
  reg  _EVAL_345;
  reg [31:0] _RAND_98;
  reg  _EVAL_346;
  reg [31:0] _RAND_99;
  reg [127:0] _EVAL_348;
  reg [127:0] _RAND_100;
  reg  _EVAL_349;
  reg [31:0] _RAND_101;
  reg  _EVAL_350;
  reg [31:0] _RAND_102;
  reg  _EVAL_352;
  reg [31:0] _RAND_103;
  reg  _EVAL_353;
  reg [31:0] _RAND_104;
  reg  _EVAL_355;
  reg [31:0] _RAND_105;
  reg  _EVAL_356;
  reg [31:0] _RAND_106;
  reg  _EVAL_358;
  reg [31:0] _RAND_107;
  reg [2:0] _EVAL_360;
  reg [31:0] _RAND_108;
  reg  _EVAL_361;
  reg [31:0] _RAND_109;
  reg  _EVAL_363;
  reg [31:0] _RAND_110;
  reg  _EVAL_365;
  reg [31:0] _RAND_111;
  reg  _EVAL_366;
  reg [31:0] _RAND_112;
  reg [4:0] _EVAL_368;
  reg [31:0] _RAND_113;
  reg  _EVAL_371;
  reg [31:0] _RAND_114;
  reg [8:0] _EVAL_372;
  reg [31:0] _RAND_115;
  reg  _EVAL_374;
  reg [31:0] _RAND_116;
  reg  _EVAL_375;
  reg [31:0] _RAND_117;
  reg  _EVAL_376;
  reg [31:0] _RAND_118;
  reg [31:0] _EVAL_377;
  reg [31:0] _RAND_119;
  reg  _EVAL_387;
  reg [31:0] _RAND_120;
  reg  _EVAL_388;
  reg [31:0] _RAND_121;
  reg  _EVAL_389;
  reg [31:0] _RAND_122;
  reg [4:0] _EVAL_390;
  reg [31:0] _RAND_123;
  reg [6:0] _EVAL_391;
  reg [31:0] _RAND_124;
  reg  _EVAL_392;
  reg [31:0] _RAND_125;
  reg [4:0] _EVAL_393;
  reg [31:0] _RAND_126;
  reg  _EVAL_398;
  reg [31:0] _RAND_127;
  reg  _EVAL_400;
  reg [31:0] _RAND_128;
  reg [6:0] _EVAL_402;
  reg [31:0] _RAND_129;
  reg  _EVAL_413;
  reg [31:0] _RAND_130;
  reg  _EVAL_414;
  reg [31:0] _RAND_131;
  reg  _EVAL_415;
  reg [31:0] _RAND_132;
  reg  _EVAL_416;
  reg [31:0] _RAND_133;
  reg [2:0] _EVAL_420;
  reg [31:0] _RAND_134;
  reg  _EVAL_421;
  reg [31:0] _RAND_135;
  reg  _EVAL_422;
  reg [31:0] _RAND_136;
  reg [4:0] _EVAL_424;
  reg [31:0] _RAND_137;
  reg [4:0] _EVAL_425;
  reg [31:0] _RAND_138;
  reg  _EVAL_426;
  reg [31:0] _RAND_139;
  reg [14:0] _EVAL_428;
  reg [31:0] _RAND_140;
  reg  _EVAL_429;
  reg [31:0] _RAND_141;
  reg  _EVAL_430;
  reg [31:0] _RAND_142;
  reg [2:0] _EVAL_431;
  reg [31:0] _RAND_143;
  reg  _EVAL_433;
  reg [31:0] _RAND_144;
  reg [127:0] _EVAL_434;
  reg [127:0] _RAND_145;
  reg  _EVAL_436;
  reg [31:0] _RAND_146;
  reg [6:0] _EVAL_439;
  reg [31:0] _RAND_147;
  reg [4:0] _EVAL_440;
  reg [31:0] _RAND_148;
  reg  _EVAL_442;
  reg [31:0] _RAND_149;
  reg  _EVAL_444;
  reg [31:0] _RAND_150;
  reg  _EVAL_445;
  reg [31:0] _RAND_151;
  reg  _EVAL_447;
  reg [31:0] _RAND_152;
  reg [1:0] _EVAL_451;
  reg [31:0] _RAND_153;
  reg  _EVAL_453;
  reg [31:0] _RAND_154;
  reg  _EVAL_455;
  reg [31:0] _RAND_155;
  reg [2:0] _EVAL_456;
  reg [31:0] _RAND_156;
  reg  _EVAL_457;
  reg [31:0] _RAND_157;
  reg  _EVAL_460;
  reg [31:0] _RAND_158;
  reg  _EVAL_461;
  reg [31:0] _RAND_159;
  reg [2:0] _EVAL_467;
  reg [31:0] _RAND_160;
  reg [6:0] _EVAL_468;
  reg [31:0] _RAND_161;
  reg  _EVAL_470;
  reg [31:0] _RAND_162;
  reg [127:0] _EVAL_471;
  reg [127:0] _RAND_163;
  reg [127:0] _EVAL_472;
  reg [127:0] _RAND_164;
  reg  _EVAL_473;
  reg [31:0] _RAND_165;
  reg [4:0] _EVAL_474;
  reg [31:0] _RAND_166;
  reg  _EVAL_475;
  reg [31:0] _RAND_167;
  reg  _EVAL_476;
  reg [31:0] _RAND_168;
  reg  _EVAL_479;
  reg [31:0] _RAND_169;
  reg  _EVAL_480;
  reg [31:0] _RAND_170;
  reg  _EVAL_482;
  reg [31:0] _RAND_171;
  reg  _EVAL_484;
  reg [31:0] _RAND_172;
  reg  _EVAL_488;
  reg [31:0] _RAND_173;
  reg  _EVAL_489;
  reg [31:0] _RAND_174;
  reg [1:0] _EVAL_490;
  reg [31:0] _RAND_175;
  reg  _EVAL_491;
  reg [31:0] _RAND_176;
  reg  _EVAL_494;
  reg [31:0] _RAND_177;
  reg  _EVAL_497;
  reg [31:0] _RAND_178;
  reg [14:0] _EVAL_498;
  reg [31:0] _RAND_179;
  reg  _EVAL_499;
  reg [31:0] _RAND_180;
  reg  _EVAL_500;
  reg [31:0] _RAND_181;
  reg  _EVAL_502;
  reg [31:0] _RAND_182;
  reg  _EVAL_504;
  reg [31:0] _RAND_183;
  reg  _EVAL_505;
  reg [31:0] _RAND_184;
  reg  _EVAL_507;
  reg [31:0] _RAND_185;
  reg  _EVAL_508;
  reg [31:0] _RAND_186;
  reg [4:0] _EVAL_509;
  reg [31:0] _RAND_187;
  reg  _EVAL_510;
  reg [31:0] _RAND_188;
  reg  _EVAL_511;
  reg [31:0] _RAND_189;
  reg [2:0] _EVAL_513;
  reg [31:0] _RAND_190;
  reg [127:0] _EVAL_515;
  reg [127:0] _RAND_191;
  reg  _EVAL_517;
  reg [31:0] _RAND_192;
  reg  _EVAL_518;
  reg [31:0] _RAND_193;
  reg  _EVAL_519;
  reg [31:0] _RAND_194;
  reg  _EVAL_521;
  reg [31:0] _RAND_195;
  reg  _EVAL_522;
  reg [31:0] _RAND_196;
  reg [127:0] _EVAL_524;
  reg [127:0] _RAND_197;
  reg  _EVAL_525;
  reg [31:0] _RAND_198;
  reg [4:0] _EVAL_527;
  reg [31:0] _RAND_199;
  reg  _EVAL_528;
  reg [31:0] _RAND_200;
  reg  _EVAL_530;
  reg [31:0] _RAND_201;
  reg  _EVAL_533;
  reg [31:0] _RAND_202;
  reg  _EVAL_534;
  reg [31:0] _RAND_203;
  reg [31:0] _EVAL_536;
  reg [31:0] _RAND_204;
  reg  _EVAL_537;
  reg [31:0] _RAND_205;
  reg [1:0] _EVAL_538;
  reg [31:0] _RAND_206;
  reg [2:0] _EVAL_541;
  reg [31:0] _RAND_207;
  reg  _EVAL_545;
  reg [31:0] _RAND_208;
  reg  _EVAL_546;
  reg [31:0] _RAND_209;
  reg  _EVAL_547;
  reg [31:0] _RAND_210;
  reg [127:0] _EVAL_548;
  reg [127:0] _RAND_211;
  reg  _EVAL_551;
  reg [31:0] _RAND_212;
  reg  _EVAL_554;
  reg [31:0] _RAND_213;
  reg  _EVAL_555;
  reg [31:0] _RAND_214;
  reg  _EVAL_556;
  reg [31:0] _RAND_215;
  reg  _EVAL_558;
  reg [31:0] _RAND_216;
  reg [2:0] _EVAL_559;
  reg [31:0] _RAND_217;
  reg  _EVAL_560;
  reg [31:0] _RAND_218;
  reg  _EVAL_561;
  reg [31:0] _RAND_219;
  reg  _EVAL_562;
  reg [31:0] _RAND_220;
  reg  _EVAL_563;
  reg [31:0] _RAND_221;
  reg  _EVAL_564;
  reg [31:0] _RAND_222;
  reg  _EVAL_565;
  reg [31:0] _RAND_223;
  reg  _EVAL_566;
  reg [31:0] _RAND_224;
  reg  _EVAL_568;
  reg [31:0] _RAND_225;
  reg [4:0] _EVAL_569;
  reg [31:0] _RAND_226;
  reg [4:0] _EVAL_571;
  reg [31:0] _RAND_227;
  reg  _EVAL_573;
  reg [31:0] _RAND_228;
  reg [4:0] _EVAL_574;
  reg [31:0] _RAND_229;
  reg [14:0] _EVAL_576;
  reg [31:0] _RAND_230;
  reg  _EVAL_579;
  reg [31:0] _RAND_231;
  reg  _EVAL_580;
  reg [31:0] _RAND_232;
  reg  _EVAL_581;
  reg [31:0] _RAND_233;
  reg  _EVAL_582;
  reg [31:0] _RAND_234;
  reg  _EVAL_584;
  reg [31:0] _RAND_235;
  reg  _EVAL_587;
  reg [31:0] _RAND_236;
  reg  _EVAL_589;
  reg [31:0] _RAND_237;
  reg  _EVAL_591;
  reg [31:0] _RAND_238;
  reg [4:0] _EVAL_593;
  reg [31:0] _RAND_239;
  reg  _EVAL_594;
  reg [31:0] _RAND_240;
  reg  _EVAL_596;
  reg [31:0] _RAND_241;
  reg  _EVAL_597;
  reg [31:0] _RAND_242;
  reg  _EVAL_598;
  reg [31:0] _RAND_243;
  reg  _EVAL_599;
  reg [31:0] _RAND_244;
  reg  _EVAL_600;
  reg [31:0] _RAND_245;
  reg  _EVAL_601;
  reg [31:0] _RAND_246;
  reg [4:0] _EVAL_602;
  reg [31:0] _RAND_247;
  reg [8:0] _EVAL_603;
  reg [31:0] _RAND_248;
  reg  _EVAL_604;
  reg [31:0] _RAND_249;
  reg  _EVAL_606;
  reg [31:0] _RAND_250;
  reg  _EVAL_607;
  reg [31:0] _RAND_251;
  reg  _EVAL_608;
  reg [31:0] _RAND_252;
  reg  _EVAL_609;
  reg [31:0] _RAND_253;
  reg  _EVAL_611;
  reg [31:0] _RAND_254;
  reg  _EVAL_612;
  reg [31:0] _RAND_255;
  reg  _EVAL_614;
  reg [31:0] _RAND_256;
  reg  _EVAL_615;
  reg [31:0] _RAND_257;
  reg  _EVAL_618;
  reg [31:0] _RAND_258;
  reg  _EVAL_619;
  reg [31:0] _RAND_259;
  reg  _EVAL_620;
  reg [31:0] _RAND_260;
  reg [2:0] _EVAL_621;
  reg [31:0] _RAND_261;
  reg  _EVAL_622;
  reg [31:0] _RAND_262;
  reg [4:0] _EVAL_623;
  reg [31:0] _RAND_263;
  reg  _EVAL_625;
  reg [31:0] _RAND_264;
  reg  _EVAL_626;
  reg [31:0] _RAND_265;
  reg  _EVAL_630;
  reg [31:0] _RAND_266;
  reg  _EVAL_633;
  reg [31:0] _RAND_267;
  reg [6:0] _EVAL_634;
  reg [31:0] _RAND_268;
  reg [4:0] _EVAL_638;
  reg [31:0] _RAND_269;
  reg  _EVAL_640;
  reg [31:0] _RAND_270;
  reg  _EVAL_644;
  reg [31:0] _RAND_271;
  reg  _EVAL_646;
  reg [31:0] _RAND_272;
  reg  _EVAL_648;
  reg [31:0] _RAND_273;
  reg  _EVAL_651;
  reg [31:0] _RAND_274;
  reg [8:0] _EVAL_653;
  reg [31:0] _RAND_275;
  reg  _EVAL_655;
  reg [31:0] _RAND_276;
  reg  _EVAL_657;
  reg [31:0] _RAND_277;
  reg  _EVAL_658;
  reg [31:0] _RAND_278;
  reg [4:0] _EVAL_661;
  reg [31:0] _RAND_279;
  reg [1:0] _EVAL_663;
  reg [31:0] _RAND_280;
  reg  _EVAL_665;
  reg [31:0] _RAND_281;
  reg [1:0] _EVAL_667;
  reg [31:0] _RAND_282;
  reg [8:0] _EVAL_668;
  reg [31:0] _RAND_283;
  reg  _EVAL_672;
  reg [31:0] _RAND_284;
  reg [3:0] _EVAL_673;
  reg [31:0] _RAND_285;
  reg [14:0] _EVAL_675;
  reg [31:0] _RAND_286;
  reg  _EVAL_681;
  reg [31:0] _RAND_287;
  reg  _EVAL_682;
  reg [31:0] _RAND_288;
  reg  _EVAL_683;
  reg [31:0] _RAND_289;
  reg  _EVAL_684;
  reg [31:0] _RAND_290;
  reg [8:0] _EVAL_685;
  reg [31:0] _RAND_291;
  reg  _EVAL_687;
  reg [31:0] _RAND_292;
  reg  _EVAL_688;
  reg [31:0] _RAND_293;
  reg  _EVAL_689;
  reg [31:0] _RAND_294;
  reg  _EVAL_692;
  reg [31:0] _RAND_295;
  reg [14:0] _EVAL_693;
  reg [31:0] _RAND_296;
  reg  _EVAL_695;
  reg [31:0] _RAND_297;
  reg  _EVAL_696;
  reg [31:0] _RAND_298;
  reg  _EVAL_697;
  reg [31:0] _RAND_299;
  reg  _EVAL_698;
  reg [31:0] _RAND_300;
  reg  _EVAL_699;
  reg [31:0] _RAND_301;
  reg  _EVAL_701;
  reg [31:0] _RAND_302;
  reg  _EVAL_702;
  reg [31:0] _RAND_303;
  reg [1:0] _EVAL_703;
  reg [31:0] _RAND_304;
  reg  _EVAL_708;
  reg [31:0] _RAND_305;
  reg  _EVAL_711;
  reg [31:0] _RAND_306;
  reg  _EVAL_714;
  reg [31:0] _RAND_307;
  reg  _EVAL_716;
  reg [31:0] _RAND_308;
  reg  _EVAL_717;
  reg [31:0] _RAND_309;
  reg  _EVAL_718;
  reg [31:0] _RAND_310;
  reg  _EVAL_719;
  reg [31:0] _RAND_311;
  reg  _EVAL_720;
  reg [31:0] _RAND_312;
  reg [2:0] _EVAL_721;
  reg [31:0] _RAND_313;
  reg  _EVAL_722;
  reg [31:0] _RAND_314;
  reg  _EVAL_723;
  reg [31:0] _RAND_315;
  reg  _EVAL_725;
  reg [31:0] _RAND_316;
  reg  _EVAL_726;
  reg [31:0] _RAND_317;
  reg  _EVAL_727;
  reg [31:0] _RAND_318;
  reg [4:0] _EVAL_728;
  reg [31:0] _RAND_319;
  reg  _EVAL_729;
  reg [31:0] _RAND_320;
  reg  _EVAL_731;
  reg [31:0] _RAND_321;
  reg  _EVAL_732;
  reg [31:0] _RAND_322;
  reg  _EVAL_734;
  reg [31:0] _RAND_323;
  reg  _EVAL_735;
  reg [31:0] _RAND_324;
  reg  _EVAL_736;
  reg [31:0] _RAND_325;
  reg  _EVAL_737;
  reg [31:0] _RAND_326;
  reg  _EVAL_738;
  reg [31:0] _RAND_327;
  reg  _EVAL_739;
  reg [31:0] _RAND_328;
  reg  _EVAL_740;
  reg [31:0] _RAND_329;
  reg  _EVAL_742;
  reg [31:0] _RAND_330;
  reg  _EVAL_743;
  reg [31:0] _RAND_331;
  reg  _EVAL_744;
  reg [31:0] _RAND_332;
  reg [4:0] _EVAL_747;
  reg [31:0] _RAND_333;
  reg [2:0] _EVAL_748;
  reg [31:0] _RAND_334;
  reg  _EVAL_750;
  reg [31:0] _RAND_335;
  reg [4:0] _EVAL_751;
  reg [31:0] _RAND_336;
  reg  _EVAL_753;
  reg [31:0] _RAND_337;
  reg [4:0] _EVAL_754;
  reg [31:0] _RAND_338;
  reg  _EVAL_756;
  reg [31:0] _RAND_339;
  reg  _EVAL_758;
  reg [31:0] _RAND_340;
  reg  _EVAL_760;
  reg [31:0] _RAND_341;
  reg  _EVAL_761;
  reg [31:0] _RAND_342;
  reg  _EVAL_762;
  reg [31:0] _RAND_343;
  reg  _EVAL_763;
  reg [31:0] _RAND_344;
  reg  _EVAL_764;
  reg [31:0] _RAND_345;
  reg  _EVAL_765;
  reg [31:0] _RAND_346;
  reg [1:0] _EVAL_768;
  reg [31:0] _RAND_347;
  reg [2:0] _EVAL_770;
  reg [31:0] _RAND_348;
  reg  _EVAL_772;
  reg [31:0] _RAND_349;
  reg  _EVAL_773;
  reg [31:0] _RAND_350;
  reg [14:0] _EVAL_774;
  reg [31:0] _RAND_351;
  reg [4:0] _EVAL_776;
  reg [31:0] _RAND_352;
  reg  _EVAL_777;
  reg [31:0] _RAND_353;
  reg  _EVAL_778;
  reg [31:0] _RAND_354;
  reg  _EVAL_780;
  reg [31:0] _RAND_355;
  reg [2:0] _EVAL_781;
  reg [31:0] _RAND_356;
  reg  _EVAL_782;
  reg [31:0] _RAND_357;
  reg  _EVAL_786;
  reg [31:0] _RAND_358;
  reg [2:0] _EVAL_787;
  reg [31:0] _RAND_359;
  reg [3:0] _EVAL_788;
  reg [31:0] _RAND_360;
  reg [6:0] _EVAL_789;
  reg [31:0] _RAND_361;
  reg  _EVAL_792;
  reg [31:0] _RAND_362;
  reg  _EVAL_793;
  reg [31:0] _RAND_363;
  reg [31:0] _EVAL_796;
  reg [31:0] _RAND_364;
  reg [2:0] _EVAL_797;
  reg [31:0] _RAND_365;
  reg  _EVAL_798;
  reg [31:0] _RAND_366;
  reg [2:0] _EVAL_799;
  reg [31:0] _RAND_367;
  reg [4:0] _EVAL_800;
  reg [31:0] _RAND_368;
  reg  _EVAL_801;
  reg [31:0] _RAND_369;
  reg  _EVAL_804;
  reg [31:0] _RAND_370;
  reg [8:0] _EVAL_805;
  reg [31:0] _RAND_371;
  reg  _EVAL_806;
  reg [31:0] _RAND_372;
  reg  _EVAL_807;
  reg [31:0] _RAND_373;
  reg  _EVAL_808;
  reg [31:0] _RAND_374;
  reg  _EVAL_809;
  reg [31:0] _RAND_375;
  reg [14:0] _EVAL_810;
  reg [31:0] _RAND_376;
  reg [8:0] _EVAL_811;
  reg [31:0] _RAND_377;
  reg [4:0] _EVAL_812;
  reg [31:0] _RAND_378;
  reg  _EVAL_815;
  reg [31:0] _RAND_379;
  reg  _EVAL_817;
  reg [31:0] _RAND_380;
  reg  _EVAL_818;
  reg [31:0] _RAND_381;
  wire  _EVAL_253;
  wire [134:0] _EVAL_383;
  wire [20:0] _EVAL_347;
  wire [34:0] _EVAL_741;
  wire [177:0] _EVAL_632;
  wire [3:0] _EVAL_298;
  wire [2:0] _EVAL_669;
  wire [3:0] _EVAL_287;
  wire  _EVAL_396;
  wire [3:0] _EVAL_226;
  wire [3:0] _EVAL_755;
  wire [2:0] _EVAL_759;
  wire  _EVAL_532;
  wire [5:0] _EVAL_492;
  wire  _EVAL_791;
  wire  _EVAL_552;
  wire  _EVAL_189;
  wire [1:0] _EVAL_575;
  wire  _EVAL_637;
  wire [134:0] _EVAL_635;
  wire  _EVAL_320;
  wire [7:0] _EVAL_319;
  wire [7:0] _EVAL_458;
  wire [7:0] _EVAL_462;
  wire  _EVAL_516;
  wire  _EVAL_629;
  wire [7:0] _EVAL_212;
  wire [6:0] _EVAL_544;
  wire  _EVAL_677;
  wire [7:0] _EVAL_469;
  wire [7:0] _EVAL_232;
  wire [7:0] _EVAL_448;
  wire  _EVAL_592;
  wire [3:0] _EVAL_220;
  wire [2:0] _EVAL_224;
  wire  _EVAL_367;
  wire  _EVAL_790;
  wire [1:0] _EVAL_803;
  wire [1:0] _EVAL_487;
  wire  _EVAL_214;
  wire [134:0] _EVAL_327;
  wire [20:0] _EVAL_293;
  wire [34:0] _EVAL_412;
  wire [177:0] _EVAL_417;
  wire  _EVAL_666;
  wire [9:0] _EVAL_570;
  wire [5:0] _EVAL_213;
  wire [11:0] _EVAL_588;
  wire [134:0] _EVAL_654;
  wire [20:0] _EVAL_769;
  wire [34:0] _EVAL_258;
  wire [177:0] _EVAL_329;
  wire [256:0] _EVAL_595;
  wire [256:0] _EVAL_671;
  wire [20:0] _EVAL_816;
  wire [20:0] _EVAL_539;
  wire [34:0] _EVAL_386;
  wire  _EVAL_674;
  wire [5:0] _EVAL_190;
  wire [5:0] _EVAL_446;
  wire [11:0] _EVAL_354;
  wire [5:0] _EVAL_680;
  wire  _EVAL_397;
  wire [9:0] _EVAL_351;
  wire [5:0] _EVAL_466;
  wire [11:0] _EVAL_266;
  wire [134:0] _EVAL_227;
  wire [177:0] _EVAL_486;
  wire [256:0] _EVAL_273;
  wire [256:0] _EVAL_265;
  wire [256:0] _EVAL_207;
  wire  _EVAL_553;
  wire  _EVAL_373;
  wire  _EVAL_705;
  wire [2:0] _EVAL_407;
  wire  _EVAL_205;
  wire [2:0] _EVAL_610;
  wire  _EVAL_463;
  wire [3:0] _EVAL_438;
  wire [9:0] _EVAL_325;
  wire [11:0] _EVAL_617;
  wire [256:0] _EVAL_283;
  wire  _EVAL_501;
  wire [9:0] _EVAL_631;
  wire  _EVAL_405;
  wire [9:0] _EVAL_642;
  wire [11:0] _EVAL_676;
  wire [134:0] _EVAL_452;
  wire [20:0] _EVAL_418;
  wire [34:0] _EVAL_493;
  wire [177:0] _EVAL_369;
  wire [256:0] _EVAL_586;
  wire [256:0] _EVAL_450;
  wire  _EVAL_549;
  wire [9:0] _EVAL_523;
  wire [11:0] _EVAL_204;
  wire [134:0] _EVAL_616;
  wire [20:0] _EVAL_730;
  wire [34:0] _EVAL_542;
  wire [177:0] _EVAL_410;
  wire [256:0] _EVAL_408;
  wire [256:0] _EVAL_529;
  wire [256:0] _EVAL_664;
  wire [34:0] _EVAL_295;
  wire [177:0] _EVAL_557;
  wire [256:0] _EVAL_590;
  wire [256:0] _EVAL_292;
  wire [256:0] _EVAL_709;
  wire  _EVAL_495;
  wire [256:0] _EVAL_659;
  wire [256:0] _EVAL_526;
  wire [9:0] _EVAL_231;
  wire [5:0] _EVAL_771;
  wire [11:0] _EVAL_656;
  wire [134:0] _EVAL_506;
  wire [20:0] _EVAL_321;
  wire [34:0] _EVAL_650;
  wire [177:0] _EVAL_464;
  wire [256:0] _EVAL_362;
  wire [256:0] _EVAL_543;
  wire [256:0] _EVAL_443;
  wire [2:0] _EVAL_641;
  wire  _EVAL_454;
  wire [3:0] _EVAL_700;
  wire [2:0] _EVAL_691;
  wire [3:0] _EVAL_357;
  wire [2:0] _EVAL_540;
  wire [3:0] _EVAL_690;
  wire [2:0] _EVAL_627;
  wire  _EVAL_710;
  wire  _EVAL_567;
  wire  _EVAL_478;
  wire [5:0] _EVAL_249;
  wire  _EVAL_193;
  wire  _EVAL_707;
  wire [9:0] _EVAL_449;
  wire [11:0] _EVAL_404;
  wire [256:0] _EVAL_314;
  wire  _EVAL_779;
  wire  _EVAL_678;
  wire [256:0] _EVAL_514;
  wire [256:0] _EVAL_712;
  wire  _EVAL_427;
  wire  _EVAL_749;
  wire  _EVAL_441;
  wire  _EVAL_238;
  wire  _EVAL_230;
  wire  _EVAL_250;
  wire  _EVAL_483;
  wire  _EVAL_724;
  wire  _EVAL_485;
  assign _EVAL_253 = _EVAL_431[0];
  assign _EVAL_383 = {_EVAL_731,_EVAL_434,_EVAL_389,_EVAL_608,_EVAL_770,_EVAL_355};
  assign _EVAL_347 = {_EVAL_538,_EVAL_675,_EVAL_309,_EVAL_718,_EVAL_763,_EVAL_200};
  assign _EVAL_741 = {_EVAL_658,_EVAL_685,_EVAL_560,_EVAL_581,_EVAL_530,_EVAL_534,_EVAL_347};
  assign _EVAL_632 = {_EVAL_597,_EVAL_415,_EVAL_727,_EVAL_604,_EVAL_257,_EVAL_353,_EVAL_383,_EVAL_741};
  assign _EVAL_298 = _EVAL_748 + 3'h1;
  assign _EVAL_669 = _EVAL_298[2:0];
  assign _EVAL_287 = _EVAL_669 + 3'h1;
  assign _EVAL_396 = _EVAL_254 == 1'h0;
  assign _EVAL_226 = _EVAL_431 - _EVAL_748;
  assign _EVAL_755 = $unsigned(_EVAL_226);
  assign _EVAL_759 = _EVAL_755[2:0];
  assign _EVAL_532 = _EVAL_759 > 3'h1;
  assign _EVAL_492 = {_EVAL_311,_EVAL_537,_EVAL_762,_EVAL_218,_EVAL_564,_EVAL_346};
  assign _EVAL_791 = _EVAL_182 & _EVAL_19;
  assign _EVAL_552 = _EVAL_56 & _EVAL_60;
  assign _EVAL_189 = _EVAL_791 & _EVAL_552;
  assign _EVAL_575 = {_EVAL_189,_EVAL_552};
  assign _EVAL_637 = _EVAL_575[1];
  assign _EVAL_635 = {_EVAL_711,_EVAL_515,_EVAL_186,_EVAL_573,_EVAL_621,_EVAL_444};
  assign _EVAL_320 = _EVAL_42 & _EVAL_94;
  assign _EVAL_319 = _EVAL_320 ? 8'hff : 8'h0;
  assign _EVAL_458 = 8'h1 << _EVAL_431;
  assign _EVAL_462 = _EVAL_319 & _EVAL_458;
  assign _EVAL_516 = _EVAL_153 & _EVAL_176;
  assign _EVAL_629 = _EVAL_516 & _EVAL_320;
  assign _EVAL_212 = _EVAL_629 ? 8'hff : 8'h0;
  assign _EVAL_544 = _EVAL_458[6:0];
  assign _EVAL_677 = _EVAL_458[7];
  assign _EVAL_469 = {_EVAL_544,_EVAL_677};
  assign _EVAL_232 = _EVAL_212 & _EVAL_469;
  assign _EVAL_448 = _EVAL_462 | _EVAL_232;
  assign _EVAL_592 = _EVAL_448[4];
  assign _EVAL_220 = {{1'd0}, _EVAL_669};
  assign _EVAL_224 = _EVAL_220[2:0];
  assign _EVAL_367 = _EVAL_748[0];
  assign _EVAL_790 = _EVAL_575[0];
  assign _EVAL_803 = {_EVAL_790,_EVAL_637};
  assign _EVAL_487 = _EVAL_367 ? _EVAL_803 : _EVAL_575;
  assign _EVAL_214 = _EVAL_487[0];
  assign _EVAL_327 = {_EVAL_533,_EVAL_348,_EVAL_473,_EVAL_374,_EVAL_260,_EVAL_278};
  assign _EVAL_293 = {_EVAL_451,_EVAL_225,_EVAL_365,_EVAL_322,_EVAL_455,_EVAL_695};
  assign _EVAL_412 = {_EVAL_508,_EVAL_603,_EVAL_818,_EVAL_626,_EVAL_555,_EVAL_612,_EVAL_293};
  assign _EVAL_417 = {_EVAL_786,_EVAL_363,_EVAL_239,_EVAL_243,_EVAL_541,_EVAL_739,_EVAL_327,_EVAL_412};
  assign _EVAL_666 = _EVAL_788[0];
  assign _EVAL_570 = {_EVAL_393,_EVAL_221,_EVAL_332,_EVAL_219,_EVAL_453,_EVAL_489};
  assign _EVAL_213 = {_EVAL_687,_EVAL_798,_EVAL_306,_EVAL_330,_EVAL_470,_EVAL_271};
  assign _EVAL_588 = {_EVAL_500,_EVAL_510,_EVAL_545,_EVAL_692,1'h0,_EVAL_447,_EVAL_213};
  assign _EVAL_654 = {_EVAL_701,_EVAL_340,_EVAL_714,_EVAL_665,_EVAL_337,_EVAL_345};
  assign _EVAL_769 = {_EVAL_490,_EVAL_810,_EVAL_318,_EVAL_246,_EVAL_248,_EVAL_806};
  assign _EVAL_258 = {_EVAL_615,_EVAL_811,_EVAL_270,_EVAL_736,_EVAL_518,_EVAL_625,_EVAL_769};
  assign _EVAL_329 = {_EVAL_202,_EVAL_601,_EVAL_808,_EVAL_554,_EVAL_467,_EVAL_723,_EVAL_654,_EVAL_258};
  assign _EVAL_595 = {_EVAL_377,_EVAL_424,_EVAL_797,_EVAL_468,_EVAL_527,_EVAL_593,_EVAL_570,_EVAL_588,_EVAL_329};
  assign _EVAL_671 = _EVAL_666 ? _EVAL_595 : 257'h0;
  assign _EVAL_816 = {_EVAL_279,_EVAL_428,_EVAL_547,_EVAL_753,_EVAL_729,_EVAL_242};
  assign _EVAL_539 = {_EVAL_663,_EVAL_693,_EVAL_237,_EVAL_491,_EVAL_494,_EVAL_807};
  assign _EVAL_386 = {_EVAL_801,_EVAL_805,_EVAL_313,_EVAL_778,_EVAL_563,_EVAL_782,_EVAL_539};
  assign _EVAL_674 = _EVAL_748 == _EVAL_431;
  assign _EVAL_190 = {_EVAL_215,_EVAL_681,_EVAL_566,_EVAL_702,_EVAL_422,_EVAL_740};
  assign _EVAL_446 = {_EVAL_594,_EVAL_619,_EVAL_484,_EVAL_398,_EVAL_505,_EVAL_528};
  assign _EVAL_354 = {_EVAL_620,_EVAL_426,_EVAL_302,_EVAL_255,1'h0,_EVAL_657,_EVAL_446};
  assign _EVAL_680 = {_EVAL_429,_EVAL_640,_EVAL_758,_EVAL_460,_EVAL_606,_EVAL_268};
  assign _EVAL_397 = _EVAL_788[1];
  assign _EVAL_351 = {_EVAL_571,_EVAL_482,_EVAL_732,_EVAL_561,_EVAL_591,_EVAL_430};
  assign _EVAL_466 = {_EVAL_720,_EVAL_648,_EVAL_288,_EVAL_717,_EVAL_488,_EVAL_684};
  assign _EVAL_266 = {_EVAL_596,_EVAL_582,_EVAL_744,_EVAL_750,1'h0,_EVAL_188,_EVAL_466};
  assign _EVAL_227 = {_EVAL_568,_EVAL_524,_EVAL_308,_EVAL_376,_EVAL_192,_EVAL_235};
  assign _EVAL_486 = {_EVAL_696,_EVAL_413,_EVAL_272,_EVAL_742,_EVAL_210,_EVAL_241,_EVAL_227,_EVAL_386};
  assign _EVAL_273 = {_EVAL_796,_EVAL_754,_EVAL_316,_EVAL_297,_EVAL_661,_EVAL_574,_EVAL_351,_EVAL_266,_EVAL_486};
  assign _EVAL_265 = _EVAL_397 ? _EVAL_273 : 257'h0;
  assign _EVAL_207 = _EVAL_671 | _EVAL_265;
  assign _EVAL_553 = _EVAL_791 == 1'h0;
  assign _EVAL_373 = _EVAL_516 == 1'h0;
  assign _EVAL_705 = _EVAL_373 ? 1'h0 : 1'h1;
  assign _EVAL_407 = {{2'd0}, _EVAL_705};
  assign _EVAL_205 = _EVAL_673[2];
  assign _EVAL_610 = _EVAL_788[2:0];
  assign _EVAL_463 = _EVAL_788[3];
  assign _EVAL_438 = {_EVAL_610,_EVAL_463};
  assign _EVAL_325 = {_EVAL_812,_EVAL_203,_EVAL_247,_EVAL_756,_EVAL_256,_EVAL_264};
  assign _EVAL_617 = {_EVAL_282,_EVAL_743,_EVAL_734,_EVAL_683,1'h0,_EVAL_358,_EVAL_190};
  assign _EVAL_283 = {_EVAL_328,_EVAL_638,_EVAL_799,_EVAL_634,_EVAL_425,_EVAL_602,_EVAL_325,_EVAL_617,_EVAL_417};
  assign _EVAL_501 = _EVAL_448[5];
  assign _EVAL_631 = {_EVAL_252,_EVAL_598,_EVAL_584,_EVAL_339,_EVAL_223,_EVAL_630};
  assign _EVAL_405 = _EVAL_673[0];
  assign _EVAL_642 = {_EVAL_747,_EVAL_618,_EVAL_315,_EVAL_525,_EVAL_817,_EVAL_229};
  assign _EVAL_676 = {_EVAL_289,_EVAL_507,_EVAL_392,_EVAL_556,1'h0,_EVAL_651,_EVAL_680};
  assign _EVAL_452 = {_EVAL_335,_EVAL_548,_EVAL_780,_EVAL_244,_EVAL_721,_EVAL_761};
  assign _EVAL_418 = {_EVAL_703,_EVAL_774,_EVAL_716,_EVAL_371,_EVAL_286,_EVAL_433};
  assign _EVAL_493 = {_EVAL_263,_EVAL_317,_EVAL_285,_EVAL_722,_EVAL_546,_EVAL_416,_EVAL_418};
  assign _EVAL_369 = {_EVAL_655,_EVAL_201,_EVAL_699,_EVAL_646,_EVAL_513,_EVAL_331,_EVAL_452,_EVAL_493};
  assign _EVAL_586 = {_EVAL_536,_EVAL_776,_EVAL_420,_EVAL_789,_EVAL_187,_EVAL_338,_EVAL_642,_EVAL_676,_EVAL_369};
  assign _EVAL_450 = _EVAL_405 ? _EVAL_586 : 257'h0;
  assign _EVAL_549 = _EVAL_673[1];
  assign _EVAL_523 = {_EVAL_751,_EVAL_442,_EVAL_558,_EVAL_436,_EVAL_352,_EVAL_356};
  assign _EVAL_204 = {_EVAL_497,_EVAL_499,_EVAL_682,_EVAL_725,1'h0,_EVAL_387,_EVAL_492};
  assign _EVAL_616 = {_EVAL_301,_EVAL_472,_EVAL_194,_EVAL_388,_EVAL_456,_EVAL_609};
  assign _EVAL_730 = {_EVAL_667,_EVAL_576,_EVAL_502,_EVAL_361,_EVAL_461,_EVAL_457};
  assign _EVAL_542 = {_EVAL_304,_EVAL_668,_EVAL_777,_EVAL_445,_EVAL_521,_EVAL_804,_EVAL_730};
  assign _EVAL_410 = {_EVAL_697,_EVAL_504,_EVAL_294,_EVAL_614,_EVAL_781,_EVAL_672,_EVAL_616,_EVAL_542};
  assign _EVAL_408 = {_EVAL_274,_EVAL_623,_EVAL_342,_EVAL_402,_EVAL_233,_EVAL_569,_EVAL_523,_EVAL_204,_EVAL_410};
  assign _EVAL_529 = _EVAL_549 ? _EVAL_408 : 257'h0;
  assign _EVAL_664 = _EVAL_450 | _EVAL_529;
  assign _EVAL_295 = {_EVAL_312,_EVAL_372,_EVAL_291,_EVAL_476,_EVAL_277,_EVAL_222,_EVAL_816};
  assign _EVAL_557 = {_EVAL_760,_EVAL_280,_EVAL_209,_EVAL_333,_EVAL_360,_EVAL_349,_EVAL_635,_EVAL_295};
  assign _EVAL_590 = {_EVAL_240,_EVAL_259,_EVAL_559,_EVAL_439,_EVAL_390,_EVAL_368,_EVAL_631,_EVAL_354,_EVAL_557};
  assign _EVAL_292 = _EVAL_205 ? _EVAL_590 : 257'h0;
  assign _EVAL_709 = _EVAL_664 | _EVAL_292;
  assign _EVAL_495 = _EVAL_788[2];
  assign _EVAL_659 = _EVAL_495 ? _EVAL_283 : 257'h0;
  assign _EVAL_526 = _EVAL_207 | _EVAL_659;
  assign _EVAL_231 = {_EVAL_728,_EVAL_519,_EVAL_688,_EVAL_323,_EVAL_793,_EVAL_517};
  assign _EVAL_771 = {_EVAL_475,_EVAL_350,_EVAL_296,_EVAL_366,_EVAL_708,_EVAL_307};
  assign _EVAL_656 = {_EVAL_765,_EVAL_600,_EVAL_809,_EVAL_599,1'h0,_EVAL_644,_EVAL_771};
  assign _EVAL_506 = {_EVAL_738,_EVAL_471,_EVAL_587,_EVAL_735,_EVAL_336,_EVAL_269};
  assign _EVAL_321 = {_EVAL_768,_EVAL_498,_EVAL_633,_EVAL_689,_EVAL_773,_EVAL_611};
  assign _EVAL_650 = {_EVAL_772,_EVAL_653,_EVAL_234,_EVAL_421,_EVAL_511,_EVAL_764,_EVAL_321};
  assign _EVAL_464 = {_EVAL_375,_EVAL_815,_EVAL_726,_EVAL_400,_EVAL_787,_EVAL_792,_EVAL_506,_EVAL_650};
  assign _EVAL_362 = {_EVAL_267,_EVAL_217,_EVAL_284,_EVAL_197,_EVAL_211,_EVAL_474,_EVAL_231,_EVAL_656,_EVAL_464};
  assign _EVAL_543 = _EVAL_463 ? _EVAL_362 : 257'h0;
  assign _EVAL_443 = _EVAL_526 | _EVAL_543;
  assign _EVAL_641 = _EVAL_673[2:0];
  assign _EVAL_454 = _EVAL_673[3];
  assign _EVAL_700 = {_EVAL_641,_EVAL_454};
  assign _EVAL_691 = _EVAL_287[2:0];
  assign _EVAL_357 = _EVAL_431 + 3'h1;
  assign _EVAL_540 = _EVAL_357[2:0];
  assign _EVAL_690 = _EVAL_540 + _EVAL_407;
  assign _EVAL_627 = _EVAL_690[2:0];
  assign _EVAL_710 = _EVAL_487[1];
  assign _EVAL_567 = _EVAL_448[3];
  assign _EVAL_478 = _EVAL_674 & _EVAL_254;
  assign _EVAL_249 = {_EVAL_589,_EVAL_414,_EVAL_622,_EVAL_551,_EVAL_562,_EVAL_199};
  assign _EVAL_193 = _EVAL_448[7];
  assign _EVAL_707 = _EVAL_448[0];
  assign _EVAL_449 = {_EVAL_509,_EVAL_579,_EVAL_698,_EVAL_522,_EVAL_580,_EVAL_737};
  assign _EVAL_404 = {_EVAL_565,_EVAL_480,_EVAL_479,_EVAL_607,1'h0,_EVAL_719,_EVAL_249};
  assign _EVAL_314 = {_EVAL_196,_EVAL_440,_EVAL_343,_EVAL_391,_EVAL_251,_EVAL_800,_EVAL_449,_EVAL_404,_EVAL_632};
  assign _EVAL_779 = _EVAL_674 & _EVAL_396;
  assign _EVAL_678 = _EVAL_779 == 1'h0;
  assign _EVAL_514 = _EVAL_454 ? _EVAL_314 : 257'h0;
  assign _EVAL_712 = _EVAL_709 | _EVAL_514;
  assign _EVAL_427 = _EVAL_553 ? 1'h0 : 1'h1;
  assign _EVAL_749 = _EVAL_705 > _EVAL_427;
  assign _EVAL_441 = _EVAL_759 < 3'h7;
  assign _EVAL_238 = _EVAL_320 & _EVAL_749;
  assign _EVAL_230 = _EVAL_320 | _EVAL_254;
  assign _EVAL_250 = _EVAL_448[6];
  assign _EVAL_483 = _EVAL_448[1];
  assign _EVAL_724 = _EVAL_448[2];
  assign _EVAL_485 = _EVAL_478 == 1'h0;
  assign _EVAL_125 = _EVAL_443[18:4];
  assign _EVAL_57 = _EVAL_712[170];
  assign _EVAL_179 = _EVAL_712[188];
  assign _EVAL_26 = _EVAL_712[189];
  assign _EVAL_52 = _EVAL_712[34];
  assign _EVAL_123 = _EVAL_712[40];
  assign _EVAL_94 = _EVAL_478 == 1'h0;
  assign _EVAL_165 = _EVAL_443[186];
  assign _EVAL_4 = _EVAL_443[170];
  assign _EVAL_176 = _EVAL_485 & _EVAL_441;
  assign _EVAL_146 = _EVAL_443[256:225];
  assign _EVAL_34 = _EVAL_443[187];
  assign _EVAL_162 = _EVAL_443[40];
  assign _EVAL_138 = _EVAL_712[187];
  assign _EVAL_145 = _EVAL_712[20:19];
  assign _EVAL_56 = _EVAL_779 == 1'h0;
  assign _EVAL_183 = _EVAL_712[219:217];
  assign _EVAL_21 = _EVAL_443[34];
  assign _EVAL_141 = _EVAL_712[224:220];
  assign _EVAL_38 = _EVAL_443[176];
  assign _EVAL_43 = _EVAL_712[182];
  assign _EVAL_93 = _EVAL_712[185];
  assign _EVAL_65 = _EVAL_443[185];
  assign _EVAL_132 = _EVAL_443[177];
  assign _EVAL_83 = _EVAL_712[21];
  assign _EVAL_2 = _EVAL_443[181];
  assign _EVAL_85 = _EVAL_712[39];
  assign _EVAL_8 = _EVAL_443[189];
  assign _EVAL_9 = _EVAL_443[224:220];
  assign _EVAL_124 = _EVAL_443[39];
  assign _EVAL_49 = _EVAL_712[186];
  assign _EVAL_69 = _EVAL_443[20:19];
  assign _EVAL_144 = _EVAL_443[183];
  assign _EVAL_96 = _EVAL_443[191];
  assign _EVAL_140 = _EVAL_712[190];
  assign _EVAL_61 = _EVAL_712[180];
  assign _EVAL_74 = _EVAL_443[209:205];
  assign _EVAL_30 = _EVAL_443[173:171];
  assign _EVAL_163 = _EVAL_443[38:36];
  assign _EVAL_20 = _EVAL_443[169];
  assign _EVAL_40 = _EVAL_712[181];
  assign _EVAL_118 = _EVAL_443[22];
  assign _EVAL_13 = _EVAL_443[199:195];
  assign _EVAL_106 = _EVAL_443[179];
  assign _EVAL_84 = _EVAL_712[179];
  assign _EVAL_24 = _EVAL_712[18:4];
  assign _EVAL_129 = _EVAL_712[216:210];
  assign _EVAL_0 = _EVAL_712[178];
  assign _EVAL_109 = _EVAL_712[204:200];
  assign _EVAL_111 = _EVAL_712[22];
  assign _EVAL_66 = _EVAL_303;
  assign _EVAL_79 = _EVAL_443[192];
  assign _EVAL_121 = _EVAL_712[192];
  assign _EVAL_98 = _EVAL_712[168:41];
  assign _EVAL_152 = _EVAL_443[168:41];
  assign _EVAL_160 = _EVAL_712[193];
  assign _EVAL_133 = _EVAL_712[199:195];
  assign _EVAL_159 = _EVAL_443[23];
  assign _EVAL_53 = _EVAL_443[178];
  assign _EVAL_45 = _EVAL_443[174];
  assign _EVAL_81 = _EVAL_712[169];
  assign _EVAL_185 = _EVAL_712[184];
  assign _EVAL_182 = _EVAL_532 | _EVAL_478;
  assign _EVAL_77 = _EVAL_712[256:225];
  assign _EVAL_17 = _EVAL_443[184];
  assign _EVAL_91 = _EVAL_712[209:205];
  assign _EVAL_70 = _EVAL_712[183];
  assign _EVAL_128 = _EVAL_712[38:36];
  assign _EVAL_59 = _EVAL_712[175];
  assign _EVAL_166 = _EVAL_443[182];
  assign _EVAL_171 = _EVAL_443[216:210];
  assign _EVAL_73 = _EVAL_443[193];
  assign _EVAL_18 = _EVAL_443[219:217];
  assign _EVAL_90 = _EVAL_712[194];
  assign _EVAL_170 = _EVAL_443[188];
  assign _EVAL_22 = _EVAL_443[175];
  assign _EVAL_67 = _EVAL_712[23];
  assign _EVAL_6 = _EVAL_712[174];
  assign _EVAL_155 = _EVAL_443[180];
  assign _EVAL_136 = _EVAL_712[191];
  assign _EVAL_134 = _EVAL_712[176];
  assign _EVAL_112 = _EVAL_443[190];
  assign _EVAL_3 = _EVAL_712[173:171];
  assign _EVAL_78 = _EVAL_748[0];
  assign _EVAL_113 = _EVAL_712[177];
  assign _EVAL_180 = _EVAL_443[21];
  assign _EVAL_27 = _EVAL_443[204:200];
  assign _EVAL_173 = _EVAL_443[194];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_187 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_188 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_192 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_194 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_196 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_197 = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_199 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_200 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_201 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_202 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_203 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_209 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_210 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_211 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_215 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_217 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_218 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_219 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_221 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_222 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_223 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_225 = _RAND_22[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_229 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_233 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_234 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_235 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_237 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_239 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_240 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_241 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_242 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_243 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_244 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_246 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_247 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_248 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_251 = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_252 = _RAND_38[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_254 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_255 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_256 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_257 = _RAND_42[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_259 = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_260 = _RAND_44[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_263 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_264 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_267 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_268 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_269 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_270 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_271 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_272 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_274 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_277 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_278 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_279 = _RAND_56[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_280 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_282 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_284 = _RAND_59[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_285 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_286 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_288 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_289 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_291 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_294 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_296 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_297 = _RAND_67[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_301 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_302 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_303 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_304 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_306 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_307 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_308 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_309 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_311 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_312 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_313 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_315 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_316 = _RAND_80[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_317 = _RAND_81[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_318 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_322 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_323 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_328 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_330 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_331 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_332 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_333 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_335 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_336 = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_337 = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_338 = _RAND_93[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_339 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {4{`RANDOM}};
  _EVAL_340 = _RAND_95[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_342 = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_343 = _RAND_97[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_345 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_346 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {4{`RANDOM}};
  _EVAL_348 = _RAND_100[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_349 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_350 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_352 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_353 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_355 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_356 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_358 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_360 = _RAND_108[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_361 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_363 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_365 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_366 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_368 = _RAND_113[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _EVAL_371 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_372 = _RAND_115[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_374 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_375 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_376 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_377 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_387 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_388 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_389 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_390 = _RAND_123[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_391 = _RAND_124[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_392 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_393 = _RAND_126[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_398 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_400 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_402 = _RAND_129[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_413 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_414 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_415 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_416 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_420 = _RAND_134[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_421 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_422 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_424 = _RAND_137[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_425 = _RAND_138[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_426 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_428 = _RAND_140[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_429 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _EVAL_430 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_431 = _RAND_143[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _EVAL_433 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {4{`RANDOM}};
  _EVAL_434 = _RAND_145[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_436 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _EVAL_439 = _RAND_147[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _EVAL_440 = _RAND_148[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _EVAL_442 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _EVAL_444 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _EVAL_445 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _EVAL_447 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _EVAL_451 = _RAND_153[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _EVAL_453 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _EVAL_455 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _EVAL_456 = _RAND_156[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _EVAL_457 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _EVAL_460 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _EVAL_461 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _EVAL_467 = _RAND_160[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _EVAL_468 = _RAND_161[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _EVAL_470 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {4{`RANDOM}};
  _EVAL_471 = _RAND_163[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {4{`RANDOM}};
  _EVAL_472 = _RAND_164[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _EVAL_473 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _EVAL_474 = _RAND_166[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _EVAL_475 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _EVAL_476 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _EVAL_479 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _EVAL_480 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _EVAL_482 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _EVAL_484 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _EVAL_488 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _EVAL_489 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _EVAL_490 = _RAND_175[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _EVAL_491 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _EVAL_494 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _EVAL_497 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _EVAL_498 = _RAND_179[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _EVAL_499 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _EVAL_500 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _EVAL_502 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _EVAL_504 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _EVAL_505 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _EVAL_507 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _EVAL_508 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _EVAL_509 = _RAND_187[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _EVAL_510 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _EVAL_511 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _EVAL_513 = _RAND_190[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {4{`RANDOM}};
  _EVAL_515 = _RAND_191[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _EVAL_517 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _EVAL_518 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _EVAL_519 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _EVAL_521 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _EVAL_522 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {4{`RANDOM}};
  _EVAL_524 = _RAND_197[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _EVAL_525 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _EVAL_527 = _RAND_199[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _EVAL_528 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _EVAL_530 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _EVAL_533 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _EVAL_534 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _EVAL_536 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _EVAL_537 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _EVAL_538 = _RAND_206[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _EVAL_541 = _RAND_207[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _EVAL_545 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _EVAL_546 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _EVAL_547 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {4{`RANDOM}};
  _EVAL_548 = _RAND_211[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _EVAL_551 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _EVAL_554 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _EVAL_555 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _EVAL_556 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _EVAL_558 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _EVAL_559 = _RAND_217[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _EVAL_560 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _EVAL_561 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _EVAL_562 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _EVAL_563 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _EVAL_564 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _EVAL_565 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _EVAL_566 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _EVAL_568 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _EVAL_569 = _RAND_226[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _EVAL_571 = _RAND_227[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _EVAL_573 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _EVAL_574 = _RAND_229[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _EVAL_576 = _RAND_230[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _EVAL_579 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _EVAL_580 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _EVAL_581 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _EVAL_582 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _EVAL_584 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _EVAL_587 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _EVAL_589 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _EVAL_591 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _EVAL_593 = _RAND_239[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _EVAL_594 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _EVAL_596 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _EVAL_597 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _EVAL_598 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _EVAL_599 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _EVAL_600 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _EVAL_601 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _EVAL_602 = _RAND_247[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _EVAL_603 = _RAND_248[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _EVAL_604 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _EVAL_606 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _EVAL_607 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _EVAL_608 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _EVAL_609 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _EVAL_611 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _EVAL_612 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _EVAL_614 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _EVAL_615 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _EVAL_618 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _EVAL_619 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _EVAL_620 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _EVAL_621 = _RAND_261[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _EVAL_622 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _EVAL_623 = _RAND_263[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _EVAL_625 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _EVAL_626 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _EVAL_630 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _EVAL_633 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _EVAL_634 = _RAND_268[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _EVAL_638 = _RAND_269[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _EVAL_640 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _EVAL_644 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _EVAL_646 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _EVAL_648 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _EVAL_651 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _EVAL_653 = _RAND_275[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _EVAL_655 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _EVAL_657 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _EVAL_658 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _EVAL_661 = _RAND_279[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _EVAL_663 = _RAND_280[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _EVAL_665 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _EVAL_667 = _RAND_282[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _EVAL_668 = _RAND_283[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _EVAL_672 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _EVAL_673 = _RAND_285[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _EVAL_675 = _RAND_286[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _EVAL_681 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _EVAL_682 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _EVAL_683 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _EVAL_684 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _EVAL_685 = _RAND_291[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _EVAL_687 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _EVAL_688 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _EVAL_689 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _EVAL_692 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _EVAL_693 = _RAND_296[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _EVAL_695 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _EVAL_696 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _EVAL_697 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _EVAL_698 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _EVAL_699 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _EVAL_701 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _EVAL_702 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _EVAL_703 = _RAND_304[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _EVAL_708 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _EVAL_711 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _EVAL_714 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _EVAL_716 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _EVAL_717 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _EVAL_718 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _EVAL_719 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _EVAL_720 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _EVAL_721 = _RAND_313[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _EVAL_722 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _EVAL_723 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _EVAL_725 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _EVAL_726 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _EVAL_727 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _EVAL_728 = _RAND_319[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _EVAL_729 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _EVAL_731 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _EVAL_732 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _EVAL_734 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _EVAL_735 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _EVAL_736 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _EVAL_737 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _EVAL_738 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _EVAL_739 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _EVAL_740 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _EVAL_742 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _EVAL_743 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _EVAL_744 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _EVAL_747 = _RAND_333[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _EVAL_748 = _RAND_334[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _EVAL_750 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _EVAL_751 = _RAND_336[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _EVAL_753 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _EVAL_754 = _RAND_338[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _EVAL_756 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _EVAL_758 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _EVAL_760 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _EVAL_761 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _EVAL_762 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _EVAL_763 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _EVAL_764 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _EVAL_765 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _EVAL_768 = _RAND_347[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _EVAL_770 = _RAND_348[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _EVAL_772 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _EVAL_773 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _EVAL_774 = _RAND_351[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _EVAL_776 = _RAND_352[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _EVAL_777 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _EVAL_778 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _EVAL_780 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _EVAL_781 = _RAND_356[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _EVAL_782 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _EVAL_786 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _EVAL_787 = _RAND_359[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _EVAL_788 = _RAND_360[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _EVAL_789 = _RAND_361[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _EVAL_792 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _EVAL_793 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _EVAL_796 = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _EVAL_797 = _RAND_365[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _EVAL_798 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _EVAL_799 = _RAND_367[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _EVAL_800 = _RAND_368[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _EVAL_801 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _EVAL_804 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _EVAL_805 = _RAND_371[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _EVAL_806 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _EVAL_807 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _EVAL_808 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _EVAL_809 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _EVAL_810 = _RAND_376[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _EVAL_811 = _RAND_377[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _EVAL_812 = _RAND_378[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _EVAL_815 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _EVAL_817 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _EVAL_818 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_32) begin
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_186 <= _EVAL_122;
      end else begin
        _EVAL_186 <= _EVAL_114;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_187 <= _EVAL_169;
      end else begin
        _EVAL_187 <= _EVAL_88;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_188 <= _EVAL_175;
      end else begin
        _EVAL_188 <= _EVAL_64;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_192 <= _EVAL_82;
      end else begin
        _EVAL_192 <= _EVAL_92;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_194 <= _EVAL_122;
      end else begin
        _EVAL_194 <= _EVAL_114;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_196 <= _EVAL_102;
      end else begin
        _EVAL_196 <= _EVAL_127;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_197 <= _EVAL_63;
      end else begin
        _EVAL_197 <= _EVAL_148;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_199 <= _EVAL_68;
      end else begin
        _EVAL_199 <= _EVAL_158;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_200 <= _EVAL_28;
      end else begin
        _EVAL_200 <= _EVAL_177;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_201 <= 1'h0;
      end else begin
        _EVAL_201 <= _EVAL_167;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_202 <= _EVAL_139;
      end else begin
        _EVAL_202 <= _EVAL_164;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_203 <= _EVAL_55;
      end else begin
        _EVAL_203 <= _EVAL_104;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_209 <= _EVAL_51;
      end else begin
        _EVAL_209 <= _EVAL_181;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_210 <= _EVAL_101;
      end else begin
        _EVAL_210 <= _EVAL_126;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_211 <= _EVAL_88;
      end else begin
        _EVAL_211 <= _EVAL_169;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_215 <= _EVAL_80;
      end else begin
        _EVAL_215 <= _EVAL_156;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_217 <= _EVAL_62;
      end else begin
        _EVAL_217 <= _EVAL_58;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_218 <= _EVAL_11;
      end else begin
        _EVAL_218 <= _EVAL_54;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_219 <= _EVAL_14;
      end else begin
        _EVAL_219 <= _EVAL_151;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_221 <= _EVAL_55;
      end else begin
        _EVAL_221 <= _EVAL_104;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_222 <= _EVAL_87;
      end else begin
        _EVAL_222 <= _EVAL_116;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_223 <= _EVAL_174;
      end else begin
        _EVAL_223 <= _EVAL_110;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_225 <= _EVAL_41;
      end else begin
        _EVAL_225 <= _EVAL_39;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_229 <= _EVAL_105;
      end else begin
        _EVAL_229 <= _EVAL_161;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_233 <= _EVAL_169;
      end else begin
        _EVAL_233 <= _EVAL_88;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_234 <= _EVAL_147;
      end else begin
        _EVAL_234 <= _EVAL_131;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_235 <= _EVAL_168;
      end else begin
        _EVAL_235 <= _EVAL_184;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_237 <= _EVAL_33;
      end else begin
        _EVAL_237 <= _EVAL_115;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_239 <= _EVAL_181;
      end else begin
        _EVAL_239 <= _EVAL_51;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_240 <= _EVAL_102;
      end else begin
        _EVAL_240 <= _EVAL_127;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_241 <= _EVAL_130;
      end else begin
        _EVAL_241 <= _EVAL_142;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_242 <= _EVAL_28;
      end else begin
        _EVAL_242 <= _EVAL_177;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_243 <= _EVAL_5;
      end else begin
        _EVAL_243 <= _EVAL_143;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_244 <= _EVAL_7;
      end else begin
        _EVAL_244 <= _EVAL_95;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_246 <= _EVAL_108;
      end else begin
        _EVAL_246 <= _EVAL_89;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_247 <= _EVAL_120;
      end else begin
        _EVAL_247 <= _EVAL_99;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_248 <= _EVAL_100;
      end else begin
        _EVAL_248 <= _EVAL_86;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_251 <= _EVAL_169;
      end else begin
        _EVAL_251 <= _EVAL_88;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_252 <= _EVAL_48;
      end else begin
        _EVAL_252 <= _EVAL_154;
      end
    end
    if (_EVAL_50) begin
      _EVAL_254 <= 1'h0;
    end else begin
      if (_EVAL_552) begin
        _EVAL_254 <= _EVAL_238;
      end else begin
        _EVAL_254 <= _EVAL_230;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_255 <= _EVAL_36;
      end else begin
        _EVAL_255 <= _EVAL;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_256 <= _EVAL_110;
      end else begin
        _EVAL_256 <= _EVAL_174;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_257 <= _EVAL_126;
      end else begin
        _EVAL_257 <= _EVAL_101;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_259 <= _EVAL_58;
      end else begin
        _EVAL_259 <= _EVAL_62;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_260 <= _EVAL_82;
      end else begin
        _EVAL_260 <= _EVAL_92;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_263 <= _EVAL_44;
      end else begin
        _EVAL_263 <= _EVAL_12;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_264 <= _EVAL_161;
      end else begin
        _EVAL_264 <= _EVAL_105;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_267 <= _EVAL_127;
      end else begin
        _EVAL_267 <= _EVAL_102;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_268 <= _EVAL_68;
      end else begin
        _EVAL_268 <= _EVAL_158;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_269 <= _EVAL_168;
      end else begin
        _EVAL_269 <= _EVAL_184;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_270 <= _EVAL_147;
      end else begin
        _EVAL_270 <= _EVAL_131;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_271 <= _EVAL_158;
      end else begin
        _EVAL_271 <= _EVAL_68;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_272 <= _EVAL_181;
      end else begin
        _EVAL_272 <= _EVAL_51;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_274 <= _EVAL_102;
      end else begin
        _EVAL_274 <= _EVAL_127;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_277 <= _EVAL_76;
      end else begin
        _EVAL_277 <= _EVAL_75;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_278 <= _EVAL_168;
      end else begin
        _EVAL_278 <= _EVAL_184;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_279 <= _EVAL_1;
      end else begin
        _EVAL_279 <= _EVAL_103;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_280 <= 1'h0;
      end else begin
        _EVAL_280 <= _EVAL_167;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_282 <= _EVAL_135;
      end else begin
        _EVAL_282 <= _EVAL_25;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_284 <= _EVAL_149;
      end else begin
        _EVAL_284 <= _EVAL_47;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_285 <= _EVAL_131;
      end else begin
        _EVAL_285 <= _EVAL_147;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_286 <= _EVAL_86;
      end else begin
        _EVAL_286 <= _EVAL_100;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_288 <= _EVAL_71;
      end else begin
        _EVAL_288 <= _EVAL_119;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_289 <= _EVAL_25;
      end else begin
        _EVAL_289 <= _EVAL_135;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_291 <= _EVAL_131;
      end else begin
        _EVAL_291 <= _EVAL_147;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_294 <= _EVAL_51;
      end else begin
        _EVAL_294 <= _EVAL_181;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_296 <= _EVAL_71;
      end else begin
        _EVAL_296 <= _EVAL_119;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_297 <= _EVAL_63;
      end else begin
        _EVAL_297 <= _EVAL_148;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_301 <= _EVAL_37;
      end else begin
        _EVAL_301 <= _EVAL_137;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_302 <= _EVAL_16;
      end else begin
        _EVAL_302 <= _EVAL_35;
      end
    end
    _EVAL_303 <= _EVAL_678 | _EVAL_42;
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_304 <= _EVAL_44;
      end else begin
        _EVAL_304 <= _EVAL_12;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_306 <= _EVAL_71;
      end else begin
        _EVAL_306 <= _EVAL_119;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_307 <= _EVAL_158;
      end else begin
        _EVAL_307 <= _EVAL_68;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_308 <= _EVAL_114;
      end else begin
        _EVAL_308 <= _EVAL_122;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_309 <= _EVAL_115;
      end else begin
        _EVAL_309 <= _EVAL_33;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_311 <= _EVAL_156;
      end else begin
        _EVAL_311 <= _EVAL_80;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_312 <= _EVAL_44;
      end else begin
        _EVAL_312 <= _EVAL_12;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_313 <= _EVAL_147;
      end else begin
        _EVAL_313 <= _EVAL_131;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_315 <= _EVAL_99;
      end else begin
        _EVAL_315 <= _EVAL_120;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_316 <= _EVAL_149;
      end else begin
        _EVAL_316 <= _EVAL_47;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_317 <= _EVAL_107;
      end else begin
        _EVAL_317 <= _EVAL_72;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_318 <= _EVAL_33;
      end else begin
        _EVAL_318 <= _EVAL_115;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_322 <= _EVAL_108;
      end else begin
        _EVAL_322 <= _EVAL_89;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_323 <= _EVAL_14;
      end else begin
        _EVAL_323 <= _EVAL_151;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_328 <= _EVAL_127;
      end else begin
        _EVAL_328 <= _EVAL_102;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_330 <= _EVAL_54;
      end else begin
        _EVAL_330 <= _EVAL_11;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_331 <= _EVAL_142;
      end else begin
        _EVAL_331 <= _EVAL_130;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_332 <= _EVAL_120;
      end else begin
        _EVAL_332 <= _EVAL_99;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_333 <= _EVAL_143;
      end else begin
        _EVAL_333 <= _EVAL_5;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_335 <= _EVAL_37;
      end else begin
        _EVAL_335 <= _EVAL_137;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_336 <= _EVAL_82;
      end else begin
        _EVAL_336 <= _EVAL_92;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_337 <= _EVAL_82;
      end else begin
        _EVAL_337 <= _EVAL_92;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_338 <= _EVAL_117;
      end else begin
        _EVAL_338 <= _EVAL_31;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_339 <= _EVAL_151;
      end else begin
        _EVAL_339 <= _EVAL_14;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_340 <= _EVAL_23;
      end else begin
        _EVAL_340 <= _EVAL_29;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_342 <= _EVAL_47;
      end else begin
        _EVAL_342 <= _EVAL_149;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_343 <= _EVAL_47;
      end else begin
        _EVAL_343 <= _EVAL_149;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_345 <= _EVAL_168;
      end else begin
        _EVAL_345 <= _EVAL_184;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_346 <= _EVAL_68;
      end else begin
        _EVAL_346 <= _EVAL_158;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_348 <= _EVAL_23;
      end else begin
        _EVAL_348 <= _EVAL_29;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_349 <= _EVAL_142;
      end else begin
        _EVAL_349 <= _EVAL_130;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_350 <= _EVAL_97;
      end else begin
        _EVAL_350 <= _EVAL_178;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_352 <= _EVAL_174;
      end else begin
        _EVAL_352 <= _EVAL_110;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_353 <= _EVAL_142;
      end else begin
        _EVAL_353 <= _EVAL_130;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_355 <= _EVAL_184;
      end else begin
        _EVAL_355 <= _EVAL_168;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_356 <= _EVAL_105;
      end else begin
        _EVAL_356 <= _EVAL_161;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_358 <= _EVAL_175;
      end else begin
        _EVAL_358 <= _EVAL_64;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_360 <= _EVAL_126;
      end else begin
        _EVAL_360 <= _EVAL_101;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_361 <= _EVAL_89;
      end else begin
        _EVAL_361 <= _EVAL_108;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_363 <= _EVAL_167;
      end else begin
        _EVAL_363 <= 1'h0;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_365 <= _EVAL_33;
      end else begin
        _EVAL_365 <= _EVAL_115;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_366 <= _EVAL_54;
      end else begin
        _EVAL_366 <= _EVAL_11;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_368 <= _EVAL_117;
      end else begin
        _EVAL_368 <= _EVAL_31;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_371 <= _EVAL_89;
      end else begin
        _EVAL_371 <= _EVAL_108;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_372 <= _EVAL_107;
      end else begin
        _EVAL_372 <= _EVAL_72;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_374 <= _EVAL_95;
      end else begin
        _EVAL_374 <= _EVAL_7;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_375 <= _EVAL_139;
      end else begin
        _EVAL_375 <= _EVAL_164;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_376 <= _EVAL_95;
      end else begin
        _EVAL_376 <= _EVAL_7;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_377 <= _EVAL_127;
      end else begin
        _EVAL_377 <= _EVAL_102;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_387 <= _EVAL_64;
      end else begin
        _EVAL_387 <= _EVAL_175;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_388 <= _EVAL_7;
      end else begin
        _EVAL_388 <= _EVAL_95;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_389 <= _EVAL_122;
      end else begin
        _EVAL_389 <= _EVAL_114;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_390 <= _EVAL_169;
      end else begin
        _EVAL_390 <= _EVAL_88;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_391 <= _EVAL_148;
      end else begin
        _EVAL_391 <= _EVAL_63;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_392 <= _EVAL_16;
      end else begin
        _EVAL_392 <= _EVAL_35;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_393 <= _EVAL_154;
      end else begin
        _EVAL_393 <= _EVAL_48;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_398 <= _EVAL_11;
      end else begin
        _EVAL_398 <= _EVAL_54;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_400 <= _EVAL_5;
      end else begin
        _EVAL_400 <= _EVAL_143;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_402 <= _EVAL_148;
      end else begin
        _EVAL_402 <= _EVAL_63;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_413 <= _EVAL_167;
      end else begin
        _EVAL_413 <= 1'h0;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_414 <= _EVAL_178;
      end else begin
        _EVAL_414 <= _EVAL_97;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_415 <= 1'h0;
      end else begin
        _EVAL_415 <= _EVAL_167;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_416 <= _EVAL_87;
      end else begin
        _EVAL_416 <= _EVAL_116;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_420 <= _EVAL_47;
      end else begin
        _EVAL_420 <= _EVAL_149;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_421 <= _EVAL_46;
      end else begin
        _EVAL_421 <= _EVAL_157;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_422 <= _EVAL_15;
      end else begin
        _EVAL_422 <= _EVAL_172;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_424 <= _EVAL_62;
      end else begin
        _EVAL_424 <= _EVAL_58;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_425 <= _EVAL_88;
      end else begin
        _EVAL_425 <= _EVAL_169;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_426 <= _EVAL_10;
      end else begin
        _EVAL_426 <= _EVAL_150;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_428 <= _EVAL_39;
      end else begin
        _EVAL_428 <= _EVAL_41;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_429 <= _EVAL_156;
      end else begin
        _EVAL_429 <= _EVAL_80;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_430 <= _EVAL_161;
      end else begin
        _EVAL_430 <= _EVAL_105;
      end
    end
    if (_EVAL_50) begin
      _EVAL_431 <= 3'h0;
    end else begin
      if (_EVAL_320) begin
        _EVAL_431 <= _EVAL_627;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_433 <= _EVAL_28;
      end else begin
        _EVAL_433 <= _EVAL_177;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_434 <= _EVAL_29;
      end else begin
        _EVAL_434 <= _EVAL_23;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_436 <= _EVAL_151;
      end else begin
        _EVAL_436 <= _EVAL_14;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_439 <= _EVAL_148;
      end else begin
        _EVAL_439 <= _EVAL_63;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_440 <= _EVAL_58;
      end else begin
        _EVAL_440 <= _EVAL_62;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_442 <= _EVAL_104;
      end else begin
        _EVAL_442 <= _EVAL_55;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_444 <= _EVAL_184;
      end else begin
        _EVAL_444 <= _EVAL_168;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_445 <= _EVAL_157;
      end else begin
        _EVAL_445 <= _EVAL_46;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_447 <= _EVAL_175;
      end else begin
        _EVAL_447 <= _EVAL_64;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_451 <= _EVAL_103;
      end else begin
        _EVAL_451 <= _EVAL_1;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_453 <= _EVAL_110;
      end else begin
        _EVAL_453 <= _EVAL_174;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_455 <= _EVAL_100;
      end else begin
        _EVAL_455 <= _EVAL_86;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_456 <= _EVAL_92;
      end else begin
        _EVAL_456 <= _EVAL_82;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_457 <= _EVAL_28;
      end else begin
        _EVAL_457 <= _EVAL_177;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_460 <= _EVAL_11;
      end else begin
        _EVAL_460 <= _EVAL_54;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_461 <= _EVAL_86;
      end else begin
        _EVAL_461 <= _EVAL_100;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_467 <= _EVAL_101;
      end else begin
        _EVAL_467 <= _EVAL_126;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_468 <= _EVAL_63;
      end else begin
        _EVAL_468 <= _EVAL_148;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_470 <= _EVAL_15;
      end else begin
        _EVAL_470 <= _EVAL_172;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_471 <= _EVAL_23;
      end else begin
        _EVAL_471 <= _EVAL_29;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_472 <= _EVAL_29;
      end else begin
        _EVAL_472 <= _EVAL_23;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_473 <= _EVAL_114;
      end else begin
        _EVAL_473 <= _EVAL_122;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_474 <= _EVAL_31;
      end else begin
        _EVAL_474 <= _EVAL_117;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_475 <= _EVAL_80;
      end else begin
        _EVAL_475 <= _EVAL_156;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_476 <= _EVAL_157;
      end else begin
        _EVAL_476 <= _EVAL_46;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_479 <= _EVAL_16;
      end else begin
        _EVAL_479 <= _EVAL_35;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_480 <= _EVAL_10;
      end else begin
        _EVAL_480 <= _EVAL_150;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_482 <= _EVAL_55;
      end else begin
        _EVAL_482 <= _EVAL_104;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_484 <= _EVAL_119;
      end else begin
        _EVAL_484 <= _EVAL_71;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_488 <= _EVAL_15;
      end else begin
        _EVAL_488 <= _EVAL_172;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_489 <= _EVAL_161;
      end else begin
        _EVAL_489 <= _EVAL_105;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_490 <= _EVAL_103;
      end else begin
        _EVAL_490 <= _EVAL_1;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_491 <= _EVAL_108;
      end else begin
        _EVAL_491 <= _EVAL_89;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_494 <= _EVAL_100;
      end else begin
        _EVAL_494 <= _EVAL_86;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_497 <= _EVAL_25;
      end else begin
        _EVAL_497 <= _EVAL_135;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_498 <= _EVAL_41;
      end else begin
        _EVAL_498 <= _EVAL_39;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_499 <= _EVAL_10;
      end else begin
        _EVAL_499 <= _EVAL_150;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_500 <= _EVAL_135;
      end else begin
        _EVAL_500 <= _EVAL_25;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_502 <= _EVAL_115;
      end else begin
        _EVAL_502 <= _EVAL_33;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_504 <= 1'h0;
      end else begin
        _EVAL_504 <= _EVAL_167;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_505 <= _EVAL_172;
      end else begin
        _EVAL_505 <= _EVAL_15;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_507 <= _EVAL_10;
      end else begin
        _EVAL_507 <= _EVAL_150;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_508 <= _EVAL_12;
      end else begin
        _EVAL_508 <= _EVAL_44;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_509 <= _EVAL_48;
      end else begin
        _EVAL_509 <= _EVAL_154;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_510 <= _EVAL_150;
      end else begin
        _EVAL_510 <= _EVAL_10;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_511 <= _EVAL_75;
      end else begin
        _EVAL_511 <= _EVAL_76;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_513 <= _EVAL_126;
      end else begin
        _EVAL_513 <= _EVAL_101;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_515 <= _EVAL_29;
      end else begin
        _EVAL_515 <= _EVAL_23;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_517 <= _EVAL_161;
      end else begin
        _EVAL_517 <= _EVAL_105;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_518 <= _EVAL_75;
      end else begin
        _EVAL_518 <= _EVAL_76;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_519 <= _EVAL_55;
      end else begin
        _EVAL_519 <= _EVAL_104;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_521 <= _EVAL_76;
      end else begin
        _EVAL_521 <= _EVAL_75;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_522 <= _EVAL_151;
      end else begin
        _EVAL_522 <= _EVAL_14;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_524 <= _EVAL_23;
      end else begin
        _EVAL_524 <= _EVAL_29;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_525 <= _EVAL_151;
      end else begin
        _EVAL_525 <= _EVAL_14;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_527 <= _EVAL_88;
      end else begin
        _EVAL_527 <= _EVAL_169;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_528 <= _EVAL_68;
      end else begin
        _EVAL_528 <= _EVAL_158;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_530 <= _EVAL_76;
      end else begin
        _EVAL_530 <= _EVAL_75;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_533 <= _EVAL_137;
      end else begin
        _EVAL_533 <= _EVAL_37;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_534 <= _EVAL_87;
      end else begin
        _EVAL_534 <= _EVAL_116;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_536 <= _EVAL_102;
      end else begin
        _EVAL_536 <= _EVAL_127;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_537 <= _EVAL_178;
      end else begin
        _EVAL_537 <= _EVAL_97;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_538 <= _EVAL_1;
      end else begin
        _EVAL_538 <= _EVAL_103;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_541 <= _EVAL_101;
      end else begin
        _EVAL_541 <= _EVAL_126;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_545 <= _EVAL_35;
      end else begin
        _EVAL_545 <= _EVAL_16;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_546 <= _EVAL_76;
      end else begin
        _EVAL_546 <= _EVAL_75;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_547 <= _EVAL_115;
      end else begin
        _EVAL_547 <= _EVAL_33;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_548 <= _EVAL_29;
      end else begin
        _EVAL_548 <= _EVAL_23;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_551 <= _EVAL_11;
      end else begin
        _EVAL_551 <= _EVAL_54;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_554 <= _EVAL_5;
      end else begin
        _EVAL_554 <= _EVAL_143;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_555 <= _EVAL_75;
      end else begin
        _EVAL_555 <= _EVAL_76;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_556 <= _EVAL_36;
      end else begin
        _EVAL_556 <= _EVAL;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_558 <= _EVAL_99;
      end else begin
        _EVAL_558 <= _EVAL_120;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_559 <= _EVAL_47;
      end else begin
        _EVAL_559 <= _EVAL_149;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_560 <= _EVAL_131;
      end else begin
        _EVAL_560 <= _EVAL_147;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_561 <= _EVAL_14;
      end else begin
        _EVAL_561 <= _EVAL_151;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_562 <= _EVAL_172;
      end else begin
        _EVAL_562 <= _EVAL_15;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_563 <= _EVAL_75;
      end else begin
        _EVAL_563 <= _EVAL_76;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_564 <= _EVAL_172;
      end else begin
        _EVAL_564 <= _EVAL_15;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_565 <= _EVAL_25;
      end else begin
        _EVAL_565 <= _EVAL_135;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_566 <= _EVAL_71;
      end else begin
        _EVAL_566 <= _EVAL_119;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_568 <= _EVAL_137;
      end else begin
        _EVAL_568 <= _EVAL_37;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_569 <= _EVAL_117;
      end else begin
        _EVAL_569 <= _EVAL_31;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_571 <= _EVAL_154;
      end else begin
        _EVAL_571 <= _EVAL_48;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_573 <= _EVAL_7;
      end else begin
        _EVAL_573 <= _EVAL_95;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_574 <= _EVAL_31;
      end else begin
        _EVAL_574 <= _EVAL_117;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_576 <= _EVAL_39;
      end else begin
        _EVAL_576 <= _EVAL_41;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_579 <= _EVAL_104;
      end else begin
        _EVAL_579 <= _EVAL_55;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_580 <= _EVAL_174;
      end else begin
        _EVAL_580 <= _EVAL_110;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_581 <= _EVAL_157;
      end else begin
        _EVAL_581 <= _EVAL_46;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_582 <= _EVAL_150;
      end else begin
        _EVAL_582 <= _EVAL_10;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_584 <= _EVAL_99;
      end else begin
        _EVAL_584 <= _EVAL_120;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_587 <= _EVAL_114;
      end else begin
        _EVAL_587 <= _EVAL_122;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_589 <= _EVAL_156;
      end else begin
        _EVAL_589 <= _EVAL_80;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_591 <= _EVAL_110;
      end else begin
        _EVAL_591 <= _EVAL_174;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_593 <= _EVAL_31;
      end else begin
        _EVAL_593 <= _EVAL_117;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_594 <= _EVAL_156;
      end else begin
        _EVAL_594 <= _EVAL_80;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_596 <= _EVAL_135;
      end else begin
        _EVAL_596 <= _EVAL_25;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_597 <= _EVAL_164;
      end else begin
        _EVAL_597 <= _EVAL_139;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_598 <= _EVAL_104;
      end else begin
        _EVAL_598 <= _EVAL_55;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_599 <= _EVAL;
      end else begin
        _EVAL_599 <= _EVAL_36;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_600 <= _EVAL_150;
      end else begin
        _EVAL_600 <= _EVAL_10;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_601 <= _EVAL_167;
      end else begin
        _EVAL_601 <= 1'h0;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_602 <= _EVAL_31;
      end else begin
        _EVAL_602 <= _EVAL_117;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_603 <= _EVAL_72;
      end else begin
        _EVAL_603 <= _EVAL_107;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_604 <= _EVAL_143;
      end else begin
        _EVAL_604 <= _EVAL_5;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_606 <= _EVAL_172;
      end else begin
        _EVAL_606 <= _EVAL_15;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_607 <= _EVAL_36;
      end else begin
        _EVAL_607 <= _EVAL;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_608 <= _EVAL_7;
      end else begin
        _EVAL_608 <= _EVAL_95;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_609 <= _EVAL_184;
      end else begin
        _EVAL_609 <= _EVAL_168;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_611 <= _EVAL_177;
      end else begin
        _EVAL_611 <= _EVAL_28;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_612 <= _EVAL_116;
      end else begin
        _EVAL_612 <= _EVAL_87;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_614 <= _EVAL_143;
      end else begin
        _EVAL_614 <= _EVAL_5;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_615 <= _EVAL_12;
      end else begin
        _EVAL_615 <= _EVAL_44;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_618 <= _EVAL_104;
      end else begin
        _EVAL_618 <= _EVAL_55;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_619 <= _EVAL_178;
      end else begin
        _EVAL_619 <= _EVAL_97;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_620 <= _EVAL_25;
      end else begin
        _EVAL_620 <= _EVAL_135;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_621 <= _EVAL_92;
      end else begin
        _EVAL_621 <= _EVAL_82;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_622 <= _EVAL_119;
      end else begin
        _EVAL_622 <= _EVAL_71;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_623 <= _EVAL_58;
      end else begin
        _EVAL_623 <= _EVAL_62;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_625 <= _EVAL_116;
      end else begin
        _EVAL_625 <= _EVAL_87;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_626 <= _EVAL_46;
      end else begin
        _EVAL_626 <= _EVAL_157;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_630 <= _EVAL_105;
      end else begin
        _EVAL_630 <= _EVAL_161;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_633 <= _EVAL_33;
      end else begin
        _EVAL_633 <= _EVAL_115;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_634 <= _EVAL_63;
      end else begin
        _EVAL_634 <= _EVAL_148;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_638 <= _EVAL_62;
      end else begin
        _EVAL_638 <= _EVAL_58;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_640 <= _EVAL_178;
      end else begin
        _EVAL_640 <= _EVAL_97;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_644 <= _EVAL_175;
      end else begin
        _EVAL_644 <= _EVAL_64;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_646 <= _EVAL_143;
      end else begin
        _EVAL_646 <= _EVAL_5;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_648 <= _EVAL_97;
      end else begin
        _EVAL_648 <= _EVAL_178;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_651 <= _EVAL_64;
      end else begin
        _EVAL_651 <= _EVAL_175;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_653 <= _EVAL_72;
      end else begin
        _EVAL_653 <= _EVAL_107;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_655 <= _EVAL_164;
      end else begin
        _EVAL_655 <= _EVAL_139;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_657 <= _EVAL_64;
      end else begin
        _EVAL_657 <= _EVAL_175;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_658 <= _EVAL_44;
      end else begin
        _EVAL_658 <= _EVAL_12;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_661 <= _EVAL_88;
      end else begin
        _EVAL_661 <= _EVAL_169;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_663 <= _EVAL_103;
      end else begin
        _EVAL_663 <= _EVAL_1;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_665 <= _EVAL_95;
      end else begin
        _EVAL_665 <= _EVAL_7;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_667 <= _EVAL_1;
      end else begin
        _EVAL_667 <= _EVAL_103;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_668 <= _EVAL_107;
      end else begin
        _EVAL_668 <= _EVAL_72;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_672 <= _EVAL_142;
      end else begin
        _EVAL_672 <= _EVAL_130;
      end
    end
    if (_EVAL_50) begin
      _EVAL_673 <= 4'h1;
    end else begin
      if (_EVAL_214) begin
        _EVAL_673 <= _EVAL_700;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_675 <= _EVAL_39;
      end else begin
        _EVAL_675 <= _EVAL_41;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_681 <= _EVAL_97;
      end else begin
        _EVAL_681 <= _EVAL_178;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_682 <= _EVAL_16;
      end else begin
        _EVAL_682 <= _EVAL_35;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_683 <= _EVAL;
      end else begin
        _EVAL_683 <= _EVAL_36;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_684 <= _EVAL_158;
      end else begin
        _EVAL_684 <= _EVAL_68;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_685 <= _EVAL_107;
      end else begin
        _EVAL_685 <= _EVAL_72;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_687 <= _EVAL_80;
      end else begin
        _EVAL_687 <= _EVAL_156;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_688 <= _EVAL_120;
      end else begin
        _EVAL_688 <= _EVAL_99;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_689 <= _EVAL_108;
      end else begin
        _EVAL_689 <= _EVAL_89;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_692 <= _EVAL;
      end else begin
        _EVAL_692 <= _EVAL_36;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_693 <= _EVAL_41;
      end else begin
        _EVAL_693 <= _EVAL_39;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_695 <= _EVAL_177;
      end else begin
        _EVAL_695 <= _EVAL_28;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_696 <= _EVAL_139;
      end else begin
        _EVAL_696 <= _EVAL_164;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_697 <= _EVAL_164;
      end else begin
        _EVAL_697 <= _EVAL_139;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_698 <= _EVAL_99;
      end else begin
        _EVAL_698 <= _EVAL_120;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_699 <= _EVAL_51;
      end else begin
        _EVAL_699 <= _EVAL_181;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_701 <= _EVAL_137;
      end else begin
        _EVAL_701 <= _EVAL_37;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_702 <= _EVAL_54;
      end else begin
        _EVAL_702 <= _EVAL_11;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_703 <= _EVAL_1;
      end else begin
        _EVAL_703 <= _EVAL_103;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_708 <= _EVAL_15;
      end else begin
        _EVAL_708 <= _EVAL_172;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_711 <= _EVAL_37;
      end else begin
        _EVAL_711 <= _EVAL_137;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_714 <= _EVAL_114;
      end else begin
        _EVAL_714 <= _EVAL_122;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_716 <= _EVAL_115;
      end else begin
        _EVAL_716 <= _EVAL_33;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_717 <= _EVAL_54;
      end else begin
        _EVAL_717 <= _EVAL_11;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_718 <= _EVAL_89;
      end else begin
        _EVAL_718 <= _EVAL_108;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_719 <= _EVAL_64;
      end else begin
        _EVAL_719 <= _EVAL_175;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_720 <= _EVAL_80;
      end else begin
        _EVAL_720 <= _EVAL_156;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_721 <= _EVAL_92;
      end else begin
        _EVAL_721 <= _EVAL_82;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_722 <= _EVAL_157;
      end else begin
        _EVAL_722 <= _EVAL_46;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_723 <= _EVAL_130;
      end else begin
        _EVAL_723 <= _EVAL_142;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_725 <= _EVAL_36;
      end else begin
        _EVAL_725 <= _EVAL;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_726 <= _EVAL_181;
      end else begin
        _EVAL_726 <= _EVAL_51;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_727 <= _EVAL_51;
      end else begin
        _EVAL_727 <= _EVAL_181;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_728 <= _EVAL_154;
      end else begin
        _EVAL_728 <= _EVAL_48;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_729 <= _EVAL_86;
      end else begin
        _EVAL_729 <= _EVAL_100;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_731 <= _EVAL_37;
      end else begin
        _EVAL_731 <= _EVAL_137;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_732 <= _EVAL_120;
      end else begin
        _EVAL_732 <= _EVAL_99;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_734 <= _EVAL_35;
      end else begin
        _EVAL_734 <= _EVAL_16;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_735 <= _EVAL_95;
      end else begin
        _EVAL_735 <= _EVAL_7;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_736 <= _EVAL_46;
      end else begin
        _EVAL_736 <= _EVAL_157;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_737 <= _EVAL_105;
      end else begin
        _EVAL_737 <= _EVAL_161;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_738 <= _EVAL_137;
      end else begin
        _EVAL_738 <= _EVAL_37;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_739 <= _EVAL_130;
      end else begin
        _EVAL_739 <= _EVAL_142;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_740 <= _EVAL_158;
      end else begin
        _EVAL_740 <= _EVAL_68;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_742 <= _EVAL_5;
      end else begin
        _EVAL_742 <= _EVAL_143;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_743 <= _EVAL_150;
      end else begin
        _EVAL_743 <= _EVAL_10;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_744 <= _EVAL_35;
      end else begin
        _EVAL_744 <= _EVAL_16;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_747 <= _EVAL_48;
      end else begin
        _EVAL_747 <= _EVAL_154;
      end
    end
    if (_EVAL_50) begin
      _EVAL_748 <= 3'h0;
    end else begin
      if (_EVAL_552) begin
        if (_EVAL_553) begin
          _EVAL_748 <= _EVAL_224;
        end else begin
          _EVAL_748 <= _EVAL_691;
        end
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_750 <= _EVAL;
      end else begin
        _EVAL_750 <= _EVAL_36;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_751 <= _EVAL_48;
      end else begin
        _EVAL_751 <= _EVAL_154;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_753 <= _EVAL_89;
      end else begin
        _EVAL_753 <= _EVAL_108;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_754 <= _EVAL_62;
      end else begin
        _EVAL_754 <= _EVAL_58;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_756 <= _EVAL_14;
      end else begin
        _EVAL_756 <= _EVAL_151;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_758 <= _EVAL_119;
      end else begin
        _EVAL_758 <= _EVAL_71;
      end
    end
    if (_EVAL_592) begin
      if (_EVAL_253) begin
        _EVAL_760 <= _EVAL_164;
      end else begin
        _EVAL_760 <= _EVAL_139;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_761 <= _EVAL_184;
      end else begin
        _EVAL_761 <= _EVAL_168;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_762 <= _EVAL_119;
      end else begin
        _EVAL_762 <= _EVAL_71;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_763 <= _EVAL_86;
      end else begin
        _EVAL_763 <= _EVAL_100;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_764 <= _EVAL_116;
      end else begin
        _EVAL_764 <= _EVAL_87;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_765 <= _EVAL_135;
      end else begin
        _EVAL_765 <= _EVAL_25;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_768 <= _EVAL_103;
      end else begin
        _EVAL_768 <= _EVAL_1;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_770 <= _EVAL_92;
      end else begin
        _EVAL_770 <= _EVAL_82;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_772 <= _EVAL_12;
      end else begin
        _EVAL_772 <= _EVAL_44;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_773 <= _EVAL_100;
      end else begin
        _EVAL_773 <= _EVAL_86;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_774 <= _EVAL_39;
      end else begin
        _EVAL_774 <= _EVAL_41;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_776 <= _EVAL_58;
      end else begin
        _EVAL_776 <= _EVAL_62;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_777 <= _EVAL_131;
      end else begin
        _EVAL_777 <= _EVAL_147;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_778 <= _EVAL_46;
      end else begin
        _EVAL_778 <= _EVAL_157;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_780 <= _EVAL_122;
      end else begin
        _EVAL_780 <= _EVAL_114;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_781 <= _EVAL_126;
      end else begin
        _EVAL_781 <= _EVAL_101;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_782 <= _EVAL_116;
      end else begin
        _EVAL_782 <= _EVAL_87;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_786 <= _EVAL_139;
      end else begin
        _EVAL_786 <= _EVAL_164;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_787 <= _EVAL_101;
      end else begin
        _EVAL_787 <= _EVAL_126;
      end
    end
    if (_EVAL_50) begin
      _EVAL_788 <= 4'h1;
    end else begin
      if (_EVAL_710) begin
        _EVAL_788 <= _EVAL_438;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_789 <= _EVAL_148;
      end else begin
        _EVAL_789 <= _EVAL_63;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_792 <= _EVAL_130;
      end else begin
        _EVAL_792 <= _EVAL_142;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_793 <= _EVAL_110;
      end else begin
        _EVAL_793 <= _EVAL_174;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_796 <= _EVAL_127;
      end else begin
        _EVAL_796 <= _EVAL_102;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_797 <= _EVAL_149;
      end else begin
        _EVAL_797 <= _EVAL_47;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_798 <= _EVAL_97;
      end else begin
        _EVAL_798 <= _EVAL_178;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_799 <= _EVAL_149;
      end else begin
        _EVAL_799 <= _EVAL_47;
      end
    end
    if (_EVAL_250) begin
      if (_EVAL_253) begin
        _EVAL_800 <= _EVAL_117;
      end else begin
        _EVAL_800 <= _EVAL_31;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_801 <= _EVAL_12;
      end else begin
        _EVAL_801 <= _EVAL_44;
      end
    end
    if (_EVAL_724) begin
      if (_EVAL_253) begin
        _EVAL_804 <= _EVAL_87;
      end else begin
        _EVAL_804 <= _EVAL_116;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_805 <= _EVAL_72;
      end else begin
        _EVAL_805 <= _EVAL_107;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_806 <= _EVAL_177;
      end else begin
        _EVAL_806 <= _EVAL_28;
      end
    end
    if (_EVAL_567) begin
      if (_EVAL_253) begin
        _EVAL_807 <= _EVAL_177;
      end else begin
        _EVAL_807 <= _EVAL_28;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_808 <= _EVAL_181;
      end else begin
        _EVAL_808 <= _EVAL_51;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_809 <= _EVAL_35;
      end else begin
        _EVAL_809 <= _EVAL_16;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_810 <= _EVAL_41;
      end else begin
        _EVAL_810 <= _EVAL_39;
      end
    end
    if (_EVAL_483) begin
      if (_EVAL_253) begin
        _EVAL_811 <= _EVAL_72;
      end else begin
        _EVAL_811 <= _EVAL_107;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_812 <= _EVAL_154;
      end else begin
        _EVAL_812 <= _EVAL_48;
      end
    end
    if (_EVAL_193) begin
      if (_EVAL_253) begin
        _EVAL_815 <= _EVAL_167;
      end else begin
        _EVAL_815 <= 1'h0;
      end
    end
    if (_EVAL_707) begin
      if (_EVAL_253) begin
        _EVAL_817 <= _EVAL_174;
      end else begin
        _EVAL_817 <= _EVAL_110;
      end
    end
    if (_EVAL_501) begin
      if (_EVAL_253) begin
        _EVAL_818 <= _EVAL_147;
      end else begin
        _EVAL_818 <= _EVAL_131;
      end
    end
  end
endmodule
