//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_18(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [63:0] _EVAL_5,
  output [31:0] _EVAL_6,
  output [1:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  output [3:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input  [7:0]  _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output [2:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23,
  input  [2:0]  _EVAL_24,
  input         _EVAL_25,
  input  [63:0] _EVAL_26,
  output [2:0]  _EVAL_27,
  output [1:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  input  [2:0]  _EVAL_30,
  input         _EVAL_31,
  input  [1:0]  _EVAL_32,
  output [63:0] _EVAL_33,
  input  [2:0]  _EVAL_34,
  input  [3:0]  _EVAL_35,
  input         _EVAL_36,
  output        _EVAL_37,
  output [3:0]  _EVAL_38,
  output [3:0]  _EVAL_39,
  input  [1:0]  _EVAL_40,
  input  [31:0] _EVAL_41,
  input  [2:0]  _EVAL_42,
  output        _EVAL_43,
  input  [31:0] _EVAL_44,
  input  [2:0]  _EVAL_45,
  input  [2:0]  _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  output [2:0]  _EVAL_49,
  output [31:0] _EVAL_50,
  output [63:0] _EVAL_51,
  output [1:0]  _EVAL_52,
  input  [1:0]  _EVAL_53,
  output [3:0]  _EVAL_54,
  input  [3:0]  _EVAL_55,
  output        _EVAL_56,
  output [1:0]  _EVAL_57,
  output [1:0]  _EVAL_58,
  output [7:0]  _EVAL_59,
  output        _EVAL_60,
  output [3:0]  _EVAL_61,
  input         _EVAL_62,
  input  [2:0]  _EVAL_63,
  input         _EVAL_64,
  input  [3:0]  _EVAL_65,
  output [1:0]  _EVAL_66,
  output        _EVAL_67,
  input  [1:0]  _EVAL_68,
  input  [2:0]  _EVAL_69,
  input  [3:0]  _EVAL_70,
  input         _EVAL_71,
  output [63:0] _EVAL_72,
  output [1:0]  _EVAL_73,
  output        _EVAL_74,
  input  [63:0] _EVAL_75,
  output [2:0]  _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output        _EVAL_79,
  output [1:0]  _EVAL_80,
  output        _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input  [3:0]  _EVAL_84,
  output [31:0] _EVAL_85,
  output [3:0]  _EVAL_86,
  output [3:0]  _EVAL_87,
  output [3:0]  _EVAL_88,
  output [63:0] _EVAL_89,
  input         _EVAL_90,
  output [31:0] _EVAL_91,
  input  [63:0] _EVAL_92,
  output [2:0]  _EVAL_93,
  output [1:0]  _EVAL_94,
  input  [3:0]  _EVAL_95,
  output        _EVAL_96,
  input         _EVAL_97,
  input         _EVAL_98,
  input  [1:0]  _EVAL_99,
  input         _EVAL_100,
  input  [31:0] _EVAL_101,
  input  [63:0] _EVAL_102,
  output        _EVAL_103,
  input         _EVAL_104,
  input  [7:0]  _EVAL_105,
  input  [1:0]  _EVAL_106,
  input         _EVAL_107
);
  wire  buffer__EVAL;
  wire [3:0] buffer__EVAL_0;
  wire [3:0] buffer__EVAL_1;
  wire [31:0] buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [31:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [63:0] buffer__EVAL_8;
  wire [31:0] buffer__EVAL_9;
  wire [7:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire [63:0] buffer__EVAL_13;
  wire [1:0] buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire [3:0] buffer__EVAL_16;
  wire [2:0] buffer__EVAL_17;
  wire [2:0] buffer__EVAL_18;
  wire [1:0] buffer__EVAL_19;
  wire [3:0] buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire [1:0] buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire [3:0] buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire [63:0] buffer__EVAL_34;
  wire [31:0] buffer__EVAL_35;
  wire [3:0] buffer__EVAL_36;
  wire  buffer__EVAL_37;
  wire [2:0] buffer__EVAL_38;
  wire [63:0] buffer__EVAL_39;
  wire [2:0] buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire [3:0] buffer__EVAL_42;
  wire [2:0] buffer__EVAL_43;
  wire [2:0] buffer__EVAL_44;
  wire [2:0] buffer__EVAL_45;
  wire [31:0] buffer__EVAL_46;
  wire [3:0] buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire [31:0] buffer__EVAL_49;
  wire  buffer__EVAL_50;
  wire [3:0] buffer__EVAL_51;
  wire  buffer__EVAL_52;
  wire  buffer__EVAL_53;
  wire [3:0] buffer__EVAL_54;
  wire [2:0] buffer__EVAL_55;
  wire [63:0] buffer__EVAL_56;
  wire  buffer__EVAL_57;
  wire  buffer__EVAL_58;
  wire  buffer__EVAL_59;
  wire [63:0] buffer__EVAL_60;
  wire  buffer__EVAL_61;
  wire  buffer__EVAL_62;
  wire [2:0] buffer__EVAL_63;
  wire [3:0] buffer__EVAL_64;
  wire [3:0] buffer__EVAL_65;
  wire  buffer__EVAL_66;
  wire [7:0] buffer__EVAL_67;
  wire [2:0] buffer__EVAL_68;
  wire [1:0] buffer__EVAL_69;
  wire  buffer__EVAL_70;
  wire  rsink__EVAL;
  wire [2:0] rsink__EVAL_0;
  wire [2:0] rsink__EVAL_1;
  wire [63:0] rsink__EVAL_2;
  wire  rsink__EVAL_3;
  wire  rsink__EVAL_4;
  wire [63:0] rsink__EVAL_5;
  wire [1:0] rsink__EVAL_6;
  wire  rsink__EVAL_7;
  wire  rsink__EVAL_8;
  wire [2:0] rsink__EVAL_9;
  wire [2:0] rsink__EVAL_10;
  wire [31:0] rsink__EVAL_11;
  wire  rsink__EVAL_12;
  wire  rsink__EVAL_13;
  wire [1:0] rsink__EVAL_14;
  wire [1:0] rsink__EVAL_15;
  wire [1:0] rsink__EVAL_16;
  wire  rsink__EVAL_17;
  wire  rsink__EVAL_18;
  wire  rsink__EVAL_19;
  wire [63:0] rsink__EVAL_20;
  wire [31:0] rsink__EVAL_21;
  wire [2:0] rsink__EVAL_22;
  wire [3:0] rsink__EVAL_23;
  wire [3:0] rsink__EVAL_24;
  wire [2:0] rsink__EVAL_25;
  wire  rsink__EVAL_26;
  wire [63:0] rsink__EVAL_27;
  wire [1:0] rsink__EVAL_28;
  wire [1:0] rsink__EVAL_29;
  wire [1:0] rsink__EVAL_30;
  wire  rsink__EVAL_31;
  wire [2:0] rsink__EVAL_32;
  wire [31:0] rsink__EVAL_33;
  wire [3:0] rsink__EVAL_34;
  wire [2:0] rsink__EVAL_35;
  wire [2:0] rsink__EVAL_36;
  wire  rsink__EVAL_37;
  wire  rsink__EVAL_38;
  wire [1:0] rsink__EVAL_39;
  wire [3:0] rsink__EVAL_40;
  wire  rsink__EVAL_41;
  wire  rsink__EVAL_42;
  wire [1:0] rsink__EVAL_43;
  wire [1:0] rsink__EVAL_44;
  wire [3:0] rsink__EVAL_45;
  wire  rsink__EVAL_46;
  wire [7:0] rsink__EVAL_47;
  wire [3:0] rsink__EVAL_48;
  wire [3:0] rsink__EVAL_49;
  wire [63:0] rsink__EVAL_50;
  wire [1:0] rsink__EVAL_51;
  wire [2:0] rsink__EVAL_52;
  wire [3:0] rsink__EVAL_53;
  wire  rsink__EVAL_54;
  wire [3:0] rsink__EVAL_55;
  wire [3:0] rsink__EVAL_56;
  wire [2:0] rsink__EVAL_57;
  wire [3:0] rsink__EVAL_58;
  wire [3:0] rsink__EVAL_59;
  wire  rsink__EVAL_60;
  wire  rsink__EVAL_61;
  wire  rsink__EVAL_62;
  wire [3:0] rsink__EVAL_63;
  wire [2:0] rsink__EVAL_64;
  wire [31:0] rsink__EVAL_65;
  wire  rsink__EVAL_66;
  wire  rsink__EVAL_67;
  wire [2:0] rsink__EVAL_68;
  wire [1:0] rsink__EVAL_69;
  wire  rsink__EVAL_70;
  wire [3:0] rsink__EVAL_71;
  wire [31:0] rsink__EVAL_72;
  wire  rsink__EVAL_73;
  wire  rsink__EVAL_74;
  wire  rsink__EVAL_75;
  wire  rsink__EVAL_76;
  wire [1:0] rsink__EVAL_77;
  wire [2:0] rsink__EVAL_78;
  wire  rsink__EVAL_79;
  wire [3:0] rsink__EVAL_80;
  wire  rsink__EVAL_81;
  wire  rsink__EVAL_82;
  wire [7:0] rsink__EVAL_83;
  wire [31:0] rsink__EVAL_84;
  wire [31:0] rsink__EVAL_85;
  wire [3:0] rsink__EVAL_86;
  wire [1:0] rsink__EVAL_87;
  wire [63:0] rsink__EVAL_88;
  wire  rsink__EVAL_89;
  wire [31:0] rsink__EVAL_90;
  wire [63:0] rsink__EVAL_91;
  wire [3:0] rsink__EVAL_92;
  wire  rsink__EVAL_93;
  wire [1:0] rsink__EVAL_94;
  wire [3:0] rsink__EVAL_95;
  wire [63:0] rsink__EVAL_96;
  wire [7:0] rsink__EVAL_97;
  wire [31:0] rsink__EVAL_98;
  wire [1:0] rsink__EVAL_99;
  wire  rsink__EVAL_100;
  wire [2:0] rsink__EVAL_101;
  wire [63:0] rsink__EVAL_102;
  wire  rsink__EVAL_103;
  wire  rsink__EVAL_104;
  wire  rsink__EVAL_105;
  wire  rsink__EVAL_106;
  wire  rsink__EVAL_107;
  wire [3:0] fixer__EVAL;
  wire [31:0] fixer__EVAL_0;
  wire [2:0] fixer__EVAL_1;
  wire [63:0] fixer__EVAL_2;
  wire  fixer__EVAL_3;
  wire [2:0] fixer__EVAL_4;
  wire [1:0] fixer__EVAL_5;
  wire  fixer__EVAL_6;
  wire [63:0] fixer__EVAL_7;
  wire  fixer__EVAL_8;
  wire  fixer__EVAL_9;
  wire  fixer__EVAL_10;
  wire [2:0] fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire  fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire [63:0] fixer__EVAL_15;
  wire  fixer__EVAL_16;
  wire [2:0] fixer__EVAL_17;
  wire  fixer__EVAL_18;
  wire  fixer__EVAL_19;
  wire  fixer__EVAL_20;
  wire [31:0] fixer__EVAL_21;
  wire [3:0] fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire [63:0] fixer__EVAL_24;
  wire [3:0] fixer__EVAL_25;
  wire  fixer__EVAL_26;
  wire [31:0] fixer__EVAL_27;
  wire [63:0] fixer__EVAL_28;
  wire  fixer__EVAL_29;
  wire [3:0] fixer__EVAL_30;
  wire  fixer__EVAL_31;
  wire [7:0] fixer__EVAL_32;
  wire [3:0] fixer__EVAL_33;
  wire [7:0] fixer__EVAL_34;
  wire [2:0] fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire [3:0] fixer__EVAL_37;
  wire [3:0] fixer__EVAL_38;
  wire [3:0] fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire [2:0] fixer__EVAL_41;
  wire  fixer__EVAL_42;
  wire [2:0] fixer__EVAL_43;
  wire  fixer__EVAL_44;
  wire  fixer__EVAL_45;
  wire [3:0] fixer__EVAL_46;
  wire [2:0] fixer__EVAL_47;
  wire [2:0] fixer__EVAL_48;
  wire [31:0] fixer__EVAL_49;
  wire [3:0] fixer__EVAL_50;
  wire  fixer__EVAL_51;
  wire  fixer__EVAL_52;
  wire [1:0] fixer__EVAL_53;
  wire  fixer__EVAL_54;
  wire  fixer__EVAL_55;
  wire  fixer__EVAL_56;
  wire  fixer__EVAL_57;
  wire [31:0] fixer__EVAL_58;
  wire  fixer__EVAL_59;
  wire [1:0] fixer__EVAL_60;
  wire  fixer__EVAL_61;
  wire [3:0] fixer__EVAL_62;
  wire [1:0] fixer__EVAL_63;
  wire [3:0] fixer__EVAL_64;
  wire  fixer__EVAL_65;
  wire [2:0] fixer__EVAL_66;
  wire [31:0] fixer__EVAL_67;
  wire  fixer__EVAL_68;
  wire [63:0] fixer__EVAL_69;
  wire  fixer__EVAL_70;
  SiFive__EVAL_4 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48),
    ._EVAL_49(buffer__EVAL_49),
    ._EVAL_50(buffer__EVAL_50),
    ._EVAL_51(buffer__EVAL_51),
    ._EVAL_52(buffer__EVAL_52),
    ._EVAL_53(buffer__EVAL_53),
    ._EVAL_54(buffer__EVAL_54),
    ._EVAL_55(buffer__EVAL_55),
    ._EVAL_56(buffer__EVAL_56),
    ._EVAL_57(buffer__EVAL_57),
    ._EVAL_58(buffer__EVAL_58),
    ._EVAL_59(buffer__EVAL_59),
    ._EVAL_60(buffer__EVAL_60),
    ._EVAL_61(buffer__EVAL_61),
    ._EVAL_62(buffer__EVAL_62),
    ._EVAL_63(buffer__EVAL_63),
    ._EVAL_64(buffer__EVAL_64),
    ._EVAL_65(buffer__EVAL_65),
    ._EVAL_66(buffer__EVAL_66),
    ._EVAL_67(buffer__EVAL_67),
    ._EVAL_68(buffer__EVAL_68),
    ._EVAL_69(buffer__EVAL_69),
    ._EVAL_70(buffer__EVAL_70)
  );
  SiFive__EVAL_17 rsink (
    ._EVAL(rsink__EVAL),
    ._EVAL_0(rsink__EVAL_0),
    ._EVAL_1(rsink__EVAL_1),
    ._EVAL_2(rsink__EVAL_2),
    ._EVAL_3(rsink__EVAL_3),
    ._EVAL_4(rsink__EVAL_4),
    ._EVAL_5(rsink__EVAL_5),
    ._EVAL_6(rsink__EVAL_6),
    ._EVAL_7(rsink__EVAL_7),
    ._EVAL_8(rsink__EVAL_8),
    ._EVAL_9(rsink__EVAL_9),
    ._EVAL_10(rsink__EVAL_10),
    ._EVAL_11(rsink__EVAL_11),
    ._EVAL_12(rsink__EVAL_12),
    ._EVAL_13(rsink__EVAL_13),
    ._EVAL_14(rsink__EVAL_14),
    ._EVAL_15(rsink__EVAL_15),
    ._EVAL_16(rsink__EVAL_16),
    ._EVAL_17(rsink__EVAL_17),
    ._EVAL_18(rsink__EVAL_18),
    ._EVAL_19(rsink__EVAL_19),
    ._EVAL_20(rsink__EVAL_20),
    ._EVAL_21(rsink__EVAL_21),
    ._EVAL_22(rsink__EVAL_22),
    ._EVAL_23(rsink__EVAL_23),
    ._EVAL_24(rsink__EVAL_24),
    ._EVAL_25(rsink__EVAL_25),
    ._EVAL_26(rsink__EVAL_26),
    ._EVAL_27(rsink__EVAL_27),
    ._EVAL_28(rsink__EVAL_28),
    ._EVAL_29(rsink__EVAL_29),
    ._EVAL_30(rsink__EVAL_30),
    ._EVAL_31(rsink__EVAL_31),
    ._EVAL_32(rsink__EVAL_32),
    ._EVAL_33(rsink__EVAL_33),
    ._EVAL_34(rsink__EVAL_34),
    ._EVAL_35(rsink__EVAL_35),
    ._EVAL_36(rsink__EVAL_36),
    ._EVAL_37(rsink__EVAL_37),
    ._EVAL_38(rsink__EVAL_38),
    ._EVAL_39(rsink__EVAL_39),
    ._EVAL_40(rsink__EVAL_40),
    ._EVAL_41(rsink__EVAL_41),
    ._EVAL_42(rsink__EVAL_42),
    ._EVAL_43(rsink__EVAL_43),
    ._EVAL_44(rsink__EVAL_44),
    ._EVAL_45(rsink__EVAL_45),
    ._EVAL_46(rsink__EVAL_46),
    ._EVAL_47(rsink__EVAL_47),
    ._EVAL_48(rsink__EVAL_48),
    ._EVAL_49(rsink__EVAL_49),
    ._EVAL_50(rsink__EVAL_50),
    ._EVAL_51(rsink__EVAL_51),
    ._EVAL_52(rsink__EVAL_52),
    ._EVAL_53(rsink__EVAL_53),
    ._EVAL_54(rsink__EVAL_54),
    ._EVAL_55(rsink__EVAL_55),
    ._EVAL_56(rsink__EVAL_56),
    ._EVAL_57(rsink__EVAL_57),
    ._EVAL_58(rsink__EVAL_58),
    ._EVAL_59(rsink__EVAL_59),
    ._EVAL_60(rsink__EVAL_60),
    ._EVAL_61(rsink__EVAL_61),
    ._EVAL_62(rsink__EVAL_62),
    ._EVAL_63(rsink__EVAL_63),
    ._EVAL_64(rsink__EVAL_64),
    ._EVAL_65(rsink__EVAL_65),
    ._EVAL_66(rsink__EVAL_66),
    ._EVAL_67(rsink__EVAL_67),
    ._EVAL_68(rsink__EVAL_68),
    ._EVAL_69(rsink__EVAL_69),
    ._EVAL_70(rsink__EVAL_70),
    ._EVAL_71(rsink__EVAL_71),
    ._EVAL_72(rsink__EVAL_72),
    ._EVAL_73(rsink__EVAL_73),
    ._EVAL_74(rsink__EVAL_74),
    ._EVAL_75(rsink__EVAL_75),
    ._EVAL_76(rsink__EVAL_76),
    ._EVAL_77(rsink__EVAL_77),
    ._EVAL_78(rsink__EVAL_78),
    ._EVAL_79(rsink__EVAL_79),
    ._EVAL_80(rsink__EVAL_80),
    ._EVAL_81(rsink__EVAL_81),
    ._EVAL_82(rsink__EVAL_82),
    ._EVAL_83(rsink__EVAL_83),
    ._EVAL_84(rsink__EVAL_84),
    ._EVAL_85(rsink__EVAL_85),
    ._EVAL_86(rsink__EVAL_86),
    ._EVAL_87(rsink__EVAL_87),
    ._EVAL_88(rsink__EVAL_88),
    ._EVAL_89(rsink__EVAL_89),
    ._EVAL_90(rsink__EVAL_90),
    ._EVAL_91(rsink__EVAL_91),
    ._EVAL_92(rsink__EVAL_92),
    ._EVAL_93(rsink__EVAL_93),
    ._EVAL_94(rsink__EVAL_94),
    ._EVAL_95(rsink__EVAL_95),
    ._EVAL_96(rsink__EVAL_96),
    ._EVAL_97(rsink__EVAL_97),
    ._EVAL_98(rsink__EVAL_98),
    ._EVAL_99(rsink__EVAL_99),
    ._EVAL_100(rsink__EVAL_100),
    ._EVAL_101(rsink__EVAL_101),
    ._EVAL_102(rsink__EVAL_102),
    ._EVAL_103(rsink__EVAL_103),
    ._EVAL_104(rsink__EVAL_104),
    ._EVAL_105(rsink__EVAL_105),
    ._EVAL_106(rsink__EVAL_106),
    ._EVAL_107(rsink__EVAL_107)
  );
  SiFive__EVAL_6 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40),
    ._EVAL_41(fixer__EVAL_41),
    ._EVAL_42(fixer__EVAL_42),
    ._EVAL_43(fixer__EVAL_43),
    ._EVAL_44(fixer__EVAL_44),
    ._EVAL_45(fixer__EVAL_45),
    ._EVAL_46(fixer__EVAL_46),
    ._EVAL_47(fixer__EVAL_47),
    ._EVAL_48(fixer__EVAL_48),
    ._EVAL_49(fixer__EVAL_49),
    ._EVAL_50(fixer__EVAL_50),
    ._EVAL_51(fixer__EVAL_51),
    ._EVAL_52(fixer__EVAL_52),
    ._EVAL_53(fixer__EVAL_53),
    ._EVAL_54(fixer__EVAL_54),
    ._EVAL_55(fixer__EVAL_55),
    ._EVAL_56(fixer__EVAL_56),
    ._EVAL_57(fixer__EVAL_57),
    ._EVAL_58(fixer__EVAL_58),
    ._EVAL_59(fixer__EVAL_59),
    ._EVAL_60(fixer__EVAL_60),
    ._EVAL_61(fixer__EVAL_61),
    ._EVAL_62(fixer__EVAL_62),
    ._EVAL_63(fixer__EVAL_63),
    ._EVAL_64(fixer__EVAL_64),
    ._EVAL_65(fixer__EVAL_65),
    ._EVAL_66(fixer__EVAL_66),
    ._EVAL_67(fixer__EVAL_67),
    ._EVAL_68(fixer__EVAL_68),
    ._EVAL_69(fixer__EVAL_69),
    ._EVAL_70(fixer__EVAL_70)
  );
  assign buffer__EVAL_55 = _EVAL_29;
  assign rsink__EVAL_63 = _EVAL_35;
  assign _EVAL_6 = buffer__EVAL_49;
  assign _EVAL_22 = buffer__EVAL_15;
  assign buffer__EVAL_50 = fixer__EVAL_55;
  assign rsink__EVAL_58 = fixer__EVAL_46;
  assign _EVAL_81 = buffer__EVAL_28;
  assign _EVAL_54 = rsink__EVAL_56;
  assign fixer__EVAL_29 = rsink__EVAL_37;
  assign buffer__EVAL_35 = _EVAL_101;
  assign fixer__EVAL_27 = rsink__EVAL_90;
  assign rsink__EVAL_76 = fixer__EVAL_6;
  assign rsink__EVAL_23 = _EVAL_10;
  assign _EVAL_76 = buffer__EVAL_38;
  assign buffer__EVAL_31 = _EVAL_0;
  assign _EVAL_38 = buffer__EVAL_42;
  assign rsink__EVAL_93 = _EVAL_18;
  assign _EVAL_57 = rsink__EVAL_94;
  assign buffer__EVAL_39 = fixer__EVAL_15;
  assign rsink__EVAL_69 = _EVAL_4;
  assign _EVAL_78 = rsink__EVAL_81;
  assign fixer__EVAL_23 = _EVAL_97;
  assign buffer__EVAL_37 = fixer__EVAL_8;
  assign fixer__EVAL_52 = buffer__EVAL_66;
  assign fixer__EVAL_65 = rsink__EVAL_70;
  assign rsink__EVAL_91 = _EVAL_102;
  assign fixer__EVAL_20 = rsink__EVAL_79;
  assign _EVAL_56 = rsink__EVAL_46;
  assign rsink__EVAL_26 = _EVAL_98;
  assign _EVAL_1 = rsink__EVAL_103;
  assign rsink__EVAL_3 = _EVAL_31;
  assign rsink__EVAL_31 = _EVAL_2;
  assign fixer__EVAL_12 = buffer__EVAL_29;
  assign buffer__EVAL_23 = fixer__EVAL_45;
  assign buffer__EVAL_44 = fixer__EVAL_35;
  assign _EVAL_87 = rsink__EVAL_92;
  assign rsink__EVAL_88 = _EVAL_5;
  assign buffer__EVAL_5 = _EVAL_71;
  assign rsink__EVAL_19 = _EVAL_64;
  assign _EVAL_48 = rsink__EVAL_61;
  assign fixer__EVAL_3 = buffer__EVAL_25;
  assign rsink__EVAL_44 = _EVAL_99;
  assign buffer__EVAL_65 = _EVAL_55;
  assign fixer__EVAL_44 = rsink__EVAL_106;
  assign rsink__EVAL_48 = _EVAL_84;
  assign _EVAL_51 = buffer__EVAL_60;
  assign _EVAL_86 = buffer__EVAL_1;
  assign fixer__EVAL_28 = buffer__EVAL_56;
  assign _EVAL_3 = rsink__EVAL_73;
  assign fixer__EVAL_47 = rsink__EVAL_1;
  assign _EVAL_93 = rsink__EVAL_68;
  assign fixer__EVAL_7 = rsink__EVAL_50;
  assign fixer__EVAL_19 = rsink__EVAL_89;
  assign rsink__EVAL_53 = _EVAL_70;
  assign _EVAL_79 = buffer__EVAL_11;
  assign rsink__EVAL_12 = _EVAL_62;
  assign buffer__EVAL_24 = fixer__EVAL_54;
  assign _EVAL_17 = rsink__EVAL_67;
  assign fixer__EVAL_59 = buffer__EVAL_12;
  assign rsink__EVAL = _EVAL_82;
  assign _EVAL_77 = rsink__EVAL_42;
  assign buffer__EVAL_27 = _EVAL_107;
  assign _EVAL_96 = rsink__EVAL_41;
  assign buffer__EVAL_0 = fixer__EVAL_33;
  assign rsink__EVAL_22 = _EVAL_45;
  assign buffer__EVAL_34 = fixer__EVAL_69;
  assign rsink__EVAL_20 = _EVAL_75;
  assign fixer__EVAL_53 = buffer__EVAL_14;
  assign _EVAL_72 = rsink__EVAL_5;
  assign rsink__EVAL_47 = _EVAL_15;
  assign rsink__EVAL_33 = _EVAL_8;
  assign fixer__EVAL_25 = buffer__EVAL_36;
  assign _EVAL_59 = buffer__EVAL_67;
  assign rsink__EVAL_30 = _EVAL_40;
  assign rsink__EVAL_17 = _EVAL_36;
  assign rsink__EVAL_38 = fixer__EVAL_42;
  assign rsink__EVAL_78 = _EVAL_34;
  assign rsink__EVAL_29 = fixer__EVAL_60;
  assign _EVAL_58 = rsink__EVAL_77;
  assign buffer__EVAL_20 = fixer__EVAL_38;
  assign _EVAL_61 = rsink__EVAL_40;
  assign rsink__EVAL_87 = _EVAL_68;
  assign buffer__EVAL_61 = fixer__EVAL_9;
  assign buffer__EVAL_8 = _EVAL_26;
  assign rsink__EVAL_57 = _EVAL_30;
  assign rsink__EVAL_98 = fixer__EVAL_0;
  assign buffer__EVAL_46 = fixer__EVAL_49;
  assign _EVAL_60 = rsink__EVAL_18;
  assign rsink__EVAL_102 = _EVAL_92;
  assign fixer__EVAL_1 = buffer__EVAL_45;
  assign rsink__EVAL_11 = _EVAL_44;
  assign _EVAL_91 = rsink__EVAL_84;
  assign fixer__EVAL_11 = rsink__EVAL_32;
  assign _EVAL_7 = rsink__EVAL_51;
  assign _EVAL_73 = rsink__EVAL_39;
  assign rsink__EVAL_100 = fixer__EVAL_16;
  assign buffer__EVAL_70 = fixer__EVAL_13;
  assign _EVAL_52 = rsink__EVAL_6;
  assign rsink__EVAL_74 = _EVAL_104;
  assign _EVAL_103 = buffer__EVAL_21;
  assign _EVAL_43 = buffer__EVAL_4;
  assign buffer__EVAL_26 = fixer__EVAL_56;
  assign _EVAL_28 = rsink__EVAL_15;
  assign rsink__EVAL_62 = fixer__EVAL_36;
  assign _EVAL_67 = buffer__EVAL_41;
  assign _EVAL_11 = buffer__EVAL_64;
  assign rsink__EVAL_28 = _EVAL_53;
  assign buffer__EVAL_18 = fixer__EVAL_66;
  assign rsink__EVAL_25 = _EVAL_24;
  assign _EVAL_49 = buffer__EVAL_43;
  assign fixer__EVAL_70 = rsink__EVAL_8;
  assign fixer__EVAL_58 = buffer__EVAL_9;
  assign rsink__EVAL_54 = _EVAL_14;
  assign _EVAL_88 = rsink__EVAL_45;
  assign rsink__EVAL_66 = _EVAL_97;
  assign fixer__EVAL_63 = buffer__EVAL_22;
  assign rsink__EVAL_64 = _EVAL_69;
  assign buffer__EVAL_6 = fixer__EVAL_67;
  assign _EVAL_27 = rsink__EVAL_101;
  assign _EVAL_94 = rsink__EVAL_99;
  assign rsink__EVAL_2 = fixer__EVAL_2;
  assign _EVAL_66 = rsink__EVAL_16;
  assign _EVAL_80 = rsink__EVAL_14;
  assign fixer__EVAL = rsink__EVAL_95;
  assign buffer__EVAL_62 = _EVAL_97;
  assign fixer__EVAL_10 = rsink__EVAL_13;
  assign _EVAL_50 = rsink__EVAL_65;
  assign fixer__EVAL_32 = rsink__EVAL_83;
  assign buffer__EVAL = _EVAL_25;
  assign buffer__EVAL_51 = _EVAL_9;
  assign buffer__EVAL_33 = fixer__EVAL_57;
  assign buffer__EVAL_17 = fixer__EVAL_4;
  assign rsink__EVAL_72 = _EVAL_41;
  assign _EVAL_85 = buffer__EVAL_2;
  assign buffer__EVAL_57 = _EVAL_83;
  assign rsink__EVAL_35 = _EVAL_46;
  assign fixer__EVAL_30 = rsink__EVAL_49;
  assign rsink__EVAL_55 = fixer__EVAL_64;
  assign fixer__EVAL_26 = buffer__EVAL_7;
  assign rsink__EVAL_82 = fixer__EVAL_68;
  assign buffer__EVAL_68 = fixer__EVAL_41;
  assign fixer__EVAL_48 = rsink__EVAL_9;
  assign fixer__EVAL_61 = rsink__EVAL_107;
  assign _EVAL_39 = buffer__EVAL_32;
  assign rsink__EVAL_97 = _EVAL_105;
  assign _EVAL_89 = buffer__EVAL_13;
  assign fixer__EVAL_43 = rsink__EVAL_0;
  assign fixer__EVAL_31 = buffer__EVAL_3;
  assign _EVAL_16 = rsink__EVAL_60;
  assign rsink__EVAL_24 = _EVAL;
  assign rsink__EVAL_105 = _EVAL_23;
  assign buffer__EVAL_53 = _EVAL_2;
  assign fixer__EVAL_40 = _EVAL_2;
  assign _EVAL_33 = rsink__EVAL_96;
  assign rsink__EVAL_71 = _EVAL_12;
  assign buffer__EVAL_69 = _EVAL_106;
  assign _EVAL_37 = rsink__EVAL_7;
  assign fixer__EVAL_39 = rsink__EVAL_80;
  assign rsink__EVAL_104 = fixer__EVAL_51;
  assign _EVAL_20 = buffer__EVAL_40;
  assign fixer__EVAL_62 = buffer__EVAL_16;
  assign _EVAL_21 = buffer__EVAL_63;
  assign fixer__EVAL_18 = buffer__EVAL_59;
  assign buffer__EVAL_52 = _EVAL_19;
  assign rsink__EVAL_85 = _EVAL_13;
  assign rsink__EVAL_43 = fixer__EVAL_5;
  assign rsink__EVAL_34 = _EVAL_65;
  assign buffer__EVAL_19 = _EVAL_32;
  assign fixer__EVAL_37 = rsink__EVAL_59;
  assign _EVAL_47 = buffer__EVAL_48;
  assign fixer__EVAL_21 = rsink__EVAL_21;
  assign buffer__EVAL_54 = fixer__EVAL_50;
  assign rsink__EVAL_86 = _EVAL_95;
  assign _EVAL_74 = buffer__EVAL_30;
  assign fixer__EVAL_24 = rsink__EVAL_27;
  assign rsink__EVAL_75 = fixer__EVAL_14;
  assign buffer__EVAL_10 = fixer__EVAL_34;
  assign rsink__EVAL_36 = _EVAL_63;
  assign buffer__EVAL_47 = fixer__EVAL_22;
  assign rsink__EVAL_10 = fixer__EVAL_17;
  assign buffer__EVAL_58 = _EVAL_100;
  assign rsink__EVAL_52 = _EVAL_42;
  assign rsink__EVAL_4 = _EVAL_90;
endmodule
