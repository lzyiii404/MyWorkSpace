//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_228_assert(
  input        _EVAL,
  input        _EVAL_0,
  input        _EVAL_2,
  input  [1:0] _EVAL_3,
  input        _EVAL_4,
  input        _EVAL_5,
  input        _EVAL_6,
  input  [1:0] _EVAL_8,
  input        _EVAL_9,
  input        _EVAL_11,
  input        _EVAL_12,
  input        _EVAL_13,
  input        _EVAL_14,
  input        _EVAL_15,
  input        _EVAL_16,
  input  [1:0] _EVAL_17,
  input  [1:0] _EVAL_19,
  input        _EVAL_21,
  input        _EVAL_22,
  input        _EVAL_23,
  input        _EVAL_24,
  input  [1:0] _EVAL_25,
  input        _EVAL_28,
  input        _EVAL_29,
  input        _EVAL_30,
  input        _EVAL_31,
  input        _EVAL_32,
  input        _EVAL_33,
  input        _EVAL_34,
  input  [1:0] _EVAL_35,
  input        _EVAL_36,
  input        _EVAL_40,
  input        _EVAL_41,
  input        _EVAL_44,
  input        _EVAL_46,
  input        _EVAL_48,
  input        _EVAL_50,
  input  [1:0] _EVAL_51,
  input        _EVAL_52,
  input        _EVAL_55,
  input  [1:0] _EVAL_56,
  input        _EVAL_58,
  input        _EVAL_226,
  input        _EVAL_116,
  input        _EVAL_79,
  input        _EVAL_306,
  input        _EVAL_237,
  input        _EVAL_242,
  input        _EVAL_180,
  input        _EVAL_311,
  input        _EVAL_74,
  input        _EVAL_201,
  input        _EVAL_302,
  input        _EVAL_258,
  input        _EVAL_304,
  input        _EVAL_315,
  input        _EVAL_178,
  input        _EVAL_235
);
  wire  _EVAL_273;
  wire  _EVAL_216;
  wire [2:0] _EVAL_210;
  wire  _EVAL_183;
  wire [2:0] _EVAL_194;
  wire  _EVAL_170;
  wire  _EVAL_143;
  wire [2:0] _EVAL_269;
  wire  _EVAL_364;
  wire  _EVAL_291;
  wire  _EVAL_350;
  wire  _EVAL_347;
  wire  _EVAL_144;
  wire  _EVAL_106;
  wire  _EVAL_145;
  wire  _EVAL_208;
  wire  _EVAL_281;
  wire  _EVAL_326;
  wire [2:0] _EVAL_150;
  wire [2:0] _EVAL_345;
  wire  _EVAL_310;
  wire [2:0] _EVAL_199;
  wire  _EVAL_265;
  wire  _EVAL_248;
  wire  _EVAL_268;
  wire  _EVAL_189;
  wire  _EVAL_322;
  wire  _EVAL_197;
  wire  _EVAL_257;
  wire  _EVAL_75;
  wire [2:0] _EVAL_329;
  wire  _EVAL_171;
  wire [2:0] _EVAL_61;
  wire  _EVAL_190;
  wire  _EVAL_275;
  wire  _EVAL_184;
  wire  _EVAL_97;
  wire  _EVAL_279;
  wire  _EVAL_134;
  wire  _EVAL_247;
  wire  _EVAL_287;
  wire  _EVAL_121;
  wire  _EVAL_238;
  wire  _EVAL_73;
  wire  _EVAL_214;
  wire  _EVAL_149;
  wire  _EVAL_80;
  wire  _EVAL_165;
  wire  _EVAL_253;
  wire  _EVAL_330;
  wire  _EVAL_179;
  wire  _EVAL_243;
  wire  _EVAL_325;
  wire  _EVAL_366;
  wire  _EVAL_369;
  wire  _EVAL_92;
  wire  _EVAL_333;
  wire  _EVAL_167;
  wire  _EVAL_154;
  wire  _EVAL_244;
  wire  _EVAL_109;
  wire  _EVAL_147;
  wire  _EVAL_60;
  wire  _EVAL_344;
  wire  _EVAL_103;
  wire  _EVAL_358;
  wire  _EVAL_117;
  wire  _EVAL_71;
  wire  _EVAL_228;
  wire  _EVAL_231;
  wire  _EVAL_108;
  wire  _EVAL_125;
  wire  _EVAL_107;
  wire  _EVAL_251;
  wire  _EVAL_159;
  wire  _EVAL_187;
  wire  _EVAL_260;
  wire  _EVAL_182;
  wire  _EVAL_319;
  wire  _EVAL_206;
  wire  _EVAL_361;
  wire  _EVAL_135;
  wire  _EVAL_163;
  wire  _EVAL_318;
  wire  _EVAL_298;
  wire  _EVAL_324;
  wire  _EVAL_356;
  wire  _EVAL_85;
  wire  _EVAL_296;
  wire  _EVAL_334;
  wire  _EVAL_227;
  wire  _EVAL_286;
  wire  _EVAL_285;
  wire  _EVAL_352;
  wire  _EVAL_207;
  wire  _EVAL_126;
  wire  _EVAL_327;
  wire  _EVAL_301;
  wire  _EVAL_78;
  wire  _EVAL_250;
  wire  _EVAL_130;
  wire  _EVAL_166;
  wire  _EVAL_177;
  wire  _EVAL_86;
  wire  _EVAL_174;
  wire  _EVAL_181;
  wire  _EVAL_198;
  wire  _EVAL_282;
  wire  _EVAL_365;
  wire  _EVAL_100;
  wire  _EVAL_66;
  wire  _EVAL_303;
  wire  _EVAL_94;
  wire  _EVAL_205;
  wire  _EVAL_215;
  wire  _EVAL_68;
  wire  _EVAL_312;
  wire  _EVAL_276;
  wire  _EVAL_164;
  wire  _EVAL_225;
  wire  _EVAL_152;
  wire  _EVAL_317;
  wire  _EVAL_127;
  wire  _EVAL_321;
  wire  _EVAL_104;
  wire  _EVAL_293;
  wire  _EVAL_133;
  wire  _EVAL_241;
  wire  _EVAL_323;
  wire  _EVAL_359;
  wire  _EVAL_234;
  wire  _EVAL_132;
  wire  _EVAL_259;
  wire  _EVAL_82;
  wire  _EVAL_292;
  wire  _EVAL_305;
  wire  _EVAL_151;
  wire  _EVAL_90;
  wire  _EVAL_267;
  wire  _EVAL_363;
  wire  _EVAL_314;
  wire  _EVAL_223;
  wire  _EVAL_270;
  wire  _EVAL_289;
  wire  _EVAL_139;
  wire  _EVAL_161;
  wire  _EVAL_354;
  wire  _EVAL_221;
  wire  _EVAL_113;
  wire  _EVAL_191;
  wire  _EVAL_255;
  wire  _EVAL_101;
  wire  _EVAL_239;
  wire  _EVAL_299;
  wire  _EVAL_362;
  wire  _EVAL_222;
  wire  _EVAL_264;
  wire  _EVAL_200;
  wire  _EVAL_368;
  wire  _EVAL_172;
  wire  _EVAL_186;
  assign _EVAL_273 = _EVAL_17 == 2'h3;
  assign _EVAL_216 = _EVAL_51 == 2'h0;
  assign _EVAL_210 = {_EVAL_30,_EVAL_4,_EVAL_22};
  assign _EVAL_183 = _EVAL_210 == 3'h5;
  assign _EVAL_194 = {_EVAL_52,_EVAL_16,_EVAL_46};
  assign _EVAL_170 = _EVAL_194 == 3'h5;
  assign _EVAL_143 = _EVAL_8 == 2'h0;
  assign _EVAL_269 = {_EVAL_13,_EVAL_23,_EVAL_33};
  assign _EVAL_364 = _EVAL_269 == 3'h3;
  assign _EVAL_291 = _EVAL_51 == 2'h1;
  assign _EVAL_350 = _EVAL_116 == 1'h0;
  assign _EVAL_347 = _EVAL_242 == 1'h0;
  assign _EVAL_144 = _EVAL_347 & _EVAL_237;
  assign _EVAL_106 = _EVAL_25 == 2'h2;
  assign _EVAL_145 = _EVAL_144 & _EVAL_106;
  assign _EVAL_208 = _EVAL_34 & _EVAL_201;
  assign _EVAL_281 = _EVAL_51 == 2'h3;
  assign _EVAL_326 = _EVAL_208 & _EVAL_281;
  assign _EVAL_150 = {_EVAL,_EVAL_28,_EVAL_21};
  assign _EVAL_345 = {_EVAL_6,_EVAL_41,_EVAL_40};
  assign _EVAL_310 = _EVAL_345 == 3'h0;
  assign _EVAL_199 = {_EVAL_2,_EVAL_50,_EVAL_15};
  assign _EVAL_265 = _EVAL_199 == 3'h3;
  assign _EVAL_248 = _EVAL_194 == 3'h7;
  assign _EVAL_268 = _EVAL_24 & _EVAL_180;
  assign _EVAL_189 = _EVAL_19 == 2'h2;
  assign _EVAL_322 = _EVAL_268 & _EVAL_189;
  assign _EVAL_197 = _EVAL_36 & _EVAL_302;
  assign _EVAL_257 = _EVAL_17 == 2'h2;
  assign _EVAL_75 = _EVAL_197 & _EVAL_257;
  assign _EVAL_329 = {_EVAL_44,_EVAL_58,_EVAL_9};
  assign _EVAL_171 = _EVAL_329 == 3'h0;
  assign _EVAL_61 = {_EVAL_14,_EVAL_0,_EVAL_12};
  assign _EVAL_190 = _EVAL_61 == 3'h1;
  assign _EVAL_275 = _EVAL_150 == 3'h1;
  assign _EVAL_184 = _EVAL_350 & _EVAL_180;
  assign _EVAL_97 = _EVAL_19 == 2'h3;
  assign _EVAL_279 = _EVAL_184 & _EVAL_97;
  assign _EVAL_134 = _EVAL_35 == 2'h0;
  assign _EVAL_247 = _EVAL_226 == 1'h0;
  assign _EVAL_287 = _EVAL_32 & _EVAL_258;
  assign _EVAL_121 = _EVAL_35 == 2'h2;
  assign _EVAL_238 = _EVAL_287 & _EVAL_121;
  assign _EVAL_73 = _EVAL_29 & _EVAL_311;
  assign _EVAL_214 = _EVAL_8 == 2'h1;
  assign _EVAL_149 = _EVAL_73 & _EVAL_214;
  assign _EVAL_80 = _EVAL_304 == 1'h0;
  assign _EVAL_165 = _EVAL_80 & _EVAL_302;
  assign _EVAL_253 = _EVAL_269 == 3'h0;
  assign _EVAL_330 = _EVAL_210 == 3'h1;
  assign _EVAL_179 = _EVAL_5 & _EVAL_79;
  assign _EVAL_243 = _EVAL_3 == 2'h2;
  assign _EVAL_325 = _EVAL_179 & _EVAL_243;
  assign _EVAL_366 = _EVAL_194 == 3'h1;
  assign _EVAL_369 = _EVAL_74 == 1'h0;
  assign _EVAL_92 = _EVAL_369 & _EVAL_311;
  assign _EVAL_333 = _EVAL_329 == 3'h3;
  assign _EVAL_167 = _EVAL_25 == 2'h3;
  assign _EVAL_154 = _EVAL_144 & _EVAL_167;
  assign _EVAL_244 = _EVAL_210 == 3'h3;
  assign _EVAL_109 = _EVAL_61 == 3'h7;
  assign _EVAL_147 = _EVAL_35 == 2'h3;
  assign _EVAL_60 = _EVAL_287 & _EVAL_147;
  assign _EVAL_344 = _EVAL_165 & _EVAL_257;
  assign _EVAL_103 = _EVAL_150 == 3'h4;
  assign _EVAL_358 = _EVAL_3 == 2'h1;
  assign _EVAL_117 = _EVAL_179 & _EVAL_358;
  assign _EVAL_71 = _EVAL_315 == 1'h0;
  assign _EVAL_228 = _EVAL_11 == 1'h0;
  assign _EVAL_231 = _EVAL_329 == 3'h7;
  assign _EVAL_108 = _EVAL_19 == 2'h1;
  assign _EVAL_125 = _EVAL_184 & _EVAL_108;
  assign _EVAL_107 = _EVAL_48 & _EVAL_237;
  assign _EVAL_251 = _EVAL_150 == 3'h3;
  assign _EVAL_159 = _EVAL_150 == 3'h5;
  assign _EVAL_187 = _EVAL_3 == 2'h3;
  assign _EVAL_260 = _EVAL_179 & _EVAL_187;
  assign _EVAL_182 = _EVAL_269 == 3'h1;
  assign _EVAL_319 = _EVAL_25 == 2'h1;
  assign _EVAL_206 = _EVAL_306 == 1'h0;
  assign _EVAL_361 = _EVAL_206 & _EVAL_79;
  assign _EVAL_135 = _EVAL_361 & _EVAL_358;
  assign _EVAL_163 = _EVAL_31 & _EVAL_178;
  assign _EVAL_318 = _EVAL_56 == 2'h2;
  assign _EVAL_298 = _EVAL_163 & _EVAL_318;
  assign _EVAL_324 = _EVAL_268 & _EVAL_108;
  assign _EVAL_356 = _EVAL_61 == 3'h4;
  assign _EVAL_85 = _EVAL_345 == 3'h4;
  assign _EVAL_296 = _EVAL_199 == 3'h4;
  assign _EVAL_334 = _EVAL_71 & _EVAL_201;
  assign _EVAL_227 = _EVAL_17 == 2'h0;
  assign _EVAL_286 = _EVAL_8 == 2'h2;
  assign _EVAL_285 = _EVAL_73 & _EVAL_286;
  assign _EVAL_352 = _EVAL_361 & _EVAL_187;
  assign _EVAL_207 = _EVAL_199 == 3'h7;
  assign _EVAL_126 = _EVAL_345 == 3'h5;
  assign _EVAL_327 = _EVAL_51 == 2'h2;
  assign _EVAL_301 = _EVAL_334 & _EVAL_327;
  assign _EVAL_78 = _EVAL_56 == 2'h1;
  assign _EVAL_250 = _EVAL_163 & _EVAL_78;
  assign _EVAL_130 = _EVAL_61 == 3'h5;
  assign _EVAL_166 = _EVAL_19 == 2'h0;
  assign _EVAL_177 = _EVAL_17 == 2'h1;
  assign _EVAL_86 = _EVAL_165 & _EVAL_177;
  assign _EVAL_174 = _EVAL_165 & _EVAL_273;
  assign _EVAL_181 = _EVAL_194 == 3'h0;
  assign _EVAL_198 = _EVAL_150 == 3'h7;
  assign _EVAL_282 = _EVAL_3 == 2'h0;
  assign _EVAL_365 = _EVAL_107 & _EVAL_319;
  assign _EVAL_100 = _EVAL_247 & _EVAL_258;
  assign _EVAL_66 = _EVAL_100 & _EVAL_121;
  assign _EVAL_303 = _EVAL_56 == 2'h3;
  assign _EVAL_94 = _EVAL_163 & _EVAL_303;
  assign _EVAL_205 = _EVAL_345 == 3'h1;
  assign _EVAL_215 = _EVAL_199 == 3'h0;
  assign _EVAL_68 = _EVAL_329 == 3'h4;
  assign _EVAL_312 = _EVAL_269 == 3'h7;
  assign _EVAL_276 = _EVAL_8 == 2'h3;
  assign _EVAL_164 = _EVAL_73 & _EVAL_276;
  assign _EVAL_225 = _EVAL_194 == 3'h3;
  assign _EVAL_152 = _EVAL_361 & _EVAL_243;
  assign _EVAL_317 = _EVAL_199 == 3'h5;
  assign _EVAL_127 = _EVAL_107 & _EVAL_106;
  assign _EVAL_321 = _EVAL_184 & _EVAL_189;
  assign _EVAL_104 = _EVAL_269 == 3'h4;
  assign _EVAL_293 = _EVAL_235 == 1'h0;
  assign _EVAL_133 = _EVAL_293 & _EVAL_178;
  assign _EVAL_241 = _EVAL_133 & _EVAL_318;
  assign _EVAL_323 = _EVAL_208 & _EVAL_327;
  assign _EVAL_359 = _EVAL_269 == 3'h5;
  assign _EVAL_234 = _EVAL_107 & _EVAL_167;
  assign _EVAL_132 = _EVAL_345 == 3'h3;
  assign _EVAL_259 = _EVAL_329 == 3'h5;
  assign _EVAL_82 = _EVAL_35 == 2'h1;
  assign _EVAL_292 = _EVAL_287 & _EVAL_82;
  assign _EVAL_305 = _EVAL_194 == 3'h4;
  assign _EVAL_151 = _EVAL_61 == 3'h3;
  assign _EVAL_90 = _EVAL_133 & _EVAL_303;
  assign _EVAL_267 = _EVAL_100 & _EVAL_82;
  assign _EVAL_363 = _EVAL_210 == 3'h4;
  assign _EVAL_314 = _EVAL_210 == 3'h0;
  assign _EVAL_223 = _EVAL_100 & _EVAL_147;
  assign _EVAL_270 = _EVAL_210 == 3'h7;
  assign _EVAL_289 = _EVAL_144 & _EVAL_319;
  assign _EVAL_139 = _EVAL_345 == 3'h7;
  assign _EVAL_161 = _EVAL_92 & _EVAL_276;
  assign _EVAL_354 = _EVAL_197 & _EVAL_273;
  assign _EVAL_221 = _EVAL_150 == 3'h0;
  assign _EVAL_113 = _EVAL_25 == 2'h0;
  assign _EVAL_191 = _EVAL_133 & _EVAL_78;
  assign _EVAL_255 = _EVAL_197 & _EVAL_177;
  assign _EVAL_101 = _EVAL_334 & _EVAL_291;
  assign _EVAL_239 = _EVAL_56 == 2'h0;
  assign _EVAL_299 = _EVAL_61 == 3'h0;
  assign _EVAL_362 = _EVAL_268 & _EVAL_97;
  assign _EVAL_222 = _EVAL_92 & _EVAL_286;
  assign _EVAL_264 = _EVAL_208 & _EVAL_291;
  assign _EVAL_200 = _EVAL_92 & _EVAL_214;
  assign _EVAL_368 = _EVAL_334 & _EVAL_281;
  assign _EVAL_172 = _EVAL_329 == 3'h1;
  assign _EVAL_186 = _EVAL_199 == 3'h1;
  always @(posedge _EVAL_55) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_327 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_363 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_362 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_354 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_358 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_366 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c803a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fa4a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d26248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635f8930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc2e5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c99191e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee41222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f742f169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab54cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b17f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fbd216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f86a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9f15ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23590644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ccaeac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7dd1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b5b278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
