//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_149(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  output [2:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [31:0] _EVAL_8,
  output [1:0]  _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  output [6:0]  _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  output [2:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [3:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  output [31:0] _EVAL_22,
  input  [6:0]  _EVAL_23,
  output [3:0]  _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output [2:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  input  [24:0] _EVAL_30,
  output        _EVAL_31,
  output [31:0] _EVAL_32,
  output        _EVAL_33,
  output [2:0]  _EVAL_34,
  output [24:0] _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input  [6:0]  _EVAL_38,
  output [6:0]  _EVAL_39,
  input  [2:0]  _EVAL_40
);
  assign _EVAL_15 = _EVAL_7;
  assign _EVAL_13 = _EVAL_23;
  assign _EVAL_28 = _EVAL_17;
  assign _EVAL_22 = _EVAL_8;
  assign _EVAL_14 = _EVAL_19;
  assign _EVAL_9 = _EVAL_12;
  assign _EVAL_31 = _EVAL_11;
  assign _EVAL_16 = _EVAL_40;
  assign _EVAL_32 = _EVAL_2;
  assign _EVAL_34 = _EVAL_0;
  assign _EVAL_10 = _EVAL_36;
  assign _EVAL_39 = _EVAL_38;
  assign _EVAL_35 = _EVAL_30;
  assign _EVAL_21 = _EVAL;
  assign _EVAL_24 = _EVAL_20;
  assign _EVAL_33 = _EVAL_6;
  assign _EVAL_4 = _EVAL_37;
  assign _EVAL_18 = _EVAL_5;
  assign _EVAL_1 = _EVAL_29;
  assign _EVAL_25 = _EVAL_26;
endmodule
