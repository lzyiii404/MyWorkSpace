//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_242(
  input  [31:0] _EVAL,
  output [31:0] _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  input  [2:0]  _EVAL_4
);
  wire  _EVAL_63;
  wire  _EVAL_165;
  wire [7:0] _EVAL_27;
  wire  _EVAL_61;
  wire [7:0] _EVAL_180;
  wire  _EVAL_13;
  wire [7:0] _EVAL_191;
  wire  _EVAL_93;
  wire [7:0] _EVAL_188;
  wire [31:0] _EVAL_154;
  wire  _EVAL_160;
  wire  _EVAL_110;
  wire [31:0] _EVAL_117;
  wire  _EVAL_236;
  wire [31:0] _EVAL_113;
  wire [31:0] _EVAL_12;
  wire [31:0] _EVAL_143;
  wire  _EVAL_16;
  wire  _EVAL_121;
  wire  _EVAL_67;
  wire  _EVAL_91;
  wire [3:0] _EVAL_183;
  wire [3:0] _EVAL_207;
  wire [2:0] _EVAL_223;
  wire [3:0] _EVAL_136;
  wire [3:0] _EVAL_187;
  wire [3:0] _EVAL_68;
  wire  _EVAL_130;
  wire  _EVAL_82;
  wire  _EVAL_150;
  wire  _EVAL_41;
  wire  _EVAL_163;
  wire  _EVAL_211;
  wire  _EVAL_166;
  wire  _EVAL_20;
  wire [3:0] _EVAL_172;
  wire [3:0] _EVAL_89;
  wire  _EVAL_218;
  wire  _EVAL_48;
  wire  _EVAL_35;
  wire  _EVAL_122;
  wire  _EVAL_153;
  wire [3:0] _EVAL_240;
  wire [3:0] _EVAL_44;
  wire  _EVAL_114;
  wire  _EVAL_14;
  wire  _EVAL_251;
  wire  _EVAL_129;
  wire  _EVAL_108;
  wire  _EVAL_175;
  wire [1:0] _EVAL_11;
  wire [1:0] _EVAL_39;
  wire [1:0] _EVAL_246;
  wire [1:0] _EVAL_126;
  wire [1:0] _EVAL_25;
  wire [1:0] _EVAL_142;
  wire [1:0] _EVAL_71;
  wire [1:0] _EVAL_45;
  wire [1:0] _EVAL_205;
  wire [3:0] _EVAL_145;
  wire [3:0] _EVAL_99;
  wire [3:0] _EVAL_158;
  wire [1:0] _EVAL_94;
  wire [3:0] _EVAL_148;
  wire  _EVAL_169;
  wire  _EVAL_203;
  wire  _EVAL_86;
  wire [1:0] _EVAL_111;
  wire [3:0] _EVAL_100;
  wire  _EVAL_212;
  wire  _EVAL_190;
  wire  _EVAL_62;
  wire [1:0] _EVAL_103;
  wire [3:0] _EVAL_214;
  wire  _EVAL_92;
  wire  _EVAL_40;
  wire  _EVAL_156;
  wire [1:0] _EVAL_244;
  wire [3:0] _EVAL_6;
  wire  _EVAL_138;
  wire  _EVAL_210;
  wire  _EVAL_49;
  wire [1:0] _EVAL_184;
  wire [3:0] _EVAL_189;
  wire  _EVAL_245;
  wire  _EVAL_197;
  wire  _EVAL_196;
  wire [1:0] _EVAL_28;
  wire [3:0] _EVAL_144;
  wire  _EVAL_42;
  wire  _EVAL_120;
  wire  _EVAL_33;
  wire [1:0] _EVAL_241;
  wire [3:0] _EVAL_185;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [1:0] _EVAL_164;
  wire [3:0] _EVAL_123;
  wire  _EVAL_112;
  wire [1:0] _EVAL_159;
  wire [3:0] _EVAL_75;
  wire  _EVAL_73;
  wire  _EVAL_235;
  wire  _EVAL_98;
  wire [1:0] _EVAL_227;
  wire [3:0] _EVAL_10;
  wire  _EVAL_30;
  wire  _EVAL_238;
  wire [1:0] _EVAL_155;
  wire [3:0] _EVAL_118;
  wire  _EVAL_194;
  wire  _EVAL_19;
  wire  _EVAL_96;
  wire [1:0] _EVAL_161;
  wire [3:0] _EVAL_87;
  wire  _EVAL_135;
  wire  _EVAL_200;
  wire  _EVAL_152;
  wire [1:0] _EVAL_219;
  wire [3:0] _EVAL_9;
  wire  _EVAL_146;
  wire  _EVAL_5;
  wire  _EVAL_206;
  wire [1:0] _EVAL_127;
  wire [3:0] _EVAL_173;
  wire  _EVAL_115;
  wire  _EVAL_182;
  wire  _EVAL_76;
  wire [1:0] _EVAL_125;
  wire [3:0] _EVAL_243;
  wire  _EVAL_131;
  wire  _EVAL_224;
  wire  _EVAL_69;
  wire [1:0] _EVAL_78;
  wire [3:0] _EVAL_34;
  wire  _EVAL_102;
  wire [7:0] _EVAL_178;
  wire [1:0] _EVAL_85;
  wire [3:0] _EVAL_177;
  wire  _EVAL_97;
  wire  _EVAL_167;
  wire  _EVAL_176;
  wire [1:0] _EVAL_107;
  wire [3:0] _EVAL_134;
  wire  _EVAL_81;
  wire  _EVAL_221;
  wire  _EVAL_60;
  wire [1:0] _EVAL_213;
  wire [3:0] _EVAL_128;
  wire  _EVAL_36;
  wire  _EVAL_8;
  wire  _EVAL_208;
  wire [1:0] _EVAL_109;
  wire [3:0] _EVAL_51;
  wire  _EVAL_174;
  wire  _EVAL_225;
  wire  _EVAL_17;
  wire [1:0] _EVAL_52;
  wire [3:0] _EVAL_79;
  wire  _EVAL_192;
  wire  _EVAL_56;
  wire [1:0] _EVAL_132;
  wire [3:0] _EVAL_18;
  wire  _EVAL_70;
  wire  _EVAL_202;
  wire  _EVAL_74;
  wire [1:0] _EVAL_77;
  wire [3:0] _EVAL_104;
  wire  _EVAL_222;
  wire  _EVAL_116;
  wire  _EVAL_43;
  wire [1:0] _EVAL_124;
  wire [3:0] _EVAL_83;
  wire  _EVAL_168;
  wire [1:0] _EVAL_84;
  wire [3:0] _EVAL_204;
  wire  _EVAL_38;
  wire  _EVAL_226;
  wire  _EVAL_209;
  wire [1:0] _EVAL_24;
  wire [3:0] _EVAL_101;
  wire  _EVAL_157;
  wire  _EVAL_21;
  wire  _EVAL_54;
  wire [1:0] _EVAL_239;
  wire [3:0] _EVAL_105;
  wire  _EVAL_15;
  wire  _EVAL_147;
  wire [1:0] _EVAL_72;
  wire [3:0] _EVAL_90;
  wire  _EVAL_64;
  wire  _EVAL_22;
  wire  _EVAL_133;
  wire [1:0] _EVAL_228;
  wire [3:0] _EVAL_181;
  wire  _EVAL_139;
  wire  _EVAL_179;
  wire  _EVAL_26;
  wire [1:0] _EVAL_249;
  wire [3:0] _EVAL_247;
  wire  _EVAL_233;
  wire  _EVAL_198;
  wire  _EVAL_193;
  wire [1:0] _EVAL_231;
  wire [3:0] _EVAL_32;
  wire  _EVAL_50;
  wire  _EVAL_106;
  wire  _EVAL_162;
  wire [1:0] _EVAL_237;
  wire [3:0] _EVAL_250;
  wire  _EVAL_220;
  wire [7:0] _EVAL_201;
  wire [15:0] _EVAL_31;
  wire [31:0] _EVAL_171;
  wire [7:0] _EVAL_186;
  wire [7:0] _EVAL_248;
  wire [7:0] _EVAL_66;
  wire [7:0] _EVAL_119;
  wire [7:0] _EVAL_58;
  wire [7:0] _EVAL_151;
  wire [7:0] _EVAL_137;
  wire [1:0] _EVAL_46;
  wire [7:0] _EVAL_170;
  wire [7:0] _EVAL_229;
  wire [7:0] _EVAL_217;
  wire [7:0] _EVAL_80;
  wire [7:0] _EVAL_234;
  wire [1:0] _EVAL_59;
  wire [7:0] _EVAL_65;
  wire [7:0] _EVAL_216;
  wire [7:0] _EVAL_149;
  wire [7:0] _EVAL_242;
  wire [7:0] _EVAL_215;
  wire [7:0] _EVAL_7;
  wire [7:0] _EVAL_95;
  wire [7:0] _EVAL_29;
  wire [7:0] _EVAL_88;
  wire [7:0] _EVAL_199;
  wire [15:0] _EVAL_37;
  wire [7:0] _EVAL_195;
  wire [1:0] _EVAL_230;
  wire [7:0] _EVAL_55;
  wire [7:0] _EVAL_57;
  wire [7:0] _EVAL_23;
  wire [7:0] _EVAL_232;
  wire [7:0] _EVAL_47;
  wire [15:0] _EVAL_252;
  assign _EVAL_63 = _EVAL_3[24];
  assign _EVAL_165 = _EVAL_1[3];
  assign _EVAL_27 = _EVAL_165 ? 8'hff : 8'h0;
  assign _EVAL_61 = _EVAL_1[2];
  assign _EVAL_180 = _EVAL_61 ? 8'hff : 8'h0;
  assign _EVAL_13 = _EVAL_1[1];
  assign _EVAL_191 = _EVAL_13 ? 8'hff : 8'h0;
  assign _EVAL_93 = _EVAL_1[0];
  assign _EVAL_188 = _EVAL_93 ? 8'hff : 8'h0;
  assign _EVAL_154 = {_EVAL_27,_EVAL_180,_EVAL_191,_EVAL_188};
  assign _EVAL_160 = _EVAL_3[10];
  assign _EVAL_110 = _EVAL_3[4];
  assign _EVAL_117 = _EVAL_154 & _EVAL_3;
  assign _EVAL_236 = _EVAL_2[2];
  assign _EVAL_113 = ~ _EVAL;
  assign _EVAL_12 = _EVAL_236 ? _EVAL : _EVAL_113;
  assign _EVAL_143 = _EVAL_117 + _EVAL_12;
  assign _EVAL_16 = _EVAL_143[31];
  assign _EVAL_121 = _EVAL_143[23];
  assign _EVAL_67 = _EVAL_143[15];
  assign _EVAL_91 = _EVAL_143[7];
  assign _EVAL_183 = {_EVAL_16,_EVAL_121,_EVAL_67,_EVAL_91};
  assign _EVAL_207 = ~ _EVAL_1;
  assign _EVAL_223 = _EVAL_207[3:1];
  assign _EVAL_136 = {1'h1,_EVAL_223};
  assign _EVAL_187 = _EVAL_1 & _EVAL_136;
  assign _EVAL_68 = _EVAL_183 & _EVAL_187;
  assign _EVAL_130 = _EVAL_68 != 4'h0;
  assign _EVAL_82 = _EVAL_130 == 1'h0;
  assign _EVAL_150 = _EVAL_3[21];
  assign _EVAL_41 = _EVAL_2[0];
  assign _EVAL_163 = _EVAL_3[31];
  assign _EVAL_211 = _EVAL_3[23];
  assign _EVAL_166 = _EVAL_3[15];
  assign _EVAL_20 = _EVAL_3[7];
  assign _EVAL_172 = {_EVAL_163,_EVAL_211,_EVAL_166,_EVAL_20};
  assign _EVAL_89 = _EVAL_172 & _EVAL_187;
  assign _EVAL_218 = _EVAL_89 != 4'h0;
  assign _EVAL_48 = _EVAL[31];
  assign _EVAL_35 = _EVAL[23];
  assign _EVAL_122 = _EVAL[15];
  assign _EVAL_153 = _EVAL[7];
  assign _EVAL_240 = {_EVAL_48,_EVAL_35,_EVAL_122,_EVAL_153};
  assign _EVAL_44 = _EVAL_240 & _EVAL_187;
  assign _EVAL_114 = _EVAL_44 != 4'h0;
  assign _EVAL_14 = _EVAL_218 == _EVAL_114;
  assign _EVAL_251 = _EVAL_2[1];
  assign _EVAL_129 = _EVAL_251 == _EVAL_218;
  assign _EVAL_108 = _EVAL_14 ? _EVAL_82 : _EVAL_129;
  assign _EVAL_175 = _EVAL_41 == _EVAL_108;
  assign _EVAL_11 = _EVAL_236 ? 2'h2 : {{1'd0}, _EVAL_175};
  assign _EVAL_39 = 3'h2 == _EVAL_4 ? _EVAL_11 : 2'h1;
  assign _EVAL_246 = 3'h3 == _EVAL_4 ? 2'h3 : _EVAL_39;
  assign _EVAL_126 = 3'h4 == _EVAL_4 ? 2'h0 : _EVAL_246;
  assign _EVAL_25 = 3'h5 == _EVAL_4 ? 2'h0 : _EVAL_126;
  assign _EVAL_142 = 3'h6 == _EVAL_4 ? 2'h0 : _EVAL_25;
  assign _EVAL_71 = 3'h7 == _EVAL_4 ? 2'h0 : _EVAL_142;
  assign _EVAL_45 = _EVAL_61 ? _EVAL_71 : 2'h0;
  assign _EVAL_205 = _EVAL_2[1:0];
  assign _EVAL_145 = 2'h1 == _EVAL_205 ? 4'he : 4'h6;
  assign _EVAL_99 = 2'h2 == _EVAL_205 ? 4'h8 : _EVAL_145;
  assign _EVAL_158 = 2'h3 == _EVAL_205 ? 4'hc : _EVAL_99;
  assign _EVAL_94 = {_EVAL_163,_EVAL_48};
  assign _EVAL_148 = _EVAL_158 >> _EVAL_94;
  assign _EVAL_169 = _EVAL_148[0];
  assign _EVAL_203 = _EVAL_3[30];
  assign _EVAL_86 = _EVAL[30];
  assign _EVAL_111 = {_EVAL_203,_EVAL_86};
  assign _EVAL_100 = _EVAL_158 >> _EVAL_111;
  assign _EVAL_212 = _EVAL_100[0];
  assign _EVAL_190 = _EVAL_3[29];
  assign _EVAL_62 = _EVAL[29];
  assign _EVAL_103 = {_EVAL_190,_EVAL_62};
  assign _EVAL_214 = _EVAL_158 >> _EVAL_103;
  assign _EVAL_92 = _EVAL_214[0];
  assign _EVAL_40 = _EVAL_3[28];
  assign _EVAL_156 = _EVAL[28];
  assign _EVAL_244 = {_EVAL_40,_EVAL_156};
  assign _EVAL_6 = _EVAL_158 >> _EVAL_244;
  assign _EVAL_138 = _EVAL_6[0];
  assign _EVAL_210 = _EVAL_3[27];
  assign _EVAL_49 = _EVAL[27];
  assign _EVAL_184 = {_EVAL_210,_EVAL_49};
  assign _EVAL_189 = _EVAL_158 >> _EVAL_184;
  assign _EVAL_245 = _EVAL_189[0];
  assign _EVAL_197 = _EVAL_3[26];
  assign _EVAL_196 = _EVAL[26];
  assign _EVAL_28 = {_EVAL_197,_EVAL_196};
  assign _EVAL_144 = _EVAL_158 >> _EVAL_28;
  assign _EVAL_42 = _EVAL_144[0];
  assign _EVAL_120 = _EVAL_3[25];
  assign _EVAL_33 = _EVAL[25];
  assign _EVAL_241 = {_EVAL_120,_EVAL_33};
  assign _EVAL_185 = _EVAL_158 >> _EVAL_241;
  assign _EVAL_140 = _EVAL_185[0];
  assign _EVAL_141 = _EVAL[24];
  assign _EVAL_164 = {_EVAL_63,_EVAL_141};
  assign _EVAL_123 = _EVAL_158 >> _EVAL_164;
  assign _EVAL_112 = _EVAL_123[0];
  assign _EVAL_159 = {_EVAL_211,_EVAL_35};
  assign _EVAL_75 = _EVAL_158 >> _EVAL_159;
  assign _EVAL_73 = _EVAL_75[0];
  assign _EVAL_235 = _EVAL_3[22];
  assign _EVAL_98 = _EVAL[22];
  assign _EVAL_227 = {_EVAL_235,_EVAL_98};
  assign _EVAL_10 = _EVAL_158 >> _EVAL_227;
  assign _EVAL_30 = _EVAL_10[0];
  assign _EVAL_238 = _EVAL[21];
  assign _EVAL_155 = {_EVAL_150,_EVAL_238};
  assign _EVAL_118 = _EVAL_158 >> _EVAL_155;
  assign _EVAL_194 = _EVAL_118[0];
  assign _EVAL_19 = _EVAL_3[20];
  assign _EVAL_96 = _EVAL[20];
  assign _EVAL_161 = {_EVAL_19,_EVAL_96};
  assign _EVAL_87 = _EVAL_158 >> _EVAL_161;
  assign _EVAL_135 = _EVAL_87[0];
  assign _EVAL_200 = _EVAL_3[19];
  assign _EVAL_152 = _EVAL[19];
  assign _EVAL_219 = {_EVAL_200,_EVAL_152};
  assign _EVAL_9 = _EVAL_158 >> _EVAL_219;
  assign _EVAL_146 = _EVAL_9[0];
  assign _EVAL_5 = _EVAL_3[18];
  assign _EVAL_206 = _EVAL[18];
  assign _EVAL_127 = {_EVAL_5,_EVAL_206};
  assign _EVAL_173 = _EVAL_158 >> _EVAL_127;
  assign _EVAL_115 = _EVAL_173[0];
  assign _EVAL_182 = _EVAL_3[17];
  assign _EVAL_76 = _EVAL[17];
  assign _EVAL_125 = {_EVAL_182,_EVAL_76};
  assign _EVAL_243 = _EVAL_158 >> _EVAL_125;
  assign _EVAL_131 = _EVAL_243[0];
  assign _EVAL_224 = _EVAL_3[16];
  assign _EVAL_69 = _EVAL[16];
  assign _EVAL_78 = {_EVAL_224,_EVAL_69};
  assign _EVAL_34 = _EVAL_158 >> _EVAL_78;
  assign _EVAL_102 = _EVAL_34[0];
  assign _EVAL_178 = {_EVAL_73,_EVAL_30,_EVAL_194,_EVAL_135,_EVAL_146,_EVAL_115,_EVAL_131,_EVAL_102};
  assign _EVAL_85 = {_EVAL_166,_EVAL_122};
  assign _EVAL_177 = _EVAL_158 >> _EVAL_85;
  assign _EVAL_97 = _EVAL_177[0];
  assign _EVAL_167 = _EVAL_3[14];
  assign _EVAL_176 = _EVAL[14];
  assign _EVAL_107 = {_EVAL_167,_EVAL_176};
  assign _EVAL_134 = _EVAL_158 >> _EVAL_107;
  assign _EVAL_81 = _EVAL_134[0];
  assign _EVAL_221 = _EVAL_3[13];
  assign _EVAL_60 = _EVAL[13];
  assign _EVAL_213 = {_EVAL_221,_EVAL_60};
  assign _EVAL_128 = _EVAL_158 >> _EVAL_213;
  assign _EVAL_36 = _EVAL_128[0];
  assign _EVAL_8 = _EVAL_3[12];
  assign _EVAL_208 = _EVAL[12];
  assign _EVAL_109 = {_EVAL_8,_EVAL_208};
  assign _EVAL_51 = _EVAL_158 >> _EVAL_109;
  assign _EVAL_174 = _EVAL_51[0];
  assign _EVAL_225 = _EVAL_3[11];
  assign _EVAL_17 = _EVAL[11];
  assign _EVAL_52 = {_EVAL_225,_EVAL_17};
  assign _EVAL_79 = _EVAL_158 >> _EVAL_52;
  assign _EVAL_192 = _EVAL_79[0];
  assign _EVAL_56 = _EVAL[10];
  assign _EVAL_132 = {_EVAL_160,_EVAL_56};
  assign _EVAL_18 = _EVAL_158 >> _EVAL_132;
  assign _EVAL_70 = _EVAL_18[0];
  assign _EVAL_202 = _EVAL_3[9];
  assign _EVAL_74 = _EVAL[9];
  assign _EVAL_77 = {_EVAL_202,_EVAL_74};
  assign _EVAL_104 = _EVAL_158 >> _EVAL_77;
  assign _EVAL_222 = _EVAL_104[0];
  assign _EVAL_116 = _EVAL_3[8];
  assign _EVAL_43 = _EVAL[8];
  assign _EVAL_124 = {_EVAL_116,_EVAL_43};
  assign _EVAL_83 = _EVAL_158 >> _EVAL_124;
  assign _EVAL_168 = _EVAL_83[0];
  assign _EVAL_84 = {_EVAL_20,_EVAL_153};
  assign _EVAL_204 = _EVAL_158 >> _EVAL_84;
  assign _EVAL_38 = _EVAL_204[0];
  assign _EVAL_226 = _EVAL_3[6];
  assign _EVAL_209 = _EVAL[6];
  assign _EVAL_24 = {_EVAL_226,_EVAL_209};
  assign _EVAL_101 = _EVAL_158 >> _EVAL_24;
  assign _EVAL_157 = _EVAL_101[0];
  assign _EVAL_21 = _EVAL_3[5];
  assign _EVAL_54 = _EVAL[5];
  assign _EVAL_239 = {_EVAL_21,_EVAL_54};
  assign _EVAL_105 = _EVAL_158 >> _EVAL_239;
  assign _EVAL_15 = _EVAL_105[0];
  assign _EVAL_147 = _EVAL[4];
  assign _EVAL_72 = {_EVAL_110,_EVAL_147};
  assign _EVAL_90 = _EVAL_158 >> _EVAL_72;
  assign _EVAL_64 = _EVAL_90[0];
  assign _EVAL_22 = _EVAL_3[3];
  assign _EVAL_133 = _EVAL[3];
  assign _EVAL_228 = {_EVAL_22,_EVAL_133};
  assign _EVAL_181 = _EVAL_158 >> _EVAL_228;
  assign _EVAL_139 = _EVAL_181[0];
  assign _EVAL_179 = _EVAL_3[2];
  assign _EVAL_26 = _EVAL[2];
  assign _EVAL_249 = {_EVAL_179,_EVAL_26};
  assign _EVAL_247 = _EVAL_158 >> _EVAL_249;
  assign _EVAL_233 = _EVAL_247[0];
  assign _EVAL_198 = _EVAL_3[1];
  assign _EVAL_193 = _EVAL[1];
  assign _EVAL_231 = {_EVAL_198,_EVAL_193};
  assign _EVAL_32 = _EVAL_158 >> _EVAL_231;
  assign _EVAL_50 = _EVAL_32[0];
  assign _EVAL_106 = _EVAL_3[0];
  assign _EVAL_162 = _EVAL[0];
  assign _EVAL_237 = {_EVAL_106,_EVAL_162};
  assign _EVAL_250 = _EVAL_158 >> _EVAL_237;
  assign _EVAL_220 = _EVAL_250[0];
  assign _EVAL_201 = {_EVAL_38,_EVAL_157,_EVAL_15,_EVAL_64,_EVAL_139,_EVAL_233,_EVAL_50,_EVAL_220};
  assign _EVAL_31 = {_EVAL_97,_EVAL_81,_EVAL_36,_EVAL_174,_EVAL_192,_EVAL_70,_EVAL_222,_EVAL_168,_EVAL_201};
  assign _EVAL_171 = {_EVAL_169,_EVAL_212,_EVAL_92,_EVAL_138,_EVAL_245,_EVAL_42,_EVAL_140,_EVAL_112,_EVAL_178,_EVAL_31};
  assign _EVAL_186 = _EVAL_171[23:16];
  assign _EVAL_248 = _EVAL_143[23:16];
  assign _EVAL_66 = _EVAL_3[23:16];
  assign _EVAL_119 = _EVAL[23:16];
  assign _EVAL_58 = 2'h1 == _EVAL_45 ? _EVAL_66 : _EVAL_119;
  assign _EVAL_151 = 2'h2 == _EVAL_45 ? _EVAL_248 : _EVAL_58;
  assign _EVAL_137 = 2'h3 == _EVAL_45 ? _EVAL_186 : _EVAL_151;
  assign _EVAL_46 = _EVAL_93 ? _EVAL_71 : 2'h0;
  assign _EVAL_170 = _EVAL_3[7:0];
  assign _EVAL_229 = _EVAL[7:0];
  assign _EVAL_217 = 2'h1 == _EVAL_46 ? _EVAL_170 : _EVAL_229;
  assign _EVAL_80 = _EVAL_143[7:0];
  assign _EVAL_234 = _EVAL_3[31:24];
  assign _EVAL_59 = _EVAL_13 ? _EVAL_71 : 2'h0;
  assign _EVAL_65 = _EVAL_171[15:8];
  assign _EVAL_216 = _EVAL_143[15:8];
  assign _EVAL_149 = _EVAL_3[15:8];
  assign _EVAL_242 = _EVAL[15:8];
  assign _EVAL_215 = 2'h1 == _EVAL_59 ? _EVAL_149 : _EVAL_242;
  assign _EVAL_7 = 2'h2 == _EVAL_59 ? _EVAL_216 : _EVAL_215;
  assign _EVAL_95 = 2'h3 == _EVAL_59 ? _EVAL_65 : _EVAL_7;
  assign _EVAL_29 = _EVAL_171[7:0];
  assign _EVAL_88 = 2'h2 == _EVAL_46 ? _EVAL_80 : _EVAL_217;
  assign _EVAL_199 = 2'h3 == _EVAL_46 ? _EVAL_29 : _EVAL_88;
  assign _EVAL_37 = {_EVAL_95,_EVAL_199};
  assign _EVAL_195 = _EVAL_171[31:24];
  assign _EVAL_230 = _EVAL_165 ? _EVAL_71 : 2'h0;
  assign _EVAL_55 = _EVAL_143[31:24];
  assign _EVAL_57 = _EVAL[31:24];
  assign _EVAL_23 = 2'h1 == _EVAL_230 ? _EVAL_234 : _EVAL_57;
  assign _EVAL_232 = 2'h2 == _EVAL_230 ? _EVAL_55 : _EVAL_23;
  assign _EVAL_47 = 2'h3 == _EVAL_230 ? _EVAL_195 : _EVAL_232;
  assign _EVAL_252 = {_EVAL_47,_EVAL_137};
  assign _EVAL_0 = {_EVAL_252,_EVAL_37};
endmodule
