//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_75(
  input         _EVAL,
  input  [7:0]  _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  output [1:0]  _EVAL_3,
  output [31:0] _EVAL_4,
  output [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  output        _EVAL_7,
  input  [31:0] _EVAL_8,
  output [7:0]  _EVAL_9,
  input         _EVAL_10,
  output [7:0]  _EVAL_11,
  input  [7:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14
);
  reg [7:0] _EVAL_18 [0:1];
  reg [31:0] _RAND_0;
  wire [7:0] _EVAL_18__EVAL_19_data;
  wire  _EVAL_18__EVAL_19_addr;
  wire [7:0] _EVAL_18__EVAL_20_data;
  wire  _EVAL_18__EVAL_20_addr;
  wire  _EVAL_18__EVAL_20_mask;
  wire  _EVAL_18__EVAL_20_en;
  reg [1:0] _EVAL_22 [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] _EVAL_22__EVAL_23_data;
  wire  _EVAL_22__EVAL_23_addr;
  wire [1:0] _EVAL_22__EVAL_24_data;
  wire  _EVAL_22__EVAL_24_addr;
  wire  _EVAL_22__EVAL_24_mask;
  wire  _EVAL_22__EVAL_24_en;
  reg [7:0] _EVAL_34 [0:1];
  reg [31:0] _RAND_2;
  wire [7:0] _EVAL_34__EVAL_35_data;
  wire  _EVAL_34__EVAL_35_addr;
  wire [7:0] _EVAL_34__EVAL_36_data;
  wire  _EVAL_34__EVAL_36_addr;
  wire  _EVAL_34__EVAL_36_mask;
  wire  _EVAL_34__EVAL_36_en;
  reg [2:0] _EVAL_41 [0:1];
  reg [31:0] _RAND_3;
  wire [2:0] _EVAL_41__EVAL_42_data;
  wire  _EVAL_41__EVAL_42_addr;
  wire [2:0] _EVAL_41__EVAL_43_data;
  wire  _EVAL_41__EVAL_43_addr;
  wire  _EVAL_41__EVAL_43_mask;
  wire  _EVAL_41__EVAL_43_en;
  reg [31:0] _EVAL_44 [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] _EVAL_44__EVAL_45_data;
  wire  _EVAL_44__EVAL_45_addr;
  wire [31:0] _EVAL_44__EVAL_46_data;
  wire  _EVAL_44__EVAL_46_addr;
  wire  _EVAL_44__EVAL_46_mask;
  wire  _EVAL_44__EVAL_46_en;
  reg  _EVAL_33;
  reg [31:0] _RAND_5;
  reg  _EVAL_38;
  reg [31:0] _RAND_6;
  reg  _EVAL_39;
  reg [31:0] _RAND_7;
  wire  _EVAL_25;
  wire  _EVAL_17;
  wire  _EVAL_30;
  wire  _EVAL_26;
  wire  _EVAL_16;
  wire  _EVAL_40;
  wire  _EVAL_28;
  wire  _EVAL_32;
  wire  _EVAL_15;
  assign _EVAL_18__EVAL_19_addr = _EVAL_33;
  assign _EVAL_18__EVAL_19_data = _EVAL_18[_EVAL_18__EVAL_19_addr];
  assign _EVAL_18__EVAL_20_data = _EVAL_0;
  assign _EVAL_18__EVAL_20_addr = _EVAL_39;
  assign _EVAL_18__EVAL_20_mask = 1'h1;
  assign _EVAL_18__EVAL_20_en = _EVAL_14 & _EVAL_10;
  assign _EVAL_22__EVAL_23_addr = _EVAL_33;
  assign _EVAL_22__EVAL_23_data = _EVAL_22[_EVAL_22__EVAL_23_addr];
  assign _EVAL_22__EVAL_24_data = _EVAL_2;
  assign _EVAL_22__EVAL_24_addr = _EVAL_39;
  assign _EVAL_22__EVAL_24_mask = 1'h1;
  assign _EVAL_22__EVAL_24_en = _EVAL_14 & _EVAL_10;
  assign _EVAL_34__EVAL_35_addr = _EVAL_33;
  assign _EVAL_34__EVAL_35_data = _EVAL_34[_EVAL_34__EVAL_35_addr];
  assign _EVAL_34__EVAL_36_data = _EVAL_12;
  assign _EVAL_34__EVAL_36_addr = _EVAL_39;
  assign _EVAL_34__EVAL_36_mask = 1'h1;
  assign _EVAL_34__EVAL_36_en = _EVAL_14 & _EVAL_10;
  assign _EVAL_41__EVAL_42_addr = _EVAL_33;
  assign _EVAL_41__EVAL_42_data = _EVAL_41[_EVAL_41__EVAL_42_addr];
  assign _EVAL_41__EVAL_43_data = _EVAL_6;
  assign _EVAL_41__EVAL_43_addr = _EVAL_39;
  assign _EVAL_41__EVAL_43_mask = 1'h1;
  assign _EVAL_41__EVAL_43_en = _EVAL_14 & _EVAL_10;
  assign _EVAL_44__EVAL_45_addr = _EVAL_33;
  assign _EVAL_44__EVAL_45_data = _EVAL_44[_EVAL_44__EVAL_45_addr];
  assign _EVAL_44__EVAL_46_data = _EVAL_8;
  assign _EVAL_44__EVAL_46_addr = _EVAL_39;
  assign _EVAL_44__EVAL_46_mask = 1'h1;
  assign _EVAL_44__EVAL_46_en = _EVAL_14 & _EVAL_10;
  assign _EVAL_25 = _EVAL_39 + 1'h1;
  assign _EVAL_17 = _EVAL_1 & _EVAL_7;
  assign _EVAL_30 = _EVAL_33 + 1'h1;
  assign _EVAL_26 = _EVAL_14 & _EVAL_10;
  assign _EVAL_16 = _EVAL_39 == _EVAL_33;
  assign _EVAL_40 = _EVAL_38 == 1'h0;
  assign _EVAL_28 = _EVAL_16 & _EVAL_40;
  assign _EVAL_32 = _EVAL_16 & _EVAL_38;
  assign _EVAL_15 = _EVAL_26 != _EVAL_17;
  assign _EVAL_4 = _EVAL_44__EVAL_45_data;
  assign _EVAL_14 = _EVAL_32 == 1'h0;
  assign _EVAL_5 = _EVAL_41__EVAL_42_data;
  assign _EVAL_9 = _EVAL_34__EVAL_35_data;
  assign _EVAL_7 = _EVAL_28 == 1'h0;
  assign _EVAL_3 = _EVAL_22__EVAL_23_data;
  assign _EVAL_11 = _EVAL_18__EVAL_19_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_18[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_22[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_34[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_41[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_44[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_33 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_38 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_39 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_13) begin
    if(_EVAL_18__EVAL_20_en & _EVAL_18__EVAL_20_mask) begin
      _EVAL_18[_EVAL_18__EVAL_20_addr] <= _EVAL_18__EVAL_20_data;
    end
    if(_EVAL_22__EVAL_24_en & _EVAL_22__EVAL_24_mask) begin
      _EVAL_22[_EVAL_22__EVAL_24_addr] <= _EVAL_22__EVAL_24_data;
    end
    if(_EVAL_34__EVAL_36_en & _EVAL_34__EVAL_36_mask) begin
      _EVAL_34[_EVAL_34__EVAL_36_addr] <= _EVAL_34__EVAL_36_data;
    end
    if(_EVAL_41__EVAL_43_en & _EVAL_41__EVAL_43_mask) begin
      _EVAL_41[_EVAL_41__EVAL_43_addr] <= _EVAL_41__EVAL_43_data;
    end
    if(_EVAL_44__EVAL_46_en & _EVAL_44__EVAL_46_mask) begin
      _EVAL_44[_EVAL_44__EVAL_46_addr] <= _EVAL_44__EVAL_46_data;
    end
    if (_EVAL) begin
      _EVAL_33 <= 1'h0;
    end else begin
      if (_EVAL_17) begin
        _EVAL_33 <= _EVAL_30;
      end
    end
    if (_EVAL) begin
      _EVAL_38 <= 1'h0;
    end else begin
      if (_EVAL_15) begin
        _EVAL_38 <= _EVAL_26;
      end
    end
    if (_EVAL) begin
      _EVAL_39 <= 1'h0;
    end else begin
      if (_EVAL_26) begin
        _EVAL_39 <= _EVAL_25;
      end
    end
  end
endmodule
