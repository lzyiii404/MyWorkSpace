//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_107_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [7:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [31:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [2:0]  _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_22;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_45;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_71;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_95;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_98;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_120;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_136;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_138;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_143;
  reg [31:0] _RAND_8;
  reg  _EVAL_144;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_183;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_202;
  reg [31:0] _RAND_11;
  reg  _EVAL_221;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_271;
  reg [31:0] _RAND_13;
  reg  _EVAL_278;
  reg [31:0] _RAND_14;
  wire  _EVAL_223;
  wire  _EVAL_195;
  wire  _EVAL_265;
  wire [1:0] _EVAL_252;
  wire [3:0] _EVAL_137;
  wire [2:0] _EVAL_214;
  wire [2:0] _EVAL_215;
  wire  _EVAL_127;
  wire  _EVAL_235;
  wire  _EVAL_158;
  wire  _EVAL_67;
  wire  _EVAL_124;
  wire  _EVAL_86;
  wire  _EVAL_115;
  wire  _EVAL_167;
  wire [12:0] _EVAL_108;
  wire [5:0] _EVAL_140;
  wire [5:0] _EVAL_267;
  wire [31:0] _EVAL_210;
  wire [32:0] _EVAL_142;
  wire  _EVAL_21;
  wire  _EVAL_152;
  wire  _EVAL_245;
  wire [12:0] _EVAL_273;
  wire [5:0] _EVAL_280;
  wire [5:0] _EVAL_250;
  wire [2:0] _EVAL_37;
  wire  _EVAL_50;
  wire  _EVAL_255;
  wire  _EVAL_128;
  wire  _EVAL_92;
  wire [2:0] _EVAL_44;
  wire [2:0] _EVAL_263;
  wire  _EVAL_26;
  wire  _EVAL_156;
  wire  _EVAL_94;
  wire  _EVAL_243;
  wire [2:0] _EVAL_111;
  wire  _EVAL_251;
  wire  _EVAL_199;
  wire  _EVAL_181;
  wire  _EVAL_87;
  wire  _EVAL_182;
  wire  _EVAL_29;
  wire  _EVAL_197;
  wire  _EVAL_177;
  wire  _EVAL_234;
  wire  _EVAL_169;
  wire [1:0] _EVAL_57;
  wire [1:0] _EVAL_194;
  wire [1:0] _EVAL_153;
  wire [1:0] _EVAL_148;
  wire  _EVAL_103;
  wire  _EVAL_135;
  wire  _EVAL_240;
  wire  _EVAL_79;
  wire  _EVAL_93;
  wire  _EVAL_72;
  wire  _EVAL_165;
  wire  _EVAL_33;
  wire  _EVAL_121;
  wire  _EVAL_157;
  wire  _EVAL_147;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_134;
  wire  _EVAL_196;
  wire  _EVAL_141;
  wire  _EVAL_62;
  wire  _EVAL_122;
  wire  _EVAL_132;
  wire  _EVAL_53;
  wire  _EVAL_75;
  wire  _EVAL_73;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_96;
  wire  _EVAL_123;
  wire [1:0] _EVAL_188;
  wire [1:0] _EVAL_227;
  wire  _EVAL_101;
  wire  _EVAL_272;
  wire  _EVAL_77;
  wire  _EVAL_261;
  wire  _EVAL_218;
  wire  _EVAL_217;
  wire  _EVAL_104;
  wire  _EVAL_206;
  wire  _EVAL_229;
  wire  _EVAL_207;
  wire  _EVAL_131;
  wire  _EVAL_40;
  wire  _EVAL_189;
  wire  _EVAL_97;
  wire  _EVAL_254;
  wire  _EVAL_220;
  wire  _EVAL_190;
  wire  _EVAL_257;
  wire  _EVAL_70;
  wire  _EVAL_239;
  wire  _EVAL_187;
  wire  _EVAL_39;
  wire  _EVAL_205;
  wire  _EVAL_52;
  wire  _EVAL_151;
  wire  _EVAL_238;
  wire [7:0] _EVAL_83;
  wire [7:0] _EVAL_24;
  wire [7:0] _EVAL_85;
  wire  _EVAL_283;
  wire  _EVAL_164;
  wire  _EVAL_244;
  wire [2:0] _EVAL_25;
  wire  _EVAL_76;
  wire  _EVAL_32;
  wire  _EVAL_213;
  wire [7:0] _EVAL_166;
  wire  _EVAL_170;
  wire  _EVAL_80;
  wire  _EVAL_224;
  wire  _EVAL_168;
  wire  _EVAL_42;
  wire  _EVAL_47;
  wire  _EVAL_246;
  wire  _EVAL_109;
  wire  _EVAL_133;
  wire  _EVAL_259;
  wire  _EVAL_91;
  wire  _EVAL_110;
  wire  _EVAL_281;
  wire  _EVAL_61;
  wire  _EVAL_262;
  wire  _EVAL_66;
  wire  _EVAL_191;
  wire  _EVAL_106;
  wire  _EVAL_41;
  wire  _EVAL_18;
  wire  _EVAL_60;
  wire  _EVAL_249;
  wire [2:0] _EVAL_242;
  wire  _EVAL_49;
  wire  _EVAL_211;
  wire  _EVAL_125;
  wire [31:0] _EVAL_216;
  wire  _EVAL_119;
  wire  _EVAL_225;
  wire  _EVAL_69;
  wire  _EVAL_58;
  wire  _EVAL_54;
  wire  _EVAL_233;
  wire  _EVAL_102;
  wire  _EVAL_117;
  wire  _EVAL_230;
  wire  _EVAL_219;
  wire [1:0] _EVAL_126;
  wire  _EVAL_84;
  wire  _EVAL_31;
  wire  _EVAL_19;
  wire  _EVAL_30;
  wire  _EVAL_178;
  wire  _EVAL_173;
  wire [31:0] _EVAL_174;
  wire [31:0] _EVAL_186;
  wire  _EVAL_46;
  wire  _EVAL_59;
  wire  _EVAL_129;
  wire  _EVAL_185;
  wire  _EVAL_82;
  wire  _EVAL_113;
  wire  _EVAL_282;
  wire  _EVAL_269;
  wire  _EVAL_208;
  wire  _EVAL_184;
  wire  _EVAL_17;
  wire  _EVAL_279;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [1:0] _EVAL_275;
  wire [1:0] _EVAL_179;
  wire  _EVAL_90;
  wire  _EVAL_116;
  wire [1:0] _EVAL_74;
  wire  _EVAL_268;
  wire  _EVAL_112;
  wire  _EVAL_100;
  wire  _EVAL_266;
  wire  _EVAL_55;
  wire  _EVAL_36;
  wire  _EVAL_231;
  wire  _EVAL_162;
  wire  _EVAL_253;
  wire  _EVAL_175;
  wire  _EVAL_27;
  wire  _EVAL_139;
  wire  _EVAL_51;
  wire  _EVAL_20;
  wire  _EVAL_68;
  wire  _EVAL_171;
  wire  _EVAL_163;
  wire  _EVAL_155;
  wire  _EVAL_209;
  wire  _EVAL_264;
  wire  _EVAL_212;
  wire  _EVAL_277;
  wire  _EVAL_236;
  wire  _EVAL_201;
  wire  _EVAL_145;
  wire  _EVAL_28;
  wire  _EVAL_180;
  wire  _EVAL_192;
  wire  _EVAL_274;
  wire  _EVAL_241;
  wire  _EVAL_154;
  wire  _EVAL_200;
  wire  _EVAL_48;
  wire  _EVAL_23;
  wire  _EVAL_78;
  wire  _EVAL_130;
  wire  _EVAL_198;
  wire  _EVAL_65;
  wire  _EVAL_256;
  wire  _EVAL_146;
  wire  _EVAL_149;
  wire  _EVAL_232;
  wire  _EVAL_159;
  wire  _EVAL_260;
  wire  _EVAL_248;
  wire  _EVAL_172;
  wire  _EVAL_64;
  wire  _EVAL_204;
  wire  _EVAL_89;
  wire  _EVAL_222;
  wire  _EVAL_114;
  wire  _EVAL_258;
  wire  _EVAL_63;
  wire  _EVAL_118;
  wire  _EVAL_38;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_223 = _EVAL_120 == 3'h0;
  assign _EVAL_195 = _EVAL_223 == 1'h0;
  assign _EVAL_265 = _EVAL_14 & _EVAL_195;
  assign _EVAL_252 = _EVAL_15[1:0];
  assign _EVAL_137 = 4'h1 << _EVAL_252;
  assign _EVAL_214 = _EVAL_137[2:0];
  assign _EVAL_215 = _EVAL_214 | 3'h1;
  assign _EVAL_127 = _EVAL_215[0];
  assign _EVAL_235 = _EVAL_5[2];
  assign _EVAL_158 = _EVAL_235 == 1'h0;
  assign _EVAL_67 = _EVAL_5[1];
  assign _EVAL_124 = _EVAL_158 & _EVAL_67;
  assign _EVAL_86 = _EVAL_5[0];
  assign _EVAL_115 = _EVAL_124 & _EVAL_86;
  assign _EVAL_167 = _EVAL_127 & _EVAL_115;
  assign _EVAL_108 = 13'h3f << _EVAL_15;
  assign _EVAL_140 = _EVAL_108[5:0];
  assign _EVAL_267 = ~ _EVAL_140;
  assign _EVAL_210 = _EVAL_5 ^ 32'h80000000;
  assign _EVAL_142 = {1'b0,$signed(_EVAL_210)};
  assign _EVAL_21 = _EVAL_235 & _EVAL_67;
  assign _EVAL_152 = _EVAL_215[2];
  assign _EVAL_245 = _EVAL_152 & _EVAL_235;
  assign _EVAL_273 = 13'h3f << _EVAL;
  assign _EVAL_280 = _EVAL_273[5:0];
  assign _EVAL_250 = ~ _EVAL_280;
  assign _EVAL_37 = _EVAL_250[5:3];
  assign _EVAL_50 = _EVAL_10 & _EVAL_13;
  assign _EVAL_255 = _EVAL_202 == 3'h0;
  assign _EVAL_128 = _EVAL_12[2];
  assign _EVAL_92 = _EVAL_128 == 1'h0;
  assign _EVAL_44 = _EVAL_267[5:3];
  assign _EVAL_263 = _EVAL_202 - 3'h1;
  assign _EVAL_26 = _EVAL_15 >= 3'h3;
  assign _EVAL_156 = _EVAL_26 | _EVAL_11;
  assign _EVAL_94 = _EVAL_156 == 1'h0;
  assign _EVAL_243 = _EVAL_45 == 3'h0;
  assign _EVAL_111 = _EVAL_45 - 3'h1;
  assign _EVAL_251 = _EVAL_152 & _EVAL_158;
  assign _EVAL_199 = _EVAL_26 | _EVAL_251;
  assign _EVAL_181 = _EVAL_215[1];
  assign _EVAL_87 = _EVAL_181 & _EVAL_124;
  assign _EVAL_182 = _EVAL_199 | _EVAL_87;
  assign _EVAL_29 = _EVAL_86 == 1'h0;
  assign _EVAL_197 = _EVAL_124 & _EVAL_29;
  assign _EVAL_177 = _EVAL_127 & _EVAL_197;
  assign _EVAL_234 = _EVAL_182 | _EVAL_177;
  assign _EVAL_169 = _EVAL_50 & _EVAL_255;
  assign _EVAL_57 = 2'h1 << _EVAL_8;
  assign _EVAL_194 = _EVAL_169 ? _EVAL_57 : 2'h0;
  assign _EVAL_153 = _EVAL_194 | _EVAL_183;
  assign _EVAL_148 = _EVAL_153 >> _EVAL_4;
  assign _EVAL_103 = _EVAL_148[0];
  assign _EVAL_135 = _EVAL_16 != 3'h0;
  assign _EVAL_240 = _EVAL_135 | _EVAL_11;
  assign _EVAL_79 = _EVAL_240 == 1'h0;
  assign _EVAL_93 = _EVAL_1 & _EVAL_14;
  assign _EVAL_72 = _EVAL_138 == 3'h0;
  assign _EVAL_165 = _EVAL_93 & _EVAL_72;
  assign _EVAL_33 = _EVAL_4 == _EVAL_278;
  assign _EVAL_121 = _EVAL_33 | _EVAL_11;
  assign _EVAL_157 = _EVAL_121 == 1'h0;
  assign _EVAL_147 = _EVAL_5 == _EVAL_271;
  assign _EVAL_150 = $signed(_EVAL_142) & $signed(-33'sh20000);
  assign _EVAL_134 = $signed(_EVAL_150);
  assign _EVAL_196 = _EVAL_67 == 1'h0;
  assign _EVAL_141 = _EVAL_158 & _EVAL_196;
  assign _EVAL_62 = _EVAL_181 & _EVAL_141;
  assign _EVAL_122 = _EVAL_199 | _EVAL_62;
  assign _EVAL_132 = _EVAL_141 & _EVAL_29;
  assign _EVAL_53 = _EVAL_127 & _EVAL_132;
  assign _EVAL_75 = _EVAL_122 | _EVAL_53;
  assign _EVAL_73 = _EVAL_7 == 1'h0;
  assign _EVAL_34 = _EVAL_73 | _EVAL_11;
  assign _EVAL_35 = _EVAL_9 == 3'h6;
  assign _EVAL_96 = _EVAL_35 == 1'h0;
  assign _EVAL_123 = _EVAL_165 & _EVAL_96;
  assign _EVAL_188 = 2'h1 << _EVAL_4;
  assign _EVAL_227 = _EVAL_123 ? _EVAL_188 : 2'h0;
  assign _EVAL_101 = _EVAL_194 != _EVAL_227;
  assign _EVAL_272 = _EVAL_194 != 2'h0;
  assign _EVAL_77 = _EVAL_272 == 1'h0;
  assign _EVAL_261 = _EVAL_101 | _EVAL_77;
  assign _EVAL_218 = _EVAL_26 | _EVAL_245;
  assign _EVAL_217 = _EVAL_181 & _EVAL_21;
  assign _EVAL_104 = _EVAL_218 | _EVAL_217;
  assign _EVAL_206 = _EVAL_21 & _EVAL_86;
  assign _EVAL_229 = _EVAL_127 & _EVAL_206;
  assign _EVAL_207 = _EVAL_104 | _EVAL_229;
  assign _EVAL_131 = _EVAL_21 & _EVAL_29;
  assign _EVAL_40 = _EVAL_127 & _EVAL_131;
  assign _EVAL_189 = _EVAL_104 | _EVAL_40;
  assign _EVAL_97 = _EVAL_235 & _EVAL_196;
  assign _EVAL_254 = _EVAL_181 & _EVAL_97;
  assign _EVAL_220 = _EVAL_218 | _EVAL_254;
  assign _EVAL_190 = _EVAL_97 & _EVAL_86;
  assign _EVAL_257 = _EVAL_127 & _EVAL_190;
  assign _EVAL_70 = _EVAL_220 | _EVAL_257;
  assign _EVAL_239 = _EVAL_97 & _EVAL_29;
  assign _EVAL_187 = _EVAL_127 & _EVAL_239;
  assign _EVAL_39 = _EVAL_220 | _EVAL_187;
  assign _EVAL_205 = _EVAL_182 | _EVAL_167;
  assign _EVAL_52 = _EVAL_141 & _EVAL_86;
  assign _EVAL_151 = _EVAL_127 & _EVAL_52;
  assign _EVAL_238 = _EVAL_122 | _EVAL_151;
  assign _EVAL_83 = {_EVAL_207,_EVAL_189,_EVAL_70,_EVAL_39,_EVAL_205,_EVAL_234,_EVAL_238,_EVAL_75};
  assign _EVAL_24 = ~ _EVAL_83;
  assign _EVAL_85 = _EVAL_2 & _EVAL_24;
  assign _EVAL_283 = _EVAL_85 == 8'h0;
  assign _EVAL_164 = _EVAL_283 | _EVAL_11;
  assign _EVAL_244 = _EVAL_16 == _EVAL_95;
  assign _EVAL_25 = _EVAL_120 - 3'h1;
  assign _EVAL_76 = _EVAL_12 == 3'h4;
  assign _EVAL_32 = _EVAL_3 == 1'h0;
  assign _EVAL_213 = _EVAL_32 | _EVAL_11;
  assign _EVAL_166 = ~ _EVAL_2;
  assign _EVAL_170 = _EVAL_166 == 8'h0;
  assign _EVAL_80 = _EVAL_170 | _EVAL_11;
  assign _EVAL_224 = plusarg_reader_out == 32'h0;
  assign _EVAL_168 = _EVAL_12 == 3'h1;
  assign _EVAL_42 = _EVAL_13 & _EVAL_168;
  assign _EVAL_47 = _EVAL_12 == _EVAL_136;
  assign _EVAL_246 = _EVAL_47 | _EVAL_11;
  assign _EVAL_109 = _EVAL_147 | _EVAL_11;
  assign _EVAL_133 = _EVAL_16 == 3'h0;
  assign _EVAL_259 = _EVAL_9 <= 3'h6;
  assign _EVAL_91 = _EVAL_259 | _EVAL_11;
  assign _EVAL_110 = $signed(_EVAL_134) == $signed(33'sh0);
  assign _EVAL_281 = _EVAL_15 <= 3'h6;
  assign _EVAL_61 = _EVAL_6 == 1'h0;
  assign _EVAL_262 = _EVAL_61 | _EVAL_11;
  assign _EVAL_66 = _EVAL_2 == _EVAL_83;
  assign _EVAL_191 = _EVAL_66 | _EVAL_11;
  assign _EVAL_106 = _EVAL_191 == 1'h0;
  assign _EVAL_41 = _EVAL_12 == 3'h2;
  assign _EVAL_18 = _EVAL_15 == _EVAL_98;
  assign _EVAL_60 = _EVAL >= 3'h3;
  assign _EVAL_249 = _EVAL_60 | _EVAL_11;
  assign _EVAL_242 = _EVAL_138 - 3'h1;
  assign _EVAL_49 = _EVAL_243 == 1'h0;
  assign _EVAL_211 = _EVAL_9 == 3'h5;
  assign _EVAL_125 = _EVAL_14 & _EVAL_211;
  assign _EVAL_216 = _EVAL_22 + 32'h1;
  assign _EVAL_119 = _EVAL_164 == 1'h0;
  assign _EVAL_225 = _EVAL_8 == _EVAL_221;
  assign _EVAL_69 = _EVAL_225 | _EVAL_11;
  assign _EVAL_58 = _EVAL_69 == 1'h0;
  assign _EVAL_54 = _EVAL_9[0];
  assign _EVAL_233 = _EVAL_12 == 3'h7;
  assign _EVAL_102 = _EVAL_13 & _EVAL_233;
  assign _EVAL_117 = _EVAL_16 <= 3'h2;
  assign _EVAL_230 = _EVAL_117 | _EVAL_11;
  assign _EVAL_219 = _EVAL_230 == 1'h0;
  assign _EVAL_126 = ~ _EVAL_227;
  assign _EVAL_84 = _EVAL_93 & _EVAL_223;
  assign _EVAL_31 = _EVAL_9 == _EVAL_71;
  assign _EVAL_19 = _EVAL_12 == 3'h3;
  assign _EVAL_30 = _EVAL_34 == 1'h0;
  assign _EVAL_178 = _EVAL_261 | _EVAL_11;
  assign _EVAL_173 = _EVAL_178 == 1'h0;
  assign _EVAL_174 = {{26'd0}, _EVAL_267};
  assign _EVAL_186 = _EVAL_5 & _EVAL_174;
  assign _EVAL_46 = _EVAL_186 == 32'h0;
  assign _EVAL_59 = _EVAL_46 | _EVAL_11;
  assign _EVAL_129 = _EVAL_281 & _EVAL_110;
  assign _EVAL_185 = _EVAL_129 | _EVAL_11;
  assign _EVAL_82 = _EVAL_185 == 1'h0;
  assign _EVAL_113 = _EVAL_103 | _EVAL_11;
  assign _EVAL_282 = _EVAL_113 == 1'h0;
  assign _EVAL_269 = _EVAL_12 == 3'h0;
  assign _EVAL_208 = _EVAL_13 & _EVAL_269;
  assign _EVAL_184 = _EVAL_16 <= 3'h4;
  assign _EVAL_17 = _EVAL_184 | _EVAL_11;
  assign _EVAL_279 = _EVAL_17 == 1'h0;
  assign _EVAL_160 = _EVAL_9 == 3'h2;
  assign _EVAL_161 = _EVAL_14 & _EVAL_160;
  assign _EVAL_275 = _EVAL_183 | _EVAL_194;
  assign _EVAL_179 = _EVAL_275 & _EVAL_126;
  assign _EVAL_90 = _EVAL_80 == 1'h0;
  assign _EVAL_116 = _EVAL_183 != 2'h0;
  assign _EVAL_74 = _EVAL_183 >> _EVAL_8;
  assign _EVAL_268 = _EVAL_74[0];
  assign _EVAL_112 = _EVAL_268 == 1'h0;
  assign _EVAL_100 = _EVAL_112 | _EVAL_11;
  assign _EVAL_266 = _EVAL_91 == 1'h0;
  assign _EVAL_55 = _EVAL_73 | _EVAL_6;
  assign _EVAL_36 = _EVAL_55 | _EVAL_11;
  assign _EVAL_231 = _EVAL_50 | _EVAL_93;
  assign _EVAL_162 = _EVAL_16 <= 3'h3;
  assign _EVAL_253 = _EVAL_162 | _EVAL_11;
  assign _EVAL_175 = _EVAL_253 == 1'h0;
  assign _EVAL_27 = _EVAL_12 == 3'h6;
  assign _EVAL_139 = _EVAL_13 & _EVAL_27;
  assign _EVAL_51 = _EVAL_249 == 1'h0;
  assign _EVAL_20 = _EVAL_13 & _EVAL_41;
  assign _EVAL_68 = _EVAL_13 & _EVAL_76;
  assign _EVAL_171 = _EVAL_11 == 1'h0;
  assign _EVAL_163 = _EVAL_262 == 1'h0;
  assign _EVAL_155 = _EVAL_13 & _EVAL_19;
  assign _EVAL_209 = _EVAL_9 == 3'h1;
  assign _EVAL_264 = _EVAL_14 & _EVAL_209;
  assign _EVAL_212 = _EVAL_9 == 3'h4;
  assign _EVAL_277 = _EVAL_14 & _EVAL_212;
  assign _EVAL_236 = _EVAL_12 == 3'h5;
  assign _EVAL_201 = _EVAL_13 & _EVAL_236;
  assign _EVAL_145 = _EVAL_246 == 1'h0;
  assign _EVAL_28 = _EVAL_9 == 3'h0;
  assign _EVAL_180 = _EVAL_13 & _EVAL_49;
  assign _EVAL_192 = _EVAL == _EVAL_143;
  assign _EVAL_274 = _EVAL_100 == 1'h0;
  assign _EVAL_241 = _EVAL_22 < plusarg_reader_out;
  assign _EVAL_154 = _EVAL_31 | _EVAL_11;
  assign _EVAL_200 = _EVAL_133 | _EVAL_11;
  assign _EVAL_48 = _EVAL_200 == 1'h0;
  assign _EVAL_23 = _EVAL_192 | _EVAL_11;
  assign _EVAL_78 = _EVAL_23 == 1'h0;
  assign _EVAL_130 = _EVAL_14 & _EVAL_28;
  assign _EVAL_198 = _EVAL_244 | _EVAL_11;
  assign _EVAL_65 = _EVAL_7 == _EVAL_144;
  assign _EVAL_256 = _EVAL_198 == 1'h0;
  assign _EVAL_146 = _EVAL_59 == 1'h0;
  assign _EVAL_149 = _EVAL_116 == 1'h0;
  assign _EVAL_232 = _EVAL_149 | _EVAL_224;
  assign _EVAL_159 = _EVAL_232 | _EVAL_241;
  assign _EVAL_260 = _EVAL_18 | _EVAL_11;
  assign _EVAL_248 = _EVAL_260 == 1'h0;
  assign _EVAL_172 = _EVAL_65 | _EVAL_11;
  assign _EVAL_64 = _EVAL_172 == 1'h0;
  assign _EVAL_204 = _EVAL_213 == 1'h0;
  assign _EVAL_89 = _EVAL_50 & _EVAL_243;
  assign _EVAL_222 = _EVAL_154 == 1'h0;
  assign _EVAL_114 = _EVAL_36 == 1'h0;
  assign _EVAL_258 = _EVAL_109 == 1'h0;
  assign _EVAL_63 = _EVAL_159 | _EVAL_11;
  assign _EVAL_118 = _EVAL_63 == 1'h0;
  assign _EVAL_38 = _EVAL_14 & _EVAL_35;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_45 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_71 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_95 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_98 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_120 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_136 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_138 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_143 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_144 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_183 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_202 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_221 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_271 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_278 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_11) begin
      _EVAL_22 <= 32'h0;
    end else begin
      if (_EVAL_231) begin
        _EVAL_22 <= 32'h0;
      end else begin
        _EVAL_22 <= _EVAL_216;
      end
    end
    if (_EVAL_11) begin
      _EVAL_45 <= 3'h0;
    end else begin
      if (_EVAL_50) begin
        if (_EVAL_243) begin
          if (_EVAL_92) begin
            _EVAL_45 <= _EVAL_44;
          end else begin
            _EVAL_45 <= 3'h0;
          end
        end else begin
          _EVAL_45 <= _EVAL_111;
        end
      end
    end
    if (_EVAL_84) begin
      _EVAL_71 <= _EVAL_9;
    end
    if (_EVAL_89) begin
      _EVAL_95 <= _EVAL_16;
    end
    if (_EVAL_89) begin
      _EVAL_98 <= _EVAL_15;
    end
    if (_EVAL_11) begin
      _EVAL_120 <= 3'h0;
    end else begin
      if (_EVAL_93) begin
        if (_EVAL_223) begin
          if (_EVAL_54) begin
            _EVAL_120 <= _EVAL_37;
          end else begin
            _EVAL_120 <= 3'h0;
          end
        end else begin
          _EVAL_120 <= _EVAL_25;
        end
      end
    end
    if (_EVAL_89) begin
      _EVAL_136 <= _EVAL_12;
    end
    if (_EVAL_11) begin
      _EVAL_138 <= 3'h0;
    end else begin
      if (_EVAL_93) begin
        if (_EVAL_72) begin
          if (_EVAL_54) begin
            _EVAL_138 <= _EVAL_37;
          end else begin
            _EVAL_138 <= 3'h0;
          end
        end else begin
          _EVAL_138 <= _EVAL_242;
        end
      end
    end
    if (_EVAL_84) begin
      _EVAL_143 <= _EVAL;
    end
    if (_EVAL_84) begin
      _EVAL_144 <= _EVAL_7;
    end
    if (_EVAL_11) begin
      _EVAL_183 <= 2'h0;
    end else begin
      _EVAL_183 <= _EVAL_179;
    end
    if (_EVAL_11) begin
      _EVAL_202 <= 3'h0;
    end else begin
      if (_EVAL_50) begin
        if (_EVAL_255) begin
          if (_EVAL_92) begin
            _EVAL_202 <= _EVAL_44;
          end else begin
            _EVAL_202 <= 3'h0;
          end
        end else begin
          _EVAL_202 <= _EVAL_263;
        end
      end
    end
    if (_EVAL_89) begin
      _EVAL_221 <= _EVAL_8;
    end
    if (_EVAL_89) begin
      _EVAL_271 <= _EVAL_5;
    end
    if (_EVAL_84) begin
      _EVAL_278 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e68bc1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfc6eadd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38c3a380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58491693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b77ed0a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66f75524)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15a284e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4a7e6a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a025fdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(777ed5de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b98c5095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9af0428)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b540c228)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5edbb95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4fcb350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97dc813c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f59560)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a207400)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ace1dbf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5f739cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(706c03e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5b49890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc2050a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53162d9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1fae00b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69e1ebdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6459485d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b14488f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6ce67f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c42c953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721dc194)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a042ba51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a56b1dd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47ecf248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9db566b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f6c7522)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c16500c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6c2de99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e707ce0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(161efcca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a78810f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c097850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad64d095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(315befc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(def89d9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aacaa672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0856b22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b0515fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ba90369)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f672c7b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3907fde7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6390e3fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(621bed34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eca7e636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e71f0aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(129714ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37082b1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a81bc1ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac7d168f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ad28b60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2651694)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(278be24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc66bfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b54d89c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7bca6d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9cdd90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
