//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_212_assert(
  input         _EVAL,
  input  [11:0] _EVAL_0,
  input  [11:0] _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [11:0] _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_23;
  reg [31:0] _RAND_0;
  reg [11:0] _EVAL_27;
  reg [31:0] _RAND_1;
  reg  _EVAL_40;
  reg [31:0] _RAND_2;
  reg  _EVAL_42;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_74;
  reg [31:0] _RAND_4;
  reg [11:0] _EVAL_98;
  reg [31:0] _RAND_5;
  reg [1:0] _EVAL_124;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_144;
  reg [31:0] _RAND_7;
  reg  _EVAL_175;
  reg [31:0] _RAND_8;
  reg [11:0] _EVAL_177;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_188;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_209;
  reg [31:0] _RAND_11;
  reg [2335:0] _EVAL_213;
  reg [2335:0] _RAND_12;
  reg [2:0] _EVAL_219;
  reg [31:0] _RAND_13;
  wire  _EVAL_168;
  wire  _EVAL_162;
  wire  _EVAL_113;
  wire  _EVAL_25;
  wire  _EVAL_150;
  wire  _EVAL_112;
  wire  _EVAL_158;
  wire  _EVAL_187;
  wire  _EVAL_159;
  wire  _EVAL_228;
  wire  _EVAL_115;
  wire  _EVAL_86;
  wire  _EVAL_135;
  wire [4095:0] _EVAL_36;
  wire [4095:0] _EVAL_205;
  wire [2335:0] _EVAL_200;
  wire [2335:0] _EVAL_194;
  wire [2335:0] _EVAL_55;
  wire  _EVAL_118;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_179;
  wire [4095:0] _EVAL_96;
  wire [4095:0] _EVAL_140;
  wire  _EVAL_75;
  wire  _EVAL_129;
  wire  _EVAL_52;
  wire  _EVAL_46;
  wire [1:0] _EVAL_131;
  wire [1:0] _EVAL_51;
  wire  _EVAL_49;
  wire  _EVAL_15;
  wire  _EVAL_178;
  wire  _EVAL_133;
  wire  _EVAL_73;
  wire [2335:0] _EVAL_214;
  wire [2335:0] _EVAL_121;
  wire [12:0] _EVAL_149;
  wire [12:0] _EVAL_45;
  wire [12:0] _EVAL_142;
  wire  _EVAL_71;
  wire  _EVAL_61;
  wire [4:0] _EVAL_81;
  wire [1:0] _EVAL_22;
  wire  _EVAL_66;
  wire  _EVAL_145;
  wire  _EVAL_198;
  wire  _EVAL_137;
  wire  _EVAL_18;
  wire  _EVAL_176;
  wire  _EVAL_220;
  wire  _EVAL_31;
  wire  _EVAL_148;
  wire  _EVAL_17;
  wire  _EVAL_180;
  wire  _EVAL_92;
  wire  _EVAL_182;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_190;
  wire  _EVAL_225;
  wire  _EVAL_216;
  wire  _EVAL_192;
  wire  _EVAL_189;
  wire [3:0] _EVAL_37;
  wire [3:0] _EVAL_89;
  wire [3:0] _EVAL_114;
  wire  _EVAL_67;
  wire  _EVAL_105;
  wire  _EVAL_127;
  wire  _EVAL_69;
  wire  _EVAL_64;
  wire  _EVAL_44;
  wire  _EVAL_157;
  wire  _EVAL_146;
  wire  _EVAL_153;
  wire  _EVAL_91;
  wire  _EVAL_53;
  wire  _EVAL_212;
  wire  _EVAL_120;
  wire  _EVAL_164;
  wire  _EVAL_125;
  wire  _EVAL_102;
  wire  _EVAL_141;
  wire  _EVAL_167;
  wire  _EVAL_38;
  wire  _EVAL_191;
  wire  _EVAL_94;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [1:0] _EVAL_147;
  wire [11:0] _EVAL_207;
  wire [11:0] _EVAL_84;
  wire  _EVAL_136;
  wire  _EVAL_199;
  wire  _EVAL_78;
  wire  _EVAL_21;
  wire  _EVAL_34;
  wire  _EVAL_184;
  wire  _EVAL_130;
  wire  _EVAL_183;
  wire  _EVAL_29;
  wire  _EVAL_155;
  wire  _EVAL_223;
  wire  _EVAL_32;
  wire  _EVAL_83;
  wire [31:0] _EVAL_231;
  wire  _EVAL_185;
  wire  _EVAL_109;
  wire  _EVAL_95;
  wire  _EVAL_171;
  wire  _EVAL_211;
  wire  _EVAL_161;
  wire  _EVAL_106;
  wire  _EVAL_206;
  wire  _EVAL_60;
  wire  _EVAL_80;
  wire [3:0] _EVAL_117;
  wire  _EVAL_122;
  wire  _EVAL_181;
  wire  _EVAL_19;
  wire  _EVAL_41;
  wire  _EVAL_85;
  wire [2335:0] _EVAL_165;
  wire  _EVAL_116;
  wire  _EVAL_229;
  wire  _EVAL_68;
  wire  _EVAL_39;
  wire  _EVAL_215;
  wire  _EVAL_143;
  wire  _EVAL_196;
  wire  _EVAL_217;
  wire  _EVAL_70;
  wire  _EVAL_108;
  wire  _EVAL_119;
  wire  _EVAL_208;
  wire  _EVAL_62;
  wire  _EVAL_103;
  wire  _EVAL_56;
  wire  _EVAL_24;
  wire  _EVAL_87;
  wire  _EVAL_77;
  wire  _EVAL_47;
  wire  _EVAL_201;
  wire  _EVAL_163;
  wire  _EVAL_134;
  wire  _EVAL_152;
  wire  _EVAL_99;
  wire  _EVAL_59;
  wire  _EVAL_110;
  wire  _EVAL_174;
  wire  _EVAL_154;
  wire  _EVAL_16;
  wire  _EVAL_156;
  wire  _EVAL_28;
  wire  _EVAL_63;
  wire  _EVAL_111;
  wire  _EVAL_166;
  wire [2335:0] _EVAL_50;
  wire  _EVAL_104;
  wire  _EVAL_210;
  wire  _EVAL_43;
  wire  _EVAL_170;
  wire  _EVAL_202;
  wire  _EVAL_76;
  wire  _EVAL_139;
  wire  _EVAL_227;
  wire  _EVAL_20;
  wire  _EVAL_126;
  wire  _EVAL_226;
  wire  _EVAL_169;
  wire  _EVAL_33;
  wire  _EVAL_65;
  wire  _EVAL_138;
  wire  _EVAL_222;
  wire  _EVAL_132;
  wire  _EVAL_72;
  wire [2335:0] _EVAL_82;
  wire  _EVAL_221;
  wire  _EVAL_224;
  wire  _EVAL_123;
  wire  _EVAL_93;
  wire  _EVAL_97;
  wire  _EVAL_193;
  wire  _EVAL_218;
  wire  _EVAL_197;
  wire  _EVAL_54;
  wire  _EVAL_90;
  wire  _EVAL_57;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_168 = _EVAL_10 <= 3'h2;
  assign _EVAL_162 = _EVAL_5 == 3'h0;
  assign _EVAL_113 = _EVAL_11 & _EVAL_162;
  assign _EVAL_25 = _EVAL_1[0];
  assign _EVAL_150 = _EVAL_213 != 2336'h0;
  assign _EVAL_112 = _EVAL_150 == 1'h0;
  assign _EVAL_158 = _EVAL_5 == 3'h5;
  assign _EVAL_187 = _EVAL_4 & _EVAL_11;
  assign _EVAL_159 = _EVAL_175 == 1'h0;
  assign _EVAL_228 = _EVAL_175 - 1'h1;
  assign _EVAL_115 = _EVAL_12 & _EVAL_9;
  assign _EVAL_86 = _EVAL_42 == 1'h0;
  assign _EVAL_135 = _EVAL_115 & _EVAL_86;
  assign _EVAL_36 = 4096'h1 << _EVAL_14;
  assign _EVAL_205 = _EVAL_135 ? _EVAL_36 : 4096'h0;
  assign _EVAL_200 = _EVAL_205[2335:0];
  assign _EVAL_194 = _EVAL_200 | _EVAL_213;
  assign _EVAL_55 = _EVAL_194 >> _EVAL_0;
  assign _EVAL_118 = _EVAL_187 & _EVAL_159;
  assign _EVAL_203 = _EVAL_5 == 3'h6;
  assign _EVAL_204 = _EVAL_203 == 1'h0;
  assign _EVAL_179 = _EVAL_118 & _EVAL_204;
  assign _EVAL_96 = 4096'h1 << _EVAL_0;
  assign _EVAL_140 = _EVAL_179 ? _EVAL_96 : 4096'h0;
  assign _EVAL_75 = _EVAL_10 <= 3'h3;
  assign _EVAL_129 = _EVAL_75 | _EVAL_3;
  assign _EVAL_52 = _EVAL_129 == 1'h0;
  assign _EVAL_46 = _EVAL_2[0];
  assign _EVAL_131 = 2'h1 << _EVAL_46;
  assign _EVAL_51 = _EVAL_131 | 2'h1;
  assign _EVAL_49 = _EVAL_51[0];
  assign _EVAL_15 = _EVAL_1[1];
  assign _EVAL_178 = _EVAL_25 == 1'h0;
  assign _EVAL_133 = _EVAL_15 & _EVAL_178;
  assign _EVAL_73 = _EVAL_49 & _EVAL_133;
  assign _EVAL_214 = _EVAL_140[2335:0];
  assign _EVAL_121 = ~ _EVAL_214;
  assign _EVAL_149 = {1'b0,$signed(_EVAL_1)};
  assign _EVAL_45 = $signed(_EVAL_149) & $signed(-13'sh1000);
  assign _EVAL_142 = $signed(_EVAL_45);
  assign _EVAL_71 = $signed(_EVAL_142) == $signed(13'sh0);
  assign _EVAL_61 = _EVAL_3 == 1'h0;
  assign _EVAL_81 = 5'h3 << _EVAL_2;
  assign _EVAL_22 = _EVAL_81[1:0];
  assign _EVAL_66 = _EVAL_23 == 1'h0;
  assign _EVAL_145 = _EVAL_0 == _EVAL_177;
  assign _EVAL_198 = _EVAL_145 | _EVAL_3;
  assign _EVAL_137 = _EVAL_2 >= 2'h2;
  assign _EVAL_18 = _EVAL_51[1];
  assign _EVAL_176 = _EVAL_18 & _EVAL_15;
  assign _EVAL_220 = _EVAL_137 | _EVAL_176;
  assign _EVAL_31 = _EVAL_15 & _EVAL_25;
  assign _EVAL_148 = _EVAL_49 & _EVAL_31;
  assign _EVAL_17 = _EVAL_220 | _EVAL_148;
  assign _EVAL_180 = _EVAL_220 | _EVAL_73;
  assign _EVAL_92 = _EVAL_15 == 1'h0;
  assign _EVAL_182 = _EVAL_18 & _EVAL_92;
  assign _EVAL_172 = _EVAL_137 | _EVAL_182;
  assign _EVAL_173 = _EVAL_92 & _EVAL_25;
  assign _EVAL_190 = _EVAL_49 & _EVAL_173;
  assign _EVAL_225 = _EVAL_172 | _EVAL_190;
  assign _EVAL_216 = _EVAL_92 & _EVAL_178;
  assign _EVAL_192 = _EVAL_49 & _EVAL_216;
  assign _EVAL_189 = _EVAL_172 | _EVAL_192;
  assign _EVAL_37 = {_EVAL_17,_EVAL_180,_EVAL_225,_EVAL_189};
  assign _EVAL_89 = ~ _EVAL_37;
  assign _EVAL_114 = _EVAL_6 & _EVAL_89;
  assign _EVAL_67 = _EVAL_114 == 4'h0;
  assign _EVAL_105 = _EVAL_67 | _EVAL_3;
  assign _EVAL_127 = _EVAL == 1'h0;
  assign _EVAL_69 = _EVAL_127 | _EVAL_3;
  assign _EVAL_64 = _EVAL_5 <= 3'h6;
  assign _EVAL_44 = _EVAL_115 | _EVAL_187;
  assign _EVAL_157 = plusarg_reader_out == 32'h0;
  assign _EVAL_146 = _EVAL_112 | _EVAL_157;
  assign _EVAL_153 = _EVAL_144 < plusarg_reader_out;
  assign _EVAL_91 = _EVAL_146 | _EVAL_153;
  assign _EVAL_53 = _EVAL_5 == 3'h1;
  assign _EVAL_212 = _EVAL_14 == _EVAL_98;
  assign _EVAL_120 = _EVAL_1 == _EVAL_27;
  assign _EVAL_164 = _EVAL_120 | _EVAL_3;
  assign _EVAL_125 = _EVAL_8 == _EVAL_219;
  assign _EVAL_102 = _EVAL_125 | _EVAL_3;
  assign _EVAL_141 = _EVAL_102 == 1'h0;
  assign _EVAL_167 = _EVAL_23 - 1'h1;
  assign _EVAL_38 = _EVAL_8 == 3'h2;
  assign _EVAL_191 = _EVAL_9 & _EVAL_38;
  assign _EVAL_94 = _EVAL_10 <= 3'h4;
  assign _EVAL_100 = _EVAL_94 | _EVAL_3;
  assign _EVAL_101 = _EVAL_100 == 1'h0;
  assign _EVAL_147 = ~ _EVAL_22;
  assign _EVAL_207 = {{10'd0}, _EVAL_147};
  assign _EVAL_84 = _EVAL_1 & _EVAL_207;
  assign _EVAL_136 = _EVAL_11 & _EVAL_53;
  assign _EVAL_199 = _EVAL_2 <= 2'h2;
  assign _EVAL_78 = _EVAL_199 & _EVAL_71;
  assign _EVAL_21 = _EVAL_168 | _EVAL_3;
  assign _EVAL_34 = _EVAL_137 | _EVAL_3;
  assign _EVAL_184 = _EVAL_34 == 1'h0;
  assign _EVAL_130 = _EVAL_8 == 3'h6;
  assign _EVAL_183 = _EVAL_9 & _EVAL_130;
  assign _EVAL_29 = _EVAL_84 == 12'h0;
  assign _EVAL_155 = _EVAL_29 | _EVAL_3;
  assign _EVAL_223 = _EVAL_155 == 1'h0;
  assign _EVAL_32 = _EVAL_10 == _EVAL_74;
  assign _EVAL_83 = _EVAL_32 | _EVAL_3;
  assign _EVAL_231 = _EVAL_144 + 32'h1;
  assign _EVAL_185 = _EVAL_2 == _EVAL_188;
  assign _EVAL_109 = _EVAL_185 | _EVAL_3;
  assign _EVAL_95 = _EVAL_109 == 1'h0;
  assign _EVAL_171 = _EVAL_212 | _EVAL_3;
  assign _EVAL_211 = _EVAL_171 == 1'h0;
  assign _EVAL_161 = _EVAL_10 == 3'h0;
  assign _EVAL_106 = _EVAL_161 | _EVAL_3;
  assign _EVAL_206 = _EVAL_40 - 1'h1;
  assign _EVAL_60 = _EVAL_69 == 1'h0;
  assign _EVAL_80 = _EVAL_64 | _EVAL_3;
  assign _EVAL_117 = ~ _EVAL_6;
  assign _EVAL_122 = _EVAL_117 == 4'h0;
  assign _EVAL_181 = _EVAL_8 == 3'h4;
  assign _EVAL_19 = _EVAL_9 & _EVAL_181;
  assign _EVAL_41 = _EVAL_40 == 1'h0;
  assign _EVAL_85 = _EVAL_14 <= 12'h91f;
  assign _EVAL_165 = _EVAL_213 >> _EVAL_14;
  assign _EVAL_116 = _EVAL_165[0];
  assign _EVAL_229 = _EVAL_116 == 1'h0;
  assign _EVAL_68 = _EVAL_229 | _EVAL_3;
  assign _EVAL_39 = _EVAL_11 & _EVAL_158;
  assign _EVAL_215 = _EVAL_187 & _EVAL_66;
  assign _EVAL_143 = _EVAL_0 <= 12'h91f;
  assign _EVAL_196 = _EVAL_143 | _EVAL_3;
  assign _EVAL_217 = _EVAL_196 == 1'h0;
  assign _EVAL_70 = _EVAL_42 - 1'h1;
  assign _EVAL_108 = _EVAL_8 == 3'h5;
  assign _EVAL_119 = _EVAL_9 & _EVAL_108;
  assign _EVAL_208 = _EVAL_5 == _EVAL_209;
  assign _EVAL_62 = _EVAL_208 | _EVAL_3;
  assign _EVAL_103 = _EVAL_62 == 1'h0;
  assign _EVAL_56 = _EVAL_8 == 3'h7;
  assign _EVAL_24 = _EVAL_7 >= 2'h2;
  assign _EVAL_87 = _EVAL_24 | _EVAL_3;
  assign _EVAL_77 = _EVAL_115 & _EVAL_41;
  assign _EVAL_47 = _EVAL_10 != 3'h0;
  assign _EVAL_201 = _EVAL_47 | _EVAL_3;
  assign _EVAL_163 = _EVAL_11 & _EVAL_203;
  assign _EVAL_134 = _EVAL_8 == 3'h3;
  assign _EVAL_152 = _EVAL_6 == _EVAL_37;
  assign _EVAL_99 = _EVAL_152 | _EVAL_3;
  assign _EVAL_59 = _EVAL_122 | _EVAL_3;
  assign _EVAL_110 = _EVAL_83 == 1'h0;
  assign _EVAL_174 = _EVAL_66 == 1'h0;
  assign _EVAL_154 = _EVAL_99 == 1'h0;
  assign _EVAL_16 = _EVAL_85 | _EVAL_3;
  assign _EVAL_156 = _EVAL_9 & _EVAL_56;
  assign _EVAL_28 = _EVAL_91 | _EVAL_3;
  assign _EVAL_63 = _EVAL_59 == 1'h0;
  assign _EVAL_111 = _EVAL_9 & _EVAL_134;
  assign _EVAL_166 = _EVAL_7 == _EVAL_124;
  assign _EVAL_50 = _EVAL_213 | _EVAL_200;
  assign _EVAL_104 = _EVAL_8 == 3'h0;
  assign _EVAL_210 = _EVAL_9 & _EVAL_104;
  assign _EVAL_43 = _EVAL_21 == 1'h0;
  assign _EVAL_170 = _EVAL_5 == 3'h2;
  assign _EVAL_202 = _EVAL_201 == 1'h0;
  assign _EVAL_76 = _EVAL_8 == 3'h1;
  assign _EVAL_139 = _EVAL_78 | _EVAL_3;
  assign _EVAL_227 = _EVAL_139 == 1'h0;
  assign _EVAL_20 = _EVAL_55[0];
  assign _EVAL_126 = _EVAL_20 | _EVAL_3;
  assign _EVAL_226 = _EVAL_80 == 1'h0;
  assign _EVAL_169 = _EVAL_28 == 1'h0;
  assign _EVAL_33 = _EVAL_198 == 1'h0;
  assign _EVAL_65 = _EVAL_5 == 3'h4;
  assign _EVAL_138 = _EVAL_11 & _EVAL_65;
  assign _EVAL_222 = _EVAL_166 | _EVAL_3;
  assign _EVAL_132 = _EVAL_222 == 1'h0;
  assign _EVAL_72 = _EVAL_11 & _EVAL_170;
  assign _EVAL_82 = _EVAL_50 & _EVAL_121;
  assign _EVAL_221 = _EVAL_164 == 1'h0;
  assign _EVAL_224 = _EVAL_16 == 1'h0;
  assign _EVAL_123 = _EVAL_106 == 1'h0;
  assign _EVAL_93 = _EVAL_105 == 1'h0;
  assign _EVAL_97 = _EVAL_68 == 1'h0;
  assign _EVAL_193 = _EVAL_9 & _EVAL_76;
  assign _EVAL_218 = _EVAL_87 == 1'h0;
  assign _EVAL_197 = _EVAL_11 & _EVAL_174;
  assign _EVAL_54 = _EVAL_41 == 1'h0;
  assign _EVAL_90 = _EVAL_9 & _EVAL_54;
  assign _EVAL_57 = _EVAL_126 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_27 = _RAND_1[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_40 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_42 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_74 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_98 = _RAND_5[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_124 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_144 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_175 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_177 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_188 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_209 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {73{`RANDOM}};
  _EVAL_213 = _RAND_12[2335:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_219 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_13) begin
    if (_EVAL_3) begin
      _EVAL_23 <= 1'h0;
    end else begin
      if (_EVAL_187) begin
        if (_EVAL_66) begin
          _EVAL_23 <= 1'h0;
        end else begin
          _EVAL_23 <= _EVAL_167;
        end
      end
    end
    if (_EVAL_77) begin
      _EVAL_27 <= _EVAL_1;
    end
    if (_EVAL_3) begin
      _EVAL_40 <= 1'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_41) begin
          _EVAL_40 <= 1'h0;
        end else begin
          _EVAL_40 <= _EVAL_206;
        end
      end
    end
    if (_EVAL_3) begin
      _EVAL_42 <= 1'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_86) begin
          _EVAL_42 <= 1'h0;
        end else begin
          _EVAL_42 <= _EVAL_70;
        end
      end
    end
    if (_EVAL_77) begin
      _EVAL_74 <= _EVAL_10;
    end
    if (_EVAL_77) begin
      _EVAL_98 <= _EVAL_14;
    end
    if (_EVAL_215) begin
      _EVAL_124 <= _EVAL_7;
    end
    if (_EVAL_3) begin
      _EVAL_144 <= 32'h0;
    end else begin
      if (_EVAL_44) begin
        _EVAL_144 <= 32'h0;
      end else begin
        _EVAL_144 <= _EVAL_231;
      end
    end
    if (_EVAL_3) begin
      _EVAL_175 <= 1'h0;
    end else begin
      if (_EVAL_187) begin
        if (_EVAL_159) begin
          _EVAL_175 <= 1'h0;
        end else begin
          _EVAL_175 <= _EVAL_228;
        end
      end
    end
    if (_EVAL_215) begin
      _EVAL_177 <= _EVAL_0;
    end
    if (_EVAL_77) begin
      _EVAL_188 <= _EVAL_2;
    end
    if (_EVAL_215) begin
      _EVAL_209 <= _EVAL_5;
    end
    if (_EVAL_3) begin
      _EVAL_213 <= 2336'h0;
    end else begin
      _EVAL_213 <= _EVAL_82;
    end
    if (_EVAL_77) begin
      _EVAL_219 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0500a6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(350e94bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e21e7ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a5e8682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8902f94b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b68efc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2adc90da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bec2bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(556b5bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(543528c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd43300a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c0d67a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28449b2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f24868b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(722a65bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(164d03cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e56f84e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eab5cbe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e6a65f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad1ff5fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b8ec99a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0fd63ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36a55aab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8424d2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1aa36530)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13c71272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c4060dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2209cb86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9ad0eb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3a5c320)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47a22de4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a132b08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f31c22c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2def4a3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5fbdd3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11178b9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc09fcdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73ce5854)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd6c1ca5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef130519)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(504f9c62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41328d28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2209e09a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43a21e74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ec32d36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbb37c7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(249f8af7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c9d8ae5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a745eaf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4795f86c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1ac052a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b00f925)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ffe2d2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b0f16ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8cd18eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a56277cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec4a6e28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d9e6f32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cacf4a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f85e734)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a45c0b66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(682da4b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4872ac31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11a4a9fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e15da5b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb18ac90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f083a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11fc701b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e74ea0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35c7693f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c34f2626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
