//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_38(
  output        _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  output [63:0] _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  output [63:0] _EVAL_11,
  input         _EVAL_12,
  output [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input  [30:0] _EVAL_17,
  input  [6:0]  _EVAL_18,
  input  [63:0] _EVAL_19,
  output [2:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  input  [6:0]  _EVAL_24,
  output        _EVAL_25,
  input  [2:0]  _EVAL_26,
  input  [2:0]  _EVAL_27,
  output        _EVAL_28,
  input  [7:0]  _EVAL_29,
  output [6:0]  _EVAL_30,
  output [6:0]  _EVAL_31,
  input  [63:0] _EVAL_32,
  output [2:0]  _EVAL_33,
  output [30:0] _EVAL_34,
  output [2:0]  _EVAL_35,
  output [7:0]  _EVAL_36
);
  assign _EVAL_34 = _EVAL_17;
  assign _EVAL_3 = _EVAL_21;
  assign _EVAL_22 = _EVAL_5;
  assign _EVAL_15 = _EVAL_10;
  assign _EVAL_28 = _EVAL_2;
  assign _EVAL_31 = _EVAL_18;
  assign _EVAL_8 = _EVAL_19;
  assign _EVAL_9 = _EVAL_4;
  assign _EVAL = _EVAL_7;
  assign _EVAL_35 = _EVAL_26;
  assign _EVAL_36 = _EVAL_29;
  assign _EVAL_11 = _EVAL_32;
  assign _EVAL_25 = _EVAL_0;
  assign _EVAL_30 = _EVAL_24;
  assign _EVAL_33 = _EVAL_14;
  assign _EVAL_23 = _EVAL_16;
  assign _EVAL_13 = _EVAL_6;
  assign _EVAL_20 = _EVAL_27;
endmodule
