//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_183(
  input  [2:0]   _EVAL,
  input  [2:0]   _EVAL_0,
  input  [2:0]   _EVAL_1,
  input  [2:0]   _EVAL_2,
  input  [2:0]   _EVAL_3,
  input  [2:0]   _EVAL_4,
  input  [2:0]   _EVAL_5,
  input  [2:0]   _EVAL_6,
  input  [2:0]   _EVAL_7,
  input  [2:0]   _EVAL_8,
  input  [2:0]   _EVAL_9,
  input  [2:0]   _EVAL_10,
  input  [2:0]   _EVAL_11,
  input  [2:0]   _EVAL_12,
  input  [2:0]   _EVAL_13,
  input  [2:0]   _EVAL_14,
  input  [2:0]   _EVAL_15,
  input  [2:0]   _EVAL_16,
  input  [2:0]   _EVAL_17,
  input  [2:0]   _EVAL_18,
  input  [2:0]   _EVAL_19,
  input  [2:0]   _EVAL_20,
  input  [2:0]   _EVAL_21,
  input  [2:0]   _EVAL_22,
  input  [2:0]   _EVAL_23,
  input  [2:0]   _EVAL_24,
  input  [2:0]   _EVAL_25,
  input  [2:0]   _EVAL_26,
  input  [2:0]   _EVAL_27,
  input  [2:0]   _EVAL_28,
  input  [2:0]   _EVAL_29,
  input  [2:0]   _EVAL_30,
  input  [2:0]   _EVAL_31,
  output [2:0]   _EVAL_32,
  input  [2:0]   _EVAL_33,
  input  [2:0]   _EVAL_34,
  input  [2:0]   _EVAL_35,
  output [6:0]   _EVAL_36,
  input  [2:0]   _EVAL_37,
  input  [2:0]   _EVAL_38,
  input  [2:0]   _EVAL_39,
  input  [2:0]   _EVAL_40,
  input  [2:0]   _EVAL_41,
  input  [2:0]   _EVAL_42,
  input  [2:0]   _EVAL_43,
  input  [2:0]   _EVAL_44,
  input  [2:0]   _EVAL_45,
  input  [2:0]   _EVAL_46,
  input  [2:0]   _EVAL_47,
  input  [2:0]   _EVAL_48,
  input  [2:0]   _EVAL_49,
  input  [2:0]   _EVAL_50,
  input  [2:0]   _EVAL_51,
  input  [2:0]   _EVAL_52,
  input  [2:0]   _EVAL_53,
  input  [2:0]   _EVAL_54,
  input  [2:0]   _EVAL_55,
  input  [2:0]   _EVAL_56,
  input  [2:0]   _EVAL_57,
  input  [2:0]   _EVAL_58,
  input  [2:0]   _EVAL_59,
  input  [2:0]   _EVAL_60,
  input  [2:0]   _EVAL_61,
  input  [2:0]   _EVAL_62,
  input  [2:0]   _EVAL_63,
  input  [2:0]   _EVAL_64,
  input  [2:0]   _EVAL_65,
  input  [2:0]   _EVAL_66,
  input  [2:0]   _EVAL_67,
  input  [2:0]   _EVAL_68,
  input  [2:0]   _EVAL_69,
  input  [2:0]   _EVAL_70,
  input  [2:0]   _EVAL_71,
  input  [2:0]   _EVAL_72,
  input  [2:0]   _EVAL_73,
  input  [2:0]   _EVAL_74,
  input  [2:0]   _EVAL_75,
  input  [2:0]   _EVAL_76,
  input  [2:0]   _EVAL_77,
  input  [2:0]   _EVAL_78,
  input  [2:0]   _EVAL_79,
  input  [2:0]   _EVAL_80,
  input  [2:0]   _EVAL_81,
  input  [2:0]   _EVAL_82,
  input  [2:0]   _EVAL_83,
  input  [2:0]   _EVAL_84,
  input  [2:0]   _EVAL_85,
  input  [2:0]   _EVAL_86,
  input  [2:0]   _EVAL_87,
  input  [2:0]   _EVAL_88,
  input  [2:0]   _EVAL_89,
  input  [2:0]   _EVAL_90,
  input  [2:0]   _EVAL_91,
  input  [2:0]   _EVAL_92,
  input  [2:0]   _EVAL_93,
  input  [2:0]   _EVAL_94,
  input  [2:0]   _EVAL_95,
  input  [2:0]   _EVAL_96,
  input  [2:0]   _EVAL_97,
  input  [2:0]   _EVAL_98,
  input  [2:0]   _EVAL_99,
  input  [2:0]   _EVAL_100,
  input  [2:0]   _EVAL_101,
  input  [2:0]   _EVAL_102,
  input  [2:0]   _EVAL_103,
  input  [2:0]   _EVAL_104,
  input  [2:0]   _EVAL_105,
  input  [2:0]   _EVAL_106,
  input  [2:0]   _EVAL_107,
  input  [2:0]   _EVAL_108,
  input  [2:0]   _EVAL_109,
  input  [2:0]   _EVAL_110,
  input  [2:0]   _EVAL_111,
  input  [2:0]   _EVAL_112,
  input  [126:0] _EVAL_113,
  input  [2:0]   _EVAL_114,
  input  [2:0]   _EVAL_115,
  input  [2:0]   _EVAL_116,
  input  [2:0]   _EVAL_117,
  input  [2:0]   _EVAL_118,
  input  [2:0]   _EVAL_119,
  input  [2:0]   _EVAL_120,
  input  [2:0]   _EVAL_121,
  input  [2:0]   _EVAL_122,
  input  [2:0]   _EVAL_123,
  input  [2:0]   _EVAL_124,
  input  [2:0]   _EVAL_125,
  input  [2:0]   _EVAL_126,
  input  [2:0]   _EVAL_127,
  input  [2:0]   _EVAL_128
);
  wire  _EVAL_595;
  wire [3:0] _EVAL_239;
  wire  _EVAL_641;
  wire [3:0] _EVAL_761;
  wire  _EVAL_862;
  wire [3:0] _EVAL_511;
  wire  _EVAL_887;
  wire [3:0] _EVAL_392;
  wire  _EVAL_203;
  wire [3:0] _EVAL_244;
  wire  _EVAL_770;
  wire [3:0] _EVAL_803;
  wire  _EVAL_702;
  wire [3:0] _EVAL_478;
  wire  _EVAL_578;
  wire [3:0] _EVAL_414;
  wire  _EVAL_886;
  wire [3:0] _EVAL_746;
  wire  _EVAL_876;
  wire [3:0] _EVAL_168;
  wire  _EVAL_514;
  wire [3:0] _EVAL_472;
  wire  _EVAL_583;
  wire [3:0] _EVAL_683;
  wire  _EVAL_192;
  wire [3:0] _EVAL_644;
  wire  _EVAL_436;
  wire [3:0] _EVAL_417;
  wire  _EVAL_486;
  wire [3:0] _EVAL_512;
  wire  _EVAL_362;
  wire [3:0] _EVAL_291;
  wire  _EVAL_539;
  wire [3:0] _EVAL_846;
  wire  _EVAL_611;
  wire [3:0] _EVAL_550;
  wire  _EVAL_198;
  wire [3:0] _EVAL_532;
  wire  _EVAL_302;
  wire [3:0] _EVAL_603;
  wire  _EVAL_468;
  wire [3:0] _EVAL_357;
  wire  _EVAL_735;
  wire [3:0] _EVAL_254;
  wire  _EVAL_855;
  wire [3:0] _EVAL_623;
  wire  _EVAL_555;
  wire [3:0] _EVAL_422;
  wire  _EVAL_758;
  wire [3:0] _EVAL_285;
  wire  _EVAL_545;
  wire [3:0] _EVAL_176;
  wire  _EVAL_666;
  wire [3:0] _EVAL_783;
  wire  _EVAL_481;
  wire [3:0] _EVAL_804;
  wire  _EVAL_820;
  wire [3:0] _EVAL_155;
  wire  _EVAL_231;
  wire [3:0] _EVAL_174;
  wire  _EVAL_727;
  wire [3:0] _EVAL_279;
  wire  _EVAL_187;
  wire [3:0] _EVAL_661;
  wire  _EVAL_301;
  wire  _EVAL_719;
  wire  _EVAL_536;
  wire [1:0] _EVAL_413;
  wire [1:0] _EVAL_567;
  wire [1:0] _EVAL_425;
  wire  _EVAL_213;
  wire [3:0] _EVAL_226;
  wire  _EVAL_299;
  wire [3:0] _EVAL_824;
  wire  _EVAL_869;
  wire [3:0] _EVAL_600;
  wire  _EVAL_310;
  wire [3:0] _EVAL_858;
  wire  _EVAL_796;
  wire [3:0] _EVAL_768;
  wire  _EVAL_703;
  wire [3:0] _EVAL_816;
  wire  _EVAL_397;
  wire  _EVAL_565;
  wire  _EVAL_247;
  wire [1:0] _EVAL_637;
  wire [1:0] _EVAL_160;
  wire [1:0] _EVAL_456;
  wire [2:0] _EVAL_151;
  wire  _EVAL_479;
  wire [3:0] _EVAL_712;
  wire  _EVAL_474;
  wire [3:0] _EVAL_706;
  wire  _EVAL_276;
  wire [3:0] _EVAL_501;
  wire  _EVAL_388;
  wire [3:0] _EVAL_724;
  wire  _EVAL_663;
  wire [3:0] _EVAL_533;
  wire  _EVAL_138;
  wire [3:0] _EVAL_483;
  wire  _EVAL_769;
  wire  _EVAL_619;
  wire [3:0] _EVAL_186;
  wire  _EVAL_348;
  wire [3:0] _EVAL_453;
  wire  _EVAL_500;
  wire [3:0] _EVAL_658;
  wire  _EVAL_609;
  wire [3:0] _EVAL_189;
  wire  _EVAL_597;
  wire [3:0] _EVAL_431;
  wire  _EVAL_224;
  wire [3:0] _EVAL_502;
  wire  _EVAL_647;
  wire [3:0] _EVAL_811;
  wire  _EVAL_343;
  wire [3:0] _EVAL_743;
  wire  _EVAL_146;
  wire [3:0] _EVAL_269;
  wire  _EVAL_467;
  wire [3:0] _EVAL_778;
  wire  _EVAL_751;
  wire [3:0] _EVAL_656;
  wire  _EVAL_335;
  wire [3:0] _EVAL_371;
  wire  _EVAL_212;
  wire [3:0] _EVAL_234;
  wire  _EVAL_708;
  wire [3:0] _EVAL_544;
  wire  _EVAL_535;
  wire  _EVAL_797;
  wire  _EVAL_713;
  wire [1:0] _EVAL_361;
  wire [1:0] _EVAL_204;
  wire [1:0] _EVAL_831;
  wire  _EVAL_798;
  wire  _EVAL_643;
  wire [1:0] _EVAL_323;
  wire [1:0] _EVAL_332;
  wire [1:0] _EVAL_372;
  wire [2:0] _EVAL_739;
  wire [2:0] _EVAL_626;
  wire [2:0] _EVAL_268;
  wire [3:0] _EVAL_284;
  wire  _EVAL_885;
  wire  _EVAL_809;
  wire [3:0] _EVAL_772;
  wire  _EVAL_274;
  wire [3:0] _EVAL_795;
  wire  _EVAL_172;
  wire [3:0] _EVAL_214;
  wire  _EVAL_494;
  wire [3:0] _EVAL_196;
  wire  _EVAL_396;
  wire [3:0] _EVAL_330;
  wire  _EVAL_318;
  wire [3:0] _EVAL_185;
  wire  _EVAL_843;
  wire [3:0] _EVAL_492;
  wire  _EVAL_732;
  wire [3:0] _EVAL_766;
  wire  _EVAL_616;
  wire [3:0] _EVAL_817;
  wire  _EVAL_564;
  wire [3:0] _EVAL_376;
  wire  _EVAL_438;
  wire [3:0] _EVAL_834;
  wire  _EVAL_257;
  wire [3:0] _EVAL_308;
  wire  _EVAL_137;
  wire [3:0] _EVAL_334;
  wire  _EVAL_744;
  wire  _EVAL_638;
  wire  _EVAL_823;
  wire [1:0] _EVAL_333;
  wire [1:0] _EVAL_684;
  wire [1:0] _EVAL_345;
  wire [2:0] _EVAL_615;
  wire [2:0] _EVAL_734;
  wire  _EVAL_755;
  wire [1:0] _EVAL_290;
  wire  _EVAL_577;
  wire [3:0] _EVAL_219;
  wire  _EVAL_738;
  wire [3:0] _EVAL_470;
  wire  _EVAL_875;
  wire  _EVAL_295;
  wire  _EVAL_840;
  wire [3:0] _EVAL_252;
  wire  _EVAL_729;
  wire [3:0] _EVAL_551;
  wire  _EVAL_801;
  wire [3:0] _EVAL_691;
  wire  _EVAL_460;
  wire [3:0] _EVAL_628;
  wire  _EVAL_433;
  wire [3:0] _EVAL_519;
  wire  _EVAL_608;
  wire [3:0] _EVAL_429;
  wire  _EVAL_584;
  wire [3:0] _EVAL_721;
  wire  _EVAL_272;
  wire [3:0] _EVAL_657;
  wire  _EVAL_704;
  wire [3:0] _EVAL_542;
  wire  _EVAL_588;
  wire [3:0] _EVAL_748;
  wire  _EVAL_182;
  wire [3:0] _EVAL_711;
  wire [3:0] _EVAL_221;
  wire  _EVAL_354;
  wire [3:0] _EVAL_307;
  wire  _EVAL_461;
  wire [3:0] _EVAL_750;
  wire  _EVAL_418;
  wire [3:0] _EVAL_482;
  wire  _EVAL_861;
  wire [3:0] _EVAL_731;
  wire  _EVAL_440;
  wire [3:0] _EVAL_140;
  wire  _EVAL_621;
  wire [3:0] _EVAL_863;
  wire  _EVAL_159;
  wire [3:0] _EVAL_312;
  wire  _EVAL_589;
  wire [3:0] _EVAL_304;
  wire  _EVAL_510;
  wire [3:0] _EVAL_437;
  wire  _EVAL_405;
  wire [3:0] _EVAL_315;
  wire  _EVAL_767;
  wire [3:0] _EVAL_813;
  wire  _EVAL_685;
  wire [3:0] _EVAL_195;
  wire  _EVAL_635;
  wire [3:0] _EVAL_166;
  wire  _EVAL_380;
  wire [3:0] _EVAL_705;
  wire  _EVAL_747;
  wire [3:0] _EVAL_549;
  wire [3:0] _EVAL_722;
  wire  _EVAL_201;
  wire [3:0] _EVAL_518;
  wire  _EVAL_849;
  wire [3:0] _EVAL_144;
  wire  _EVAL_242;
  wire [3:0] _EVAL_851;
  wire [3:0] _EVAL_391;
  wire  _EVAL_799;
  wire [3:0] _EVAL_507;
  wire  _EVAL_505;
  wire [3:0] _EVAL_826;
  wire  _EVAL_350;
  wire [3:0] _EVAL_618;
  wire  _EVAL_401;
  wire [3:0] _EVAL_864;
  wire  _EVAL_452;
  wire [3:0] _EVAL_415;
  wire  _EVAL_590;
  wire [3:0] _EVAL_802;
  wire [3:0] _EVAL_668;
  wire  _EVAL_416;
  wire [3:0] _EVAL_856;
  wire  _EVAL_464;
  wire [3:0] _EVAL_614;
  wire  _EVAL_419;
  wire [3:0] _EVAL_873;
  wire  _EVAL_435;
  wire [3:0] _EVAL_650;
  wire  _EVAL_591;
  wire [3:0] _EVAL_206;
  wire  _EVAL_374;
  wire  _EVAL_726;
  wire [3:0] _EVAL_692;
  wire  _EVAL_136;
  wire [3:0] _EVAL_161;
  wire  _EVAL_366;
  wire  _EVAL_541;
  wire [3:0] _EVAL_181;
  wire  _EVAL_884;
  wire [3:0] _EVAL_728;
  wire  _EVAL_717;
  wire [3:0] _EVAL_844;
  wire  _EVAL_485;
  wire [3:0] _EVAL_303;
  wire  _EVAL_612;
  wire [3:0] _EVAL_516;
  wire  _EVAL_720;
  wire [3:0] _EVAL_458;
  wire  _EVAL_130;
  wire [3:0] _EVAL_378;
  wire  _EVAL_465;
  wire  _EVAL_496;
  wire [3:0] _EVAL_693;
  wire  _EVAL_853;
  wire [3:0] _EVAL_359;
  wire  _EVAL_207;
  wire  _EVAL_249;
  wire [1:0] _EVAL_367;
  wire [1:0] _EVAL_232;
  wire  _EVAL_349;
  wire [3:0] _EVAL_227;
  wire  _EVAL_527;
  wire [3:0] _EVAL_636;
  wire  _EVAL_449;
  wire  _EVAL_819;
  wire [1:0] _EVAL_548;
  wire  _EVAL_753;
  wire [3:0] _EVAL_558;
  wire  _EVAL_593;
  wire [3:0] _EVAL_373;
  wire  _EVAL_845;
  wire  _EVAL_408;
  wire  _EVAL_287;
  wire [3:0] _EVAL_278;
  wire  _EVAL_789;
  wire [3:0] _EVAL_356;
  wire  _EVAL_723;
  wire [3:0] _EVAL_673;
  wire  _EVAL_205;
  wire [3:0] _EVAL_211;
  wire  _EVAL_807;
  wire [3:0] _EVAL_531;
  wire  _EVAL_877;
  wire [3:0] _EVAL_521;
  wire  _EVAL_792;
  wire [3:0] _EVAL_286;
  wire  _EVAL_439;
  wire  _EVAL_363;
  wire [1:0] _EVAL_605;
  wire [1:0] _EVAL_170;
  wire [1:0] _EVAL_407;
  wire  _EVAL_522;
  wire [3:0] _EVAL_382;
  wire  _EVAL_183;
  wire [3:0] _EVAL_336;
  wire  _EVAL_830;
  wire [1:0] _EVAL_774;
  wire [1:0] _EVAL_471;
  wire  _EVAL_157;
  wire  _EVAL_175;
  wire [3:0] _EVAL_760;
  wire  _EVAL_594;
  wire [3:0] _EVAL_457;
  wire  _EVAL_640;
  wire  _EVAL_338;
  wire [3:0] _EVAL_570;
  wire  _EVAL_282;
  wire [3:0] _EVAL_553;
  wire  _EVAL_675;
  wire [3:0] _EVAL_859;
  wire  _EVAL_569;
  wire [3:0] _EVAL_520;
  wire [3:0] _EVAL_523;
  wire  _EVAL_848;
  wire [3:0] _EVAL_572;
  wire  _EVAL_718;
  wire [3:0] _EVAL_534;
  wire  _EVAL_169;
  wire [3:0] _EVAL_665;
  wire  _EVAL_543;
  wire [3:0] _EVAL_385;
  wire  _EVAL_484;
  wire [3:0] _EVAL_678;
  wire [3:0] _EVAL_446;
  wire  _EVAL_686;
  wire [3:0] _EVAL_375;
  wire  _EVAL_765;
  wire  _EVAL_699;
  wire  _EVAL_725;
  wire [1:0] _EVAL_629;
  wire [1:0] _EVAL_624;
  wire [1:0] _EVAL_800;
  wire  _EVAL_681;
  wire [1:0] _EVAL_208;
  wire [2:0] _EVAL_489;
  wire [2:0] _EVAL_561;
  wire [2:0] _EVAL_131;
  wire [3:0] _EVAL_781;
  wire  _EVAL_360;
  wire [3:0] _EVAL_680;
  wire  _EVAL_230;
  wire [3:0] _EVAL_676;
  wire  _EVAL_381;
  wire  _EVAL_707;
  wire  _EVAL_222;
  wire [3:0] _EVAL_164;
  wire  _EVAL_347;
  wire [3:0] _EVAL_495;
  wire  _EVAL_216;
  wire [3:0] _EVAL_390;
  wire  _EVAL_808;
  wire [3:0] _EVAL_370;
  wire  _EVAL_810;
  wire [3:0] _EVAL_313;
  wire  _EVAL_412;
  wire [3:0] _EVAL_342;
  wire  _EVAL_253;
  wire [3:0] _EVAL_364;
  wire [3:0] _EVAL_402;
  wire  _EVAL_822;
  wire [3:0] _EVAL_424;
  wire  _EVAL_135;
  wire [3:0] _EVAL_794;
  wire  _EVAL_710;
  wire [3:0] _EVAL_818;
  wire  _EVAL_190;
  wire [3:0] _EVAL_870;
  wire  _EVAL_630;
  wire  _EVAL_837;
  wire  _EVAL_610;
  wire [1:0] _EVAL_141;
  wire [1:0] _EVAL_672;
  wire [1:0] _EVAL_358;
  wire  _EVAL_627;
  wire  _EVAL_236;
  wire [1:0] _EVAL_517;
  wire [1:0] _EVAL_223;
  wire [1:0] _EVAL_503;
  wire [2:0] _EVAL_814;
  wire [2:0] _EVAL_882;
  wire [2:0] _EVAL_754;
  wire [3:0] _EVAL_445;
  wire  _EVAL_733;
  wire [3:0] _EVAL_574;
  wire  _EVAL_776;
  wire [3:0] _EVAL_184;
  wire  _EVAL_283;
  wire [3:0] _EVAL_607;
  wire  _EVAL_188;
  wire [3:0] _EVAL_229;
  wire  _EVAL_759;
  wire [3:0] _EVAL_689;
  wire  _EVAL_568;
  wire [3:0] _EVAL_156;
  wire  _EVAL_653;
  wire  _EVAL_506;
  wire  _EVAL_669;
  wire [1:0] _EVAL_162;
  wire [1:0] _EVAL_455;
  wire [1:0] _EVAL_697;
  wire [2:0] _EVAL_632;
  wire  _EVAL_339;
  wire [3:0] _EVAL_173;
  wire  _EVAL_745;
  wire [3:0] _EVAL_690;
  wire  _EVAL_426;
  wire [3:0] _EVAL_762;
  wire  _EVAL_275;
  wire [3:0] _EVAL_880;
  wire  _EVAL_280;
  wire [3:0] _EVAL_200;
  wire  _EVAL_322;
  wire [3:0] _EVAL_298;
  wire  _EVAL_599;
  wire [3:0] _EVAL_134;
  wire  _EVAL_580;
  wire [3:0] _EVAL_601;
  wire [3:0] _EVAL_294;
  wire  _EVAL_777;
  wire [3:0] _EVAL_659;
  wire  _EVAL_617;
  wire [3:0] _EVAL_827;
  wire  _EVAL_582;
  wire [3:0] _EVAL_368;
  wire  _EVAL_441;
  wire [3:0] _EVAL_444;
  wire  _EVAL_639;
  wire  _EVAL_488;
  wire  _EVAL_649;
  wire [1:0] _EVAL_490;
  wire [1:0] _EVAL_327;
  wire [1:0] _EVAL_874;
  wire  _EVAL_326;
  wire  _EVAL_825;
  wire [1:0] _EVAL_145;
  wire [1:0] _EVAL_821;
  wire [1:0] _EVAL_317;
  wire [2:0] _EVAL_592;
  wire [2:0] _EVAL_694;
  wire [2:0] _EVAL_409;
  wire [3:0] _EVAL_238;
  wire [3:0] _EVAL_805;
  wire  _EVAL_682;
  wire  _EVAL_386;
  wire [1:0] _EVAL_566;
  wire  _EVAL_475;
  wire [3:0] _EVAL_540;
  wire  _EVAL_153;
  wire [3:0] _EVAL_379;
  wire  _EVAL_251;
  wire [3:0] _EVAL_293;
  wire [3:0] _EVAL_421;
  wire  _EVAL_749;
  wire  _EVAL_258;
  wire [3:0] _EVAL_480;
  wire [3:0] _EVAL_191;
  wire  _EVAL_604;
  wire  _EVAL_847;
  wire [1:0] _EVAL_316;
  wire [1:0] _EVAL_526;
  wire  _EVAL_218;
  wire [1:0] _EVAL_714;
  wire  _EVAL_560;
  wire [3:0] _EVAL_281;
  wire  _EVAL_812;
  wire [3:0] _EVAL_448;
  wire  _EVAL_833;
  wire [3:0] _EVAL_498;
  wire  _EVAL_842;
  wire [1:0] _EVAL_394;
  wire [1:0] _EVAL_554;
  wire  _EVAL_319;
  wire  _EVAL_642;
  wire [1:0] _EVAL_233;
  wire [1:0] _EVAL_670;
  wire [1:0] _EVAL_340;
  wire [2:0] _EVAL_152;
  wire [2:0] _EVAL_194;
  wire [2:0] _EVAL_865;
  wire [3:0] _EVAL_756;
  wire [3:0] _EVAL_557;
  wire [3:0] _EVAL_406;
  wire  _EVAL_255;
  wire [3:0] _EVAL_598;
  wire [3:0] _EVAL_868;
  wire [3:0] _EVAL_369;
  wire  _EVAL_351;
  wire [3:0] _EVAL_147;
  wire [3:0] _EVAL_645;
  wire  _EVAL_305;
  wire [3:0] _EVAL_587;
  wire  _EVAL_337;
  wire [3:0] _EVAL_149;
  wire [3:0] _EVAL_881;
  wire [1:0] _EVAL_210;
  wire  _EVAL_736;
  wire  _EVAL_353;
  wire [3:0] _EVAL_384;
  wire  _EVAL_871;
  wire [3:0] _EVAL_241;
  wire  _EVAL_377;
  wire [3:0] _EVAL_434;
  wire [3:0] _EVAL_259;
  wire  _EVAL_698;
  wire [3:0] _EVAL_508;
  wire  _EVAL_466;
  wire [3:0] _EVAL_243;
  wire  _EVAL_423;
  wire [3:0] _EVAL_139;
  wire  _EVAL_428;
  wire [3:0] _EVAL_306;
  wire [3:0] _EVAL_791;
  wire  _EVAL_784;
  wire [3:0] _EVAL_606;
  wire  _EVAL_193;
  wire [3:0] _EVAL_651;
  wire  _EVAL_404;
  wire [3:0] _EVAL_576;
  wire  _EVAL_430;
  wire [1:0] _EVAL_835;
  wire [1:0] _EVAL_631;
  wire [1:0] _EVAL_742;
  wire  _EVAL_829;
  wire  _EVAL_432;
  wire [1:0] _EVAL_447;
  wire [1:0] _EVAL_469;
  wire [1:0] _EVAL_709;
  wire [2:0] _EVAL_158;
  wire [2:0] _EVAL_395;
  wire [2:0] _EVAL_477;
  wire [3:0] _EVAL_493;
  wire  _EVAL_142;
  wire [3:0] _EVAL_537;
  wire  _EVAL_410;
  wire [3:0] _EVAL_786;
  wire  _EVAL_248;
  wire  _EVAL_393;
  wire [3:0] _EVAL_559;
  wire  _EVAL_646;
  wire [3:0] _EVAL_546;
  wire  _EVAL_552;
  wire [3:0] _EVAL_562;
  wire [3:0] _EVAL_165;
  wire  _EVAL_365;
  wire [3:0] _EVAL_613;
  wire  _EVAL_220;
  wire [3:0] _EVAL_513;
  wire  _EVAL_491;
  wire [3:0] _EVAL_883;
  wire [3:0] _EVAL_538;
  wire  _EVAL_509;
  wire [3:0] _EVAL_267;
  wire [3:0] _EVAL_443;
  wire  _EVAL_459;
  wire [3:0] _EVAL_741;
  wire [3:0] _EVAL_237;
  wire  _EVAL_266;
  wire [3:0] _EVAL_524;
  wire  _EVAL_217;
  wire [3:0] _EVAL_177;
  wire [3:0] _EVAL_771;
  wire  _EVAL_163;
  wire [3:0] _EVAL_815;
  wire [3:0] _EVAL_806;
  wire  _EVAL_775;
  wire [3:0] _EVAL_579;
  wire  _EVAL_178;
  wire [3:0] _EVAL_715;
  wire  _EVAL_752;
  wire [3:0] _EVAL_264;
  wire  _EVAL_504;
  wire [3:0] _EVAL_850;
  wire [3:0] _EVAL_150;
  wire  _EVAL_399;
  wire [3:0] _EVAL_225;
  wire  _EVAL_344;
  wire [3:0] _EVAL_320;
  wire  _EVAL_857;
  wire [3:0] _EVAL_648;
  wire [3:0] _EVAL_620;
  wire  _EVAL_154;
  wire [3:0] _EVAL_660;
  wire  _EVAL_581;
  wire [3:0] _EVAL_737;
  wire  _EVAL_695;
  wire [3:0] _EVAL_528;
  wire  _EVAL_260;
  wire  _EVAL_171;
  wire [1:0] _EVAL_785;
  wire  _EVAL_625;
  wire  _EVAL_787;
  wire [1:0] _EVAL_270;
  wire [1:0] _EVAL_228;
  wire [1:0] _EVAL_838;
  wire [2:0] _EVAL_790;
  wire [2:0] _EVAL_573;
  wire [2:0] _EVAL_389;
  wire [3:0] _EVAL_398;
  wire [3:0] _EVAL_586;
  wire [2:0] _EVAL_454;
  wire [2:0] _EVAL_383;
  wire [3:0] _EVAL_263;
  wire [3:0] _EVAL_209;
  wire [4:0] _EVAL_314;
  wire [4:0] _EVAL_215;
  wire [4:0] _EVAL_297;
  wire  _EVAL_701;
  wire  _EVAL_476;
  wire [1:0] _EVAL_289;
  wire [1:0] _EVAL_256;
  wire [1:0] _EVAL_324;
  wire  _EVAL_841;
  wire  _EVAL_879;
  wire [1:0] _EVAL_547;
  wire [1:0] _EVAL_866;
  wire [1:0] _EVAL_730;
  wire [2:0] _EVAL_296;
  wire [2:0] _EVAL_411;
  wire [2:0] _EVAL_129;
  wire [3:0] _EVAL_167;
  wire  _EVAL_288;
  wire  _EVAL_652;
  wire [1:0] _EVAL_878;
  wire [1:0] _EVAL_860;
  wire [1:0] _EVAL_355;
  wire  _EVAL_199;
  wire  _EVAL_245;
  wire [1:0] _EVAL_265;
  wire [1:0] _EVAL_832;
  wire [1:0] _EVAL_442;
  wire [2:0] _EVAL_262;
  wire [2:0] _EVAL_667;
  wire [2:0] _EVAL_180;
  wire  _EVAL_292;
  wire  _EVAL_328;
  wire [1:0] _EVAL_773;
  wire [1:0] _EVAL_836;
  wire [1:0] _EVAL_311;
  wire  _EVAL_387;
  wire [1:0] _EVAL_487;
  wire [2:0] _EVAL_240;
  wire [2:0] _EVAL_451;
  wire [2:0] _EVAL_329;
  wire [3:0] _EVAL_757;
  wire [3:0] _EVAL_346;
  wire [3:0] _EVAL_674;
  wire [4:0] _EVAL_246;
  wire [4:0] _EVAL_664;
  wire [4:0] _EVAL_450;
  wire [5:0] _EVAL_852;
  wire [5:0] _EVAL_321;
  wire [5:0] _EVAL_197;
  wire [6:0] _EVAL_872;
  wire [6:0] _EVAL_716;
  wire  _EVAL_679;
  wire  _EVAL_497;
  wire [1:0] _EVAL_602;
  wire [1:0] _EVAL_427;
  wire [1:0] _EVAL_400;
  wire  _EVAL_261;
  wire  _EVAL_499;
  wire [1:0] _EVAL_525;
  wire [1:0] _EVAL_331;
  wire [1:0] _EVAL_854;
  wire [2:0] _EVAL_839;
  wire [2:0] _EVAL_341;
  wire [2:0] _EVAL_688;
  wire [3:0] _EVAL_596;
  wire  _EVAL_700;
  wire [1:0] _EVAL_634;
  wire [1:0] _EVAL_788;
  wire  _EVAL_740;
  wire  _EVAL_132;
  wire [1:0] _EVAL_529;
  wire [1:0] _EVAL_780;
  wire [1:0] _EVAL_654;
  wire [2:0] _EVAL_133;
  wire [2:0] _EVAL_782;
  wire [2:0] _EVAL_571;
  wire [3:0] _EVAL_622;
  wire [3:0] _EVAL_202;
  wire  _EVAL_655;
  wire  _EVAL_463;
  wire [1:0] _EVAL_763;
  wire [1:0] _EVAL_696;
  wire [1:0] _EVAL_352;
  wire  _EVAL_530;
  wire [1:0] _EVAL_277;
  wire [1:0] _EVAL_273;
  wire [2:0] _EVAL_179;
  wire [2:0] _EVAL_687;
  wire [2:0] _EVAL_779;
  wire [3:0] _EVAL_473;
  wire [3:0] _EVAL_677;
  wire [4:0] _EVAL_793;
  wire [4:0] _EVAL_515;
  wire [4:0] _EVAL_271;
  wire [5:0] _EVAL_309;
  wire [5:0] _EVAL_462;
  wire  _EVAL_828;
  wire [1:0] _EVAL_867;
  wire [3:0] _EVAL_671;
  wire  _EVAL_585;
  wire [3:0] _EVAL_420;
  wire [3:0] _EVAL_148;
  wire  _EVAL_633;
  wire [2:0] _EVAL_662;
  wire [3:0] _EVAL_300;
  wire [3:0] _EVAL_888;
  wire [2:0] _EVAL_556;
  wire [2:0] _EVAL_403;
  wire [3:0] _EVAL_143;
  wire [3:0] _EVAL_575;
  wire [4:0] _EVAL_563;
  wire [4:0] _EVAL_764;
  wire [4:0] _EVAL_325;
  wire [5:0] _EVAL_235;
  wire [3:0] _EVAL_250;
  assign _EVAL_595 = _EVAL_113[87];
  assign _EVAL_239 = {_EVAL_595,_EVAL_39};
  assign _EVAL_641 = _EVAL_113[88];
  assign _EVAL_761 = {_EVAL_641,_EVAL_120};
  assign _EVAL_862 = _EVAL_239 >= _EVAL_761;
  assign _EVAL_511 = _EVAL_862 ? _EVAL_239 : _EVAL_761;
  assign _EVAL_887 = _EVAL_113[89];
  assign _EVAL_392 = {_EVAL_887,_EVAL_23};
  assign _EVAL_203 = _EVAL_113[90];
  assign _EVAL_244 = {_EVAL_203,_EVAL_92};
  assign _EVAL_770 = _EVAL_392 >= _EVAL_244;
  assign _EVAL_803 = _EVAL_770 ? _EVAL_392 : _EVAL_244;
  assign _EVAL_702 = _EVAL_511 >= _EVAL_803;
  assign _EVAL_478 = _EVAL_702 ? _EVAL_511 : _EVAL_803;
  assign _EVAL_578 = _EVAL_113[91];
  assign _EVAL_414 = {_EVAL_578,_EVAL_27};
  assign _EVAL_886 = _EVAL_113[92];
  assign _EVAL_746 = {_EVAL_886,_EVAL_91};
  assign _EVAL_876 = _EVAL_414 >= _EVAL_746;
  assign _EVAL_168 = _EVAL_876 ? _EVAL_414 : _EVAL_746;
  assign _EVAL_514 = _EVAL_113[93];
  assign _EVAL_472 = {_EVAL_514,_EVAL_75};
  assign _EVAL_583 = _EVAL_113[94];
  assign _EVAL_683 = {_EVAL_583,_EVAL_53};
  assign _EVAL_192 = _EVAL_472 >= _EVAL_683;
  assign _EVAL_644 = _EVAL_192 ? _EVAL_472 : _EVAL_683;
  assign _EVAL_436 = _EVAL_168 >= _EVAL_644;
  assign _EVAL_417 = _EVAL_436 ? _EVAL_168 : _EVAL_644;
  assign _EVAL_486 = _EVAL_478 >= _EVAL_417;
  assign _EVAL_512 = _EVAL_486 ? _EVAL_478 : _EVAL_417;
  assign _EVAL_362 = _EVAL_113[39];
  assign _EVAL_291 = {_EVAL_362,_EVAL_124};
  assign _EVAL_539 = _EVAL_113[40];
  assign _EVAL_846 = {_EVAL_539,_EVAL_50};
  assign _EVAL_611 = _EVAL_291 >= _EVAL_846;
  assign _EVAL_550 = _EVAL_611 ? _EVAL_291 : _EVAL_846;
  assign _EVAL_198 = _EVAL_113[54];
  assign _EVAL_532 = {_EVAL_198,_EVAL_24};
  assign _EVAL_302 = _EVAL_113[0];
  assign _EVAL_603 = {_EVAL_302,_EVAL_95};
  assign _EVAL_468 = 4'h8 >= _EVAL_603;
  assign _EVAL_357 = _EVAL_468 ? 4'h8 : _EVAL_603;
  assign _EVAL_735 = _EVAL_113[1];
  assign _EVAL_254 = {_EVAL_735,_EVAL_21};
  assign _EVAL_855 = _EVAL_113[2];
  assign _EVAL_623 = {_EVAL_855,_EVAL_55};
  assign _EVAL_555 = _EVAL_254 >= _EVAL_623;
  assign _EVAL_422 = _EVAL_555 ? _EVAL_254 : _EVAL_623;
  assign _EVAL_758 = _EVAL_357 >= _EVAL_422;
  assign _EVAL_285 = _EVAL_758 ? _EVAL_357 : _EVAL_422;
  assign _EVAL_545 = _EVAL_113[3];
  assign _EVAL_176 = {_EVAL_545,_EVAL_103};
  assign _EVAL_666 = _EVAL_113[4];
  assign _EVAL_783 = {_EVAL_666,_EVAL_108};
  assign _EVAL_481 = _EVAL_176 >= _EVAL_783;
  assign _EVAL_804 = _EVAL_481 ? _EVAL_176 : _EVAL_783;
  assign _EVAL_820 = _EVAL_113[5];
  assign _EVAL_155 = {_EVAL_820,_EVAL_48};
  assign _EVAL_231 = _EVAL_113[6];
  assign _EVAL_174 = {_EVAL_231,_EVAL_101};
  assign _EVAL_727 = _EVAL_155 >= _EVAL_174;
  assign _EVAL_279 = _EVAL_727 ? _EVAL_155 : _EVAL_174;
  assign _EVAL_187 = _EVAL_804 >= _EVAL_279;
  assign _EVAL_661 = _EVAL_187 ? _EVAL_804 : _EVAL_279;
  assign _EVAL_301 = _EVAL_285 >= _EVAL_661;
  assign _EVAL_719 = _EVAL_468 ? 1'h0 : 1'h1;
  assign _EVAL_536 = _EVAL_555 ? 1'h0 : 1'h1;
  assign _EVAL_413 = {{1'd0}, _EVAL_536};
  assign _EVAL_567 = 2'h2 | _EVAL_413;
  assign _EVAL_425 = _EVAL_758 ? {{1'd0}, _EVAL_719} : _EVAL_567;
  assign _EVAL_213 = _EVAL_113[19];
  assign _EVAL_226 = {_EVAL_213,_EVAL_81};
  assign _EVAL_299 = _EVAL_113[20];
  assign _EVAL_824 = {_EVAL_299,_EVAL_96};
  assign _EVAL_869 = _EVAL_226 >= _EVAL_824;
  assign _EVAL_600 = _EVAL_869 ? _EVAL_226 : _EVAL_824;
  assign _EVAL_310 = _EVAL_113[21];
  assign _EVAL_858 = {_EVAL_310,_EVAL_76};
  assign _EVAL_796 = _EVAL_113[22];
  assign _EVAL_768 = {_EVAL_796,_EVAL_6};
  assign _EVAL_703 = _EVAL_858 >= _EVAL_768;
  assign _EVAL_816 = _EVAL_703 ? _EVAL_858 : _EVAL_768;
  assign _EVAL_397 = _EVAL_600 >= _EVAL_816;
  assign _EVAL_565 = _EVAL_869 ? 1'h0 : 1'h1;
  assign _EVAL_247 = _EVAL_703 ? 1'h0 : 1'h1;
  assign _EVAL_637 = {{1'd0}, _EVAL_247};
  assign _EVAL_160 = 2'h2 | _EVAL_637;
  assign _EVAL_456 = _EVAL_397 ? {{1'd0}, _EVAL_565} : _EVAL_160;
  assign _EVAL_151 = {{1'd0}, _EVAL_456};
  assign _EVAL_479 = _EVAL_113[15];
  assign _EVAL_712 = {_EVAL_479,_EVAL_47};
  assign _EVAL_474 = _EVAL_113[16];
  assign _EVAL_706 = {_EVAL_474,_EVAL_35};
  assign _EVAL_276 = _EVAL_712 >= _EVAL_706;
  assign _EVAL_501 = _EVAL_276 ? _EVAL_712 : _EVAL_706;
  assign _EVAL_388 = _EVAL_113[17];
  assign _EVAL_724 = {_EVAL_388,_EVAL_67};
  assign _EVAL_663 = _EVAL_113[18];
  assign _EVAL_533 = {_EVAL_663,_EVAL_97};
  assign _EVAL_138 = _EVAL_724 >= _EVAL_533;
  assign _EVAL_483 = _EVAL_138 ? _EVAL_724 : _EVAL_533;
  assign _EVAL_769 = _EVAL_501 >= _EVAL_483;
  assign _EVAL_619 = _EVAL_113[71];
  assign _EVAL_186 = {_EVAL_619,_EVAL_89};
  assign _EVAL_348 = _EVAL_113[72];
  assign _EVAL_453 = {_EVAL_348,_EVAL_102};
  assign _EVAL_500 = _EVAL_186 >= _EVAL_453;
  assign _EVAL_658 = _EVAL_500 ? _EVAL_186 : _EVAL_453;
  assign _EVAL_609 = _EVAL_113[73];
  assign _EVAL_189 = {_EVAL_609,_EVAL_59};
  assign _EVAL_597 = _EVAL_113[74];
  assign _EVAL_431 = {_EVAL_597,_EVAL_51};
  assign _EVAL_224 = _EVAL_189 >= _EVAL_431;
  assign _EVAL_502 = _EVAL_224 ? _EVAL_189 : _EVAL_431;
  assign _EVAL_647 = _EVAL_658 >= _EVAL_502;
  assign _EVAL_811 = _EVAL_647 ? _EVAL_658 : _EVAL_502;
  assign _EVAL_343 = _EVAL_113[75];
  assign _EVAL_743 = {_EVAL_343,_EVAL_63};
  assign _EVAL_146 = _EVAL_113[76];
  assign _EVAL_269 = {_EVAL_146,_EVAL_64};
  assign _EVAL_467 = _EVAL_743 >= _EVAL_269;
  assign _EVAL_778 = _EVAL_467 ? _EVAL_743 : _EVAL_269;
  assign _EVAL_751 = _EVAL_113[77];
  assign _EVAL_656 = {_EVAL_751,_EVAL_1};
  assign _EVAL_335 = _EVAL_113[78];
  assign _EVAL_371 = {_EVAL_335,_EVAL_44};
  assign _EVAL_212 = _EVAL_656 >= _EVAL_371;
  assign _EVAL_234 = _EVAL_212 ? _EVAL_656 : _EVAL_371;
  assign _EVAL_708 = _EVAL_778 >= _EVAL_234;
  assign _EVAL_544 = _EVAL_708 ? _EVAL_778 : _EVAL_234;
  assign _EVAL_535 = _EVAL_811 >= _EVAL_544;
  assign _EVAL_797 = _EVAL_500 ? 1'h0 : 1'h1;
  assign _EVAL_713 = _EVAL_224 ? 1'h0 : 1'h1;
  assign _EVAL_361 = {{1'd0}, _EVAL_713};
  assign _EVAL_204 = 2'h2 | _EVAL_361;
  assign _EVAL_831 = _EVAL_647 ? {{1'd0}, _EVAL_797} : _EVAL_204;
  assign _EVAL_798 = _EVAL_467 ? 1'h0 : 1'h1;
  assign _EVAL_643 = _EVAL_212 ? 1'h0 : 1'h1;
  assign _EVAL_323 = {{1'd0}, _EVAL_643};
  assign _EVAL_332 = 2'h2 | _EVAL_323;
  assign _EVAL_372 = _EVAL_708 ? {{1'd0}, _EVAL_798} : _EVAL_332;
  assign _EVAL_739 = {{1'd0}, _EVAL_372};
  assign _EVAL_626 = 3'h4 | _EVAL_739;
  assign _EVAL_268 = _EVAL_535 ? {{1'd0}, _EVAL_831} : _EVAL_626;
  assign _EVAL_284 = {{1'd0}, _EVAL_268};
  assign _EVAL_885 = _EVAL_113[57];
  assign _EVAL_809 = _EVAL_113[47];
  assign _EVAL_772 = {_EVAL_809,_EVAL_119};
  assign _EVAL_274 = _EVAL_113[48];
  assign _EVAL_795 = {_EVAL_274,_EVAL_100};
  assign _EVAL_172 = _EVAL_772 >= _EVAL_795;
  assign _EVAL_214 = _EVAL_172 ? _EVAL_772 : _EVAL_795;
  assign _EVAL_494 = _EVAL_113[49];
  assign _EVAL_196 = {_EVAL_494,_EVAL_122};
  assign _EVAL_396 = _EVAL_113[50];
  assign _EVAL_330 = {_EVAL_396,_EVAL_98};
  assign _EVAL_318 = _EVAL_196 >= _EVAL_330;
  assign _EVAL_185 = _EVAL_318 ? _EVAL_196 : _EVAL_330;
  assign _EVAL_843 = _EVAL_214 >= _EVAL_185;
  assign _EVAL_492 = _EVAL_843 ? _EVAL_214 : _EVAL_185;
  assign _EVAL_732 = _EVAL_113[51];
  assign _EVAL_766 = {_EVAL_732,_EVAL_77};
  assign _EVAL_616 = _EVAL_113[52];
  assign _EVAL_817 = {_EVAL_616,_EVAL_116};
  assign _EVAL_564 = _EVAL_766 >= _EVAL_817;
  assign _EVAL_376 = _EVAL_564 ? _EVAL_766 : _EVAL_817;
  assign _EVAL_438 = _EVAL_113[53];
  assign _EVAL_834 = {_EVAL_438,_EVAL_11};
  assign _EVAL_257 = _EVAL_834 >= _EVAL_532;
  assign _EVAL_308 = _EVAL_257 ? _EVAL_834 : _EVAL_532;
  assign _EVAL_137 = _EVAL_376 >= _EVAL_308;
  assign _EVAL_334 = _EVAL_137 ? _EVAL_376 : _EVAL_308;
  assign _EVAL_744 = _EVAL_492 >= _EVAL_334;
  assign _EVAL_638 = _EVAL_481 ? 1'h0 : 1'h1;
  assign _EVAL_823 = _EVAL_727 ? 1'h0 : 1'h1;
  assign _EVAL_333 = {{1'd0}, _EVAL_823};
  assign _EVAL_684 = 2'h2 | _EVAL_333;
  assign _EVAL_345 = _EVAL_187 ? {{1'd0}, _EVAL_638} : _EVAL_684;
  assign _EVAL_615 = {{1'd0}, _EVAL_345};
  assign _EVAL_734 = 3'h4 | _EVAL_615;
  assign _EVAL_755 = _EVAL_257 ? 1'h0 : 1'h1;
  assign _EVAL_290 = {{1'd0}, _EVAL_755};
  assign _EVAL_577 = _EVAL_113[37];
  assign _EVAL_219 = {_EVAL_577,_EVAL_121};
  assign _EVAL_738 = _EVAL_113[38];
  assign _EVAL_470 = {_EVAL_738,_EVAL_61};
  assign _EVAL_875 = _EVAL_219 >= _EVAL_470;
  assign _EVAL_295 = _EVAL_113[61];
  assign _EVAL_840 = _EVAL_113[101];
  assign _EVAL_252 = {_EVAL_840,_EVAL_73};
  assign _EVAL_729 = _EVAL_113[31];
  assign _EVAL_551 = {_EVAL_729,_EVAL_117};
  assign _EVAL_801 = _EVAL_113[32];
  assign _EVAL_691 = {_EVAL_801,_EVAL_125};
  assign _EVAL_460 = _EVAL_551 >= _EVAL_691;
  assign _EVAL_628 = _EVAL_460 ? _EVAL_551 : _EVAL_691;
  assign _EVAL_433 = _EVAL_113[33];
  assign _EVAL_519 = {_EVAL_433,_EVAL_111};
  assign _EVAL_608 = _EVAL_113[34];
  assign _EVAL_429 = {_EVAL_608,_EVAL_90};
  assign _EVAL_584 = _EVAL_519 >= _EVAL_429;
  assign _EVAL_721 = _EVAL_584 ? _EVAL_519 : _EVAL_429;
  assign _EVAL_272 = _EVAL_628 >= _EVAL_721;
  assign _EVAL_657 = _EVAL_272 ? _EVAL_628 : _EVAL_721;
  assign _EVAL_704 = _EVAL_113[35];
  assign _EVAL_542 = {_EVAL_704,_EVAL_58};
  assign _EVAL_588 = _EVAL_113[36];
  assign _EVAL_748 = {_EVAL_588,_EVAL_60};
  assign _EVAL_182 = _EVAL_542 >= _EVAL_748;
  assign _EVAL_711 = _EVAL_182 ? _EVAL_542 : _EVAL_748;
  assign _EVAL_221 = _EVAL_875 ? _EVAL_219 : _EVAL_470;
  assign _EVAL_354 = _EVAL_711 >= _EVAL_221;
  assign _EVAL_307 = _EVAL_354 ? _EVAL_711 : _EVAL_221;
  assign _EVAL_461 = _EVAL_657 >= _EVAL_307;
  assign _EVAL_750 = _EVAL_461 ? _EVAL_657 : _EVAL_307;
  assign _EVAL_418 = _EVAL_113[41];
  assign _EVAL_482 = {_EVAL_418,_EVAL_42};
  assign _EVAL_861 = _EVAL_113[42];
  assign _EVAL_731 = {_EVAL_861,_EVAL_79};
  assign _EVAL_440 = _EVAL_482 >= _EVAL_731;
  assign _EVAL_140 = _EVAL_440 ? _EVAL_482 : _EVAL_731;
  assign _EVAL_621 = _EVAL_550 >= _EVAL_140;
  assign _EVAL_863 = _EVAL_621 ? _EVAL_550 : _EVAL_140;
  assign _EVAL_159 = _EVAL_113[43];
  assign _EVAL_312 = {_EVAL_159,_EVAL_4};
  assign _EVAL_589 = _EVAL_113[44];
  assign _EVAL_304 = {_EVAL_589,_EVAL_93};
  assign _EVAL_510 = _EVAL_312 >= _EVAL_304;
  assign _EVAL_437 = _EVAL_510 ? _EVAL_312 : _EVAL_304;
  assign _EVAL_405 = _EVAL_113[45];
  assign _EVAL_315 = {_EVAL_405,_EVAL_115};
  assign _EVAL_767 = _EVAL_113[46];
  assign _EVAL_813 = {_EVAL_767,_EVAL_118};
  assign _EVAL_685 = _EVAL_315 >= _EVAL_813;
  assign _EVAL_195 = _EVAL_685 ? _EVAL_315 : _EVAL_813;
  assign _EVAL_635 = _EVAL_437 >= _EVAL_195;
  assign _EVAL_166 = _EVAL_635 ? _EVAL_437 : _EVAL_195;
  assign _EVAL_380 = _EVAL_863 >= _EVAL_166;
  assign _EVAL_705 = _EVAL_380 ? _EVAL_863 : _EVAL_166;
  assign _EVAL_747 = _EVAL_750 >= _EVAL_705;
  assign _EVAL_549 = _EVAL_747 ? _EVAL_750 : _EVAL_705;
  assign _EVAL_722 = _EVAL_744 ? _EVAL_492 : _EVAL_334;
  assign _EVAL_201 = _EVAL_113[55];
  assign _EVAL_518 = {_EVAL_201,_EVAL_8};
  assign _EVAL_849 = _EVAL_113[56];
  assign _EVAL_144 = {_EVAL_849,_EVAL_71};
  assign _EVAL_242 = _EVAL_518 >= _EVAL_144;
  assign _EVAL_851 = _EVAL_242 ? _EVAL_518 : _EVAL_144;
  assign _EVAL_391 = {_EVAL_885,_EVAL_78};
  assign _EVAL_799 = _EVAL_113[58];
  assign _EVAL_507 = {_EVAL_799,_EVAL_84};
  assign _EVAL_505 = _EVAL_391 >= _EVAL_507;
  assign _EVAL_826 = _EVAL_505 ? _EVAL_391 : _EVAL_507;
  assign _EVAL_350 = _EVAL_851 >= _EVAL_826;
  assign _EVAL_618 = _EVAL_350 ? _EVAL_851 : _EVAL_826;
  assign _EVAL_401 = _EVAL_113[59];
  assign _EVAL_864 = {_EVAL_401,_EVAL_33};
  assign _EVAL_452 = _EVAL_113[60];
  assign _EVAL_415 = {_EVAL_452,_EVAL_5};
  assign _EVAL_590 = _EVAL_864 >= _EVAL_415;
  assign _EVAL_802 = _EVAL_590 ? _EVAL_864 : _EVAL_415;
  assign _EVAL_668 = {_EVAL_295,_EVAL_105};
  assign _EVAL_416 = _EVAL_113[62];
  assign _EVAL_856 = {_EVAL_416,_EVAL_31};
  assign _EVAL_464 = _EVAL_668 >= _EVAL_856;
  assign _EVAL_614 = _EVAL_464 ? _EVAL_668 : _EVAL_856;
  assign _EVAL_419 = _EVAL_802 >= _EVAL_614;
  assign _EVAL_873 = _EVAL_419 ? _EVAL_802 : _EVAL_614;
  assign _EVAL_435 = _EVAL_618 >= _EVAL_873;
  assign _EVAL_650 = _EVAL_435 ? _EVAL_618 : _EVAL_873;
  assign _EVAL_591 = _EVAL_722 >= _EVAL_650;
  assign _EVAL_206 = _EVAL_591 ? _EVAL_722 : _EVAL_650;
  assign _EVAL_374 = _EVAL_549 >= _EVAL_206;
  assign _EVAL_726 = _EVAL_113[107];
  assign _EVAL_692 = {_EVAL_726,_EVAL_30};
  assign _EVAL_136 = _EVAL_113[108];
  assign _EVAL_161 = {_EVAL_136,_EVAL_86};
  assign _EVAL_366 = _EVAL_692 >= _EVAL_161;
  assign _EVAL_541 = _EVAL_113[115];
  assign _EVAL_181 = {_EVAL_541,_EVAL_127};
  assign _EVAL_884 = _EVAL_113[116];
  assign _EVAL_728 = {_EVAL_884,_EVAL_126};
  assign _EVAL_717 = _EVAL_181 >= _EVAL_728;
  assign _EVAL_844 = _EVAL_717 ? _EVAL_181 : _EVAL_728;
  assign _EVAL_485 = _EVAL_113[117];
  assign _EVAL_303 = {_EVAL_485,_EVAL_10};
  assign _EVAL_612 = _EVAL_113[118];
  assign _EVAL_516 = {_EVAL_612,_EVAL};
  assign _EVAL_720 = _EVAL_303 >= _EVAL_516;
  assign _EVAL_458 = _EVAL_720 ? _EVAL_303 : _EVAL_516;
  assign _EVAL_130 = _EVAL_844 >= _EVAL_458;
  assign _EVAL_378 = _EVAL_130 ? _EVAL_844 : _EVAL_458;
  assign _EVAL_465 = _EVAL_113[26];
  assign _EVAL_496 = _EVAL_113[29];
  assign _EVAL_693 = {_EVAL_496,_EVAL_52};
  assign _EVAL_853 = _EVAL_113[30];
  assign _EVAL_359 = {_EVAL_853,_EVAL_16};
  assign _EVAL_207 = _EVAL_693 >= _EVAL_359;
  assign _EVAL_249 = _EVAL_207 ? 1'h0 : 1'h1;
  assign _EVAL_367 = {{1'd0}, _EVAL_249};
  assign _EVAL_232 = 2'h2 | _EVAL_367;
  assign _EVAL_349 = _EVAL_113[125];
  assign _EVAL_227 = {_EVAL_349,_EVAL_70};
  assign _EVAL_527 = _EVAL_113[126];
  assign _EVAL_636 = {_EVAL_527,_EVAL_72};
  assign _EVAL_449 = _EVAL_227 >= _EVAL_636;
  assign _EVAL_819 = _EVAL_449 ? 1'h0 : 1'h1;
  assign _EVAL_548 = {{1'd0}, _EVAL_819};
  assign _EVAL_753 = _EVAL_113[79];
  assign _EVAL_558 = {_EVAL_753,_EVAL_7};
  assign _EVAL_593 = _EVAL_113[80];
  assign _EVAL_373 = {_EVAL_593,_EVAL_22};
  assign _EVAL_845 = _EVAL_558 >= _EVAL_373;
  assign _EVAL_408 = _EVAL_845 ? 1'h0 : 1'h1;
  assign _EVAL_287 = _EVAL_113[70];
  assign _EVAL_278 = {_EVAL_287,_EVAL_128};
  assign _EVAL_789 = _EVAL_113[97];
  assign _EVAL_356 = {_EVAL_789,_EVAL_18};
  assign _EVAL_723 = _EVAL_113[98];
  assign _EVAL_673 = {_EVAL_723,_EVAL_68};
  assign _EVAL_205 = _EVAL_356 >= _EVAL_673;
  assign _EVAL_211 = _EVAL_845 ? _EVAL_558 : _EVAL_373;
  assign _EVAL_807 = _EVAL_113[81];
  assign _EVAL_531 = {_EVAL_807,_EVAL_57};
  assign _EVAL_877 = _EVAL_113[82];
  assign _EVAL_521 = {_EVAL_877,_EVAL_13};
  assign _EVAL_792 = _EVAL_531 >= _EVAL_521;
  assign _EVAL_286 = _EVAL_792 ? _EVAL_531 : _EVAL_521;
  assign _EVAL_439 = _EVAL_211 >= _EVAL_286;
  assign _EVAL_363 = _EVAL_792 ? 1'h0 : 1'h1;
  assign _EVAL_605 = {{1'd0}, _EVAL_363};
  assign _EVAL_170 = 2'h2 | _EVAL_605;
  assign _EVAL_407 = _EVAL_439 ? {{1'd0}, _EVAL_408} : _EVAL_170;
  assign _EVAL_522 = _EVAL_113[102];
  assign _EVAL_382 = {_EVAL_522,_EVAL_74};
  assign _EVAL_183 = _EVAL_252 >= _EVAL_382;
  assign _EVAL_336 = _EVAL_183 ? _EVAL_252 : _EVAL_382;
  assign _EVAL_830 = _EVAL_138 ? 1'h0 : 1'h1;
  assign _EVAL_774 = {{1'd0}, _EVAL_830};
  assign _EVAL_471 = 2'h2 | _EVAL_774;
  assign _EVAL_157 = _EVAL_113[69];
  assign _EVAL_175 = _EVAL_113[11];
  assign _EVAL_760 = {_EVAL_175,_EVAL_99};
  assign _EVAL_594 = _EVAL_113[12];
  assign _EVAL_457 = {_EVAL_594,_EVAL_12};
  assign _EVAL_640 = _EVAL_760 >= _EVAL_457;
  assign _EVAL_338 = _EVAL_113[23];
  assign _EVAL_570 = {_EVAL_338,_EVAL_123};
  assign _EVAL_282 = _EVAL_113[24];
  assign _EVAL_553 = {_EVAL_282,_EVAL_26};
  assign _EVAL_675 = _EVAL_570 >= _EVAL_553;
  assign _EVAL_859 = _EVAL_675 ? _EVAL_570 : _EVAL_553;
  assign _EVAL_569 = _EVAL_113[25];
  assign _EVAL_520 = {_EVAL_569,_EVAL_62};
  assign _EVAL_523 = {_EVAL_465,_EVAL_37};
  assign _EVAL_848 = _EVAL_520 >= _EVAL_523;
  assign _EVAL_572 = _EVAL_848 ? _EVAL_520 : _EVAL_523;
  assign _EVAL_718 = _EVAL_859 >= _EVAL_572;
  assign _EVAL_534 = _EVAL_718 ? _EVAL_859 : _EVAL_572;
  assign _EVAL_169 = _EVAL_113[27];
  assign _EVAL_665 = {_EVAL_169,_EVAL_82};
  assign _EVAL_543 = _EVAL_113[28];
  assign _EVAL_385 = {_EVAL_543,_EVAL_2};
  assign _EVAL_484 = _EVAL_665 >= _EVAL_385;
  assign _EVAL_678 = _EVAL_484 ? _EVAL_665 : _EVAL_385;
  assign _EVAL_446 = _EVAL_207 ? _EVAL_693 : _EVAL_359;
  assign _EVAL_686 = _EVAL_678 >= _EVAL_446;
  assign _EVAL_375 = _EVAL_686 ? _EVAL_678 : _EVAL_446;
  assign _EVAL_765 = _EVAL_534 >= _EVAL_375;
  assign _EVAL_699 = _EVAL_675 ? 1'h0 : 1'h1;
  assign _EVAL_725 = _EVAL_848 ? 1'h0 : 1'h1;
  assign _EVAL_629 = {{1'd0}, _EVAL_725};
  assign _EVAL_624 = 2'h2 | _EVAL_629;
  assign _EVAL_800 = _EVAL_718 ? {{1'd0}, _EVAL_699} : _EVAL_624;
  assign _EVAL_681 = _EVAL_484 ? 1'h0 : 1'h1;
  assign _EVAL_208 = _EVAL_686 ? {{1'd0}, _EVAL_681} : _EVAL_232;
  assign _EVAL_489 = {{1'd0}, _EVAL_208};
  assign _EVAL_561 = 3'h4 | _EVAL_489;
  assign _EVAL_131 = _EVAL_765 ? {{1'd0}, _EVAL_800} : _EVAL_561;
  assign _EVAL_781 = {{1'd0}, _EVAL_131};
  assign _EVAL_360 = _EVAL_113[111];
  assign _EVAL_680 = {_EVAL_360,_EVAL_106};
  assign _EVAL_230 = _EVAL_113[112];
  assign _EVAL_676 = {_EVAL_230,_EVAL_29};
  assign _EVAL_381 = _EVAL_680 >= _EVAL_676;
  assign _EVAL_707 = _EVAL_113[66];
  assign _EVAL_222 = _EVAL_113[7];
  assign _EVAL_164 = {_EVAL_222,_EVAL_9};
  assign _EVAL_347 = _EVAL_113[8];
  assign _EVAL_495 = {_EVAL_347,_EVAL_104};
  assign _EVAL_216 = _EVAL_164 >= _EVAL_495;
  assign _EVAL_390 = _EVAL_216 ? _EVAL_164 : _EVAL_495;
  assign _EVAL_808 = _EVAL_113[9];
  assign _EVAL_370 = {_EVAL_808,_EVAL_94};
  assign _EVAL_810 = _EVAL_113[10];
  assign _EVAL_313 = {_EVAL_810,_EVAL_19};
  assign _EVAL_412 = _EVAL_370 >= _EVAL_313;
  assign _EVAL_342 = _EVAL_412 ? _EVAL_370 : _EVAL_313;
  assign _EVAL_253 = _EVAL_390 >= _EVAL_342;
  assign _EVAL_364 = _EVAL_253 ? _EVAL_390 : _EVAL_342;
  assign _EVAL_402 = _EVAL_640 ? _EVAL_760 : _EVAL_457;
  assign _EVAL_822 = _EVAL_113[13];
  assign _EVAL_424 = {_EVAL_822,_EVAL_15};
  assign _EVAL_135 = _EVAL_113[14];
  assign _EVAL_794 = {_EVAL_135,_EVAL_40};
  assign _EVAL_710 = _EVAL_424 >= _EVAL_794;
  assign _EVAL_818 = _EVAL_710 ? _EVAL_424 : _EVAL_794;
  assign _EVAL_190 = _EVAL_402 >= _EVAL_818;
  assign _EVAL_870 = _EVAL_190 ? _EVAL_402 : _EVAL_818;
  assign _EVAL_630 = _EVAL_364 >= _EVAL_870;
  assign _EVAL_837 = _EVAL_216 ? 1'h0 : 1'h1;
  assign _EVAL_610 = _EVAL_412 ? 1'h0 : 1'h1;
  assign _EVAL_141 = {{1'd0}, _EVAL_610};
  assign _EVAL_672 = 2'h2 | _EVAL_141;
  assign _EVAL_358 = _EVAL_253 ? {{1'd0}, _EVAL_837} : _EVAL_672;
  assign _EVAL_627 = _EVAL_640 ? 1'h0 : 1'h1;
  assign _EVAL_236 = _EVAL_710 ? 1'h0 : 1'h1;
  assign _EVAL_517 = {{1'd0}, _EVAL_236};
  assign _EVAL_223 = 2'h2 | _EVAL_517;
  assign _EVAL_503 = _EVAL_190 ? {{1'd0}, _EVAL_627} : _EVAL_223;
  assign _EVAL_814 = {{1'd0}, _EVAL_503};
  assign _EVAL_882 = 3'h4 | _EVAL_814;
  assign _EVAL_754 = _EVAL_630 ? {{1'd0}, _EVAL_358} : _EVAL_882;
  assign _EVAL_445 = {{1'd0}, _EVAL_754};
  assign _EVAL_733 = _EVAL_113[83];
  assign _EVAL_574 = {_EVAL_733,_EVAL_65};
  assign _EVAL_776 = _EVAL_113[84];
  assign _EVAL_184 = {_EVAL_776,_EVAL_66};
  assign _EVAL_283 = _EVAL_574 >= _EVAL_184;
  assign _EVAL_607 = _EVAL_283 ? _EVAL_574 : _EVAL_184;
  assign _EVAL_188 = _EVAL_113[85];
  assign _EVAL_229 = {_EVAL_188,_EVAL_25};
  assign _EVAL_759 = _EVAL_113[86];
  assign _EVAL_689 = {_EVAL_759,_EVAL_49};
  assign _EVAL_568 = _EVAL_229 >= _EVAL_689;
  assign _EVAL_156 = _EVAL_568 ? _EVAL_229 : _EVAL_689;
  assign _EVAL_653 = _EVAL_607 >= _EVAL_156;
  assign _EVAL_506 = _EVAL_283 ? 1'h0 : 1'h1;
  assign _EVAL_669 = _EVAL_568 ? 1'h0 : 1'h1;
  assign _EVAL_162 = {{1'd0}, _EVAL_669};
  assign _EVAL_455 = 2'h2 | _EVAL_162;
  assign _EVAL_697 = _EVAL_653 ? {{1'd0}, _EVAL_506} : _EVAL_455;
  assign _EVAL_632 = {{1'd0}, _EVAL_697};
  assign _EVAL_339 = _EVAL_113[95];
  assign _EVAL_173 = {_EVAL_339,_EVAL_17};
  assign _EVAL_745 = _EVAL_113[103];
  assign _EVAL_690 = {_EVAL_745,_EVAL_109};
  assign _EVAL_426 = _EVAL_113[104];
  assign _EVAL_762 = {_EVAL_426,_EVAL_107};
  assign _EVAL_275 = _EVAL_690 >= _EVAL_762;
  assign _EVAL_880 = _EVAL_275 ? _EVAL_690 : _EVAL_762;
  assign _EVAL_280 = _EVAL_113[105];
  assign _EVAL_200 = {_EVAL_280,_EVAL_69};
  assign _EVAL_322 = _EVAL_113[106];
  assign _EVAL_298 = {_EVAL_322,_EVAL_114};
  assign _EVAL_599 = _EVAL_200 >= _EVAL_298;
  assign _EVAL_134 = _EVAL_599 ? _EVAL_200 : _EVAL_298;
  assign _EVAL_580 = _EVAL_880 >= _EVAL_134;
  assign _EVAL_601 = _EVAL_580 ? _EVAL_880 : _EVAL_134;
  assign _EVAL_294 = _EVAL_366 ? _EVAL_692 : _EVAL_161;
  assign _EVAL_777 = _EVAL_113[109];
  assign _EVAL_659 = {_EVAL_777,_EVAL_38};
  assign _EVAL_617 = _EVAL_113[110];
  assign _EVAL_827 = {_EVAL_617,_EVAL_85};
  assign _EVAL_582 = _EVAL_659 >= _EVAL_827;
  assign _EVAL_368 = _EVAL_582 ? _EVAL_659 : _EVAL_827;
  assign _EVAL_441 = _EVAL_294 >= _EVAL_368;
  assign _EVAL_444 = _EVAL_441 ? _EVAL_294 : _EVAL_368;
  assign _EVAL_639 = _EVAL_601 >= _EVAL_444;
  assign _EVAL_488 = _EVAL_275 ? 1'h0 : 1'h1;
  assign _EVAL_649 = _EVAL_599 ? 1'h0 : 1'h1;
  assign _EVAL_490 = {{1'd0}, _EVAL_649};
  assign _EVAL_327 = 2'h2 | _EVAL_490;
  assign _EVAL_874 = _EVAL_580 ? {{1'd0}, _EVAL_488} : _EVAL_327;
  assign _EVAL_326 = _EVAL_366 ? 1'h0 : 1'h1;
  assign _EVAL_825 = _EVAL_582 ? 1'h0 : 1'h1;
  assign _EVAL_145 = {{1'd0}, _EVAL_825};
  assign _EVAL_821 = 2'h2 | _EVAL_145;
  assign _EVAL_317 = _EVAL_441 ? {{1'd0}, _EVAL_326} : _EVAL_821;
  assign _EVAL_592 = {{1'd0}, _EVAL_317};
  assign _EVAL_694 = 3'h4 | _EVAL_592;
  assign _EVAL_409 = _EVAL_639 ? {{1'd0}, _EVAL_874} : _EVAL_694;
  assign _EVAL_238 = {{1'd0}, _EVAL_409};
  assign _EVAL_805 = 4'h8 | _EVAL_238;
  assign _EVAL_682 = _EVAL_862 ? 1'h0 : 1'h1;
  assign _EVAL_386 = _EVAL_584 ? 1'h0 : 1'h1;
  assign _EVAL_566 = {{1'd0}, _EVAL_386};
  assign _EVAL_475 = _EVAL_113[123];
  assign _EVAL_540 = {_EVAL_475,_EVAL_88};
  assign _EVAL_153 = _EVAL_113[124];
  assign _EVAL_379 = {_EVAL_153,_EVAL_46};
  assign _EVAL_251 = _EVAL_540 >= _EVAL_379;
  assign _EVAL_293 = _EVAL_251 ? _EVAL_540 : _EVAL_379;
  assign _EVAL_421 = _EVAL_449 ? _EVAL_227 : _EVAL_636;
  assign _EVAL_749 = _EVAL_293 >= _EVAL_421;
  assign _EVAL_258 = _EVAL_113[65];
  assign _EVAL_480 = {_EVAL_258,_EVAL_56};
  assign _EVAL_191 = {_EVAL_707,_EVAL_110};
  assign _EVAL_604 = _EVAL_480 >= _EVAL_191;
  assign _EVAL_847 = _EVAL_604 ? 1'h0 : 1'h1;
  assign _EVAL_316 = {{1'd0}, _EVAL_847};
  assign _EVAL_526 = 2'h2 | _EVAL_316;
  assign _EVAL_218 = _EVAL_505 ? 1'h0 : 1'h1;
  assign _EVAL_714 = {{1'd0}, _EVAL_218};
  assign _EVAL_560 = _EVAL_113[113];
  assign _EVAL_281 = {_EVAL_560,_EVAL_112};
  assign _EVAL_812 = _EVAL_113[114];
  assign _EVAL_448 = {_EVAL_812,_EVAL_54};
  assign _EVAL_833 = _EVAL_281 >= _EVAL_448;
  assign _EVAL_498 = _EVAL_833 ? _EVAL_281 : _EVAL_448;
  assign _EVAL_842 = _EVAL_242 ? 1'h0 : 1'h1;
  assign _EVAL_394 = 2'h2 | _EVAL_714;
  assign _EVAL_554 = _EVAL_350 ? {{1'd0}, _EVAL_842} : _EVAL_394;
  assign _EVAL_319 = _EVAL_590 ? 1'h0 : 1'h1;
  assign _EVAL_642 = _EVAL_464 ? 1'h0 : 1'h1;
  assign _EVAL_233 = {{1'd0}, _EVAL_642};
  assign _EVAL_670 = 2'h2 | _EVAL_233;
  assign _EVAL_340 = _EVAL_419 ? {{1'd0}, _EVAL_319} : _EVAL_670;
  assign _EVAL_152 = {{1'd0}, _EVAL_340};
  assign _EVAL_194 = 3'h4 | _EVAL_152;
  assign _EVAL_865 = _EVAL_435 ? {{1'd0}, _EVAL_554} : _EVAL_194;
  assign _EVAL_756 = {{1'd0}, _EVAL_865};
  assign _EVAL_557 = _EVAL_301 ? _EVAL_285 : _EVAL_661;
  assign _EVAL_406 = _EVAL_630 ? _EVAL_364 : _EVAL_870;
  assign _EVAL_255 = _EVAL_557 >= _EVAL_406;
  assign _EVAL_598 = _EVAL_255 ? _EVAL_557 : _EVAL_406;
  assign _EVAL_868 = _EVAL_769 ? _EVAL_501 : _EVAL_483;
  assign _EVAL_369 = _EVAL_397 ? _EVAL_600 : _EVAL_816;
  assign _EVAL_351 = _EVAL_868 >= _EVAL_369;
  assign _EVAL_147 = _EVAL_351 ? _EVAL_868 : _EVAL_369;
  assign _EVAL_645 = _EVAL_765 ? _EVAL_534 : _EVAL_375;
  assign _EVAL_305 = _EVAL_147 >= _EVAL_645;
  assign _EVAL_587 = _EVAL_305 ? _EVAL_147 : _EVAL_645;
  assign _EVAL_337 = _EVAL_598 >= _EVAL_587;
  assign _EVAL_149 = _EVAL_337 ? _EVAL_598 : _EVAL_587;
  assign _EVAL_881 = _EVAL_653 ? _EVAL_607 : _EVAL_156;
  assign _EVAL_210 = 2'h2 | _EVAL_548;
  assign _EVAL_736 = _EVAL_113[96];
  assign _EVAL_353 = _EVAL_113[63];
  assign _EVAL_384 = {_EVAL_353,_EVAL_14};
  assign _EVAL_871 = _EVAL_113[64];
  assign _EVAL_241 = {_EVAL_871,_EVAL_20};
  assign _EVAL_377 = _EVAL_384 >= _EVAL_241;
  assign _EVAL_434 = _EVAL_377 ? _EVAL_384 : _EVAL_241;
  assign _EVAL_259 = _EVAL_604 ? _EVAL_480 : _EVAL_191;
  assign _EVAL_698 = _EVAL_434 >= _EVAL_259;
  assign _EVAL_508 = _EVAL_698 ? _EVAL_434 : _EVAL_259;
  assign _EVAL_466 = _EVAL_113[67];
  assign _EVAL_243 = {_EVAL_466,_EVAL_87};
  assign _EVAL_423 = _EVAL_113[68];
  assign _EVAL_139 = {_EVAL_423,_EVAL_3};
  assign _EVAL_428 = _EVAL_243 >= _EVAL_139;
  assign _EVAL_306 = _EVAL_428 ? _EVAL_243 : _EVAL_139;
  assign _EVAL_791 = {_EVAL_157,_EVAL_34};
  assign _EVAL_784 = _EVAL_791 >= _EVAL_278;
  assign _EVAL_606 = _EVAL_784 ? _EVAL_791 : _EVAL_278;
  assign _EVAL_193 = _EVAL_306 >= _EVAL_606;
  assign _EVAL_651 = _EVAL_193 ? _EVAL_306 : _EVAL_606;
  assign _EVAL_404 = _EVAL_508 >= _EVAL_651;
  assign _EVAL_576 = _EVAL_404 ? _EVAL_508 : _EVAL_651;
  assign _EVAL_430 = _EVAL_770 ? 1'h0 : 1'h1;
  assign _EVAL_835 = {{1'd0}, _EVAL_430};
  assign _EVAL_631 = 2'h2 | _EVAL_835;
  assign _EVAL_742 = _EVAL_702 ? {{1'd0}, _EVAL_682} : _EVAL_631;
  assign _EVAL_829 = _EVAL_876 ? 1'h0 : 1'h1;
  assign _EVAL_432 = _EVAL_192 ? 1'h0 : 1'h1;
  assign _EVAL_447 = {{1'd0}, _EVAL_432};
  assign _EVAL_469 = 2'h2 | _EVAL_447;
  assign _EVAL_709 = _EVAL_436 ? {{1'd0}, _EVAL_829} : _EVAL_469;
  assign _EVAL_158 = {{1'd0}, _EVAL_709};
  assign _EVAL_395 = 3'h4 | _EVAL_158;
  assign _EVAL_477 = _EVAL_486 ? {{1'd0}, _EVAL_742} : _EVAL_395;
  assign _EVAL_493 = {{1'd0}, _EVAL_477};
  assign _EVAL_142 = _EVAL_113[99];
  assign _EVAL_537 = {_EVAL_142,_EVAL_28};
  assign _EVAL_410 = _EVAL_113[100];
  assign _EVAL_786 = {_EVAL_410,_EVAL_83};
  assign _EVAL_248 = _EVAL_537 >= _EVAL_786;
  assign _EVAL_393 = _EVAL_113[119];
  assign _EVAL_559 = {_EVAL_393,_EVAL_0};
  assign _EVAL_646 = _EVAL_113[121];
  assign _EVAL_546 = _EVAL_535 ? _EVAL_811 : _EVAL_544;
  assign _EVAL_552 = _EVAL_576 >= _EVAL_546;
  assign _EVAL_562 = _EVAL_552 ? _EVAL_576 : _EVAL_546;
  assign _EVAL_165 = _EVAL_439 ? _EVAL_211 : _EVAL_286;
  assign _EVAL_365 = _EVAL_165 >= _EVAL_881;
  assign _EVAL_613 = _EVAL_365 ? _EVAL_165 : _EVAL_881;
  assign _EVAL_220 = _EVAL_613 >= _EVAL_512;
  assign _EVAL_513 = _EVAL_220 ? _EVAL_613 : _EVAL_512;
  assign _EVAL_491 = _EVAL_562 >= _EVAL_513;
  assign _EVAL_883 = _EVAL_491 ? _EVAL_562 : _EVAL_513;
  assign _EVAL_538 = {_EVAL_736,_EVAL_43};
  assign _EVAL_509 = _EVAL_173 >= _EVAL_538;
  assign _EVAL_267 = _EVAL_509 ? _EVAL_173 : _EVAL_538;
  assign _EVAL_443 = _EVAL_205 ? _EVAL_356 : _EVAL_673;
  assign _EVAL_459 = _EVAL_267 >= _EVAL_443;
  assign _EVAL_741 = _EVAL_459 ? _EVAL_267 : _EVAL_443;
  assign _EVAL_237 = _EVAL_248 ? _EVAL_537 : _EVAL_786;
  assign _EVAL_266 = _EVAL_237 >= _EVAL_336;
  assign _EVAL_524 = _EVAL_266 ? _EVAL_237 : _EVAL_336;
  assign _EVAL_217 = _EVAL_741 >= _EVAL_524;
  assign _EVAL_177 = _EVAL_217 ? _EVAL_741 : _EVAL_524;
  assign _EVAL_771 = _EVAL_639 ? _EVAL_601 : _EVAL_444;
  assign _EVAL_163 = _EVAL_177 >= _EVAL_771;
  assign _EVAL_815 = _EVAL_163 ? _EVAL_177 : _EVAL_771;
  assign _EVAL_806 = _EVAL_381 ? _EVAL_680 : _EVAL_676;
  assign _EVAL_775 = _EVAL_806 >= _EVAL_498;
  assign _EVAL_579 = _EVAL_775 ? _EVAL_806 : _EVAL_498;
  assign _EVAL_178 = _EVAL_579 >= _EVAL_378;
  assign _EVAL_715 = _EVAL_178 ? _EVAL_579 : _EVAL_378;
  assign _EVAL_752 = _EVAL_113[120];
  assign _EVAL_264 = {_EVAL_752,_EVAL_41};
  assign _EVAL_504 = _EVAL_559 >= _EVAL_264;
  assign _EVAL_850 = _EVAL_504 ? _EVAL_559 : _EVAL_264;
  assign _EVAL_150 = {_EVAL_646,_EVAL_80};
  assign _EVAL_399 = _EVAL_113[122];
  assign _EVAL_225 = {_EVAL_399,_EVAL_45};
  assign _EVAL_344 = _EVAL_150 >= _EVAL_225;
  assign _EVAL_320 = _EVAL_344 ? _EVAL_150 : _EVAL_225;
  assign _EVAL_857 = _EVAL_850 >= _EVAL_320;
  assign _EVAL_648 = _EVAL_857 ? _EVAL_850 : _EVAL_320;
  assign _EVAL_620 = _EVAL_749 ? _EVAL_293 : _EVAL_421;
  assign _EVAL_154 = _EVAL_648 >= _EVAL_620;
  assign _EVAL_660 = _EVAL_154 ? _EVAL_648 : _EVAL_620;
  assign _EVAL_581 = _EVAL_715 >= _EVAL_660;
  assign _EVAL_737 = _EVAL_581 ? _EVAL_715 : _EVAL_660;
  assign _EVAL_695 = _EVAL_815 >= _EVAL_737;
  assign _EVAL_528 = _EVAL_695 ? _EVAL_815 : _EVAL_737;
  assign _EVAL_260 = _EVAL_883 >= _EVAL_528;
  assign _EVAL_171 = _EVAL_377 ? 1'h0 : 1'h1;
  assign _EVAL_785 = _EVAL_698 ? {{1'd0}, _EVAL_171} : _EVAL_526;
  assign _EVAL_625 = _EVAL_428 ? 1'h0 : 1'h1;
  assign _EVAL_787 = _EVAL_784 ? 1'h0 : 1'h1;
  assign _EVAL_270 = {{1'd0}, _EVAL_787};
  assign _EVAL_228 = 2'h2 | _EVAL_270;
  assign _EVAL_838 = _EVAL_193 ? {{1'd0}, _EVAL_625} : _EVAL_228;
  assign _EVAL_790 = {{1'd0}, _EVAL_838};
  assign _EVAL_573 = 3'h4 | _EVAL_790;
  assign _EVAL_389 = _EVAL_404 ? {{1'd0}, _EVAL_785} : _EVAL_573;
  assign _EVAL_398 = 4'h8 | _EVAL_284;
  assign _EVAL_586 = _EVAL_552 ? {{1'd0}, _EVAL_389} : _EVAL_398;
  assign _EVAL_454 = 3'h4 | _EVAL_632;
  assign _EVAL_383 = _EVAL_365 ? {{1'd0}, _EVAL_407} : _EVAL_454;
  assign _EVAL_263 = 4'h8 | _EVAL_493;
  assign _EVAL_209 = _EVAL_220 ? {{1'd0}, _EVAL_383} : _EVAL_263;
  assign _EVAL_314 = {{1'd0}, _EVAL_209};
  assign _EVAL_215 = 5'h10 | _EVAL_314;
  assign _EVAL_297 = _EVAL_491 ? {{1'd0}, _EVAL_586} : _EVAL_215;
  assign _EVAL_701 = _EVAL_509 ? 1'h0 : 1'h1;
  assign _EVAL_476 = _EVAL_205 ? 1'h0 : 1'h1;
  assign _EVAL_289 = {{1'd0}, _EVAL_476};
  assign _EVAL_256 = 2'h2 | _EVAL_289;
  assign _EVAL_324 = _EVAL_459 ? {{1'd0}, _EVAL_701} : _EVAL_256;
  assign _EVAL_841 = _EVAL_248 ? 1'h0 : 1'h1;
  assign _EVAL_879 = _EVAL_183 ? 1'h0 : 1'h1;
  assign _EVAL_547 = {{1'd0}, _EVAL_879};
  assign _EVAL_866 = 2'h2 | _EVAL_547;
  assign _EVAL_730 = _EVAL_266 ? {{1'd0}, _EVAL_841} : _EVAL_866;
  assign _EVAL_296 = {{1'd0}, _EVAL_730};
  assign _EVAL_411 = 3'h4 | _EVAL_296;
  assign _EVAL_129 = _EVAL_217 ? {{1'd0}, _EVAL_324} : _EVAL_411;
  assign _EVAL_167 = _EVAL_163 ? {{1'd0}, _EVAL_129} : _EVAL_805;
  assign _EVAL_288 = _EVAL_381 ? 1'h0 : 1'h1;
  assign _EVAL_652 = _EVAL_833 ? 1'h0 : 1'h1;
  assign _EVAL_878 = {{1'd0}, _EVAL_652};
  assign _EVAL_860 = 2'h2 | _EVAL_878;
  assign _EVAL_355 = _EVAL_775 ? {{1'd0}, _EVAL_288} : _EVAL_860;
  assign _EVAL_199 = _EVAL_717 ? 1'h0 : 1'h1;
  assign _EVAL_245 = _EVAL_720 ? 1'h0 : 1'h1;
  assign _EVAL_265 = {{1'd0}, _EVAL_245};
  assign _EVAL_832 = 2'h2 | _EVAL_265;
  assign _EVAL_442 = _EVAL_130 ? {{1'd0}, _EVAL_199} : _EVAL_832;
  assign _EVAL_262 = {{1'd0}, _EVAL_442};
  assign _EVAL_667 = 3'h4 | _EVAL_262;
  assign _EVAL_180 = _EVAL_178 ? {{1'd0}, _EVAL_355} : _EVAL_667;
  assign _EVAL_292 = _EVAL_504 ? 1'h0 : 1'h1;
  assign _EVAL_328 = _EVAL_344 ? 1'h0 : 1'h1;
  assign _EVAL_773 = {{1'd0}, _EVAL_328};
  assign _EVAL_836 = 2'h2 | _EVAL_773;
  assign _EVAL_311 = _EVAL_857 ? {{1'd0}, _EVAL_292} : _EVAL_836;
  assign _EVAL_387 = _EVAL_251 ? 1'h0 : 1'h1;
  assign _EVAL_487 = _EVAL_749 ? {{1'd0}, _EVAL_387} : _EVAL_210;
  assign _EVAL_240 = {{1'd0}, _EVAL_487};
  assign _EVAL_451 = 3'h4 | _EVAL_240;
  assign _EVAL_329 = _EVAL_154 ? {{1'd0}, _EVAL_311} : _EVAL_451;
  assign _EVAL_757 = {{1'd0}, _EVAL_329};
  assign _EVAL_346 = 4'h8 | _EVAL_757;
  assign _EVAL_674 = _EVAL_581 ? {{1'd0}, _EVAL_180} : _EVAL_346;
  assign _EVAL_246 = {{1'd0}, _EVAL_674};
  assign _EVAL_664 = 5'h10 | _EVAL_246;
  assign _EVAL_450 = _EVAL_695 ? {{1'd0}, _EVAL_167} : _EVAL_664;
  assign _EVAL_852 = {{1'd0}, _EVAL_450};
  assign _EVAL_321 = 6'h20 | _EVAL_852;
  assign _EVAL_197 = _EVAL_260 ? {{1'd0}, _EVAL_297} : _EVAL_321;
  assign _EVAL_872 = {{1'd0}, _EVAL_197};
  assign _EVAL_716 = 7'h40 | _EVAL_872;
  assign _EVAL_679 = _EVAL_611 ? 1'h0 : 1'h1;
  assign _EVAL_497 = _EVAL_440 ? 1'h0 : 1'h1;
  assign _EVAL_602 = {{1'd0}, _EVAL_497};
  assign _EVAL_427 = 2'h2 | _EVAL_602;
  assign _EVAL_400 = _EVAL_621 ? {{1'd0}, _EVAL_679} : _EVAL_427;
  assign _EVAL_261 = _EVAL_510 ? 1'h0 : 1'h1;
  assign _EVAL_499 = _EVAL_685 ? 1'h0 : 1'h1;
  assign _EVAL_525 = {{1'd0}, _EVAL_499};
  assign _EVAL_331 = 2'h2 | _EVAL_525;
  assign _EVAL_854 = _EVAL_635 ? {{1'd0}, _EVAL_261} : _EVAL_331;
  assign _EVAL_839 = {{1'd0}, _EVAL_854};
  assign _EVAL_341 = 3'h4 | _EVAL_839;
  assign _EVAL_688 = _EVAL_380 ? {{1'd0}, _EVAL_400} : _EVAL_341;
  assign _EVAL_596 = {{1'd0}, _EVAL_688};
  assign _EVAL_700 = _EVAL_460 ? 1'h0 : 1'h1;
  assign _EVAL_634 = 2'h2 | _EVAL_566;
  assign _EVAL_788 = _EVAL_272 ? {{1'd0}, _EVAL_700} : _EVAL_634;
  assign _EVAL_740 = _EVAL_182 ? 1'h0 : 1'h1;
  assign _EVAL_132 = _EVAL_875 ? 1'h0 : 1'h1;
  assign _EVAL_529 = {{1'd0}, _EVAL_132};
  assign _EVAL_780 = 2'h2 | _EVAL_529;
  assign _EVAL_654 = _EVAL_354 ? {{1'd0}, _EVAL_740} : _EVAL_780;
  assign _EVAL_133 = {{1'd0}, _EVAL_654};
  assign _EVAL_782 = 3'h4 | _EVAL_133;
  assign _EVAL_571 = _EVAL_461 ? {{1'd0}, _EVAL_788} : _EVAL_782;
  assign _EVAL_622 = 4'h8 | _EVAL_596;
  assign _EVAL_202 = _EVAL_747 ? {{1'd0}, _EVAL_571} : _EVAL_622;
  assign _EVAL_655 = _EVAL_172 ? 1'h0 : 1'h1;
  assign _EVAL_463 = _EVAL_318 ? 1'h0 : 1'h1;
  assign _EVAL_763 = {{1'd0}, _EVAL_463};
  assign _EVAL_696 = 2'h2 | _EVAL_763;
  assign _EVAL_352 = _EVAL_843 ? {{1'd0}, _EVAL_655} : _EVAL_696;
  assign _EVAL_530 = _EVAL_564 ? 1'h0 : 1'h1;
  assign _EVAL_277 = 2'h2 | _EVAL_290;
  assign _EVAL_273 = _EVAL_137 ? {{1'd0}, _EVAL_530} : _EVAL_277;
  assign _EVAL_179 = {{1'd0}, _EVAL_273};
  assign _EVAL_687 = 3'h4 | _EVAL_179;
  assign _EVAL_779 = _EVAL_744 ? {{1'd0}, _EVAL_352} : _EVAL_687;
  assign _EVAL_473 = 4'h8 | _EVAL_756;
  assign _EVAL_677 = _EVAL_591 ? {{1'd0}, _EVAL_779} : _EVAL_473;
  assign _EVAL_793 = {{1'd0}, _EVAL_677};
  assign _EVAL_515 = 5'h10 | _EVAL_793;
  assign _EVAL_271 = _EVAL_374 ? {{1'd0}, _EVAL_202} : _EVAL_515;
  assign _EVAL_309 = {{1'd0}, _EVAL_271};
  assign _EVAL_462 = 6'h20 | _EVAL_309;
  assign _EVAL_828 = _EVAL_276 ? 1'h0 : 1'h1;
  assign _EVAL_867 = _EVAL_769 ? {{1'd0}, _EVAL_828} : _EVAL_471;
  assign _EVAL_671 = _EVAL_374 ? _EVAL_549 : _EVAL_206;
  assign _EVAL_585 = _EVAL_149 >= _EVAL_671;
  assign _EVAL_420 = _EVAL_585 ? _EVAL_149 : _EVAL_671;
  assign _EVAL_148 = _EVAL_260 ? _EVAL_883 : _EVAL_528;
  assign _EVAL_633 = _EVAL_420 >= _EVAL_148;
  assign _EVAL_662 = _EVAL_301 ? {{1'd0}, _EVAL_425} : _EVAL_734;
  assign _EVAL_300 = 4'h8 | _EVAL_445;
  assign _EVAL_888 = _EVAL_255 ? {{1'd0}, _EVAL_662} : _EVAL_300;
  assign _EVAL_556 = 3'h4 | _EVAL_151;
  assign _EVAL_403 = _EVAL_351 ? {{1'd0}, _EVAL_867} : _EVAL_556;
  assign _EVAL_143 = 4'h8 | _EVAL_781;
  assign _EVAL_575 = _EVAL_305 ? {{1'd0}, _EVAL_403} : _EVAL_143;
  assign _EVAL_563 = {{1'd0}, _EVAL_575};
  assign _EVAL_764 = 5'h10 | _EVAL_563;
  assign _EVAL_325 = _EVAL_337 ? {{1'd0}, _EVAL_888} : _EVAL_764;
  assign _EVAL_235 = _EVAL_585 ? {{1'd0}, _EVAL_325} : _EVAL_462;
  assign _EVAL_250 = _EVAL_633 ? _EVAL_420 : _EVAL_148;
  assign _EVAL_32 = _EVAL_250[2:0];
  assign _EVAL_36 = _EVAL_633 ? {{1'd0}, _EVAL_235} : _EVAL_716;
endmodule
