//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_33_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_7,
  input  [3:0]  _EVAL_11,
  input         _EVAL_13,
  input         _EVAL_15,
  input         _EVAL_19,
  input         _EVAL_34,
  input  [2:0]  _EVAL_39,
  input  [6:0]  _EVAL_41,
  input  [30:0] _EVAL_43,
  input         _EVAL_48,
  input         _EVAL_54,
  input  [2:0]  _EVAL_58,
  input         _EVAL_103,
  input  [3:0]  _EVAL_128,
  input  [3:0]  _EVAL_158,
  input  [2:0]  _EVAL_209,
  input         _EVAL_212,
  input  [3:0]  _EVAL_252,
  input         _EVAL_299,
  input  [3:0]  _EVAL_377,
  input         _EVAL_141,
  input         _EVAL_177,
  input         _EVAL_333,
  input         _EVAL_429,
  input         _EVAL_87,
  input         _EVAL_329,
  input         _EVAL_253,
  input         _EVAL_243,
  input         _EVAL_108,
  input         _EVAL_283,
  input         _EVAL_139,
  input         _EVAL_191,
  input         _EVAL_439,
  input         _EVAL_152,
  input         _EVAL_181,
  input  [6:0]  _EVAL_277,
  input         _EVAL_77,
  input         _EVAL_278,
  input         _EVAL_385,
  input         _EVAL_349,
  input         _EVAL_322,
  input         _EVAL_327,
  input  [2:0]  _EVAL_208,
  input  [6:0]  _EVAL_389,
  input  [2:0]  _EVAL_79,
  input         _EVAL_86
);
  wire  TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire [6:0] TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [6:0] TLMonitor__EVAL_7;
  wire [30:0] TLMonitor__EVAL_8;
  wire [2:0] TLMonitor__EVAL_9;
  wire [2:0] TLMonitor__EVAL_10;
  wire [3:0] TLMonitor__EVAL_11;
  wire [2:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire  TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire  _EVAL_437;
  wire  _EVAL_297;
  wire  _EVAL_438;
  wire  _EVAL_132;
  wire  _EVAL_325;
  wire  _EVAL_425;
  wire  _EVAL_106;
  wire  _EVAL_271;
  wire  _EVAL_417;
  wire  _EVAL_237;
  wire  _EVAL_376;
  wire  _EVAL_60;
  wire  _EVAL_127;
  wire  _EVAL_224;
  wire  _EVAL_272;
  wire  _EVAL_233;
  wire  _EVAL_405;
  wire  _EVAL_248;
  wire  _EVAL_140;
  wire  _EVAL_228;
  wire  _EVAL_451;
  wire  _EVAL_358;
  wire  _EVAL_207;
  wire  _EVAL_411;
  wire  _EVAL_375;
  wire  _EVAL_460;
  wire  _EVAL_75;
  wire  _EVAL_213;
  wire  _EVAL_368;
  wire  _EVAL_188;
  wire  _EVAL_372;
  wire  _EVAL_265;
  wire  _EVAL_67;
  wire  _EVAL_122;
  wire  _EVAL_149;
  wire  _EVAL_96;
  wire  _EVAL_174;
  wire  _EVAL_104;
  wire  _EVAL_249;
  wire  _EVAL_260;
  wire  _EVAL_159;
  wire  _EVAL_198;
  wire  _EVAL_354;
  wire  _EVAL_453;
  wire  _EVAL_231;
  wire  _EVAL_98;
  wire  _EVAL_84;
  wire  _EVAL_214;
  wire  _EVAL_367;
  wire  _EVAL_323;
  wire  _EVAL_348;
  wire  _EVAL_217;
  wire  _EVAL_68;
  wire  _EVAL_245;
  wire  _EVAL_221;
  wire  _EVAL_173;
  wire  _EVAL_65;
  wire  _EVAL_257;
  wire  _EVAL_114;
  wire  _EVAL_381;
  wire  _EVAL_412;
  wire  _EVAL_176;
  wire  _EVAL_167;
  wire  _EVAL_80;
  wire  _EVAL_219;
  wire  _EVAL_150;
  wire  _EVAL_193;
  wire  _EVAL_102;
  wire  _EVAL_218;
  wire  _EVAL_107;
  wire  _EVAL_361;
  wire  _EVAL_61;
  wire  _EVAL_115;
  wire  _EVAL_246;
  wire  _EVAL_130;
  wire  _EVAL_269;
  wire  _EVAL_318;
  SiFive__EVAL_30_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16)
  );
  assign _EVAL_437 = _EVAL_177 == 1'h0;
  assign _EVAL_297 = _EVAL_377 != 4'h8;
  assign _EVAL_438 = _EVAL_437 | _EVAL_297;
  assign _EVAL_132 = _EVAL_438 | _EVAL_15;
  assign _EVAL_325 = _EVAL_132 == 1'h0;
  assign _EVAL_425 = _EVAL_87 == 1'h0;
  assign _EVAL_106 = _EVAL_252 != 4'h8;
  assign _EVAL_271 = _EVAL_425 | _EVAL_106;
  assign _EVAL_417 = _EVAL_271 | _EVAL_15;
  assign _EVAL_237 = _EVAL_329 == 1'h0;
  assign _EVAL_376 = _EVAL_128 != 4'h0;
  assign _EVAL_60 = _EVAL_237 | _EVAL_376;
  assign _EVAL_127 = _EVAL_108 == 1'h0;
  assign _EVAL_224 = _EVAL_139 == 1'h0;
  assign _EVAL_272 = _EVAL_209 != 3'h0;
  assign _EVAL_233 = _EVAL_224 | _EVAL_272;
  assign _EVAL_405 = _EVAL_233 | _EVAL_15;
  assign _EVAL_248 = _EVAL_405 == 1'h0;
  assign _EVAL_140 = _EVAL_377 != 4'h0;
  assign _EVAL_228 = _EVAL_152 == 1'h0;
  assign _EVAL_451 = _EVAL_253 == 1'h0;
  assign _EVAL_358 = _EVAL_128 != 4'h8;
  assign _EVAL_207 = _EVAL_451 | _EVAL_358;
  assign _EVAL_411 = _EVAL_243 == 1'h0;
  assign _EVAL_375 = _EVAL_158 != 4'h8;
  assign _EVAL_460 = _EVAL_411 | _EVAL_375;
  assign _EVAL_75 = _EVAL_460 | _EVAL_15;
  assign _EVAL_213 = _EVAL_439 == 1'h0;
  assign _EVAL_368 = _EVAL_212 != 1'h1;
  assign _EVAL_188 = _EVAL_213 | _EVAL_368;
  assign _EVAL_372 = _EVAL_188 | _EVAL_15;
  assign _EVAL_265 = _EVAL_77 == 1'h0;
  assign _EVAL_67 = _EVAL_265 | _EVAL_140;
  assign _EVAL_122 = _EVAL_67 | _EVAL_15;
  assign _EVAL_149 = _EVAL_122 == 1'h0;
  assign _EVAL_96 = _EVAL_278 == 1'h0;
  assign _EVAL_174 = _EVAL_299 != 1'h1;
  assign _EVAL_104 = _EVAL_96 | _EVAL_174;
  assign _EVAL_249 = _EVAL_104 | _EVAL_15;
  assign _EVAL_260 = _EVAL_385 == 1'h0;
  assign _EVAL_159 = _EVAL_252 != 4'h0;
  assign _EVAL_198 = _EVAL_260 | _EVAL_159;
  assign _EVAL_354 = _EVAL_349 == 1'h0;
  assign _EVAL_453 = _EVAL_354 | _EVAL_212;
  assign _EVAL_231 = _EVAL_429 == 1'h0;
  assign _EVAL_98 = _EVAL_231 | _EVAL_299;
  assign _EVAL_84 = _EVAL_98 | _EVAL_15;
  assign _EVAL_214 = _EVAL_84 == 1'h0;
  assign _EVAL_367 = _EVAL_322 == 1'h0;
  assign _EVAL_323 = _EVAL_367 | _EVAL_103;
  assign _EVAL_348 = _EVAL_60 | _EVAL_15;
  assign _EVAL_217 = _EVAL_348 == 1'h0;
  assign _EVAL_68 = _EVAL_75 == 1'h0;
  assign _EVAL_245 = _EVAL_198 | _EVAL_15;
  assign _EVAL_221 = _EVAL_181 == 1'h0;
  assign _EVAL_173 = _EVAL_103 != 1'h1;
  assign _EVAL_65 = _EVAL_221 | _EVAL_173;
  assign _EVAL_257 = _EVAL_158 != 4'h0;
  assign _EVAL_114 = _EVAL_127 | _EVAL_257;
  assign _EVAL_381 = _EVAL_114 | _EVAL_15;
  assign _EVAL_412 = _EVAL_381 == 1'h0;
  assign _EVAL_176 = _EVAL_249 == 1'h0;
  assign _EVAL_167 = _EVAL_209 != 3'h7;
  assign _EVAL_80 = _EVAL_228 | _EVAL_167;
  assign _EVAL_219 = _EVAL_245 == 1'h0;
  assign _EVAL_150 = _EVAL_80 | _EVAL_15;
  assign _EVAL_193 = _EVAL_65 | _EVAL_15;
  assign _EVAL_102 = _EVAL_193 == 1'h0;
  assign _EVAL_218 = _EVAL_372 == 1'h0;
  assign _EVAL_107 = _EVAL_207 | _EVAL_15;
  assign _EVAL_361 = _EVAL_323 | _EVAL_15;
  assign _EVAL_61 = _EVAL_361 == 1'h0;
  assign _EVAL_115 = _EVAL_107 == 1'h0;
  assign _EVAL_246 = _EVAL_453 | _EVAL_15;
  assign _EVAL_130 = _EVAL_246 == 1'h0;
  assign _EVAL_269 = _EVAL_150 == 1'h0;
  assign _EVAL_318 = _EVAL_417 == 1'h0;
  assign TLMonitor__EVAL_16 = _EVAL_333 ? _EVAL_327 : 1'h0;
  assign TLMonitor__EVAL_10 = _EVAL_39;
  assign TLMonitor__EVAL_6 = _EVAL_19;
  assign TLMonitor__EVAL = _EVAL_333 ? _EVAL_191 : _EVAL_86;
  assign TLMonitor__EVAL_12 = _EVAL_333 ? 3'h1 : 3'h0;
  assign TLMonitor__EVAL_14 = _EVAL_13;
  assign TLMonitor__EVAL_3 = _EVAL_7;
  assign TLMonitor__EVAL_1 = _EVAL_333 ? _EVAL : _EVAL_48;
  assign TLMonitor__EVAL_8 = _EVAL_43;
  assign TLMonitor__EVAL_13 = _EVAL_15;
  assign TLMonitor__EVAL_5 = _EVAL_41;
  assign TLMonitor__EVAL_9 = _EVAL_58;
  assign TLMonitor__EVAL_11 = _EVAL_11;
  assign TLMonitor__EVAL_15 = _EVAL_141 & _EVAL_283;
  assign TLMonitor__EVAL_2 = _EVAL_333 ? _EVAL_208 : _EVAL_79;
  assign TLMonitor__EVAL_4 = _EVAL_54;
  assign TLMonitor__EVAL_7 = _EVAL_333 ? _EVAL_389 : _EVAL_277;
  assign TLMonitor__EVAL_0 = _EVAL_34;
  always @(posedge _EVAL_54) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6634d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e96417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
