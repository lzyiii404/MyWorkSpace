//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_122(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [1:0]  _EVAL_3,
  output        _EVAL_4,
  output [1:0]  _EVAL_5,
  input  [6:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  output [29:0] _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  output [3:0]  _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  output [31:0] _EVAL_19,
  input         _EVAL_20,
  input  [6:0]  _EVAL_21,
  output [6:0]  _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output [3:0]  _EVAL_25,
  input         _EVAL_26,
  input  [29:0] _EVAL_27,
  output [31:0] _EVAL_28,
  input  [3:0]  _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  output [6:0]  _EVAL_33,
  output        _EVAL_34,
  output [3:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  input  [3:0]  _EVAL_37,
  input         _EVAL_38,
  input  [31:0] _EVAL_39,
  input  [2:0]  _EVAL_40
);
  reg [2:0] _EVAL_41;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_46;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_53;
  reg [31:0] _RAND_2;
  reg [5:0] _EVAL_54;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_88;
  reg [31:0] _RAND_4;
  reg  _EVAL_128;
  reg [31:0] _RAND_5;
  reg [29:0] _EVAL_130;
  reg [31:0] _RAND_6;
  reg [6:0] _EVAL_176;
  reg [31:0] _RAND_7;
  reg  _EVAL_262;
  reg [31:0] _RAND_8;
  reg  _EVAL_273;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_298;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_299;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_312;
  reg [31:0] _RAND_12;
  reg  _EVAL_327;
  reg [31:0] _RAND_13;
  reg  _EVAL_368;
  reg [31:0] _RAND_14;
  reg [3:0] _EVAL_394;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_402;
  reg [31:0] _RAND_16;
  wire  _EVAL_348;
  wire [1:0] _EVAL_435;
  wire [2:0] _EVAL_114;
  wire  _EVAL_265;
  wire  _EVAL_439;
  wire  _EVAL_155;
  wire [1:0] _EVAL_178;
  wire [3:0] _EVAL_307;
  wire  _EVAL_48;
  wire  _EVAL_177;
  wire  _EVAL_99;
  wire  _EVAL_405;
  wire  _EVAL_329;
  wire  _EVAL_264;
  wire  _EVAL_416;
  wire  _EVAL_425;
  wire  _EVAL_444;
  wire  _EVAL_76;
  wire  _EVAL_140;
  wire  _EVAL_304;
  wire  _EVAL_52;
  wire [29:0] _EVAL_430;
  wire [30:0] _EVAL_212;
  wire [30:0] _EVAL_75;
  wire [30:0] _EVAL_144;
  wire  _EVAL_228;
  wire [29:0] _EVAL_68;
  wire [30:0] _EVAL_452;
  wire [30:0] _EVAL_183;
  wire [30:0] _EVAL_162;
  wire  _EVAL_384;
  wire  _EVAL_168;
  wire  _EVAL_214;
  wire  _EVAL_106;
  wire  _EVAL_352;
  wire  _EVAL_198;
  wire  _EVAL_283;
  wire  _EVAL_375;
  wire  _EVAL_236;
  wire [1:0] _EVAL_401;
  wire [2:0] _EVAL_119;
  wire [1:0] _EVAL_80;
  wire [1:0] _EVAL_388;
  wire [2:0] _EVAL_163;
  wire [1:0] _EVAL_284;
  wire [1:0] _EVAL_81;
  wire  _EVAL_72;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_279;
  wire  _EVAL_87;
  wire  _EVAL_440;
  wire  _EVAL_453;
  wire  _EVAL_121;
  wire  _EVAL_126;
  wire  _EVAL_377;
  wire  _EVAL_175;
  wire  _EVAL_325;
  wire  _EVAL_445;
  wire  _EVAL_373;
  wire [3:0] _EVAL_446;
  wire [3:0] _EVAL_266;
  wire [2:0] _EVAL_259;
  wire [3:0] _EVAL_256;
  wire [3:0] _EVAL_105;
  wire [3:0] _EVAL_196;
  wire [3:0] _EVAL_448;
  wire [4:0] _EVAL_393;
  wire [3:0] _EVAL_240;
  wire [4:0] _EVAL_152;
  wire [3:0] _EVAL_172;
  wire [3:0] _EVAL_267;
  wire [5:0] _EVAL_142;
  wire [3:0] _EVAL_79;
  wire [3:0] _EVAL_367;
  wire  _EVAL_56;
  wire  _EVAL_213;
  wire  _EVAL_255;
  wire [1:0] _EVAL_109;
  wire  _EVAL_277;
  wire  _EVAL_363;
  wire  _EVAL_409;
  wire  _EVAL_231;
  wire  _EVAL_138;
  wire  _EVAL_417;
  wire [1:0] _EVAL_245;
  wire [3:0] _EVAL_376;
  wire  _EVAL_62;
  wire  _EVAL_171;
  wire [1:0] _EVAL_252;
  wire [3:0] _EVAL_195;
  wire  _EVAL_167;
  wire  _EVAL_282;
  wire  _EVAL_64;
  wire  _EVAL_156;
  wire [1:0] _EVAL_47;
  wire  _EVAL_258;
  wire  _EVAL_151;
  wire  _EVAL_60;
  wire  _EVAL_449;
  wire  _EVAL_451;
  wire [3:0] _EVAL_50;
  wire [3:0] _EVAL_441;
  wire  _EVAL_428;
  wire  _EVAL_408;
  wire  _EVAL_173;
  wire [1:0] _EVAL_410;
  wire  _EVAL_386;
  wire  _EVAL_235;
  wire  _EVAL_129;
  wire [1:0] _EVAL_349;
  wire [3:0] _EVAL_170;
  wire  _EVAL_92;
  wire  _EVAL_45;
  wire  _EVAL_334;
  wire [22:0] _EVAL_357;
  wire [7:0] _EVAL_51;
  wire [7:0] _EVAL_225;
  wire [5:0] _EVAL_74;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_320;
  wire  _EVAL_174;
  wire  _EVAL_274;
  wire [5:0] _EVAL_339;
  wire [5:0] _EVAL_455;
  wire  _EVAL_355;
  wire  _EVAL_397;
  wire [1:0] _EVAL_341;
  wire [3:0] _EVAL_165;
  wire  _EVAL_362;
  wire [2:0] _EVAL_281;
  wire  _EVAL_261;
  wire  _EVAL_276;
  wire  _EVAL_100;
  wire [1:0] _EVAL_238;
  wire [3:0] _EVAL_331;
  wire  _EVAL_94;
  wire  _EVAL_422;
  wire  _EVAL_250;
  wire  _EVAL_280;
  wire  _EVAL_118;
  wire  _EVAL_104;
  wire [7:0] _EVAL_292;
  wire  _EVAL_420;
  wire [7:0] _EVAL_319;
  wire  _EVAL_189;
  wire [7:0] _EVAL_147;
  wire  _EVAL_103;
  wire [7:0] _EVAL_137;
  wire [31:0] _EVAL_407;
  wire [31:0] _EVAL_318;
  wire  _EVAL_434;
  wire [7:0] _EVAL_101;
  wire  _EVAL_188;
  wire [7:0] _EVAL_44;
  wire  _EVAL_223;
  wire [7:0] _EVAL_57;
  wire [7:0] _EVAL_169;
  wire [31:0] _EVAL_447;
  wire [31:0] _EVAL_316;
  wire  _EVAL_239;
  wire [31:0] _EVAL_396;
  wire [4:0] _EVAL_233;
  wire [3:0] _EVAL_197;
  wire [4:0] _EVAL_66;
  wire [3:0] _EVAL_346;
  wire [3:0] _EVAL_153;
  wire [5:0] _EVAL_356;
  wire [3:0] _EVAL_55;
  wire [3:0] _EVAL_326;
  wire  _EVAL_458;
  wire [7:0] _EVAL_350;
  wire  _EVAL_49;
  wire [7:0] _EVAL_414;
  wire  _EVAL_260;
  wire [7:0] _EVAL_359;
  wire  _EVAL_110;
  wire [7:0] _EVAL_303;
  wire [31:0] _EVAL_86;
  wire [31:0] _EVAL_310;
  wire [31:0] _EVAL_323;
  wire [31:0] _EVAL_215;
  wire [31:0] _EVAL_395;
  wire  _EVAL_131;
  wire [22:0] _EVAL_457;
  wire [7:0] _EVAL_371;
  wire  _EVAL_297;
  wire [1:0] _EVAL_125;
  wire  _EVAL_220;
  wire  _EVAL_436;
  wire  _EVAL_324;
  wire  _EVAL_379;
  wire  _EVAL_290;
  wire  _EVAL_450;
  wire  _EVAL_221;
  wire  _EVAL_124;
  wire  _EVAL_313;
  wire  _EVAL_248;
  wire  _EVAL_432;
  wire  _EVAL_166;
  wire [1:0] _EVAL_161;
  wire  _EVAL_460;
  wire [1:0] _EVAL_263;
  wire [3:0] _EVAL_95;
  wire  _EVAL_205;
  wire  _EVAL_70;
  wire [1:0] _EVAL_365;
  wire [3:0] _EVAL_187;
  wire  _EVAL_180;
  wire  _EVAL_257;
  wire [1:0] _EVAL_433;
  wire [3:0] _EVAL_226;
  wire  _EVAL_73;
  wire  _EVAL_333;
  wire [1:0] _EVAL_275;
  wire [3:0] _EVAL_421;
  wire  _EVAL_400;
  wire [3:0] _EVAL_201;
  wire  _EVAL_443;
  wire [3:0] _EVAL_360;
  wire  _EVAL_65;
  wire [3:0] _EVAL_314;
  wire  _EVAL_102;
  wire [3:0] _EVAL_438;
  wire  _EVAL_383;
  wire  _EVAL_111;
  wire  _EVAL_157;
  wire [1:0] _EVAL_192;
  wire [3:0] _EVAL_202;
  wire  _EVAL_286;
  wire [1:0] _EVAL_200;
  wire [3:0] _EVAL_154;
  wire  _EVAL_454;
  wire  _EVAL_305;
  wire  _EVAL_302;
  wire [1:0] _EVAL_296;
  wire [3:0] _EVAL_251;
  wire  _EVAL_399;
  wire  _EVAL_387;
  wire  _EVAL_193;
  wire [1:0] _EVAL_123;
  wire [3:0] _EVAL_224;
  wire  _EVAL_77;
  wire  _EVAL_403;
  wire [1:0] _EVAL_97;
  wire [3:0] _EVAL_269;
  wire  _EVAL_158;
  wire  _EVAL_271;
  wire [1:0] _EVAL_229;
  wire [3:0] _EVAL_404;
  wire  _EVAL_308;
  wire  _EVAL_364;
  wire  _EVAL_218;
  wire [1:0] _EVAL_160;
  wire [3:0] _EVAL_372;
  wire  _EVAL_419;
  wire [7:0] _EVAL_84;
  wire [1:0] _EVAL_69;
  wire [3:0] _EVAL_242;
  wire  _EVAL_342;
  wire  _EVAL_391;
  wire  _EVAL_217;
  wire [1:0] _EVAL_164;
  wire [3:0] _EVAL_61;
  wire  _EVAL_423;
  wire  _EVAL_83;
  wire  _EVAL_317;
  wire [1:0] _EVAL_429;
  wire [3:0] _EVAL_254;
  wire  _EVAL_456;
  wire  _EVAL_115;
  wire [3:0] _EVAL_134;
  wire  _EVAL_148;
  wire  _EVAL_322;
  wire  _EVAL_415;
  wire [1:0] _EVAL_190;
  wire [3:0] _EVAL_358;
  wire  _EVAL_431;
  wire  _EVAL_90;
  wire [1:0] _EVAL_389;
  wire [3:0] _EVAL_340;
  wire  _EVAL_203;
  wire  _EVAL_122;
  wire  _EVAL_347;
  wire [1:0] _EVAL_361;
  wire [3:0] _EVAL_232;
  wire  _EVAL_335;
  wire  _EVAL_78;
  wire [1:0] _EVAL_207;
  wire [3:0] _EVAL_234;
  wire  _EVAL_59;
  wire  _EVAL_442;
  wire  _EVAL_288;
  wire [1:0] _EVAL_390;
  wire [3:0] _EVAL_427;
  wire  _EVAL_146;
  wire  _EVAL_332;
  wire  _EVAL_133;
  wire [1:0] _EVAL_398;
  wire [3:0] _EVAL_413;
  wire  _EVAL_150;
  wire  _EVAL_344;
  wire  _EVAL_353;
  wire [1:0] _EVAL_241;
  wire [3:0] _EVAL_306;
  wire  _EVAL_462;
  wire [7:0] _EVAL_243;
  wire [15:0] _EVAL_437;
  wire [31:0] _EVAL_108;
  wire [31:0] _EVAL_209;
  wire [31:0] _EVAL_315;
  wire [31:0] _EVAL_143;
  wire [7:0] _EVAL_378;
  wire [5:0] _EVAL_211;
  wire [5:0] _EVAL_204;
  wire  _EVAL_321;
  wire [1:0] _EVAL_424;
  wire [1:0] _EVAL_96;
  wire  _EVAL_222;
  wire  _EVAL_291;
  wire  _EVAL_184;
  wire  _EVAL_345;
  wire  _EVAL_210;
  wire  _EVAL_244;
  wire  _EVAL_186;
  wire  _EVAL_149;
  wire  _EVAL_380;
  wire  _EVAL_385;
  wire  _EVAL_366;
  wire  _EVAL_268;
  wire  _EVAL_370;
  wire  _EVAL_43;
  wire  _EVAL_116;
  wire  _EVAL_42;
  wire  _EVAL_107;
  wire  _EVAL_270;
  wire  _EVAL_295;
  wire  _EVAL_330;
  wire  _EVAL_351;
  wire [2:0] _EVAL_112;
  wire [83:0] _EVAL_117;
  wire  _EVAL_336;
  wire  _EVAL_369;
  wire  _EVAL_278;
  wire  _EVAL_411;
  wire  _EVAL_253;
  wire  _EVAL_301;
  wire  _EVAL_392;
  wire  _EVAL_459;
  wire  _EVAL_141;
  wire  _EVAL_294;
  wire  _EVAL_93;
  wire  _EVAL_199;
  wire  _EVAL_289;
  wire [83:0] _EVAL_328;
  wire [83:0] _EVAL_309;
  wire  _EVAL_412;
  wire [83:0] _EVAL_132;
  wire [83:0] _EVAL_381;
  wire  _EVAL_237;
  wire  _EVAL_139;
  wire  _EVAL_206;
  assign _EVAL_348 = _EVAL_46[21];
  assign _EVAL_435 = _EVAL_14[1:0];
  assign _EVAL_114 = {{1'd0}, _EVAL_435};
  assign _EVAL_265 = 3'h2 == _EVAL_114;
  assign _EVAL_439 = _EVAL_46[6];
  assign _EVAL_155 = _EVAL_312[6];
  assign _EVAL_178 = {_EVAL_439,_EVAL_155};
  assign _EVAL_307 = _EVAL_299 >> _EVAL_178;
  assign _EVAL_48 = _EVAL_307[0];
  assign _EVAL_177 = _EVAL_88 == 2'h0;
  assign _EVAL_99 = _EVAL_176 == _EVAL_6;
  assign _EVAL_405 = _EVAL_88 != 2'h0;
  assign _EVAL_329 = _EVAL_99 & _EVAL_405;
  assign _EVAL_264 = _EVAL_12 == 3'h1;
  assign _EVAL_416 = _EVAL_298 == 6'h0;
  assign _EVAL_425 = _EVAL_88 == 2'h3;
  assign _EVAL_444 = _EVAL_88 == 2'h2;
  assign _EVAL_76 = _EVAL_425 | _EVAL_444;
  assign _EVAL_140 = _EVAL_76 == 1'h0;
  assign _EVAL_304 = _EVAL_40 == 3'h3;
  assign _EVAL_52 = _EVAL_13 <= 4'h2;
  assign _EVAL_430 = _EVAL_27 ^ 30'h1000;
  assign _EVAL_212 = {1'b0,$signed(_EVAL_430)};
  assign _EVAL_75 = $signed(_EVAL_212) & $signed(31'sh2b101000);
  assign _EVAL_144 = $signed(_EVAL_75);
  assign _EVAL_228 = $signed(_EVAL_144) == $signed(31'sh0);
  assign _EVAL_68 = _EVAL_27 ^ 30'h1100000;
  assign _EVAL_452 = {1'b0,$signed(_EVAL_68)};
  assign _EVAL_183 = $signed(_EVAL_452) & $signed(31'sh2b100000);
  assign _EVAL_162 = $signed(_EVAL_183);
  assign _EVAL_384 = $signed(_EVAL_162) == $signed(31'sh0);
  assign _EVAL_168 = _EVAL_228 | _EVAL_384;
  assign _EVAL_214 = _EVAL_52 & _EVAL_168;
  assign _EVAL_106 = _EVAL_40 == 3'h2;
  assign _EVAL_352 = _EVAL_106 ? _EVAL_214 : 1'h1;
  assign _EVAL_198 = _EVAL_304 ? _EVAL_214 : _EVAL_352;
  assign _EVAL_283 = _EVAL_198 | _EVAL_177;
  assign _EVAL_375 = _EVAL_140 & _EVAL_283;
  assign _EVAL_236 = _EVAL_2 & _EVAL_375;
  assign _EVAL_401 = {_EVAL_236,_EVAL_444};
  assign _EVAL_119 = {_EVAL_401, 1'h0};
  assign _EVAL_80 = _EVAL_119[1:0];
  assign _EVAL_388 = _EVAL_401 | _EVAL_80;
  assign _EVAL_163 = {_EVAL_388, 1'h0};
  assign _EVAL_284 = _EVAL_163[1:0];
  assign _EVAL_81 = ~ _EVAL_284;
  assign _EVAL_72 = _EVAL_81[0];
  assign _EVAL_246 = _EVAL_416 ? _EVAL_72 : _EVAL_327;
  assign _EVAL_247 = _EVAL_26 & _EVAL_246;
  assign _EVAL_279 = _EVAL_247 & _EVAL_444;
  assign _EVAL_87 = _EVAL_81[1];
  assign _EVAL_440 = _EVAL_416 ? _EVAL_87 : _EVAL_368;
  assign _EVAL_453 = _EVAL_26 & _EVAL_440;
  assign _EVAL_121 = _EVAL_453 & _EVAL_236;
  assign _EVAL_126 = _EVAL_198 == 1'h0;
  assign _EVAL_377 = _EVAL_121 & _EVAL_126;
  assign _EVAL_175 = _EVAL_46[31];
  assign _EVAL_325 = _EVAL_46[23];
  assign _EVAL_445 = _EVAL_46[15];
  assign _EVAL_373 = _EVAL_46[7];
  assign _EVAL_446 = {_EVAL_175,_EVAL_325,_EVAL_445,_EVAL_373};
  assign _EVAL_266 = ~ _EVAL_394;
  assign _EVAL_259 = _EVAL_394[3:1];
  assign _EVAL_256 = {{1'd0}, _EVAL_259};
  assign _EVAL_105 = _EVAL_266 | _EVAL_256;
  assign _EVAL_196 = ~ _EVAL_105;
  assign _EVAL_448 = _EVAL_446 & _EVAL_196;
  assign _EVAL_393 = {_EVAL_448, 1'h0};
  assign _EVAL_240 = _EVAL_393[3:0];
  assign _EVAL_152 = {_EVAL_240, 1'h0};
  assign _EVAL_172 = _EVAL_152[3:0];
  assign _EVAL_267 = _EVAL_240 | _EVAL_172;
  assign _EVAL_142 = {_EVAL_267, 2'h0};
  assign _EVAL_79 = _EVAL_142[3:0];
  assign _EVAL_367 = _EVAL_267 | _EVAL_79;
  assign _EVAL_56 = _EVAL_367[0];
  assign _EVAL_213 = _EVAL_46[11];
  assign _EVAL_255 = _EVAL_312[11];
  assign _EVAL_109 = {_EVAL_213,_EVAL_255};
  assign _EVAL_277 = _EVAL_46[12];
  assign _EVAL_363 = _EVAL_444 | _EVAL_236;
  assign _EVAL_409 = _EVAL_72 & _EVAL_444;
  assign _EVAL_231 = _EVAL_87 & _EVAL_236;
  assign _EVAL_138 = _EVAL_46[22];
  assign _EVAL_417 = _EVAL_312[22];
  assign _EVAL_245 = {_EVAL_138,_EVAL_417};
  assign _EVAL_376 = _EVAL_299 >> _EVAL_245;
  assign _EVAL_62 = _EVAL_46[24];
  assign _EVAL_171 = _EVAL_312[24];
  assign _EVAL_252 = {_EVAL_62,_EVAL_171};
  assign _EVAL_195 = _EVAL_299 >> _EVAL_252;
  assign _EVAL_167 = _EVAL_195[0];
  assign _EVAL_282 = _EVAL_376[0];
  assign _EVAL_64 = _EVAL_46[28];
  assign _EVAL_156 = _EVAL_312[28];
  assign _EVAL_47 = {_EVAL_64,_EVAL_156};
  assign _EVAL_258 = _EVAL_402[0];
  assign _EVAL_151 = _EVAL_312[31];
  assign _EVAL_60 = _EVAL_312[23];
  assign _EVAL_449 = _EVAL_312[15];
  assign _EVAL_451 = _EVAL_312[7];
  assign _EVAL_50 = {_EVAL_151,_EVAL_60,_EVAL_449,_EVAL_451};
  assign _EVAL_441 = _EVAL_50 & _EVAL_196;
  assign _EVAL_428 = _EVAL_312[2];
  assign _EVAL_408 = _EVAL_46[29];
  assign _EVAL_173 = _EVAL_312[29];
  assign _EVAL_410 = {_EVAL_408,_EVAL_173};
  assign _EVAL_386 = _EVAL_329 & _EVAL_264;
  assign _EVAL_235 = _EVAL_46[8];
  assign _EVAL_129 = _EVAL_312[8];
  assign _EVAL_349 = {_EVAL_235,_EVAL_129};
  assign _EVAL_170 = _EVAL_299 >> _EVAL_349;
  assign _EVAL_92 = _EVAL_416 & _EVAL_26;
  assign _EVAL_45 = _EVAL_40[2];
  assign _EVAL_334 = _EVAL_45 == 1'h0;
  assign _EVAL_357 = 23'hff << _EVAL_13;
  assign _EVAL_51 = _EVAL_357[7:0];
  assign _EVAL_225 = ~ _EVAL_51;
  assign _EVAL_74 = _EVAL_225[7:2];
  assign _EVAL_179 = _EVAL_327 ? _EVAL_444 : 1'h0;
  assign _EVAL_181 = _EVAL_368 ? _EVAL_236 : 1'h0;
  assign _EVAL_320 = _EVAL_179 | _EVAL_181;
  assign _EVAL_174 = _EVAL_416 ? _EVAL_363 : _EVAL_320;
  assign _EVAL_274 = _EVAL_26 & _EVAL_174;
  assign _EVAL_339 = {{5'd0}, _EVAL_274};
  assign _EVAL_455 = _EVAL_298 - _EVAL_339;
  assign _EVAL_355 = _EVAL_46[30];
  assign _EVAL_397 = _EVAL_312[30];
  assign _EVAL_341 = {_EVAL_355,_EVAL_397};
  assign _EVAL_165 = _EVAL_299 >> _EVAL_341;
  assign _EVAL_362 = _EVAL_165[0];
  assign _EVAL_281 = _EVAL_126 ? 3'h0 : _EVAL_14;
  assign _EVAL_261 = _EVAL_46[27];
  assign _EVAL_276 = _EVAL_46[4];
  assign _EVAL_100 = _EVAL_46[2];
  assign _EVAL_238 = {_EVAL_100,_EVAL_428};
  assign _EVAL_331 = _EVAL_299 >> _EVAL_238;
  assign _EVAL_94 = _EVAL_331[0];
  assign _EVAL_422 = _EVAL_312[18];
  assign _EVAL_250 = _EVAL_41[0];
  assign _EVAL_280 = _EVAL_54 == 6'h0;
  assign _EVAL_118 = _EVAL_280 & _EVAL_264;
  assign _EVAL_104 = _EVAL_394[3];
  assign _EVAL_292 = _EVAL_104 ? 8'hff : 8'h0;
  assign _EVAL_420 = _EVAL_394[2];
  assign _EVAL_319 = _EVAL_420 ? 8'hff : 8'h0;
  assign _EVAL_189 = _EVAL_394[1];
  assign _EVAL_147 = _EVAL_189 ? 8'hff : 8'h0;
  assign _EVAL_103 = _EVAL_394[0];
  assign _EVAL_137 = _EVAL_103 ? 8'hff : 8'h0;
  assign _EVAL_407 = {_EVAL_292,_EVAL_319,_EVAL_147,_EVAL_137};
  assign _EVAL_318 = _EVAL_46 & _EVAL_407;
  assign _EVAL_434 = _EVAL_367[3];
  assign _EVAL_101 = _EVAL_434 ? 8'hff : 8'h0;
  assign _EVAL_188 = _EVAL_367[2];
  assign _EVAL_44 = _EVAL_188 ? 8'hff : 8'h0;
  assign _EVAL_223 = _EVAL_367[1];
  assign _EVAL_57 = _EVAL_223 ? 8'hff : 8'h0;
  assign _EVAL_169 = _EVAL_56 ? 8'hff : 8'h0;
  assign _EVAL_447 = {_EVAL_101,_EVAL_44,_EVAL_57,_EVAL_169};
  assign _EVAL_316 = _EVAL_318 | _EVAL_447;
  assign _EVAL_239 = _EVAL_41[2];
  assign _EVAL_396 = _EVAL_312 & _EVAL_407;
  assign _EVAL_233 = {_EVAL_441, 1'h0};
  assign _EVAL_197 = _EVAL_233[3:0];
  assign _EVAL_66 = {_EVAL_197, 1'h0};
  assign _EVAL_346 = _EVAL_66[3:0];
  assign _EVAL_153 = _EVAL_197 | _EVAL_346;
  assign _EVAL_356 = {_EVAL_153, 2'h0};
  assign _EVAL_55 = _EVAL_356[3:0];
  assign _EVAL_326 = _EVAL_153 | _EVAL_55;
  assign _EVAL_458 = _EVAL_326[3];
  assign _EVAL_350 = _EVAL_458 ? 8'hff : 8'h0;
  assign _EVAL_49 = _EVAL_326[2];
  assign _EVAL_414 = _EVAL_49 ? 8'hff : 8'h0;
  assign _EVAL_260 = _EVAL_326[1];
  assign _EVAL_359 = _EVAL_260 ? 8'hff : 8'h0;
  assign _EVAL_110 = _EVAL_326[0];
  assign _EVAL_303 = _EVAL_110 ? 8'hff : 8'h0;
  assign _EVAL_86 = {_EVAL_350,_EVAL_414,_EVAL_359,_EVAL_303};
  assign _EVAL_310 = _EVAL_396 | _EVAL_86;
  assign _EVAL_323 = ~ _EVAL_310;
  assign _EVAL_215 = _EVAL_239 ? _EVAL_310 : _EVAL_323;
  assign _EVAL_395 = _EVAL_316 + _EVAL_215;
  assign _EVAL_131 = 3'h3 == _EVAL_114;
  assign _EVAL_457 = 23'hff << _EVAL_37;
  assign _EVAL_371 = _EVAL_457[7:0];
  assign _EVAL_297 = _EVAL_312[27];
  assign _EVAL_125 = {_EVAL_261,_EVAL_297};
  assign _EVAL_220 = _EVAL_46[17];
  assign _EVAL_436 = _EVAL_316[31];
  assign _EVAL_324 = _EVAL_310[31];
  assign _EVAL_379 = _EVAL_436 == _EVAL_324;
  assign _EVAL_290 = _EVAL_395[31];
  assign _EVAL_450 = _EVAL_290 == 1'h0;
  assign _EVAL_221 = _EVAL_41[1];
  assign _EVAL_124 = _EVAL_221 == _EVAL_436;
  assign _EVAL_313 = _EVAL_379 ? _EVAL_450 : _EVAL_124;
  assign _EVAL_248 = _EVAL_250 == _EVAL_313;
  assign _EVAL_432 = _EVAL_46[26];
  assign _EVAL_166 = _EVAL_312[26];
  assign _EVAL_161 = {_EVAL_432,_EVAL_166};
  assign _EVAL_460 = _EVAL_312[12];
  assign _EVAL_263 = {_EVAL_277,_EVAL_460};
  assign _EVAL_95 = _EVAL_299 >> _EVAL_263;
  assign _EVAL_205 = _EVAL_46[9];
  assign _EVAL_70 = _EVAL_312[9];
  assign _EVAL_365 = {_EVAL_205,_EVAL_70};
  assign _EVAL_187 = _EVAL_299 >> _EVAL_365;
  assign _EVAL_180 = _EVAL_187[0];
  assign _EVAL_257 = _EVAL_312[21];
  assign _EVAL_433 = {_EVAL_348,_EVAL_257};
  assign _EVAL_226 = _EVAL_299 >> _EVAL_433;
  assign _EVAL_73 = _EVAL_226[0];
  assign _EVAL_333 = _EVAL_53[0];
  assign _EVAL_275 = {_EVAL_175,_EVAL_151};
  assign _EVAL_421 = _EVAL_299 >> _EVAL_275;
  assign _EVAL_400 = _EVAL_421[0];
  assign _EVAL_201 = _EVAL_299 >> _EVAL_410;
  assign _EVAL_443 = _EVAL_201[0];
  assign _EVAL_360 = _EVAL_299 >> _EVAL_47;
  assign _EVAL_65 = _EVAL_360[0];
  assign _EVAL_314 = _EVAL_299 >> _EVAL_125;
  assign _EVAL_102 = _EVAL_314[0];
  assign _EVAL_438 = _EVAL_299 >> _EVAL_161;
  assign _EVAL_383 = _EVAL_438[0];
  assign _EVAL_111 = _EVAL_46[25];
  assign _EVAL_157 = _EVAL_312[25];
  assign _EVAL_192 = {_EVAL_111,_EVAL_157};
  assign _EVAL_202 = _EVAL_299 >> _EVAL_192;
  assign _EVAL_286 = _EVAL_202[0];
  assign _EVAL_200 = {_EVAL_325,_EVAL_60};
  assign _EVAL_154 = _EVAL_299 >> _EVAL_200;
  assign _EVAL_454 = _EVAL_154[0];
  assign _EVAL_305 = _EVAL_46[20];
  assign _EVAL_302 = _EVAL_312[20];
  assign _EVAL_296 = {_EVAL_305,_EVAL_302};
  assign _EVAL_251 = _EVAL_299 >> _EVAL_296;
  assign _EVAL_399 = _EVAL_251[0];
  assign _EVAL_387 = _EVAL_46[19];
  assign _EVAL_193 = _EVAL_312[19];
  assign _EVAL_123 = {_EVAL_387,_EVAL_193};
  assign _EVAL_224 = _EVAL_299 >> _EVAL_123;
  assign _EVAL_77 = _EVAL_224[0];
  assign _EVAL_403 = _EVAL_46[18];
  assign _EVAL_97 = {_EVAL_403,_EVAL_422};
  assign _EVAL_269 = _EVAL_299 >> _EVAL_97;
  assign _EVAL_158 = _EVAL_269[0];
  assign _EVAL_271 = _EVAL_312[17];
  assign _EVAL_229 = {_EVAL_220,_EVAL_271};
  assign _EVAL_404 = _EVAL_299 >> _EVAL_229;
  assign _EVAL_308 = _EVAL_404[0];
  assign _EVAL_364 = _EVAL_46[16];
  assign _EVAL_218 = _EVAL_312[16];
  assign _EVAL_160 = {_EVAL_364,_EVAL_218};
  assign _EVAL_372 = _EVAL_299 >> _EVAL_160;
  assign _EVAL_419 = _EVAL_372[0];
  assign _EVAL_84 = {_EVAL_454,_EVAL_282,_EVAL_73,_EVAL_399,_EVAL_77,_EVAL_158,_EVAL_308,_EVAL_419};
  assign _EVAL_69 = {_EVAL_445,_EVAL_449};
  assign _EVAL_242 = _EVAL_299 >> _EVAL_69;
  assign _EVAL_342 = _EVAL_242[0];
  assign _EVAL_391 = _EVAL_46[14];
  assign _EVAL_217 = _EVAL_312[14];
  assign _EVAL_164 = {_EVAL_391,_EVAL_217};
  assign _EVAL_61 = _EVAL_299 >> _EVAL_164;
  assign _EVAL_423 = _EVAL_61[0];
  assign _EVAL_83 = _EVAL_46[13];
  assign _EVAL_317 = _EVAL_312[13];
  assign _EVAL_429 = {_EVAL_83,_EVAL_317};
  assign _EVAL_254 = _EVAL_299 >> _EVAL_429;
  assign _EVAL_456 = _EVAL_254[0];
  assign _EVAL_115 = _EVAL_95[0];
  assign _EVAL_134 = _EVAL_299 >> _EVAL_109;
  assign _EVAL_148 = _EVAL_134[0];
  assign _EVAL_322 = _EVAL_46[10];
  assign _EVAL_415 = _EVAL_312[10];
  assign _EVAL_190 = {_EVAL_322,_EVAL_415};
  assign _EVAL_358 = _EVAL_299 >> _EVAL_190;
  assign _EVAL_431 = _EVAL_358[0];
  assign _EVAL_90 = _EVAL_170[0];
  assign _EVAL_389 = {_EVAL_373,_EVAL_451};
  assign _EVAL_340 = _EVAL_299 >> _EVAL_389;
  assign _EVAL_203 = _EVAL_340[0];
  assign _EVAL_122 = _EVAL_46[5];
  assign _EVAL_347 = _EVAL_312[5];
  assign _EVAL_361 = {_EVAL_122,_EVAL_347};
  assign _EVAL_232 = _EVAL_299 >> _EVAL_361;
  assign _EVAL_335 = _EVAL_232[0];
  assign _EVAL_78 = _EVAL_312[4];
  assign _EVAL_207 = {_EVAL_276,_EVAL_78};
  assign _EVAL_234 = _EVAL_299 >> _EVAL_207;
  assign _EVAL_59 = _EVAL_234[0];
  assign _EVAL_442 = _EVAL_46[3];
  assign _EVAL_288 = _EVAL_312[3];
  assign _EVAL_390 = {_EVAL_442,_EVAL_288};
  assign _EVAL_427 = _EVAL_299 >> _EVAL_390;
  assign _EVAL_146 = _EVAL_427[0];
  assign _EVAL_332 = _EVAL_46[1];
  assign _EVAL_133 = _EVAL_312[1];
  assign _EVAL_398 = {_EVAL_332,_EVAL_133};
  assign _EVAL_413 = _EVAL_299 >> _EVAL_398;
  assign _EVAL_150 = _EVAL_413[0];
  assign _EVAL_344 = _EVAL_46[0];
  assign _EVAL_353 = _EVAL_312[0];
  assign _EVAL_241 = {_EVAL_344,_EVAL_353};
  assign _EVAL_306 = _EVAL_299 >> _EVAL_241;
  assign _EVAL_462 = _EVAL_306[0];
  assign _EVAL_243 = {_EVAL_203,_EVAL_48,_EVAL_335,_EVAL_59,_EVAL_146,_EVAL_94,_EVAL_150,_EVAL_462};
  assign _EVAL_437 = {_EVAL_342,_EVAL_423,_EVAL_456,_EVAL_115,_EVAL_148,_EVAL_431,_EVAL_180,_EVAL_90,_EVAL_243};
  assign _EVAL_108 = {_EVAL_400,_EVAL_362,_EVAL_443,_EVAL_65,_EVAL_102,_EVAL_383,_EVAL_286,_EVAL_167,_EVAL_84,_EVAL_437};
  assign _EVAL_209 = _EVAL_248 ? _EVAL_46 : _EVAL_312;
  assign _EVAL_315 = _EVAL_239 ? _EVAL_395 : _EVAL_209;
  assign _EVAL_143 = _EVAL_333 ? _EVAL_108 : _EVAL_315;
  assign _EVAL_378 = ~ _EVAL_371;
  assign _EVAL_211 = _EVAL_378[7:2];
  assign _EVAL_204 = _EVAL_54 - 6'h1;
  assign _EVAL_321 = _EVAL_118 & _EVAL_329;
  assign _EVAL_424 = 2'h1 << _EVAL_258;
  assign _EVAL_96 = _EVAL_424 | 2'h1;
  assign _EVAL_222 = _EVAL_96[1];
  assign _EVAL_291 = _EVAL_23 | _EVAL_321;
  assign _EVAL_184 = _EVAL_291 & _EVAL_17;
  assign _EVAL_345 = _EVAL_12[0];
  assign _EVAL_210 = 3'h1 == _EVAL_114;
  assign _EVAL_244 = 3'h0 == _EVAL_114;
  assign _EVAL_186 = _EVAL_130[1];
  assign _EVAL_149 = _EVAL_186 == 1'h0;
  assign _EVAL_380 = _EVAL_130[0];
  assign _EVAL_385 = _EVAL_149 & _EVAL_380;
  assign _EVAL_366 = _EVAL_402 >= 4'h2;
  assign _EVAL_268 = _EVAL_222 & _EVAL_186;
  assign _EVAL_370 = _EVAL_366 | _EVAL_268;
  assign _EVAL_43 = _EVAL_96[0];
  assign _EVAL_116 = _EVAL_186 & _EVAL_380;
  assign _EVAL_42 = _EVAL_43 & _EVAL_116;
  assign _EVAL_107 = _EVAL_370 | _EVAL_42;
  assign _EVAL_270 = _EVAL_416 ? _EVAL_409 : _EVAL_327;
  assign _EVAL_295 = _EVAL_12 == 3'h0;
  assign _EVAL_330 = _EVAL_280 & _EVAL_295;
  assign _EVAL_351 = _EVAL_321 == 1'h0;
  assign _EVAL_112 = _EVAL_126 ? 3'h4 : _EVAL_40;
  assign _EVAL_117 = {_EVAL_112,_EVAL_281,_EVAL_13,_EVAL_21,_EVAL_27,_EVAL_29,_EVAL_39,_EVAL_32};
  assign _EVAL_336 = _EVAL_380 == 1'h0;
  assign _EVAL_369 = _EVAL_222 & _EVAL_149;
  assign _EVAL_278 = _EVAL_366 | _EVAL_369;
  assign _EVAL_411 = _EVAL_43 & _EVAL_385;
  assign _EVAL_253 = _EVAL_278 | _EVAL_411;
  assign _EVAL_301 = _EVAL_330 & _EVAL_329;
  assign _EVAL_392 = _EVAL_186 & _EVAL_336;
  assign _EVAL_459 = _EVAL_43 & _EVAL_392;
  assign _EVAL_141 = _EVAL_370 | _EVAL_459;
  assign _EVAL_294 = _EVAL_149 & _EVAL_336;
  assign _EVAL_93 = _EVAL_43 & _EVAL_294;
  assign _EVAL_199 = _EVAL_278 | _EVAL_93;
  assign _EVAL_289 = _EVAL_262 | _EVAL_128;
  assign _EVAL_328 = {6'h0,_EVAL_402,_EVAL_176,_EVAL_130,_EVAL_107,_EVAL_141,_EVAL_253,_EVAL_199,_EVAL_143,_EVAL_289};
  assign _EVAL_309 = _EVAL_270 ? _EVAL_328 : 84'h0;
  assign _EVAL_412 = _EVAL_416 ? _EVAL_231 : _EVAL_368;
  assign _EVAL_132 = _EVAL_412 ? _EVAL_117 : 84'h0;
  assign _EVAL_381 = _EVAL_309 | _EVAL_132;
  assign _EVAL_237 = _EVAL_128 | _EVAL_20;
  assign _EVAL_139 = _EVAL_184 & _EVAL_280;
  assign _EVAL_206 = _EVAL_273 | _EVAL_20;
  assign _EVAL = _EVAL_416 ? _EVAL_363 : _EVAL_320;
  assign _EVAL_28 = _EVAL_381[32:1];
  assign _EVAL_34 = _EVAL_453 & _EVAL_375;
  assign _EVAL_22 = _EVAL_6;
  assign _EVAL_18 = _EVAL_381[83:81];
  assign _EVAL_19 = _EVAL_301 ? _EVAL_312 : _EVAL_0;
  assign _EVAL_25 = _EVAL_381[36:33];
  assign _EVAL_31 = _EVAL_301 ? _EVAL_206 : _EVAL_20;
  assign _EVAL_4 = _EVAL_381[0];
  assign _EVAL_24 = _EVAL_17 & _EVAL_351;
  assign _EVAL_11 = _EVAL_381[66:37];
  assign _EVAL_10 = _EVAL_23 | _EVAL_321;
  assign _EVAL_15 = _EVAL_381[77:74];
  assign _EVAL_35 = _EVAL_37;
  assign _EVAL_9 = _EVAL_301 ? _EVAL_237 : _EVAL_7;
  assign _EVAL_33 = _EVAL_381[73:67];
  assign _EVAL_16 = _EVAL_301 ? 3'h1 : _EVAL_12;
  assign _EVAL_36 = _EVAL_381[80:78];
  assign _EVAL_30 = _EVAL_38;
  assign _EVAL_5 = _EVAL_3;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_41 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_46 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_53 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_54 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_88 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_128 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_130 = _RAND_6[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_176 = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_262 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_273 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_298 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_299 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_312 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_327 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_368 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_394 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_402 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_8) begin
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_41 <= _EVAL_14;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_46 <= _EVAL_39;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_53 <= _EVAL_40;
      end
    end
    if (_EVAL_1) begin
      _EVAL_54 <= 6'h0;
    end else begin
      if (_EVAL_184) begin
        if (_EVAL_280) begin
          if (_EVAL_345) begin
            _EVAL_54 <= _EVAL_211;
          end else begin
            _EVAL_54 <= 6'h0;
          end
        end else begin
          _EVAL_54 <= _EVAL_204;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_88 <= 2'h0;
    end else begin
      if (_EVAL_139) begin
        if (_EVAL_329) begin
          if (_EVAL_264) begin
            _EVAL_88 <= 2'h2;
          end else begin
            _EVAL_88 <= 2'h0;
          end
        end else begin
          if (_EVAL_279) begin
            if (_EVAL_444) begin
              _EVAL_88 <= 2'h1;
            end else begin
              if (_EVAL_377) begin
                if (_EVAL_177) begin
                  _EVAL_88 <= 2'h3;
                end
              end
            end
          end else begin
            if (_EVAL_377) begin
              if (_EVAL_177) begin
                _EVAL_88 <= 2'h3;
              end
            end
          end
        end
      end else begin
        if (_EVAL_279) begin
          if (_EVAL_444) begin
            _EVAL_88 <= 2'h1;
          end else begin
            if (_EVAL_377) begin
              if (_EVAL_177) begin
                _EVAL_88 <= 2'h3;
              end
            end
          end
        end else begin
          if (_EVAL_377) begin
            if (_EVAL_177) begin
              _EVAL_88 <= 2'h3;
            end
          end
        end
      end
    end
    if (_EVAL_139) begin
      if (_EVAL_386) begin
        _EVAL_128 <= _EVAL_7;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_130 <= _EVAL_27;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_176 <= _EVAL_21;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_262 <= _EVAL_32;
      end
    end
    if (_EVAL_139) begin
      if (_EVAL_386) begin
        _EVAL_273 <= _EVAL_20;
      end
    end
    if (_EVAL_1) begin
      _EVAL_298 <= 6'h0;
    end else begin
      if (_EVAL_92) begin
        if (_EVAL_231) begin
          if (_EVAL_334) begin
            _EVAL_298 <= _EVAL_74;
          end else begin
            _EVAL_298 <= 6'h0;
          end
        end else begin
          _EVAL_298 <= 6'h0;
        end
      end else begin
        _EVAL_298 <= _EVAL_455;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        if (_EVAL_265) begin
          _EVAL_299 <= 4'h8;
        end else begin
          if (_EVAL_210) begin
            _EVAL_299 <= 4'he;
          end else begin
            if (_EVAL_244) begin
              _EVAL_299 <= 4'h6;
            end else begin
              if (_EVAL_131) begin
                _EVAL_299 <= 4'hc;
              end else begin
                _EVAL_299 <= 4'h0;
              end
            end
          end
        end
      end
    end
    if (_EVAL_139) begin
      if (_EVAL_386) begin
        _EVAL_312 <= _EVAL_0;
      end
    end
    if (_EVAL_1) begin
      _EVAL_327 <= 1'h0;
    end else begin
      if (_EVAL_416) begin
        _EVAL_327 <= _EVAL_409;
      end
    end
    if (_EVAL_1) begin
      _EVAL_368 <= 1'h0;
    end else begin
      if (_EVAL_416) begin
        _EVAL_368 <= _EVAL_231;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_394 <= _EVAL_29;
      end
    end
    if (_EVAL_377) begin
      if (_EVAL_177) begin
        _EVAL_402 <= _EVAL_13;
      end
    end
  end
endmodule
