//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_138_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [6:0]  _EVAL_8,
  input  [6:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [11:0] _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_16;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_40;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_58;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_69;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_82;
  reg [31:0] _RAND_4;
  reg [72:0] _EVAL_110;
  reg [95:0] _RAND_5;
  reg [3:0] _EVAL_130;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_166;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_170;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_190;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_199;
  reg [31:0] _RAND_10;
  reg [11:0] _EVAL_212;
  reg [31:0] _RAND_11;
  reg [6:0] _EVAL_217;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_253;
  reg [31:0] _RAND_13;
  wire  _EVAL_80;
  wire  _EVAL_275;
  wire  _EVAL_185;
  wire [127:0] _EVAL_123;
  wire [127:0] _EVAL_270;
  wire [72:0] _EVAL_148;
  wire [72:0] _EVAL_36;
  wire  _EVAL_86;
  wire  _EVAL_153;
  wire [12:0] _EVAL_226;
  wire [12:0] _EVAL_124;
  wire [12:0] _EVAL_18;
  wire  _EVAL_76;
  wire [1:0] _EVAL_223;
  wire [1:0] _EVAL_102;
  wire  _EVAL_98;
  wire  _EVAL_232;
  wire  _EVAL_158;
  wire  _EVAL_260;
  wire  _EVAL_122;
  wire  _EVAL_222;
  wire  _EVAL_244;
  wire  _EVAL_35;
  wire  _EVAL_181;
  wire [12:0] _EVAL_257;
  wire [5:0] _EVAL_281;
  wire [5:0] _EVAL_156;
  wire [3:0] _EVAL_31;
  wire [3:0] _EVAL_163;
  wire  _EVAL_135;
  wire [72:0] _EVAL_96;
  wire  _EVAL_127;
  wire [3:0] _EVAL_20;
  wire  _EVAL_107;
  wire  _EVAL_220;
  wire  _EVAL_140;
  wire  _EVAL_178;
  wire  _EVAL_26;
  wire  _EVAL_41;
  wire  _EVAL_173;
  wire  _EVAL_189;
  wire  _EVAL_90;
  wire [127:0] _EVAL_228;
  wire [127:0] _EVAL_192;
  wire [72:0] _EVAL_33;
  wire [72:0] _EVAL_131;
  wire [72:0] _EVAL_245;
  wire  _EVAL_57;
  wire  _EVAL_63;
  wire  _EVAL_93;
  wire [12:0] _EVAL_105;
  wire [5:0] _EVAL_74;
  wire [5:0] _EVAL_143;
  wire [3:0] _EVAL_94;
  wire  _EVAL_225;
  wire  _EVAL_115;
  wire  _EVAL_265;
  wire  _EVAL_277;
  wire  _EVAL_171;
  wire  _EVAL_29;
  wire [3:0] _EVAL_121;
  wire  _EVAL_43;
  wire  _EVAL_237;
  wire  _EVAL_262;
  wire  _EVAL_120;
  wire [2:0] _EVAL_219;
  wire  _EVAL_70;
  wire  _EVAL_133;
  wire  _EVAL_271;
  wire  _EVAL_188;
  wire  _EVAL_206;
  wire  _EVAL_37;
  wire [11:0] _EVAL_224;
  wire  _EVAL_162;
  wire  _EVAL_81;
  wire  _EVAL_75;
  wire  _EVAL_118;
  wire  _EVAL_150;
  wire  _EVAL_112;
  wire  _EVAL_195;
  wire  _EVAL_243;
  wire  _EVAL_83;
  wire [3:0] _EVAL_230;
  wire  _EVAL_272;
  wire  _EVAL_183;
  wire  _EVAL_106;
  wire  _EVAL_154;
  wire  _EVAL_269;
  wire  _EVAL_136;
  wire  _EVAL_149;
  wire  _EVAL_78;
  wire  _EVAL_177;
  wire  _EVAL_210;
  wire [3:0] _EVAL_128;
  wire  _EVAL_160;
  wire  _EVAL_276;
  wire  _EVAL_55;
  wire  _EVAL_200;
  wire  _EVAL_137;
  wire [72:0] _EVAL_205;
  wire [72:0] _EVAL_215;
  wire  _EVAL_236;
  wire [2:0] _EVAL_203;
  wire  _EVAL_97;
  wire  _EVAL_155;
  wire  _EVAL_175;
  wire  _EVAL_103;
  wire  _EVAL_64;
  wire  _EVAL_66;
  wire  _EVAL_22;
  wire [3:0] _EVAL_184;
  wire  _EVAL_25;
  wire  _EVAL_45;
  wire  _EVAL_208;
  wire  _EVAL_179;
  wire  _EVAL_68;
  wire  _EVAL_258;
  wire  _EVAL_176;
  wire  _EVAL_207;
  wire  _EVAL_111;
  wire  _EVAL_15;
  wire  _EVAL_62;
  wire  _EVAL_172;
  wire  _EVAL_39;
  wire [3:0] _EVAL_246;
  wire [3:0] _EVAL_72;
  wire [3:0] _EVAL_233;
  wire  _EVAL_255;
  wire  _EVAL_221;
  wire  _EVAL_202;
  wire  _EVAL_250;
  wire  _EVAL_235;
  wire  _EVAL_201;
  wire  _EVAL_231;
  wire  _EVAL_251;
  wire  _EVAL_32;
  wire  _EVAL_95;
  wire  _EVAL_254;
  wire  _EVAL_248;
  wire  _EVAL_216;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_100;
  wire  _EVAL_213;
  wire  _EVAL_99;
  wire  _EVAL_168;
  wire  _EVAL_193;
  wire  _EVAL_108;
  wire  _EVAL_234;
  wire  _EVAL_141;
  wire  _EVAL_187;
  wire [31:0] _EVAL_264;
  wire  _EVAL_214;
  wire  _EVAL_266;
  wire  _EVAL_89;
  wire  _EVAL_92;
  wire  _EVAL_267;
  wire  _EVAL_278;
  wire  _EVAL_60;
  wire  _EVAL_268;
  wire  _EVAL_165;
  wire  _EVAL_52;
  wire  _EVAL_71;
  wire  _EVAL_67;
  wire  _EVAL_238;
  wire  _EVAL_144;
  wire  _EVAL_61;
  wire  _EVAL_42;
  wire  _EVAL_125;
  wire  _EVAL_116;
  wire  _EVAL_145;
  wire  _EVAL_138;
  wire  _EVAL_24;
  wire [3:0] _EVAL_54;
  wire [11:0] _EVAL_139;
  wire  _EVAL_252;
  wire  _EVAL_240;
  wire  _EVAL_279;
  wire  _EVAL_247;
  wire  _EVAL_142;
  wire  _EVAL_53;
  wire  _EVAL_84;
  wire  _EVAL_164;
  wire  _EVAL_132;
  wire  _EVAL_157;
  wire  _EVAL_134;
  wire  _EVAL_241;
  wire  _EVAL_227;
  wire  _EVAL_28;
  wire  _EVAL_147;
  wire  _EVAL_49;
  wire  _EVAL_114;
  wire  _EVAL_151;
  wire  _EVAL_249;
  wire  _EVAL_119;
  wire  _EVAL_196;
  wire  _EVAL_101;
  wire  _EVAL_129;
  wire  _EVAL_242;
  wire  _EVAL_263;
  wire  _EVAL_50;
  wire  _EVAL_79;
  wire  _EVAL_146;
  wire  _EVAL_229;
  wire  _EVAL_44;
  wire  _EVAL_186;
  wire  _EVAL_46;
  wire  _EVAL_159;
  wire  _EVAL_73;
  wire  _EVAL_197;
  wire  _EVAL_259;
  wire  _EVAL_34;
  wire  _EVAL_169;
  wire  _EVAL_51;
  wire  _EVAL_19;
  wire  _EVAL_91;
  wire  _EVAL_109;
  wire  _EVAL_191;
  wire  _EVAL_180;
  wire  _EVAL_113;
  wire  _EVAL_21;
  wire  _EVAL_23;
  wire  _EVAL_182;
  wire  _EVAL_104;
  wire  _EVAL_261;
  wire  _EVAL_88;
  wire  _EVAL_77;
  wire  _EVAL_152;
  wire  _EVAL_167;
  wire  _EVAL_198;
  wire  _EVAL_256;
  wire  _EVAL_273;
  wire  _EVAL_280;
  wire  _EVAL_30;
  wire  _EVAL_126;
  wire  _EVAL_117;
  wire  _EVAL_194;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_80 = _EVAL & _EVAL_6;
  assign _EVAL_275 = _EVAL_130 == 4'h0;
  assign _EVAL_185 = _EVAL_80 & _EVAL_275;
  assign _EVAL_123 = 128'h1 << _EVAL_9;
  assign _EVAL_270 = _EVAL_185 ? _EVAL_123 : 128'h0;
  assign _EVAL_148 = _EVAL_270[72:0];
  assign _EVAL_36 = _EVAL_110 | _EVAL_148;
  assign _EVAL_86 = _EVAL_2 == _EVAL_170;
  assign _EVAL_153 = _EVAL_86 | _EVAL_13;
  assign _EVAL_226 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_124 = $signed(_EVAL_226) & $signed(-13'sh1000);
  assign _EVAL_18 = $signed(_EVAL_124);
  assign _EVAL_76 = _EVAL_2[0];
  assign _EVAL_223 = 2'h1 << _EVAL_76;
  assign _EVAL_102 = _EVAL_223 | 2'h1;
  assign _EVAL_98 = _EVAL_102[0];
  assign _EVAL_232 = _EVAL_12[1];
  assign _EVAL_158 = _EVAL_232 == 1'h0;
  assign _EVAL_260 = _EVAL_12[0];
  assign _EVAL_122 = _EVAL_260 == 1'h0;
  assign _EVAL_222 = _EVAL_158 & _EVAL_122;
  assign _EVAL_244 = _EVAL_98 & _EVAL_222;
  assign _EVAL_35 = _EVAL_5[2];
  assign _EVAL_181 = _EVAL_35 == 1'h0;
  assign _EVAL_257 = 13'h3f << _EVAL_2;
  assign _EVAL_281 = _EVAL_257[5:0];
  assign _EVAL_156 = ~ _EVAL_281;
  assign _EVAL_31 = _EVAL_156[5:2];
  assign _EVAL_163 = _EVAL_130 - 4'h1;
  assign _EVAL_135 = _EVAL_5 == 3'h3;
  assign _EVAL_96 = _EVAL_110 >> _EVAL_9;
  assign _EVAL_127 = _EVAL_96[0];
  assign _EVAL_20 = _EVAL_8[6:3];
  assign _EVAL_107 = _EVAL_20 == 4'h2;
  assign _EVAL_220 = _EVAL_2 >= 3'h2;
  assign _EVAL_140 = _EVAL_220 | _EVAL_13;
  assign _EVAL_178 = _EVAL_4 & _EVAL_3;
  assign _EVAL_26 = _EVAL_58 == 4'h0;
  assign _EVAL_41 = _EVAL_178 & _EVAL_26;
  assign _EVAL_173 = _EVAL_0 == 3'h6;
  assign _EVAL_189 = _EVAL_173 == 1'h0;
  assign _EVAL_90 = _EVAL_41 & _EVAL_189;
  assign _EVAL_228 = 128'h1 << _EVAL_8;
  assign _EVAL_192 = _EVAL_90 ? _EVAL_228 : 128'h0;
  assign _EVAL_33 = _EVAL_192[72:0];
  assign _EVAL_131 = ~ _EVAL_33;
  assign _EVAL_245 = _EVAL_36 & _EVAL_131;
  assign _EVAL_57 = $signed(_EVAL_18) == $signed(13'sh0);
  assign _EVAL_63 = _EVAL_1 >= 3'h2;
  assign _EVAL_93 = _EVAL_0[0];
  assign _EVAL_105 = 13'h3f << _EVAL_1;
  assign _EVAL_74 = _EVAL_105[5:0];
  assign _EVAL_143 = ~ _EVAL_74;
  assign _EVAL_94 = _EVAL_143[5:2];
  assign _EVAL_225 = _EVAL_0 == 3'h0;
  assign _EVAL_115 = _EVAL_9 == 7'h40;
  assign _EVAL_265 = 3'h6 == _EVAL_2;
  assign _EVAL_277 = _EVAL_115 ? _EVAL_265 : 1'h0;
  assign _EVAL_171 = _EVAL_277 | _EVAL_13;
  assign _EVAL_29 = _EVAL_69 == 4'h0;
  assign _EVAL_121 = _EVAL_69 - 4'h1;
  assign _EVAL_43 = _EVAL_5 == 3'h2;
  assign _EVAL_237 = _EVAL_6 & _EVAL_43;
  assign _EVAL_262 = _EVAL_232 & _EVAL_260;
  assign _EVAL_120 = _EVAL_98 & _EVAL_262;
  assign _EVAL_219 = _EVAL_8[2:0];
  assign _EVAL_70 = 3'h1 <= _EVAL_219;
  assign _EVAL_133 = _EVAL_9 == _EVAL_217;
  assign _EVAL_271 = _EVAL_133 | _EVAL_13;
  assign _EVAL_188 = _EVAL_127 == 1'h0;
  assign _EVAL_206 = _EVAL_188 | _EVAL_13;
  assign _EVAL_37 = _EVAL_206 == 1'h0;
  assign _EVAL_224 = {{6'd0}, _EVAL_156};
  assign _EVAL_162 = plusarg_reader_out == 32'h0;
  assign _EVAL_81 = _EVAL_190 == 4'h0;
  assign _EVAL_75 = _EVAL_81 == 1'h0;
  assign _EVAL_118 = _EVAL_102[1];
  assign _EVAL_150 = _EVAL_118 & _EVAL_158;
  assign _EVAL_112 = _EVAL_220 | _EVAL_150;
  assign _EVAL_195 = _EVAL_158 & _EVAL_260;
  assign _EVAL_243 = _EVAL_98 & _EVAL_195;
  assign _EVAL_83 = _EVAL_112 | _EVAL_243;
  assign _EVAL_230 = _EVAL_58 - 4'h1;
  assign _EVAL_272 = _EVAL_0 == 3'h1;
  assign _EVAL_183 = _EVAL_3 & _EVAL_272;
  assign _EVAL_106 = _EVAL_11 == 1'h0;
  assign _EVAL_154 = _EVAL_8 == 7'h48;
  assign _EVAL_269 = _EVAL_110 != 73'h0;
  assign _EVAL_136 = _EVAL_269 == 1'h0;
  assign _EVAL_149 = _EVAL_136 | _EVAL_162;
  assign _EVAL_78 = _EVAL_0 == 3'h5;
  assign _EVAL_177 = _EVAL_8 == 7'h40;
  assign _EVAL_210 = _EVAL_20 == 4'h3;
  assign _EVAL_128 = _EVAL_9[6:3];
  assign _EVAL_160 = _EVAL_29 == 1'h0;
  assign _EVAL_276 = _EVAL_6 & _EVAL_160;
  assign _EVAL_55 = _EVAL_118 & _EVAL_232;
  assign _EVAL_200 = _EVAL_220 | _EVAL_55;
  assign _EVAL_137 = _EVAL_200 | _EVAL_120;
  assign _EVAL_205 = _EVAL_148 | _EVAL_110;
  assign _EVAL_215 = _EVAL_205 >> _EVAL_8;
  assign _EVAL_236 = _EVAL_215[0];
  assign _EVAL_203 = _EVAL_9[2:0];
  assign _EVAL_97 = _EVAL_0 <= 3'h6;
  assign _EVAL_155 = _EVAL_97 | _EVAL_13;
  assign _EVAL_175 = _EVAL_5 == 3'h5;
  assign _EVAL_103 = _EVAL_8 == _EVAL_40;
  assign _EVAL_64 = _EVAL_6 & _EVAL_135;
  assign _EVAL_66 = _EVAL_106 | _EVAL_13;
  assign _EVAL_22 = _EVAL_66 == 1'h0;
  assign _EVAL_184 = ~ _EVAL_7;
  assign _EVAL_25 = _EVAL_14 <= 3'h4;
  assign _EVAL_45 = _EVAL_25 | _EVAL_13;
  assign _EVAL_208 = _EVAL_5 == 3'h7;
  assign _EVAL_179 = _EVAL_6 & _EVAL_208;
  assign _EVAL_68 = _EVAL_140 == 1'h0;
  assign _EVAL_258 = _EVAL_14 <= 3'h2;
  assign _EVAL_176 = _EVAL_14 <= 3'h3;
  assign _EVAL_207 = _EVAL_176 | _EVAL_13;
  assign _EVAL_111 = _EVAL_207 == 1'h0;
  assign _EVAL_15 = _EVAL_232 & _EVAL_122;
  assign _EVAL_62 = _EVAL_98 & _EVAL_15;
  assign _EVAL_172 = _EVAL_200 | _EVAL_62;
  assign _EVAL_39 = _EVAL_112 | _EVAL_244;
  assign _EVAL_246 = {_EVAL_137,_EVAL_172,_EVAL_83,_EVAL_39};
  assign _EVAL_72 = ~ _EVAL_246;
  assign _EVAL_233 = _EVAL_7 & _EVAL_72;
  assign _EVAL_255 = _EVAL_233 == 4'h0;
  assign _EVAL_221 = _EVAL_255 | _EVAL_13;
  assign _EVAL_202 = _EVAL_1 == _EVAL_82;
  assign _EVAL_250 = _EVAL_202 | _EVAL_13;
  assign _EVAL_235 = _EVAL_5 == 3'h6;
  assign _EVAL_201 = _EVAL_6 & _EVAL_235;
  assign _EVAL_231 = _EVAL_80 & _EVAL_29;
  assign _EVAL_251 = _EVAL_154 | _EVAL_177;
  assign _EVAL_32 = _EVAL_20 == 4'h8;
  assign _EVAL_95 = _EVAL_32 & _EVAL_70;
  assign _EVAL_254 = _EVAL_251 | _EVAL_95;
  assign _EVAL_248 = _EVAL_8 == 7'h20;
  assign _EVAL_216 = _EVAL_254 | _EVAL_248;
  assign _EVAL_47 = _EVAL_20 == 4'h0;
  assign _EVAL_48 = _EVAL_216 | _EVAL_47;
  assign _EVAL_100 = _EVAL_20 == 4'h1;
  assign _EVAL_213 = _EVAL_48 | _EVAL_100;
  assign _EVAL_99 = _EVAL_213 | _EVAL_107;
  assign _EVAL_168 = _EVAL_99 | _EVAL_210;
  assign _EVAL_193 = _EVAL_168 | _EVAL_13;
  assign _EVAL_108 = _EVAL_63 | _EVAL_13;
  assign _EVAL_234 = _EVAL_45 == 1'h0;
  assign _EVAL_141 = _EVAL_155 == 1'h0;
  assign _EVAL_187 = _EVAL_80 | _EVAL_178;
  assign _EVAL_264 = _EVAL_166 + 32'h1;
  assign _EVAL_214 = _EVAL_9 == 7'h48;
  assign _EVAL_266 = _EVAL_214 | _EVAL_115;
  assign _EVAL_89 = _EVAL_128 == 4'h8;
  assign _EVAL_92 = 3'h1 <= _EVAL_203;
  assign _EVAL_267 = _EVAL_89 & _EVAL_92;
  assign _EVAL_278 = _EVAL_266 | _EVAL_267;
  assign _EVAL_60 = _EVAL_9 == 7'h20;
  assign _EVAL_268 = _EVAL_278 | _EVAL_60;
  assign _EVAL_165 = _EVAL_128 == 4'h0;
  assign _EVAL_52 = _EVAL_268 | _EVAL_165;
  assign _EVAL_71 = _EVAL_128 == 4'h1;
  assign _EVAL_67 = _EVAL_52 | _EVAL_71;
  assign _EVAL_238 = _EVAL_128 == 4'h2;
  assign _EVAL_144 = _EVAL_67 | _EVAL_238;
  assign _EVAL_61 = _EVAL_171 == 1'h0;
  assign _EVAL_42 = _EVAL_166 < plusarg_reader_out;
  assign _EVAL_125 = _EVAL_6 & _EVAL_175;
  assign _EVAL_116 = _EVAL_12 == _EVAL_212;
  assign _EVAL_145 = _EVAL_116 | _EVAL_13;
  assign _EVAL_138 = _EVAL_145 == 1'h0;
  assign _EVAL_24 = _EVAL_128 == 4'h3;
  assign _EVAL_54 = _EVAL_190 - 4'h1;
  assign _EVAL_139 = _EVAL_12 & _EVAL_224;
  assign _EVAL_252 = _EVAL_139 == 12'h0;
  assign _EVAL_240 = _EVAL_252 | _EVAL_13;
  assign _EVAL_279 = _EVAL_240 == 1'h0;
  assign _EVAL_247 = _EVAL_13 == 1'h0;
  assign _EVAL_142 = _EVAL_149 | _EVAL_42;
  assign _EVAL_53 = _EVAL_142 | _EVAL_13;
  assign _EVAL_84 = _EVAL_184 == 4'h0;
  assign _EVAL_164 = _EVAL_236 | _EVAL_13;
  assign _EVAL_132 = _EVAL_258 | _EVAL_13;
  assign _EVAL_157 = _EVAL_132 == 1'h0;
  assign _EVAL_134 = _EVAL_14 == _EVAL_199;
  assign _EVAL_241 = _EVAL_134 | _EVAL_13;
  assign _EVAL_227 = _EVAL_241 == 1'h0;
  assign _EVAL_28 = _EVAL_5 == 3'h0;
  assign _EVAL_147 = _EVAL_6 & _EVAL_28;
  assign _EVAL_49 = _EVAL_5 == _EVAL_253;
  assign _EVAL_114 = _EVAL_49 | _EVAL_13;
  assign _EVAL_151 = _EVAL_103 | _EVAL_13;
  assign _EVAL_249 = _EVAL_151 == 1'h0;
  assign _EVAL_119 = _EVAL_0 == 3'h4;
  assign _EVAL_196 = _EVAL_3 & _EVAL_119;
  assign _EVAL_101 = _EVAL_144 | _EVAL_24;
  assign _EVAL_129 = _EVAL_101 | _EVAL_13;
  assign _EVAL_242 = _EVAL_2 <= 3'h6;
  assign _EVAL_263 = _EVAL_242 & _EVAL_57;
  assign _EVAL_50 = _EVAL_3 & _EVAL_75;
  assign _EVAL_79 = _EVAL_14 != 3'h0;
  assign _EVAL_146 = _EVAL_79 | _EVAL_13;
  assign _EVAL_229 = _EVAL_7 == _EVAL_246;
  assign _EVAL_44 = _EVAL_229 | _EVAL_13;
  assign _EVAL_186 = _EVAL_44 == 1'h0;
  assign _EVAL_46 = _EVAL_114 == 1'h0;
  assign _EVAL_159 = _EVAL_221 == 1'h0;
  assign _EVAL_73 = _EVAL_5 == 3'h1;
  assign _EVAL_197 = _EVAL_263 | _EVAL_13;
  assign _EVAL_259 = _EVAL_271 == 1'h0;
  assign _EVAL_34 = _EVAL_250 == 1'h0;
  assign _EVAL_169 = _EVAL_0 == _EVAL_16;
  assign _EVAL_51 = _EVAL_0 == 3'h2;
  assign _EVAL_19 = _EVAL_3 & _EVAL_51;
  assign _EVAL_91 = _EVAL_169 | _EVAL_13;
  assign _EVAL_109 = _EVAL_14 == 3'h0;
  assign _EVAL_191 = _EVAL_109 | _EVAL_13;
  assign _EVAL_180 = _EVAL_191 == 1'h0;
  assign _EVAL_113 = _EVAL_164 == 1'h0;
  assign _EVAL_21 = _EVAL_129 == 1'h0;
  assign _EVAL_23 = _EVAL_178 & _EVAL_81;
  assign _EVAL_182 = _EVAL_3 & _EVAL_78;
  assign _EVAL_104 = _EVAL_5 == 3'h4;
  assign _EVAL_261 = _EVAL_6 & _EVAL_104;
  assign _EVAL_88 = _EVAL_53 == 1'h0;
  assign _EVAL_77 = _EVAL_153 == 1'h0;
  assign _EVAL_152 = _EVAL_84 | _EVAL_13;
  assign _EVAL_167 = _EVAL_152 == 1'h0;
  assign _EVAL_198 = _EVAL_146 == 1'h0;
  assign _EVAL_256 = _EVAL_193 == 1'h0;
  assign _EVAL_273 = _EVAL_3 & _EVAL_173;
  assign _EVAL_280 = _EVAL_108 == 1'h0;
  assign _EVAL_30 = _EVAL_3 & _EVAL_225;
  assign _EVAL_126 = _EVAL_197 == 1'h0;
  assign _EVAL_117 = _EVAL_91 == 1'h0;
  assign _EVAL_194 = _EVAL_6 & _EVAL_73;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_16 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_40 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_58 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_69 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_82 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  _EVAL_110 = _RAND_5[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_130 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_166 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_170 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_190 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_199 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_212 = _RAND_11[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_217 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_253 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_10) begin
    if (_EVAL_23) begin
      _EVAL_16 <= _EVAL_0;
    end
    if (_EVAL_23) begin
      _EVAL_40 <= _EVAL_8;
    end
    if (_EVAL_13) begin
      _EVAL_58 <= 4'h0;
    end else begin
      if (_EVAL_178) begin
        if (_EVAL_26) begin
          if (_EVAL_93) begin
            _EVAL_58 <= _EVAL_94;
          end else begin
            _EVAL_58 <= 4'h0;
          end
        end else begin
          _EVAL_58 <= _EVAL_230;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_69 <= 4'h0;
    end else begin
      if (_EVAL_80) begin
        if (_EVAL_29) begin
          if (_EVAL_181) begin
            _EVAL_69 <= _EVAL_31;
          end else begin
            _EVAL_69 <= 4'h0;
          end
        end else begin
          _EVAL_69 <= _EVAL_121;
        end
      end
    end
    if (_EVAL_23) begin
      _EVAL_82 <= _EVAL_1;
    end
    if (_EVAL_13) begin
      _EVAL_110 <= 73'h0;
    end else begin
      _EVAL_110 <= _EVAL_245;
    end
    if (_EVAL_13) begin
      _EVAL_130 <= 4'h0;
    end else begin
      if (_EVAL_80) begin
        if (_EVAL_275) begin
          if (_EVAL_181) begin
            _EVAL_130 <= _EVAL_31;
          end else begin
            _EVAL_130 <= 4'h0;
          end
        end else begin
          _EVAL_130 <= _EVAL_163;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_166 <= 32'h0;
    end else begin
      if (_EVAL_187) begin
        _EVAL_166 <= 32'h0;
      end else begin
        _EVAL_166 <= _EVAL_264;
      end
    end
    if (_EVAL_231) begin
      _EVAL_170 <= _EVAL_2;
    end
    if (_EVAL_13) begin
      _EVAL_190 <= 4'h0;
    end else begin
      if (_EVAL_178) begin
        if (_EVAL_81) begin
          if (_EVAL_93) begin
            _EVAL_190 <= _EVAL_94;
          end else begin
            _EVAL_190 <= 4'h0;
          end
        end else begin
          _EVAL_190 <= _EVAL_54;
        end
      end
    end
    if (_EVAL_231) begin
      _EVAL_199 <= _EVAL_14;
    end
    if (_EVAL_231) begin
      _EVAL_212 <= _EVAL_12;
    end
    if (_EVAL_231) begin
      _EVAL_217 <= _EVAL_9;
    end
    if (_EVAL_231) begin
      _EVAL_253 <= _EVAL_5;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3bcee72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4f3d28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18a7364c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b7188d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29317591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67472586)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a85a3fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b44e85bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f49a9c4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b3587d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(894ebfd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e46fda66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b66c415d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daaaa63a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(488ed1b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2349f4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f85a74c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36f2212b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7544076d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55b521b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad31f79f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31df0777)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(151c3079)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(441a7ec4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3521201d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3899f7a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f33abd86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e246004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7579b359)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1074c9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f812a499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2321987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f771b3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5a79c24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a1c6a33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbcc9481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73c19bb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdef24fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da39d438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e320fcce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb3d189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0d1b1f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44b2d735)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a29ea69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e4664b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8a87908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff701874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f5031f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ce2edf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(244c9019)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d04bf07a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15a8da5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43c1baa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e08b29c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77e323e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b35391d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57862079)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47aeb1f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(433e5fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c102e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e29d0512)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(242d1183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b302ee8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94dc3a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac87238d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1bca6b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff1b8cc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd793072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baff2ca5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2d0c707)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2077470e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
