//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_292(
  input         _EVAL,
  input         _EVAL_0,
  input  [32:0] _EVAL_1,
  output        _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [32:0] _EVAL_5,
  input  [32:0] _EVAL_6,
  output [4:0]  _EVAL_7,
  output [32:0] _EVAL_8
);
  wire  mulAddRecFNToRaw_postMul__EVAL;
  wire [4:0] mulAddRecFNToRaw_postMul__EVAL_0;
  wire  mulAddRecFNToRaw_postMul__EVAL_1;
  wire  mulAddRecFNToRaw_postMul__EVAL_2;
  wire  mulAddRecFNToRaw_postMul__EVAL_3;
  wire  mulAddRecFNToRaw_postMul__EVAL_4;
  wire  mulAddRecFNToRaw_postMul__EVAL_5;
  wire  mulAddRecFNToRaw_postMul__EVAL_6;
  wire [9:0] mulAddRecFNToRaw_postMul__EVAL_7;
  wire  mulAddRecFNToRaw_postMul__EVAL_8;
  wire  mulAddRecFNToRaw_postMul__EVAL_9;
  wire [48:0] mulAddRecFNToRaw_postMul__EVAL_10;
  wire [9:0] mulAddRecFNToRaw_postMul__EVAL_11;
  wire  mulAddRecFNToRaw_postMul__EVAL_12;
  wire [25:0] mulAddRecFNToRaw_postMul__EVAL_13;
  wire  mulAddRecFNToRaw_postMul__EVAL_14;
  wire  mulAddRecFNToRaw_postMul__EVAL_15;
  wire [2:0] mulAddRecFNToRaw_postMul__EVAL_16;
  wire  mulAddRecFNToRaw_postMul__EVAL_17;
  wire [26:0] mulAddRecFNToRaw_postMul__EVAL_18;
  wire  mulAddRecFNToRaw_postMul__EVAL_19;
  wire  mulAddRecFNToRaw_postMul__EVAL_20;
  wire  mulAddRecFNToRaw_postMul__EVAL_21;
  wire  mulAddRecFNToRaw_postMul__EVAL_22;
  wire  mulAddRecFNToRaw_postMul__EVAL_23;
  wire [32:0] roundRawFNToRecFN__EVAL;
  wire [9:0] roundRawFNToRecFN__EVAL_0;
  wire  roundRawFNToRecFN__EVAL_1;
  wire [2:0] roundRawFNToRecFN__EVAL_2;
  wire  roundRawFNToRecFN__EVAL_3;
  wire [4:0] roundRawFNToRecFN__EVAL_4;
  wire  roundRawFNToRecFN__EVAL_5;
  wire [26:0] roundRawFNToRecFN__EVAL_6;
  wire  roundRawFNToRecFN__EVAL_7;
  wire  roundRawFNToRecFN__EVAL_8;
  wire  roundRawFNToRecFN__EVAL_9;
  wire [32:0] mulAddRecFNToRaw_preMul__EVAL;
  wire  mulAddRecFNToRaw_preMul__EVAL_0;
  wire [23:0] mulAddRecFNToRaw_preMul__EVAL_1;
  wire [25:0] mulAddRecFNToRaw_preMul__EVAL_2;
  wire  mulAddRecFNToRaw_preMul__EVAL_3;
  wire  mulAddRecFNToRaw_preMul__EVAL_4;
  wire  mulAddRecFNToRaw_preMul__EVAL_5;
  wire [32:0] mulAddRecFNToRaw_preMul__EVAL_6;
  wire  mulAddRecFNToRaw_preMul__EVAL_7;
  wire [4:0] mulAddRecFNToRaw_preMul__EVAL_8;
  wire  mulAddRecFNToRaw_preMul__EVAL_9;
  wire [23:0] mulAddRecFNToRaw_preMul__EVAL_10;
  wire  mulAddRecFNToRaw_preMul__EVAL_11;
  wire  mulAddRecFNToRaw_preMul__EVAL_12;
  wire [47:0] mulAddRecFNToRaw_preMul__EVAL_13;
  wire  mulAddRecFNToRaw_preMul__EVAL_14;
  wire  mulAddRecFNToRaw_preMul__EVAL_15;
  wire  mulAddRecFNToRaw_preMul__EVAL_16;
  wire [32:0] mulAddRecFNToRaw_preMul__EVAL_17;
  wire  mulAddRecFNToRaw_preMul__EVAL_18;
  wire  mulAddRecFNToRaw_preMul__EVAL_19;
  wire [9:0] mulAddRecFNToRaw_preMul__EVAL_20;
  reg  _EVAL_9;
  reg [31:0] _RAND_0;
  reg  _EVAL_10;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_11;
  reg [31:0] _RAND_2;
  reg  _EVAL_13;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_14;
  reg [31:0] _RAND_4;
  reg [26:0] _EVAL_15;
  reg [31:0] _RAND_5;
  reg  _EVAL_16;
  reg [31:0] _RAND_6;
  reg  _EVAL_17;
  reg [31:0] _RAND_7;
  reg  _EVAL_19;
  reg [31:0] _RAND_8;
  reg [25:0] _EVAL_20;
  reg [31:0] _RAND_9;
  reg [9:0] _EVAL_21;
  reg [31:0] _RAND_10;
  reg  _EVAL_22;
  reg [31:0] _RAND_11;
  reg  _EVAL_23;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_24;
  reg [31:0] _RAND_13;
  reg  _EVAL_25;
  reg [31:0] _RAND_14;
  reg  _EVAL_26;
  reg [31:0] _RAND_15;
  reg  _EVAL_27;
  reg [31:0] _RAND_16;
  reg [2:0] _EVAL_28;
  reg [31:0] _RAND_17;
  reg  _EVAL_29;
  reg [31:0] _RAND_18;
  reg  _EVAL_30;
  reg [31:0] _RAND_19;
  reg  _EVAL_31;
  reg [31:0] _RAND_20;
  reg  _EVAL_32;
  reg [31:0] _RAND_21;
  reg  _EVAL_33;
  reg [31:0] _RAND_22;
  reg  _EVAL_34;
  reg [31:0] _RAND_23;
  reg  _EVAL_35;
  reg [31:0] _RAND_24;
  reg [48:0] _EVAL_36;
  reg [63:0] _RAND_25;
  reg  _EVAL_37;
  reg [31:0] _RAND_26;
  reg  _EVAL_38;
  reg [31:0] _RAND_27;
  reg [9:0] _EVAL_39;
  reg [31:0] _RAND_28;
  wire [47:0] _EVAL_18;
  wire [48:0] _EVAL_12;
  SiFive__EVAL_289 mulAddRecFNToRaw_postMul (
    ._EVAL(mulAddRecFNToRaw_postMul__EVAL),
    ._EVAL_0(mulAddRecFNToRaw_postMul__EVAL_0),
    ._EVAL_1(mulAddRecFNToRaw_postMul__EVAL_1),
    ._EVAL_2(mulAddRecFNToRaw_postMul__EVAL_2),
    ._EVAL_3(mulAddRecFNToRaw_postMul__EVAL_3),
    ._EVAL_4(mulAddRecFNToRaw_postMul__EVAL_4),
    ._EVAL_5(mulAddRecFNToRaw_postMul__EVAL_5),
    ._EVAL_6(mulAddRecFNToRaw_postMul__EVAL_6),
    ._EVAL_7(mulAddRecFNToRaw_postMul__EVAL_7),
    ._EVAL_8(mulAddRecFNToRaw_postMul__EVAL_8),
    ._EVAL_9(mulAddRecFNToRaw_postMul__EVAL_9),
    ._EVAL_10(mulAddRecFNToRaw_postMul__EVAL_10),
    ._EVAL_11(mulAddRecFNToRaw_postMul__EVAL_11),
    ._EVAL_12(mulAddRecFNToRaw_postMul__EVAL_12),
    ._EVAL_13(mulAddRecFNToRaw_postMul__EVAL_13),
    ._EVAL_14(mulAddRecFNToRaw_postMul__EVAL_14),
    ._EVAL_15(mulAddRecFNToRaw_postMul__EVAL_15),
    ._EVAL_16(mulAddRecFNToRaw_postMul__EVAL_16),
    ._EVAL_17(mulAddRecFNToRaw_postMul__EVAL_17),
    ._EVAL_18(mulAddRecFNToRaw_postMul__EVAL_18),
    ._EVAL_19(mulAddRecFNToRaw_postMul__EVAL_19),
    ._EVAL_20(mulAddRecFNToRaw_postMul__EVAL_20),
    ._EVAL_21(mulAddRecFNToRaw_postMul__EVAL_21),
    ._EVAL_22(mulAddRecFNToRaw_postMul__EVAL_22),
    ._EVAL_23(mulAddRecFNToRaw_postMul__EVAL_23)
  );
  SiFive__EVAL_291 roundRawFNToRecFN (
    ._EVAL(roundRawFNToRecFN__EVAL),
    ._EVAL_0(roundRawFNToRecFN__EVAL_0),
    ._EVAL_1(roundRawFNToRecFN__EVAL_1),
    ._EVAL_2(roundRawFNToRecFN__EVAL_2),
    ._EVAL_3(roundRawFNToRecFN__EVAL_3),
    ._EVAL_4(roundRawFNToRecFN__EVAL_4),
    ._EVAL_5(roundRawFNToRecFN__EVAL_5),
    ._EVAL_6(roundRawFNToRecFN__EVAL_6),
    ._EVAL_7(roundRawFNToRecFN__EVAL_7),
    ._EVAL_8(roundRawFNToRecFN__EVAL_8),
    ._EVAL_9(roundRawFNToRecFN__EVAL_9)
  );
  SiFive__EVAL_288 mulAddRecFNToRaw_preMul (
    ._EVAL(mulAddRecFNToRaw_preMul__EVAL),
    ._EVAL_0(mulAddRecFNToRaw_preMul__EVAL_0),
    ._EVAL_1(mulAddRecFNToRaw_preMul__EVAL_1),
    ._EVAL_2(mulAddRecFNToRaw_preMul__EVAL_2),
    ._EVAL_3(mulAddRecFNToRaw_preMul__EVAL_3),
    ._EVAL_4(mulAddRecFNToRaw_preMul__EVAL_4),
    ._EVAL_5(mulAddRecFNToRaw_preMul__EVAL_5),
    ._EVAL_6(mulAddRecFNToRaw_preMul__EVAL_6),
    ._EVAL_7(mulAddRecFNToRaw_preMul__EVAL_7),
    ._EVAL_8(mulAddRecFNToRaw_preMul__EVAL_8),
    ._EVAL_9(mulAddRecFNToRaw_preMul__EVAL_9),
    ._EVAL_10(mulAddRecFNToRaw_preMul__EVAL_10),
    ._EVAL_11(mulAddRecFNToRaw_preMul__EVAL_11),
    ._EVAL_12(mulAddRecFNToRaw_preMul__EVAL_12),
    ._EVAL_13(mulAddRecFNToRaw_preMul__EVAL_13),
    ._EVAL_14(mulAddRecFNToRaw_preMul__EVAL_14),
    ._EVAL_15(mulAddRecFNToRaw_preMul__EVAL_15),
    ._EVAL_16(mulAddRecFNToRaw_preMul__EVAL_16),
    ._EVAL_17(mulAddRecFNToRaw_preMul__EVAL_17),
    ._EVAL_18(mulAddRecFNToRaw_preMul__EVAL_18),
    ._EVAL_19(mulAddRecFNToRaw_preMul__EVAL_19),
    ._EVAL_20(mulAddRecFNToRaw_preMul__EVAL_20)
  );
  assign _EVAL_18 = mulAddRecFNToRaw_preMul__EVAL_1 * mulAddRecFNToRaw_preMul__EVAL_10;
  assign _EVAL_12 = _EVAL_18 + mulAddRecFNToRaw_preMul__EVAL_13;
  assign mulAddRecFNToRaw_postMul__EVAL_22 = _EVAL_37;
  assign mulAddRecFNToRaw_postMul__EVAL_10 = _EVAL_36;
  assign roundRawFNToRecFN__EVAL_9 = _EVAL_13;
  assign mulAddRecFNToRaw_postMul__EVAL_23 = _EVAL_23;
  assign roundRawFNToRecFN__EVAL_1 = _EVAL_38;
  assign roundRawFNToRecFN__EVAL_3 = _EVAL_29;
  assign _EVAL_7 = roundRawFNToRecFN__EVAL_4;
  assign mulAddRecFNToRaw_preMul__EVAL_17 = _EVAL_5;
  assign mulAddRecFNToRaw_postMul__EVAL_20 = _EVAL_32;
  assign roundRawFNToRecFN__EVAL_8 = 1'h0;
  assign mulAddRecFNToRaw_postMul__EVAL_19 = _EVAL_31;
  assign mulAddRecFNToRaw_postMul__EVAL_1 = _EVAL_30;
  assign mulAddRecFNToRaw_postMul__EVAL_5 = _EVAL_34;
  assign mulAddRecFNToRaw_postMul__EVAL = _EVAL_25;
  assign mulAddRecFNToRaw_postMul__EVAL_0 = _EVAL_24;
  assign mulAddRecFNToRaw_postMul__EVAL_17 = _EVAL_35;
  assign _EVAL_2 = _EVAL_16;
  assign mulAddRecFNToRaw_postMul__EVAL_21 = _EVAL_33;
  assign mulAddRecFNToRaw_postMul__EVAL_7 = _EVAL_21;
  assign mulAddRecFNToRaw_preMul__EVAL = _EVAL_1;
  assign mulAddRecFNToRaw_postMul__EVAL_16 = _EVAL_11;
  assign mulAddRecFNToRaw_postMul__EVAL_2 = _EVAL_27;
  assign _EVAL_8 = roundRawFNToRecFN__EVAL;
  assign mulAddRecFNToRaw_postMul__EVAL_3 = _EVAL_17;
  assign roundRawFNToRecFN__EVAL_2 = _EVAL_14;
  assign mulAddRecFNToRaw_postMul__EVAL_14 = _EVAL_22;
  assign roundRawFNToRecFN__EVAL_6 = _EVAL_15;
  assign mulAddRecFNToRaw_postMul__EVAL_13 = _EVAL_20;
  assign mulAddRecFNToRaw_preMul__EVAL_6 = _EVAL_6;
  assign roundRawFNToRecFN__EVAL_0 = _EVAL_39;
  assign roundRawFNToRecFN__EVAL_7 = _EVAL_26;
  assign roundRawFNToRecFN__EVAL_5 = _EVAL_19;
  assign mulAddRecFNToRaw_postMul__EVAL_4 = _EVAL_10;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_9 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_10 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_11 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_13 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_14 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_15 = _RAND_5[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_16 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_17 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_19 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_20 = _RAND_9[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_21 = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_22 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_23 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_24 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_25 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_26 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_27 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_28 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_29 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_30 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_31 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_32 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_33 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_34 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_35 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _EVAL_36 = _RAND_25[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_37 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_38 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_39 = _RAND_28[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL) begin
    if (_EVAL_4) begin
      _EVAL_9 <= 1'h0;
    end else begin
      _EVAL_9 <= _EVAL_0;
    end
    if (_EVAL_0) begin
      _EVAL_10 <= mulAddRecFNToRaw_preMul__EVAL_3;
    end
    if (_EVAL_0) begin
      _EVAL_11 <= _EVAL_3;
    end
    if (_EVAL_9) begin
      _EVAL_13 <= mulAddRecFNToRaw_postMul__EVAL_9;
    end
    if (_EVAL_9) begin
      _EVAL_14 <= _EVAL_28;
    end
    if (_EVAL_9) begin
      _EVAL_15 <= mulAddRecFNToRaw_postMul__EVAL_18;
    end
    if (_EVAL_4) begin
      _EVAL_16 <= 1'h0;
    end else begin
      _EVAL_16 <= _EVAL_9;
    end
    if (_EVAL_0) begin
      _EVAL_17 <= mulAddRecFNToRaw_preMul__EVAL_18;
    end
    if (_EVAL_9) begin
      _EVAL_19 <= mulAddRecFNToRaw_postMul__EVAL_12;
    end
    if (_EVAL_0) begin
      _EVAL_20 <= mulAddRecFNToRaw_preMul__EVAL_2;
    end
    if (_EVAL_0) begin
      _EVAL_21 <= mulAddRecFNToRaw_preMul__EVAL_20;
    end
    if (_EVAL_0) begin
      _EVAL_22 <= mulAddRecFNToRaw_preMul__EVAL_7;
    end
    if (_EVAL_0) begin
      _EVAL_23 <= mulAddRecFNToRaw_preMul__EVAL_11;
    end
    if (_EVAL_0) begin
      _EVAL_24 <= mulAddRecFNToRaw_preMul__EVAL_8;
    end
    if (_EVAL_0) begin
      _EVAL_25 <= mulAddRecFNToRaw_preMul__EVAL_12;
    end
    if (_EVAL_9) begin
      _EVAL_26 <= mulAddRecFNToRaw_postMul__EVAL_8;
    end
    if (_EVAL_0) begin
      _EVAL_27 <= mulAddRecFNToRaw_preMul__EVAL_19;
    end
    if (_EVAL_0) begin
      _EVAL_28 <= _EVAL_3;
    end
    if (_EVAL_9) begin
      _EVAL_29 <= mulAddRecFNToRaw_postMul__EVAL_6;
    end
    if (_EVAL_0) begin
      _EVAL_30 <= mulAddRecFNToRaw_preMul__EVAL_4;
    end
    if (_EVAL_0) begin
      _EVAL_31 <= mulAddRecFNToRaw_preMul__EVAL_5;
    end
    if (_EVAL_0) begin
      _EVAL_32 <= mulAddRecFNToRaw_preMul__EVAL_14;
    end
    if (_EVAL_0) begin
      _EVAL_33 <= mulAddRecFNToRaw_preMul__EVAL_9;
    end
    if (_EVAL_0) begin
      _EVAL_34 <= mulAddRecFNToRaw_preMul__EVAL_15;
    end
    if (_EVAL_0) begin
      _EVAL_35 <= mulAddRecFNToRaw_preMul__EVAL_0;
    end
    if (_EVAL_0) begin
      _EVAL_36 <= _EVAL_12;
    end
    if (_EVAL_0) begin
      _EVAL_37 <= mulAddRecFNToRaw_preMul__EVAL_16;
    end
    if (_EVAL_9) begin
      _EVAL_38 <= mulAddRecFNToRaw_postMul__EVAL_15;
    end
    if (_EVAL_9) begin
      _EVAL_39 <= mulAddRecFNToRaw_postMul__EVAL_11;
    end
  end
endmodule
