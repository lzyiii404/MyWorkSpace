//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_147(
  input         _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  output [2:0]  _EVAL_3,
  input  [31:0] _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  output        _EVAL_7,
  input  [3:0]  _EVAL_8,
  output        _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [6:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output [31:0] _EVAL_18,
  output [1:0]  _EVAL_19,
  output [24:0] _EVAL_20,
  input  [2:0]  _EVAL_21,
  output        _EVAL_22,
  output [2:0]  _EVAL_23,
  input         _EVAL_24,
  input  [31:0] _EVAL_25,
  input  [31:0] _EVAL_26,
  output        _EVAL_27,
  output [3:0]  _EVAL_28,
  output [1:0]  _EVAL_29,
  input         _EVAL_30,
  output [2:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  output        _EVAL_33,
  input  [2:0]  _EVAL_34,
  output [1:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  input  [6:0]  _EVAL_37,
  output [6:0]  _EVAL_38,
  output [2:0]  _EVAL_39,
  input  [2:0]  _EVAL_40,
  output [2:0]  _EVAL_41,
  output        _EVAL_42,
  input  [6:0]  _EVAL_43,
  input  [24:0] _EVAL_44,
  output [24:0] _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  output [31:0] _EVAL_48,
  output [2:0]  _EVAL_49,
  input         _EVAL_50,
  output [6:0]  _EVAL_51,
  input  [1:0]  _EVAL_52,
  input         _EVAL_53,
  output [3:0]  _EVAL_54,
  output        _EVAL_55,
  output [6:0]  _EVAL_56,
  input  [2:0]  _EVAL_57,
  output [31:0] _EVAL_58,
  input  [1:0]  _EVAL_59,
  input         _EVAL_60
);
  wire [6:0] RationalCrossingSink__EVAL;
  wire [1:0] RationalCrossingSink__EVAL_0;
  wire  RationalCrossingSink__EVAL_1;
  wire  RationalCrossingSink__EVAL_2;
  wire [6:0] RationalCrossingSink__EVAL_3;
  wire  RationalCrossingSink__EVAL_4;
  wire [31:0] RationalCrossingSink__EVAL_5;
  wire  RationalCrossingSink__EVAL_6;
  wire  RationalCrossingSink__EVAL_7;
  wire  RationalCrossingSink__EVAL_8;
  wire  RationalCrossingSink__EVAL_9;
  wire  RationalCrossingSink__EVAL_10;
  wire  RationalCrossingSink__EVAL_11;
  wire  RationalCrossingSink__EVAL_12;
  wire  RationalCrossingSink__EVAL_13;
  wire  RationalCrossingSink__EVAL_14;
  wire [2:0] RationalCrossingSink__EVAL_15;
  wire  RationalCrossingSink__EVAL_16;
  wire [1:0] RationalCrossingSink__EVAL_17;
  wire [31:0] RationalCrossingSink__EVAL_18;
  wire [31:0] RationalCrossingSink__EVAL_19;
  wire [2:0] RationalCrossingSink__EVAL_20;
  wire [6:0] RationalCrossingSink__EVAL_21;
  wire  RationalCrossingSink__EVAL_22;
  wire [2:0] RationalCrossingSink__EVAL_23;
  wire [1:0] RationalCrossingSink__EVAL_24;
  wire [2:0] RationalCrossingSink__EVAL_25;
  wire [2:0] RationalCrossingSink__EVAL_26;
  wire [1:0] RationalCrossingSink__EVAL_27;
  wire [1:0] RationalCrossingSink__EVAL_28;
  wire [2:0] RationalCrossingSink__EVAL_29;
  wire  RationalCrossingSink__EVAL_30;
  wire [2:0] RationalCrossingSource__EVAL;
  wire [1:0] RationalCrossingSource__EVAL_0;
  wire [2:0] RationalCrossingSource__EVAL_1;
  wire [6:0] RationalCrossingSource__EVAL_2;
  wire [31:0] RationalCrossingSource__EVAL_3;
  wire [6:0] RationalCrossingSource__EVAL_4;
  wire  RationalCrossingSource__EVAL_5;
  wire [6:0] RationalCrossingSource__EVAL_6;
  wire [2:0] RationalCrossingSource__EVAL_7;
  wire [2:0] RationalCrossingSource__EVAL_8;
  wire [24:0] RationalCrossingSource__EVAL_9;
  wire  RationalCrossingSource__EVAL_10;
  wire [2:0] RationalCrossingSource__EVAL_11;
  wire [3:0] RationalCrossingSource__EVAL_12;
  wire  RationalCrossingSource__EVAL_13;
  wire [1:0] RationalCrossingSource__EVAL_14;
  wire [24:0] RationalCrossingSource__EVAL_15;
  wire [24:0] RationalCrossingSource__EVAL_16;
  wire [2:0] RationalCrossingSource__EVAL_17;
  wire [2:0] RationalCrossingSource__EVAL_18;
  wire [31:0] RationalCrossingSource__EVAL_19;
  wire  RationalCrossingSource__EVAL_20;
  wire  RationalCrossingSource__EVAL_21;
  wire [3:0] RationalCrossingSource__EVAL_22;
  wire  RationalCrossingSource__EVAL_23;
  wire  RationalCrossingSource__EVAL_24;
  wire [2:0] RationalCrossingSource__EVAL_25;
  wire [3:0] RationalCrossingSource__EVAL_26;
  wire  RationalCrossingSource__EVAL_27;
  wire [2:0] RationalCrossingSource__EVAL_28;
  wire [31:0] RationalCrossingSource__EVAL_29;
  wire  RationalCrossingSource__EVAL_30;
  SiFive__EVAL_146 RationalCrossingSink (
    ._EVAL(RationalCrossingSink__EVAL),
    ._EVAL_0(RationalCrossingSink__EVAL_0),
    ._EVAL_1(RationalCrossingSink__EVAL_1),
    ._EVAL_2(RationalCrossingSink__EVAL_2),
    ._EVAL_3(RationalCrossingSink__EVAL_3),
    ._EVAL_4(RationalCrossingSink__EVAL_4),
    ._EVAL_5(RationalCrossingSink__EVAL_5),
    ._EVAL_6(RationalCrossingSink__EVAL_6),
    ._EVAL_7(RationalCrossingSink__EVAL_7),
    ._EVAL_8(RationalCrossingSink__EVAL_8),
    ._EVAL_9(RationalCrossingSink__EVAL_9),
    ._EVAL_10(RationalCrossingSink__EVAL_10),
    ._EVAL_11(RationalCrossingSink__EVAL_11),
    ._EVAL_12(RationalCrossingSink__EVAL_12),
    ._EVAL_13(RationalCrossingSink__EVAL_13),
    ._EVAL_14(RationalCrossingSink__EVAL_14),
    ._EVAL_15(RationalCrossingSink__EVAL_15),
    ._EVAL_16(RationalCrossingSink__EVAL_16),
    ._EVAL_17(RationalCrossingSink__EVAL_17),
    ._EVAL_18(RationalCrossingSink__EVAL_18),
    ._EVAL_19(RationalCrossingSink__EVAL_19),
    ._EVAL_20(RationalCrossingSink__EVAL_20),
    ._EVAL_21(RationalCrossingSink__EVAL_21),
    ._EVAL_22(RationalCrossingSink__EVAL_22),
    ._EVAL_23(RationalCrossingSink__EVAL_23),
    ._EVAL_24(RationalCrossingSink__EVAL_24),
    ._EVAL_25(RationalCrossingSink__EVAL_25),
    ._EVAL_26(RationalCrossingSink__EVAL_26),
    ._EVAL_27(RationalCrossingSink__EVAL_27),
    ._EVAL_28(RationalCrossingSink__EVAL_28),
    ._EVAL_29(RationalCrossingSink__EVAL_29),
    ._EVAL_30(RationalCrossingSink__EVAL_30)
  );
  SiFive__EVAL_144 RationalCrossingSource (
    ._EVAL(RationalCrossingSource__EVAL),
    ._EVAL_0(RationalCrossingSource__EVAL_0),
    ._EVAL_1(RationalCrossingSource__EVAL_1),
    ._EVAL_2(RationalCrossingSource__EVAL_2),
    ._EVAL_3(RationalCrossingSource__EVAL_3),
    ._EVAL_4(RationalCrossingSource__EVAL_4),
    ._EVAL_5(RationalCrossingSource__EVAL_5),
    ._EVAL_6(RationalCrossingSource__EVAL_6),
    ._EVAL_7(RationalCrossingSource__EVAL_7),
    ._EVAL_8(RationalCrossingSource__EVAL_8),
    ._EVAL_9(RationalCrossingSource__EVAL_9),
    ._EVAL_10(RationalCrossingSource__EVAL_10),
    ._EVAL_11(RationalCrossingSource__EVAL_11),
    ._EVAL_12(RationalCrossingSource__EVAL_12),
    ._EVAL_13(RationalCrossingSource__EVAL_13),
    ._EVAL_14(RationalCrossingSource__EVAL_14),
    ._EVAL_15(RationalCrossingSource__EVAL_15),
    ._EVAL_16(RationalCrossingSource__EVAL_16),
    ._EVAL_17(RationalCrossingSource__EVAL_17),
    ._EVAL_18(RationalCrossingSource__EVAL_18),
    ._EVAL_19(RationalCrossingSource__EVAL_19),
    ._EVAL_20(RationalCrossingSource__EVAL_20),
    ._EVAL_21(RationalCrossingSource__EVAL_21),
    ._EVAL_22(RationalCrossingSource__EVAL_22),
    ._EVAL_23(RationalCrossingSource__EVAL_23),
    ._EVAL_24(RationalCrossingSource__EVAL_24),
    ._EVAL_25(RationalCrossingSource__EVAL_25),
    ._EVAL_26(RationalCrossingSource__EVAL_26),
    ._EVAL_27(RationalCrossingSource__EVAL_27),
    ._EVAL_28(RationalCrossingSource__EVAL_28),
    ._EVAL_29(RationalCrossingSource__EVAL_29),
    ._EVAL_30(RationalCrossingSource__EVAL_30)
  );
  assign _EVAL_16 = RationalCrossingSink__EVAL_25;
  assign RationalCrossingSink__EVAL_30 = _EVAL;
  assign _EVAL_20 = RationalCrossingSource__EVAL_9;
  assign RationalCrossingSource__EVAL_0 = _EVAL_6;
  assign RationalCrossingSink__EVAL_5 = _EVAL_25;
  assign RationalCrossingSource__EVAL_23 = _EVAL_46;
  assign _EVAL_48 = RationalCrossingSource__EVAL_29;
  assign RationalCrossingSink__EVAL_11 = _EVAL_5;
  assign RationalCrossingSink__EVAL_16 = _EVAL_17;
  assign RationalCrossingSource__EVAL_15 = _EVAL_44;
  assign RationalCrossingSink__EVAL_28 = _EVAL_10;
  assign _EVAL_29 = RationalCrossingSink__EVAL_17;
  assign _EVAL_41 = RationalCrossingSource__EVAL_11;
  assign _EVAL_36 = RationalCrossingSource__EVAL_8;
  assign _EVAL_15 = RationalCrossingSource__EVAL_30;
  assign RationalCrossingSink__EVAL_6 = _EVAL_24;
  assign RationalCrossingSource__EVAL_27 = _EVAL_24;
  assign _EVAL_38 = RationalCrossingSource__EVAL_6;
  assign _EVAL_27 = RationalCrossingSource__EVAL_13;
  assign RationalCrossingSink__EVAL_29 = _EVAL_34;
  assign _EVAL_19 = RationalCrossingSource__EVAL_14;
  assign _EVAL_22 = RationalCrossingSink__EVAL_14;
  assign RationalCrossingSource__EVAL_19 = _EVAL_26;
  assign _EVAL_35 = RationalCrossingSink__EVAL_24;
  assign RationalCrossingSink__EVAL = _EVAL_43;
  assign RationalCrossingSink__EVAL_0 = _EVAL_59;
  assign RationalCrossingSource__EVAL_1 = _EVAL_32;
  assign RationalCrossingSource__EVAL_12 = _EVAL_8;
  assign _EVAL_51 = RationalCrossingSource__EVAL_2;
  assign _EVAL_9 = RationalCrossingSink__EVAL_8;
  assign _EVAL_31 = RationalCrossingSink__EVAL_15;
  assign RationalCrossingSink__EVAL_12 = _EVAL_0;
  assign RationalCrossingSink__EVAL_26 = _EVAL_40;
  assign RationalCrossingSink__EVAL_9 = _EVAL_30;
  assign _EVAL_56 = RationalCrossingSink__EVAL_21;
  assign RationalCrossingSink__EVAL_22 = _EVAL_2;
  assign _EVAL_45 = RationalCrossingSource__EVAL_16;
  assign RationalCrossingSink__EVAL_13 = _EVAL_50;
  assign _EVAL_3 = RationalCrossingSource__EVAL_7;
  assign RationalCrossingSource__EVAL_18 = _EVAL_12;
  assign _EVAL_49 = RationalCrossingSource__EVAL_17;
  assign _EVAL_14 = RationalCrossingSink__EVAL_10;
  assign RationalCrossingSink__EVAL_27 = _EVAL_52;
  assign RationalCrossingSource__EVAL_4 = _EVAL_11;
  assign _EVAL_58 = RationalCrossingSource__EVAL_3;
  assign RationalCrossingSink__EVAL_2 = _EVAL_47;
  assign RationalCrossingSink__EVAL_19 = _EVAL_4;
  assign RationalCrossingSink__EVAL_3 = _EVAL_37;
  assign _EVAL_54 = RationalCrossingSource__EVAL_22;
  assign RationalCrossingSource__EVAL_20 = _EVAL;
  assign _EVAL_39 = RationalCrossingSource__EVAL;
  assign RationalCrossingSink__EVAL_20 = _EVAL_1;
  assign RationalCrossingSource__EVAL_24 = _EVAL_13;
  assign _EVAL_42 = RationalCrossingSource__EVAL_5;
  assign _EVAL_23 = RationalCrossingSource__EVAL_28;
  assign _EVAL_18 = RationalCrossingSink__EVAL_18;
  assign _EVAL_33 = RationalCrossingSink__EVAL_7;
  assign RationalCrossingSink__EVAL_23 = _EVAL_57;
  assign RationalCrossingSource__EVAL_21 = _EVAL_53;
  assign RationalCrossingSource__EVAL_25 = _EVAL_21;
  assign _EVAL_7 = RationalCrossingSource__EVAL_10;
  assign _EVAL_28 = RationalCrossingSource__EVAL_26;
  assign RationalCrossingSink__EVAL_4 = _EVAL_60;
  assign _EVAL_55 = RationalCrossingSink__EVAL_1;
endmodule
