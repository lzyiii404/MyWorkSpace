//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_96_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  input         _EVAL_11,
  input  [7:0]  _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_22;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_40;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_47;
  reg [31:0] _RAND_2;
  reg  _EVAL_50;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_124;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_128;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_139;
  reg [31:0] _RAND_6;
  reg  _EVAL_169;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_172;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_185;
  reg [31:0] _RAND_9;
  reg [31:0] _EVAL_244;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_249;
  reg [31:0] _RAND_11;
  reg  _EVAL_257;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_262;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_269;
  reg [31:0] _RAND_14;
  wire  _EVAL_205;
  wire [1:0] _EVAL_141;
  wire [3:0] _EVAL_196;
  wire [2:0] _EVAL_184;
  wire [2:0] _EVAL_95;
  wire  _EVAL_122;
  wire  _EVAL_116;
  wire  _EVAL_250;
  wire  _EVAL_146;
  wire  _EVAL_110;
  wire  _EVAL_263;
  wire  _EVAL_236;
  wire  _EVAL_63;
  wire  _EVAL_271;
  wire  _EVAL_254;
  wire  _EVAL_154;
  wire  _EVAL_27;
  wire  _EVAL_25;
  wire  _EVAL_82;
  wire  _EVAL_157;
  wire  _EVAL_38;
  wire  _EVAL_77;
  wire [1:0] _EVAL_24;
  wire [1:0] _EVAL_30;
  wire [1:0] _EVAL_219;
  wire [1:0] _EVAL_170;
  wire  _EVAL_255;
  wire  _EVAL_224;
  wire  _EVAL_86;
  wire  _EVAL_94;
  wire  _EVAL_256;
  wire  _EVAL_214;
  wire  _EVAL_117;
  wire  _EVAL_207;
  wire  _EVAL_57;
  wire  _EVAL_189;
  wire  _EVAL_140;
  wire  _EVAL_174;
  wire  _EVAL_156;
  wire  _EVAL_119;
  wire [31:0] _EVAL_162;
  wire [32:0] _EVAL_155;
  wire [32:0] _EVAL_29;
  wire [12:0] _EVAL_52;
  wire [5:0] _EVAL_267;
  wire [5:0] _EVAL_131;
  wire [2:0] _EVAL_26;
  wire  _EVAL_100;
  wire  _EVAL_167;
  wire  _EVAL_144;
  wire  _EVAL_106;
  wire  _EVAL_251;
  wire  _EVAL_268;
  wire  _EVAL_83;
  wire [31:0] _EVAL_164;
  wire [31:0] _EVAL_217;
  wire  _EVAL_134;
  wire  _EVAL_81;
  wire  _EVAL_148;
  wire  _EVAL_278;
  wire  _EVAL_109;
  wire  _EVAL_213;
  wire  _EVAL_151;
  wire  _EVAL_274;
  wire  _EVAL_143;
  wire  _EVAL_49;
  wire  _EVAL_136;
  wire  _EVAL_135;
  wire [1:0] _EVAL_101;
  wire [1:0] _EVAL_152;
  wire  _EVAL_186;
  wire [12:0] _EVAL_48;
  wire [5:0] _EVAL_105;
  wire [5:0] _EVAL_175;
  wire [2:0] _EVAL_17;
  wire  _EVAL_264;
  wire  _EVAL_177;
  wire  _EVAL_191;
  wire  _EVAL_266;
  wire  _EVAL_190;
  wire  _EVAL_80;
  wire  _EVAL_243;
  wire  _EVAL_61;
  wire  _EVAL_234;
  wire  _EVAL_142;
  wire  _EVAL_273;
  wire  _EVAL_64;
  wire  _EVAL_69;
  wire [7:0] _EVAL_253;
  wire  _EVAL_112;
  wire  _EVAL_178;
  wire  _EVAL_129;
  wire  _EVAL_212;
  wire [32:0] _EVAL_92;
  wire  _EVAL_78;
  wire  _EVAL_259;
  wire  _EVAL_79;
  wire  _EVAL_195;
  wire  _EVAL_132;
  wire  _EVAL_280;
  wire  _EVAL_147;
  wire  _EVAL_235;
  wire  _EVAL_130;
  wire  _EVAL_23;
  wire  _EVAL_173;
  wire  _EVAL_171;
  wire  _EVAL_62;
  wire  _EVAL_206;
  wire  _EVAL_19;
  wire  _EVAL_67;
  wire  _EVAL_229;
  wire  _EVAL_261;
  wire  _EVAL_265;
  wire  _EVAL_179;
  wire  _EVAL_222;
  wire  _EVAL_187;
  wire  _EVAL_59;
  wire  _EVAL_211;
  wire  _EVAL_36;
  wire  _EVAL_56;
  wire  _EVAL_123;
  wire  _EVAL_209;
  wire  _EVAL_281;
  wire  _EVAL_176;
  wire  _EVAL_242;
  wire  _EVAL_65;
  wire  _EVAL_193;
  wire  _EVAL_272;
  wire  _EVAL_85;
  wire  _EVAL_283;
  wire  _EVAL_201;
  wire [7:0] _EVAL_197;
  wire [7:0] _EVAL_192;
  wire [7:0] _EVAL_125;
  wire  _EVAL_99;
  wire  _EVAL_188;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_34;
  wire  _EVAL_210;
  wire  _EVAL_220;
  wire  _EVAL_102;
  wire  _EVAL_248;
  wire  _EVAL_113;
  wire  _EVAL_183;
  wire  _EVAL_89;
  wire  _EVAL_161;
  wire  _EVAL_90;
  wire  _EVAL_163;
  wire  _EVAL_73;
  wire  _EVAL_28;
  wire  _EVAL_74;
  wire  _EVAL_194;
  wire  _EVAL_226;
  wire  _EVAL_111;
  wire  _EVAL_43;
  wire  _EVAL_133;
  wire  _EVAL_104;
  wire  _EVAL_252;
  wire  _EVAL_198;
  wire  _EVAL_228;
  wire [2:0] _EVAL_223;
  wire  _EVAL_182;
  wire [1:0] _EVAL_165;
  wire  _EVAL_42;
  wire  _EVAL_120;
  wire  _EVAL_159;
  wire  _EVAL_70;
  wire [2:0] _EVAL_240;
  wire  _EVAL_66;
  wire  _EVAL_45;
  wire  _EVAL_246;
  wire  _EVAL_20;
  wire  _EVAL_44;
  wire [31:0] _EVAL_115;
  wire  _EVAL_160;
  wire  _EVAL_279;
  wire  _EVAL_166;
  wire  _EVAL_239;
  wire  _EVAL_153;
  wire  _EVAL_276;
  wire  _EVAL_208;
  wire  _EVAL_137;
  wire  _EVAL_84;
  wire  _EVAL_275;
  wire  _EVAL_96;
  wire  _EVAL_258;
  wire [1:0] _EVAL_18;
  wire [1:0] _EVAL_230;
  wire [1:0] _EVAL_37;
  wire  _EVAL_181;
  wire  _EVAL_75;
  wire  _EVAL_260;
  wire  _EVAL_46;
  wire  _EVAL_277;
  wire  _EVAL_233;
  wire  _EVAL_282;
  wire  _EVAL_31;
  wire [2:0] _EVAL_158;
  wire  _EVAL_221;
  wire  _EVAL_21;
  wire  _EVAL_216;
  wire  _EVAL_232;
  wire  _EVAL_145;
  wire  _EVAL_87;
  wire  _EVAL_41;
  wire  _EVAL_76;
  wire  _EVAL_150;
  wire  _EVAL_60;
  wire  _EVAL_35;
  wire  _EVAL_138;
  wire  _EVAL_71;
  wire [2:0] _EVAL_91;
  wire  _EVAL_93;
  wire  _EVAL_241;
  wire  _EVAL_72;
  wire  _EVAL_58;
  wire  _EVAL_39;
  wire  _EVAL_202;
  wire  _EVAL_97;
  wire  _EVAL_227;
  wire  _EVAL_55;
  wire  _EVAL_118;
  wire  _EVAL_32;
  wire  _EVAL_126;
  wire  _EVAL_231;
  wire  _EVAL_53;
  wire  _EVAL_103;
  wire  _EVAL_168;
  wire  _EVAL_68;
  wire  _EVAL_270;
  wire  _EVAL_245;
  wire  _EVAL_114;
  wire  _EVAL_88;
  wire  _EVAL_204;
  wire  _EVAL_218;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_205 = _EVAL_7 >= 3'h3;
  assign _EVAL_141 = _EVAL_7[1:0];
  assign _EVAL_196 = 4'h1 << _EVAL_141;
  assign _EVAL_184 = _EVAL_196[2:0];
  assign _EVAL_95 = _EVAL_184 | 3'h1;
  assign _EVAL_122 = _EVAL_95[2];
  assign _EVAL_116 = _EVAL_10[2];
  assign _EVAL_250 = _EVAL_116 == 1'h0;
  assign _EVAL_146 = _EVAL_122 & _EVAL_250;
  assign _EVAL_110 = _EVAL_205 | _EVAL_146;
  assign _EVAL_263 = _EVAL_95[1];
  assign _EVAL_236 = _EVAL_10[1];
  assign _EVAL_63 = _EVAL_250 & _EVAL_236;
  assign _EVAL_271 = _EVAL_263 & _EVAL_63;
  assign _EVAL_254 = _EVAL_110 | _EVAL_271;
  assign _EVAL_154 = _EVAL_3 <= 3'h6;
  assign _EVAL_27 = _EVAL_7 == _EVAL_185;
  assign _EVAL_25 = _EVAL_27 | _EVAL_8;
  assign _EVAL_82 = _EVAL_25 == 1'h0;
  assign _EVAL_157 = _EVAL_15 & _EVAL_5;
  assign _EVAL_38 = _EVAL_47 == 3'h0;
  assign _EVAL_77 = _EVAL_157 & _EVAL_38;
  assign _EVAL_24 = 2'h1 << _EVAL_1;
  assign _EVAL_30 = _EVAL_77 ? _EVAL_24 : 2'h0;
  assign _EVAL_219 = _EVAL_30 | _EVAL_249;
  assign _EVAL_170 = _EVAL_219 >> _EVAL_11;
  assign _EVAL_255 = _EVAL_95[0];
  assign _EVAL_224 = _EVAL_236 == 1'h0;
  assign _EVAL_86 = _EVAL_116 & _EVAL_224;
  assign _EVAL_94 = _EVAL_10[0];
  assign _EVAL_256 = _EVAL_86 & _EVAL_94;
  assign _EVAL_214 = _EVAL_255 & _EVAL_256;
  assign _EVAL_117 = _EVAL_6 == 1'h0;
  assign _EVAL_207 = _EVAL_117 | _EVAL;
  assign _EVAL_57 = _EVAL_6 == _EVAL_169;
  assign _EVAL_189 = _EVAL_14[2];
  assign _EVAL_140 = _EVAL_189 == 1'h0;
  assign _EVAL_174 = _EVAL_14 == 3'h2;
  assign _EVAL_156 = _EVAL_4 == _EVAL_124;
  assign _EVAL_119 = _EVAL_3 == 3'h4;
  assign _EVAL_162 = _EVAL_10 ^ 32'h80000000;
  assign _EVAL_155 = {1'b0,$signed(_EVAL_162)};
  assign _EVAL_29 = $signed(_EVAL_155) & $signed(-33'sh20000);
  assign _EVAL_52 = 13'h3f << _EVAL_7;
  assign _EVAL_267 = _EVAL_52[5:0];
  assign _EVAL_131 = ~ _EVAL_267;
  assign _EVAL_26 = _EVAL_131[5:3];
  assign _EVAL_100 = _EVAL == 1'h0;
  assign _EVAL_167 = _EVAL_100 | _EVAL_8;
  assign _EVAL_144 = _EVAL_3 == 3'h0;
  assign _EVAL_106 = _EVAL_1 == _EVAL_50;
  assign _EVAL_251 = _EVAL_106 | _EVAL_8;
  assign _EVAL_268 = _EVAL_94 == 1'h0;
  assign _EVAL_83 = _EVAL_63 & _EVAL_268;
  assign _EVAL_164 = {{26'd0}, _EVAL_131};
  assign _EVAL_217 = _EVAL_10 & _EVAL_164;
  assign _EVAL_134 = _EVAL_217 == 32'h0;
  assign _EVAL_81 = _EVAL_134 | _EVAL_8;
  assign _EVAL_148 = _EVAL_81 == 1'h0;
  assign _EVAL_278 = _EVAL_63 & _EVAL_94;
  assign _EVAL_109 = _EVAL_4 >= 3'h3;
  assign _EVAL_213 = _EVAL_109 | _EVAL_8;
  assign _EVAL_151 = _EVAL_9 & _EVAL_16;
  assign _EVAL_274 = _EVAL_139 == 3'h0;
  assign _EVAL_143 = _EVAL_151 & _EVAL_274;
  assign _EVAL_49 = _EVAL_3 == 3'h6;
  assign _EVAL_136 = _EVAL_49 == 1'h0;
  assign _EVAL_135 = _EVAL_143 & _EVAL_136;
  assign _EVAL_101 = 2'h1 << _EVAL_11;
  assign _EVAL_152 = _EVAL_135 ? _EVAL_101 : 2'h0;
  assign _EVAL_186 = _EVAL_3[0];
  assign _EVAL_48 = 13'h3f << _EVAL_4;
  assign _EVAL_105 = _EVAL_48[5:0];
  assign _EVAL_175 = ~ _EVAL_105;
  assign _EVAL_17 = _EVAL_175[5:3];
  assign _EVAL_264 = _EVAL_172 == 3'h0;
  assign _EVAL_177 = _EVAL_157 & _EVAL_264;
  assign _EVAL_191 = _EVAL_14 == 3'h4;
  assign _EVAL_266 = _EVAL_13 == 1'h0;
  assign _EVAL_190 = _EVAL_266 | _EVAL_8;
  assign _EVAL_80 = _EVAL_2 == _EVAL_22;
  assign _EVAL_243 = _EVAL_80 | _EVAL_8;
  assign _EVAL_61 = _EVAL_243 == 1'h0;
  assign _EVAL_234 = _EVAL_86 & _EVAL_268;
  assign _EVAL_142 = _EVAL_255 & _EVAL_234;
  assign _EVAL_273 = _EVAL_116 & _EVAL_236;
  assign _EVAL_64 = _EVAL_273 & _EVAL_268;
  assign _EVAL_69 = _EVAL_255 & _EVAL_64;
  assign _EVAL_253 = ~ _EVAL_12;
  assign _EVAL_112 = _EVAL_253 == 8'h0;
  assign _EVAL_178 = _EVAL_2 <= 3'h2;
  assign _EVAL_129 = _EVAL_178 | _EVAL_8;
  assign _EVAL_212 = _EVAL_129 == 1'h0;
  assign _EVAL_92 = $signed(_EVAL_29);
  assign _EVAL_78 = _EVAL_11 == _EVAL_257;
  assign _EVAL_259 = _EVAL_78 | _EVAL_8;
  assign _EVAL_79 = _EVAL_250 & _EVAL_224;
  assign _EVAL_195 = _EVAL_2 <= 3'h3;
  assign _EVAL_132 = _EVAL_30 != 2'h0;
  assign _EVAL_280 = _EVAL_132 == 1'h0;
  assign _EVAL_147 = _EVAL_14 == 3'h7;
  assign _EVAL_235 = _EVAL_30 != _EVAL_152;
  assign _EVAL_130 = _EVAL_263 & _EVAL_79;
  assign _EVAL_23 = _EVAL_122 & _EVAL_116;
  assign _EVAL_173 = _EVAL_205 | _EVAL_8;
  assign _EVAL_171 = _EVAL_3 == _EVAL_269;
  assign _EVAL_62 = _EVAL_171 | _EVAL_8;
  assign _EVAL_206 = _EVAL_62 == 1'h0;
  assign _EVAL_19 = _EVAL_14 == 3'h5;
  assign _EVAL_67 = _EVAL_110 | _EVAL_130;
  assign _EVAL_229 = _EVAL_79 & _EVAL_94;
  assign _EVAL_261 = _EVAL_255 & _EVAL_229;
  assign _EVAL_265 = _EVAL_67 | _EVAL_261;
  assign _EVAL_179 = _EVAL_255 & _EVAL_83;
  assign _EVAL_222 = _EVAL_205 | _EVAL_23;
  assign _EVAL_187 = _EVAL_263 & _EVAL_273;
  assign _EVAL_59 = _EVAL_222 | _EVAL_187;
  assign _EVAL_211 = _EVAL_273 & _EVAL_94;
  assign _EVAL_36 = _EVAL_255 & _EVAL_211;
  assign _EVAL_56 = _EVAL_59 | _EVAL_36;
  assign _EVAL_123 = _EVAL_59 | _EVAL_69;
  assign _EVAL_209 = _EVAL_263 & _EVAL_86;
  assign _EVAL_281 = _EVAL_222 | _EVAL_209;
  assign _EVAL_176 = _EVAL_281 | _EVAL_214;
  assign _EVAL_242 = _EVAL_281 | _EVAL_142;
  assign _EVAL_65 = _EVAL_255 & _EVAL_278;
  assign _EVAL_193 = _EVAL_254 | _EVAL_65;
  assign _EVAL_272 = _EVAL_254 | _EVAL_179;
  assign _EVAL_85 = _EVAL_79 & _EVAL_268;
  assign _EVAL_283 = _EVAL_255 & _EVAL_85;
  assign _EVAL_201 = _EVAL_67 | _EVAL_283;
  assign _EVAL_197 = {_EVAL_56,_EVAL_123,_EVAL_176,_EVAL_242,_EVAL_193,_EVAL_272,_EVAL_265,_EVAL_201};
  assign _EVAL_192 = ~ _EVAL_197;
  assign _EVAL_125 = _EVAL_12 & _EVAL_192;
  assign _EVAL_99 = _EVAL_125 == 8'h0;
  assign _EVAL_188 = _EVAL_99 | _EVAL_8;
  assign _EVAL_237 = _EVAL_213 == 1'h0;
  assign _EVAL_238 = _EVAL_14 == _EVAL_128;
  assign _EVAL_34 = _EVAL_238 | _EVAL_8;
  assign _EVAL_210 = _EVAL_34 == 1'h0;
  assign _EVAL_220 = _EVAL_14 == 3'h6;
  assign _EVAL_102 = _EVAL_5 & _EVAL_220;
  assign _EVAL_248 = _EVAL_156 | _EVAL_8;
  assign _EVAL_113 = _EVAL_248 == 1'h0;
  assign _EVAL_183 = _EVAL_7 <= 3'h6;
  assign _EVAL_89 = $signed(_EVAL_92) == $signed(33'sh0);
  assign _EVAL_161 = _EVAL_183 & _EVAL_89;
  assign _EVAL_90 = _EVAL_161 | _EVAL_8;
  assign _EVAL_163 = _EVAL_90 == 1'h0;
  assign _EVAL_73 = _EVAL_10 == _EVAL_244;
  assign _EVAL_28 = _EVAL_16 & _EVAL_119;
  assign _EVAL_74 = _EVAL_235 | _EVAL_280;
  assign _EVAL_194 = _EVAL_74 | _EVAL_8;
  assign _EVAL_226 = _EVAL_194 == 1'h0;
  assign _EVAL_111 = _EVAL_3 == 3'h5;
  assign _EVAL_43 = _EVAL_5 & _EVAL_19;
  assign _EVAL_133 = _EVAL_2 != 3'h0;
  assign _EVAL_104 = _EVAL_133 | _EVAL_8;
  assign _EVAL_252 = _EVAL_104 == 1'h0;
  assign _EVAL_198 = _EVAL_264 == 1'h0;
  assign _EVAL_228 = _EVAL_5 & _EVAL_198;
  assign _EVAL_223 = _EVAL_172 - 3'h1;
  assign _EVAL_182 = _EVAL_170[0];
  assign _EVAL_165 = _EVAL_249 >> _EVAL_1;
  assign _EVAL_42 = _EVAL_165[0];
  assign _EVAL_120 = _EVAL_42 == 1'h0;
  assign _EVAL_159 = _EVAL_120 | _EVAL_8;
  assign _EVAL_70 = _EVAL_40 == 3'h0;
  assign _EVAL_240 = _EVAL_40 - 3'h1;
  assign _EVAL_66 = plusarg_reader_out == 32'h0;
  assign _EVAL_45 = _EVAL_195 | _EVAL_8;
  assign _EVAL_246 = _EVAL_45 == 1'h0;
  assign _EVAL_20 = _EVAL_14 == 3'h1;
  assign _EVAL_44 = _EVAL_14 == 3'h0;
  assign _EVAL_115 = _EVAL_262 + 32'h1;
  assign _EVAL_160 = _EVAL_173 == 1'h0;
  assign _EVAL_279 = _EVAL_249 != 2'h0;
  assign _EVAL_166 = _EVAL_279 == 1'h0;
  assign _EVAL_239 = _EVAL_166 | _EVAL_66;
  assign _EVAL_153 = _EVAL_262 < plusarg_reader_out;
  assign _EVAL_276 = _EVAL_239 | _EVAL_153;
  assign _EVAL_208 = _EVAL_276 | _EVAL_8;
  assign _EVAL_137 = _EVAL_208 == 1'h0;
  assign _EVAL_84 = _EVAL_182 | _EVAL_8;
  assign _EVAL_275 = _EVAL_84 == 1'h0;
  assign _EVAL_96 = _EVAL_154 | _EVAL_8;
  assign _EVAL_258 = _EVAL_96 == 1'h0;
  assign _EVAL_18 = _EVAL_249 | _EVAL_30;
  assign _EVAL_230 = ~ _EVAL_152;
  assign _EVAL_37 = _EVAL_18 & _EVAL_230;
  assign _EVAL_181 = _EVAL_207 | _EVAL_8;
  assign _EVAL_75 = _EVAL_181 == 1'h0;
  assign _EVAL_260 = _EVAL_3 == 3'h1;
  assign _EVAL_46 = _EVAL_14 == 3'h3;
  assign _EVAL_277 = _EVAL_2 == 3'h0;
  assign _EVAL_233 = _EVAL_277 | _EVAL_8;
  assign _EVAL_282 = _EVAL_233 == 1'h0;
  assign _EVAL_31 = _EVAL_16 & _EVAL_49;
  assign _EVAL_158 = _EVAL_47 - 3'h1;
  assign _EVAL_221 = _EVAL_57 | _EVAL_8;
  assign _EVAL_21 = _EVAL_221 == 1'h0;
  assign _EVAL_216 = _EVAL_5 & _EVAL_44;
  assign _EVAL_232 = _EVAL_2 <= 3'h4;
  assign _EVAL_145 = _EVAL_12 == _EVAL_197;
  assign _EVAL_87 = _EVAL_73 | _EVAL_8;
  assign _EVAL_41 = _EVAL_117 | _EVAL_8;
  assign _EVAL_76 = _EVAL_41 == 1'h0;
  assign _EVAL_150 = _EVAL_5 & _EVAL_46;
  assign _EVAL_60 = _EVAL_167 == 1'h0;
  assign _EVAL_35 = _EVAL_5 & _EVAL_191;
  assign _EVAL_138 = _EVAL_3 == 3'h2;
  assign _EVAL_71 = _EVAL_16 & _EVAL_138;
  assign _EVAL_91 = _EVAL_139 - 3'h1;
  assign _EVAL_93 = _EVAL_251 == 1'h0;
  assign _EVAL_241 = _EVAL_112 | _EVAL_8;
  assign _EVAL_72 = _EVAL_241 == 1'h0;
  assign _EVAL_58 = _EVAL_16 & _EVAL_260;
  assign _EVAL_39 = _EVAL_232 | _EVAL_8;
  assign _EVAL_202 = _EVAL_8 == 1'h0;
  assign _EVAL_97 = _EVAL_159 == 1'h0;
  assign _EVAL_227 = _EVAL_190 == 1'h0;
  assign _EVAL_55 = _EVAL_157 | _EVAL_151;
  assign _EVAL_118 = _EVAL_145 | _EVAL_8;
  assign _EVAL_32 = _EVAL_5 & _EVAL_147;
  assign _EVAL_126 = _EVAL_39 == 1'h0;
  assign _EVAL_231 = _EVAL_259 == 1'h0;
  assign _EVAL_53 = _EVAL_118 == 1'h0;
  assign _EVAL_103 = _EVAL_87 == 1'h0;
  assign _EVAL_168 = _EVAL_70 == 1'h0;
  assign _EVAL_68 = _EVAL_16 & _EVAL_168;
  assign _EVAL_270 = _EVAL_16 & _EVAL_111;
  assign _EVAL_245 = _EVAL_5 & _EVAL_20;
  assign _EVAL_114 = _EVAL_151 & _EVAL_70;
  assign _EVAL_88 = _EVAL_5 & _EVAL_174;
  assign _EVAL_204 = _EVAL_188 == 1'h0;
  assign _EVAL_218 = _EVAL_16 & _EVAL_144;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_40 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_47 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_50 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_124 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_128 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_139 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_169 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_172 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_185 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_244 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_249 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_257 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_262 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_269 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_177) begin
      _EVAL_22 <= _EVAL_2;
    end
    if (_EVAL_8) begin
      _EVAL_40 <= 3'h0;
    end else begin
      if (_EVAL_151) begin
        if (_EVAL_70) begin
          if (_EVAL_186) begin
            _EVAL_40 <= _EVAL_17;
          end else begin
            _EVAL_40 <= 3'h0;
          end
        end else begin
          _EVAL_40 <= _EVAL_240;
        end
      end
    end
    if (_EVAL_8) begin
      _EVAL_47 <= 3'h0;
    end else begin
      if (_EVAL_157) begin
        if (_EVAL_38) begin
          if (_EVAL_140) begin
            _EVAL_47 <= _EVAL_26;
          end else begin
            _EVAL_47 <= 3'h0;
          end
        end else begin
          _EVAL_47 <= _EVAL_158;
        end
      end
    end
    if (_EVAL_177) begin
      _EVAL_50 <= _EVAL_1;
    end
    if (_EVAL_114) begin
      _EVAL_124 <= _EVAL_4;
    end
    if (_EVAL_177) begin
      _EVAL_128 <= _EVAL_14;
    end
    if (_EVAL_8) begin
      _EVAL_139 <= 3'h0;
    end else begin
      if (_EVAL_151) begin
        if (_EVAL_274) begin
          if (_EVAL_186) begin
            _EVAL_139 <= _EVAL_17;
          end else begin
            _EVAL_139 <= 3'h0;
          end
        end else begin
          _EVAL_139 <= _EVAL_91;
        end
      end
    end
    if (_EVAL_114) begin
      _EVAL_169 <= _EVAL_6;
    end
    if (_EVAL_8) begin
      _EVAL_172 <= 3'h0;
    end else begin
      if (_EVAL_157) begin
        if (_EVAL_264) begin
          if (_EVAL_140) begin
            _EVAL_172 <= _EVAL_26;
          end else begin
            _EVAL_172 <= 3'h0;
          end
        end else begin
          _EVAL_172 <= _EVAL_223;
        end
      end
    end
    if (_EVAL_177) begin
      _EVAL_185 <= _EVAL_7;
    end
    if (_EVAL_177) begin
      _EVAL_244 <= _EVAL_10;
    end
    if (_EVAL_8) begin
      _EVAL_249 <= 2'h0;
    end else begin
      _EVAL_249 <= _EVAL_37;
    end
    if (_EVAL_114) begin
      _EVAL_257 <= _EVAL_11;
    end
    if (_EVAL_8) begin
      _EVAL_262 <= 32'h0;
    end else begin
      if (_EVAL_55) begin
        _EVAL_262 <= 32'h0;
      end else begin
        _EVAL_262 <= _EVAL_115;
      end
    end
    if (_EVAL_114) begin
      _EVAL_269 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a06ded2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d76eb22d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c337960)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ef3002e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903b7d90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3935710)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6a598be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1057ef2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1bd71fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec9379f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ad77dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a2e0a00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cd658ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d710224e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b251817)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa69b0ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d408c0a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(240d1035)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fadb5151)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13e4113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b6a6aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48a17114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79d96399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8adaad9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccbefb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b3ab547)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cb9961d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cfafc7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e307c24f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eff63031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fc5e871)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9645df2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59886bad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f14dd24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbcd2ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb36814f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f761b56b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(860f7d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3c080c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(139b6cd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5d34a34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95822163)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7393617)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5ab3cad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3270a85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2f7b7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cee8acb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ff36632)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ffbe1d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a53efa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1da79672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(640968fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68a71cfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec2e4c1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66337432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9b89cec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31465f35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f2ffd45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(409bc1cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(423b0965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be01676a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6314659d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a97401d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97d6c362)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3543bdbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91cfae7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
