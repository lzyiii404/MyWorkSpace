//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_265_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [7:0]  _EVAL_1,
  input  [3:0]  _EVAL_2,
  input         _EVAL_3,
  input  [31:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input  [3:0]  _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input  [3:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [3:0]  _EVAL_25,
  input  [3:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [2:0]  _EVAL_28,
  input         _EVAL_29,
  input  [1:0]  _EVAL_30,
  input  [1:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  input         _EVAL_33
);
  wire [31:0] plusarg_reader_out;
  reg [31:0] _EVAL_82;
  reg [31:0] _RAND_0;
  reg [8:0] _EVAL_100;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_113;
  reg [31:0] _RAND_2;
  reg [4:0] _EVAL_120;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_133;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_138;
  reg [31:0] _RAND_5;
  reg [31:0] _EVAL_149;
  reg [31:0] _RAND_6;
  reg  _EVAL_150;
  reg [31:0] _RAND_7;
  reg [4:0] _EVAL_159;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_219;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_252;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_255;
  reg [31:0] _RAND_11;
  reg [1:0] _EVAL_280;
  reg [31:0] _RAND_12;
  reg [4:0] _EVAL_356;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_358;
  reg [31:0] _RAND_14;
  reg [31:0] _EVAL_407;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_415;
  reg [31:0] _RAND_16;
  reg [3:0] _EVAL_417;
  reg [31:0] _RAND_17;
  reg [2:0] _EVAL_424;
  reg [31:0] _RAND_18;
  reg  _EVAL_425;
  reg [31:0] _RAND_19;
  reg [4:0] _EVAL_447;
  reg [31:0] _RAND_20;
  reg [3:0] _EVAL_499;
  reg [31:0] _RAND_21;
  reg [1:0] _EVAL_540;
  reg [31:0] _RAND_22;
  reg [3:0] _EVAL_543;
  reg [31:0] _RAND_23;
  reg [1:0] _EVAL_548;
  reg [31:0] _RAND_24;
  reg [31:0] _EVAL_559;
  reg [31:0] _RAND_25;
  reg [3:0] _EVAL_568;
  reg [31:0] _RAND_26;
  reg [4:0] _EVAL_669;
  reg [31:0] _RAND_27;
  wire [31:0] _EVAL_471;
  wire [32:0] _EVAL_398;
  wire  _EVAL_61;
  wire [1:0] _EVAL_221;
  wire [3:0] _EVAL_522;
  wire [2:0] _EVAL_551;
  wire [2:0] _EVAL_655;
  wire  _EVAL_641;
  wire  _EVAL_194;
  wire  _EVAL_182;
  wire  _EVAL_224;
  wire  _EVAL_315;
  wire  _EVAL_464;
  wire  _EVAL_328;
  wire  _EVAL_592;
  wire  _EVAL_591;
  wire  _EVAL_364;
  wire  _EVAL_176;
  wire  _EVAL_55;
  wire  _EVAL_590;
  wire  _EVAL_177;
  wire  _EVAL_154;
  wire  _EVAL_222;
  wire [31:0] _EVAL_426;
  wire [32:0] _EVAL_186;
  wire [32:0] _EVAL_560;
  wire [32:0] _EVAL_405;
  wire  _EVAL_112;
  wire [4:0] _EVAL_497;
  wire [4:0] _EVAL_171;
  wire [31:0] _EVAL_203;
  wire [32:0] _EVAL_501;
  wire  _EVAL_505;
  wire  _EVAL_68;
  wire [4:0] _EVAL_365;
  wire  _EVAL_429;
  wire [15:0] _EVAL_310;
  wire [31:0] _EVAL_309;
  wire [32:0] _EVAL_508;
  wire [32:0] _EVAL_193;
  wire [31:0] _EVAL_498;
  wire [32:0] _EVAL_466;
  wire [32:0] _EVAL_452;
  wire [32:0] _EVAL_545;
  wire  _EVAL_156;
  wire [7:0] _EVAL_279;
  wire  _EVAL_187;
  wire  _EVAL_173;
  wire  _EVAL_293;
  wire  _EVAL_596;
  wire  _EVAL_51;
  wire  _EVAL_250;
  wire [2:0] _EVAL_401;
  wire  _EVAL_262;
  wire  _EVAL_66;
  wire  _EVAL_136;
  wire  _EVAL_605;
  wire  _EVAL_645;
  wire  _EVAL_146;
  wire  _EVAL_496;
  wire  _EVAL_103;
  wire  _EVAL_403;
  wire  _EVAL_244;
  wire  _EVAL_384;
  wire [31:0] _EVAL_406;
  wire [32:0] _EVAL_649;
  wire [31:0] _EVAL_316;
  wire [32:0] _EVAL_75;
  wire [32:0] _EVAL_614;
  wire [32:0] _EVAL_230;
  wire  _EVAL_95;
  wire  _EVAL_671;
  wire  _EVAL_395;
  wire  _EVAL_312;
  wire  _EVAL_142;
  wire  _EVAL_518;
  wire [32:0] _EVAL_330;
  wire [32:0] _EVAL_491;
  wire  _EVAL_477;
  wire  _EVAL_123;
  wire  _EVAL_143;
  wire  _EVAL_313;
  wire  _EVAL_132;
  wire [2:0] _EVAL_663;
  wire  _EVAL_368;
  wire  _EVAL_300;
  wire  _EVAL_492;
  wire [31:0] _EVAL_168;
  wire  _EVAL_167;
  wire  _EVAL_190;
  wire  _EVAL_295;
  wire  _EVAL_134;
  wire  _EVAL_342;
  wire  _EVAL_191;
  wire  _EVAL_227;
  wire  _EVAL_170;
  wire  _EVAL_377;
  wire [2:0] _EVAL_117;
  wire  _EVAL_211;
  wire  _EVAL_660;
  wire  _EVAL_239;
  wire  _EVAL_306;
  wire  _EVAL_412;
  wire [31:0] _EVAL_420;
  wire [32:0] _EVAL_620;
  wire [32:0] _EVAL_135;
  wire [31:0] _EVAL_566;
  wire [32:0] _EVAL_616;
  wire [32:0] _EVAL_258;
  wire  _EVAL_593;
  wire  _EVAL_114;
  wire [32:0] _EVAL_72;
  wire [32:0] _EVAL_352;
  wire  _EVAL_261;
  wire [31:0] _EVAL_436;
  wire [32:0] _EVAL_353;
  wire [32:0] _EVAL_608;
  wire [32:0] _EVAL_390;
  wire  _EVAL_670;
  wire  _EVAL_348;
  wire [31:0] _EVAL_571;
  wire [32:0] _EVAL_58;
  wire [32:0] _EVAL_236;
  wire [32:0] _EVAL_77;
  wire  _EVAL_525;
  wire  _EVAL_169;
  wire [32:0] _EVAL_585;
  wire [32:0] _EVAL_277;
  wire [32:0] _EVAL_611;
  wire  _EVAL_440;
  wire  _EVAL_465;
  wire [31:0] _EVAL_428;
  wire [32:0] _EVAL_533;
  wire [32:0] _EVAL_122;
  wire [32:0] _EVAL_198;
  wire  _EVAL_598;
  wire  _EVAL_232;
  wire [31:0] _EVAL_85;
  wire [32:0] _EVAL_205;
  wire [32:0] _EVAL_438;
  wire [32:0] _EVAL_263;
  wire  _EVAL_504;
  wire  _EVAL_480;
  wire [31:0] _EVAL_153;
  wire [32:0] _EVAL_386;
  wire [32:0] _EVAL_521;
  wire [32:0] _EVAL_346;
  wire  _EVAL_409;
  wire [31:0] _EVAL_242;
  wire [32:0] _EVAL_38;
  wire [32:0] _EVAL_381;
  wire [32:0] _EVAL_513;
  wire  _EVAL_619;
  wire  _EVAL_208;
  wire  _EVAL_642;
  wire  _EVAL_319;
  wire  _EVAL_90;
  wire  _EVAL_345;
  wire  _EVAL_128;
  wire [31:0] _EVAL_254;
  wire [32:0] _EVAL_536;
  wire [32:0] _EVAL_520;
  wire [32:0] _EVAL_298;
  wire  _EVAL_527;
  wire  _EVAL_229;
  wire  _EVAL_638;
  wire  _EVAL_147;
  wire  _EVAL_237;
  wire [15:0] _EVAL_288;
  wire [8:0] _EVAL_481;
  wire [8:0] _EVAL_524;
  wire [8:0] _EVAL_212;
  wire  _EVAL_247;
  wire  _EVAL_383;
  wire  _EVAL_558;
  wire  _EVAL_333;
  wire  _EVAL_582;
  wire  _EVAL_493;
  wire  _EVAL_450;
  wire  _EVAL_63;
  wire  _EVAL_245;
  wire  _EVAL_656;
  wire  _EVAL_324;
  wire  _EVAL_549;
  wire  _EVAL_53;
  wire  _EVAL_165;
  wire  _EVAL_334;
  wire  _EVAL_296;
  wire  _EVAL_217;
  wire  _EVAL_375;
  wire  _EVAL_256;
  wire  _EVAL_484;
  wire  _EVAL_35;
  wire  _EVAL_98;
  wire  _EVAL_290;
  wire  _EVAL_88;
  wire  _EVAL_209;
  wire  _EVAL_363;
  wire  _EVAL_93;
  wire  _EVAL_284;
  wire  _EVAL_60;
  wire  _EVAL_609;
  wire  _EVAL_160;
  wire  _EVAL_583;
  wire  _EVAL_397;
  wire  _EVAL_422;
  wire  _EVAL_577;
  wire  _EVAL_535;
  wire  _EVAL_228;
  wire [7:0] _EVAL_216;
  wire  _EVAL_486;
  wire [31:0] _EVAL_652;
  wire [32:0] _EVAL_42;
  wire [32:0] _EVAL_574;
  wire [32:0] _EVAL_335;
  wire  _EVAL_91;
  wire [31:0] _EVAL_151;
  wire [32:0] _EVAL_271;
  wire [32:0] _EVAL_597;
  wire [32:0] _EVAL_378;
  wire  _EVAL_601;
  wire  _EVAL_538;
  wire [31:0] _EVAL_99;
  wire [32:0] _EVAL_241;
  wire [32:0] _EVAL_139;
  wire [32:0] _EVAL_512;
  wire  _EVAL_530;
  wire  _EVAL_529;
  wire [31:0] _EVAL_624;
  wire [32:0] _EVAL_305;
  wire [32:0] _EVAL_651;
  wire [32:0] _EVAL_410;
  wire  _EVAL_371;
  wire  _EVAL_78;
  wire  _EVAL_650;
  wire [32:0] _EVAL_192;
  wire [32:0] _EVAL_131;
  wire  _EVAL_373;
  wire  _EVAL_400;
  wire [32:0] _EVAL_565;
  wire  _EVAL_623;
  wire  _EVAL_489;
  wire [31:0] _EVAL_109;
  wire [32:0] _EVAL_391;
  wire [32:0] _EVAL_468;
  wire [32:0] _EVAL_157;
  wire  _EVAL_562;
  wire  _EVAL_202;
  wire [31:0] _EVAL_528;
  wire [32:0] _EVAL_627;
  wire [32:0] _EVAL_188;
  wire [32:0] _EVAL_526;
  wire  _EVAL_259;
  wire  _EVAL_637;
  wire [22:0] _EVAL_64;
  wire [7:0] _EVAL_661;
  wire [7:0] _EVAL_654;
  wire [31:0] _EVAL_49;
  wire  _EVAL_71;
  wire  _EVAL_276;
  wire  _EVAL_369;
  wire [31:0] _EVAL_411;
  wire  _EVAL_441;
  wire  _EVAL_226;
  wire [4:0] _EVAL_327;
  wire [4:0] _EVAL_653;
  wire  _EVAL_546;
  wire  _EVAL_515;
  wire  _EVAL_569;
  wire  _EVAL_201;
  wire [22:0] _EVAL_588;
  wire [7:0] _EVAL_482;
  wire [7:0] _EVAL_59;
  wire [4:0] _EVAL_200;
  wire [4:0] _EVAL_451;
  wire  _EVAL_382;
  wire [31:0] _EVAL_349;
  wire [32:0] _EVAL_459;
  wire [32:0] _EVAL_97;
  wire [32:0] _EVAL_286;
  wire [32:0] _EVAL_523;
  wire  _EVAL_622;
  wire [32:0] _EVAL_189;
  wire [32:0] _EVAL_632;
  wire [32:0] _EVAL_336;
  wire  _EVAL_243;
  wire  _EVAL_266;
  wire [31:0] _EVAL_467;
  wire [32:0] _EVAL_423;
  wire [32:0] _EVAL_602;
  wire [32:0] _EVAL_69;
  wire  _EVAL_268;
  wire  _EVAL_476;
  wire  _EVAL_444;
  wire  _EVAL_488;
  wire  _EVAL_248;
  wire  _EVAL_607;
  wire [32:0] _EVAL_70;
  wire [32:0] _EVAL_446;
  wire [32:0] _EVAL_351;
  wire  _EVAL_267;
  wire  _EVAL_129;
  wire [32:0] _EVAL_618;
  wire [32:0] _EVAL_270;
  wire  _EVAL_119;
  wire  _EVAL_197;
  wire  _EVAL_394;
  wire  _EVAL_218;
  wire  _EVAL_347;
  wire  _EVAL_615;
  wire [31:0] _EVAL_257;
  wire [32:0] _EVAL_195;
  wire [32:0] _EVAL_463;
  wire [32:0] _EVAL_174;
  wire  _EVAL_238;
  wire  _EVAL_240;
  wire  _EVAL_572;
  wire  _EVAL_556;
  wire [8:0] _EVAL_166;
  wire  _EVAL_121;
  wire  _EVAL_547;
  wire  _EVAL_399;
  wire  _EVAL_517;
  wire  _EVAL_393;
  wire  _EVAL_339;
  wire  _EVAL_502;
  wire [31:0] _EVAL_667;
  wire  _EVAL_617;
  wire  _EVAL_635;
  wire  _EVAL_291;
  wire  _EVAL_647;
  wire  _EVAL_273;
  wire  _EVAL_367;
  wire  _EVAL_272;
  wire  _EVAL_478;
  wire [15:0] _EVAL_325;
  wire [15:0] _EVAL_372;
  wire [8:0] _EVAL_299;
  wire  _EVAL_265;
  wire  _EVAL_289;
  wire  _EVAL_111;
  wire  _EVAL_460;
  wire  _EVAL_323;
  wire [1:0] _EVAL_595;
  wire [1:0] _EVAL_673;
  wire [1:0] _EVAL_457;
  wire  _EVAL_124;
  wire  _EVAL_308;
  wire  _EVAL_433;
  wire  _EVAL_118;
  wire  _EVAL_340;
  wire  _EVAL_81;
  wire  _EVAL_303;
  wire  _EVAL_606;
  wire  _EVAL_552;
  wire  _EVAL_662;
  wire  _EVAL_152;
  wire  _EVAL_294;
  wire  _EVAL_374;
  wire  _EVAL_302;
  wire  _EVAL_102;
  wire  _EVAL_251;
  wire  _EVAL_648;
  wire  _EVAL_115;
  wire  _EVAL_475;
  wire  _EVAL_292;
  wire  _EVAL_50;
  wire  _EVAL_387;
  wire  _EVAL_360;
  wire  _EVAL_207;
  wire  _EVAL_233;
  wire [1:0] _EVAL_65;
  wire  _EVAL_39;
  wire  _EVAL_483;
  wire  _EVAL_79;
  wire  _EVAL_332;
  wire  _EVAL_567;
  wire [7:0] _EVAL_494;
  wire [7:0] _EVAL_532;
  wire [4:0] _EVAL_214;
  wire  _EVAL_500;
  wire  _EVAL_84;
  wire  _EVAL_231;
  wire  _EVAL_137;
  wire  _EVAL_626;
  wire  _EVAL_534;
  wire  _EVAL_140;
  wire  _EVAL_80;
  wire  _EVAL_180;
  wire  _EVAL_220;
  wire  _EVAL_580;
  wire [22:0] _EVAL_34;
  wire  _EVAL_264;
  wire  _EVAL_495;
  wire  _EVAL_223;
  wire  _EVAL_430;
  wire  _EVAL_454;
  wire  _EVAL_92;
  wire  _EVAL_89;
  wire  _EVAL_665;
  wire  _EVAL_281;
  wire [7:0] _EVAL_631;
  wire [7:0] _EVAL_664;
  wire [31:0] _EVAL_603;
  wire [31:0] _EVAL_449;
  wire  _EVAL_636;
  wire  _EVAL_155;
  wire  _EVAL_414;
  wire  _EVAL_613;
  wire  _EVAL_474;
  wire  _EVAL_235;
  wire [4:0] _EVAL_301;
  wire  _EVAL_490;
  wire [32:0] _EVAL_76;
  wire  _EVAL_196;
  wire  _EVAL_573;
  wire [32:0] _EVAL_341;
  wire  _EVAL_234;
  wire  _EVAL_304;
  wire  _EVAL_321;
  wire  _EVAL_544;
  wire  _EVAL_634;
  wire  _EVAL_589;
  wire  _EVAL_621;
  wire  _EVAL_594;
  wire [1:0] _EVAL_519;
  wire [1:0] _EVAL_659;
  wire [1:0] _EVAL_396;
  wire [1:0] _EVAL_107;
  wire  _EVAL_269;
  wire  _EVAL_511;
  wire  _EVAL_470;
  wire  _EVAL_110;
  wire  _EVAL_178;
  wire  _EVAL_437;
  wire  _EVAL_311;
  wire  _EVAL_542;
  wire  _EVAL_96;
  wire  _EVAL_317;
  wire  _EVAL_432;
  wire  _EVAL_604;
  wire  _EVAL_408;
  wire  _EVAL_473;
  wire  _EVAL_625;
  wire  _EVAL_599;
  wire  _EVAL_581;
  wire  _EVAL_145;
  wire  _EVAL_507;
  wire  _EVAL_162;
  wire  _EVAL_388;
  wire  _EVAL_366;
  wire  _EVAL_350;
  wire  _EVAL_541;
  wire [8:0] _EVAL_56;
  wire  _EVAL_314;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_40;
  wire  _EVAL_586;
  wire  _EVAL_164;
  wire  _EVAL_179;
  wire  _EVAL_41;
  wire  _EVAL_297;
  wire  _EVAL_359;
  wire  _EVAL_668;
  wire  _EVAL_287;
  wire  _EVAL_52;
  wire  _EVAL_445;
  wire  _EVAL_329;
  wire  _EVAL_326;
  wire  _EVAL_37;
  wire  _EVAL_628;
  wire  _EVAL_357;
  wire  _EVAL_561;
  wire  _EVAL_225;
  wire  _EVAL_62;
  wire  _EVAL_285;
  wire  _EVAL_657;
  wire  _EVAL_362;
  wire  _EVAL_579;
  wire [8:0] _EVAL_54;
  wire [8:0] _EVAL_338;
  wire  _EVAL_469;
  wire  _EVAL_439;
  wire  _EVAL_537;
  wire  _EVAL_105;
  wire  _EVAL_630;
  wire  _EVAL_610;
  wire  _EVAL_74;
  wire  _EVAL_215;
  wire [1:0] _EVAL_514;
  wire [1:0] _EVAL_600;
  wire  _EVAL_204;
  wire [31:0] _EVAL_307;
  wire  _EVAL_44;
  wire  _EVAL_318;
  wire  _EVAL_646;
  wire  _EVAL_404;
  wire  _EVAL_343;
  wire  _EVAL_419;
  wire  _EVAL_45;
  wire  _EVAL_175;
  wire  _EVAL_503;
  wire  _EVAL_392;
  wire  _EVAL_101;
  wire  _EVAL_418;
  wire  _EVAL_413;
  wire  _EVAL_106;
  wire  _EVAL_427;
  wire  _EVAL_184;
  wire  _EVAL_86;
  wire  _EVAL_354;
  wire  _EVAL_564;
  wire  _EVAL_434;
  wire  _EVAL_672;
  wire  _EVAL_278;
  wire  _EVAL_148;
  wire  _EVAL_163;
  wire  _EVAL_555;
  wire  _EVAL_385;
  wire  _EVAL_553;
  wire  _EVAL_104;
  wire  _EVAL_344;
  wire  _EVAL_36;
  wire  _EVAL_510;
  wire  _EVAL_246;
  wire  _EVAL_563;
  wire  _EVAL_506;
  wire  _EVAL_260;
  wire  _EVAL_253;
  wire  _EVAL_361;
  wire  _EVAL_87;
  wire  _EVAL_472;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_43;
  wire  _EVAL_640;
  wire  _EVAL_570;
  wire  _EVAL_479;
  wire  _EVAL_275;
  wire  _EVAL_57;
  wire  _EVAL_639;
  wire  _EVAL_127;
  wire  _EVAL_575;
  wire  _EVAL_584;
  wire  _EVAL_587;
  wire  _EVAL_456;
  wire  _EVAL_509;
  wire  _EVAL_380;
  wire  _EVAL_402;
  wire  _EVAL_578;
  wire  _EVAL_370;
  wire  _EVAL_487;
  wire  _EVAL_629;
  wire  _EVAL_458;
  wire  _EVAL_199;
  wire  _EVAL_462;
  wire  _EVAL_108;
  wire  _EVAL_322;
  wire  _EVAL_144;
  wire  _EVAL_443;
  wire  _EVAL_274;
  wire [4:0] _EVAL_181;
  wire  _EVAL_376;
  wire  _EVAL_185;
  wire  _EVAL_658;
  wire  _EVAL_94;
  wire  _EVAL_206;
  wire  _EVAL_83;
  wire  _EVAL_337;
  wire  _EVAL_633;
  wire  _EVAL_158;
  wire  _EVAL_213;
  wire  _EVAL_130;
  wire  _EVAL_435;
  wire  _EVAL_485;
  wire  _EVAL_421;
  wire  _EVAL_442;
  wire  _EVAL_666;
  wire  _EVAL_431;
  wire  _EVAL_73;
  wire  _EVAL_516;
  wire  _EVAL_141;
  wire  _EVAL_455;
  wire  _EVAL_183;
  wire  _EVAL_550;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_471 = _EVAL_4 ^ 32'h1800000;
  assign _EVAL_398 = {1'b0,$signed(_EVAL_471)};
  assign _EVAL_61 = _EVAL_19 >= 4'h3;
  assign _EVAL_221 = _EVAL_19[1:0];
  assign _EVAL_522 = 4'h1 << _EVAL_221;
  assign _EVAL_551 = _EVAL_522[2:0];
  assign _EVAL_655 = _EVAL_551 | 3'h1;
  assign _EVAL_641 = _EVAL_655[2];
  assign _EVAL_194 = _EVAL_27[2];
  assign _EVAL_182 = _EVAL_194 == 1'h0;
  assign _EVAL_224 = _EVAL_641 & _EVAL_182;
  assign _EVAL_315 = _EVAL_61 | _EVAL_224;
  assign _EVAL_464 = _EVAL_655[1];
  assign _EVAL_328 = _EVAL_27[1];
  assign _EVAL_592 = _EVAL_328 == 1'h0;
  assign _EVAL_591 = _EVAL_182 & _EVAL_592;
  assign _EVAL_364 = _EVAL_464 & _EVAL_591;
  assign _EVAL_176 = _EVAL_315 | _EVAL_364;
  assign _EVAL_55 = _EVAL_655[0];
  assign _EVAL_590 = _EVAL_27[0];
  assign _EVAL_177 = _EVAL_591 & _EVAL_590;
  assign _EVAL_154 = _EVAL_55 & _EVAL_177;
  assign _EVAL_222 = _EVAL_176 | _EVAL_154;
  assign _EVAL_426 = _EVAL_12 ^ 32'h2000000;
  assign _EVAL_186 = {1'b0,$signed(_EVAL_426)};
  assign _EVAL_560 = $signed(_EVAL_186) & $signed(-33'sh10000);
  assign _EVAL_405 = $signed(_EVAL_560);
  assign _EVAL_112 = $signed(_EVAL_405) == $signed(33'sh0);
  assign _EVAL_497 = _EVAL_159 - 5'h1;
  assign _EVAL_171 = _EVAL_358 - 5'h1;
  assign _EVAL_203 = _EVAL_27 ^ 32'h3000;
  assign _EVAL_501 = {1'b0,$signed(_EVAL_203)};
  assign _EVAL_505 = _EVAL_13 == 3'h6;
  assign _EVAL_68 = _EVAL_22 >= 4'h3;
  assign _EVAL_365 = _EVAL_356 - 5'h1;
  assign _EVAL_429 = _EVAL_28 == 3'h2;
  assign _EVAL_310 = 16'h1 << _EVAL_25;
  assign _EVAL_309 = _EVAL_4 ^ 32'h2000000;
  assign _EVAL_508 = {1'b0,$signed(_EVAL_309)};
  assign _EVAL_193 = $signed(_EVAL_508) & $signed(-33'sh10000);
  assign _EVAL_498 = _EVAL_27 ^ 32'h80000000;
  assign _EVAL_466 = {1'b0,$signed(_EVAL_498)};
  assign _EVAL_452 = $signed(_EVAL_466) & $signed(-33'sh20000);
  assign _EVAL_545 = $signed(_EVAL_452);
  assign _EVAL_156 = $signed(_EVAL_545) == $signed(33'sh0);
  assign _EVAL_279 = ~ _EVAL_1;
  assign _EVAL_187 = _EVAL_279 == 8'h0;
  assign _EVAL_173 = _EVAL_15 == 4'h8;
  assign _EVAL_293 = _EVAL_15 == 4'h0;
  assign _EVAL_596 = _EVAL_173 | _EVAL_293;
  assign _EVAL_51 = _EVAL_15[3:3];
  assign _EVAL_250 = _EVAL_51 == 1'h0;
  assign _EVAL_401 = _EVAL_15[2:0];
  assign _EVAL_262 = 3'h1 <= _EVAL_401;
  assign _EVAL_66 = _EVAL_250 & _EVAL_262;
  assign _EVAL_136 = _EVAL_596 | _EVAL_66;
  assign _EVAL_605 = _EVAL_136 | _EVAL_0;
  assign _EVAL_645 = _EVAL_605 == 1'h0;
  assign _EVAL_146 = _EVAL_18 == 1'h0;
  assign _EVAL_496 = _EVAL_146 | _EVAL_0;
  assign _EVAL_103 = _EVAL_496 == 1'h0;
  assign _EVAL_403 = _EVAL_8 & _EVAL_16;
  assign _EVAL_244 = _EVAL_669 == 5'h0;
  assign _EVAL_384 = _EVAL_403 & _EVAL_244;
  assign _EVAL_406 = _EVAL_4 ^ 32'h4000;
  assign _EVAL_649 = {1'b0,$signed(_EVAL_406)};
  assign _EVAL_316 = _EVAL_4 ^ 32'h40000000;
  assign _EVAL_75 = {1'b0,$signed(_EVAL_316)};
  assign _EVAL_614 = $signed(_EVAL_75) & $signed(-33'sh2000);
  assign _EVAL_230 = $signed(_EVAL_614);
  assign _EVAL_95 = _EVAL_146 | _EVAL_33;
  assign _EVAL_671 = _EVAL_12 == _EVAL_559;
  assign _EVAL_395 = _EVAL_671 | _EVAL_0;
  assign _EVAL_312 = _EVAL_395 == 1'h0;
  assign _EVAL_142 = _EVAL_194 & _EVAL_592;
  assign _EVAL_518 = _EVAL_142 & _EVAL_590;
  assign _EVAL_330 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_491 = $signed(_EVAL_649) & $signed(-33'sh1000);
  assign _EVAL_477 = _EVAL_25 == 4'h8;
  assign _EVAL_123 = _EVAL_25 == 4'h0;
  assign _EVAL_143 = _EVAL_477 | _EVAL_123;
  assign _EVAL_313 = _EVAL_25[3:3];
  assign _EVAL_132 = _EVAL_313 == 1'h0;
  assign _EVAL_663 = _EVAL_25[2:0];
  assign _EVAL_368 = 3'h1 <= _EVAL_663;
  assign _EVAL_300 = _EVAL_132 & _EVAL_368;
  assign _EVAL_492 = _EVAL_143 | _EVAL_300;
  assign _EVAL_168 = _EVAL_4 ^ 32'h80000000;
  assign _EVAL_167 = _EVAL_31 == 2'h0;
  assign _EVAL_190 = _EVAL_167 | _EVAL_0;
  assign _EVAL_295 = _EVAL_190 == 1'h0;
  assign _EVAL_134 = _EVAL_19 <= 4'h8;
  assign _EVAL_342 = _EVAL_2 == 4'h8;
  assign _EVAL_191 = _EVAL_2 == 4'h0;
  assign _EVAL_227 = _EVAL_342 | _EVAL_191;
  assign _EVAL_170 = _EVAL_2[3:3];
  assign _EVAL_377 = _EVAL_170 == 1'h0;
  assign _EVAL_117 = _EVAL_2[2:0];
  assign _EVAL_211 = 3'h1 <= _EVAL_117;
  assign _EVAL_660 = _EVAL_377 & _EVAL_211;
  assign _EVAL_239 = _EVAL_227 | _EVAL_660;
  assign _EVAL_306 = _EVAL_239 | _EVAL_0;
  assign _EVAL_412 = _EVAL_306 == 1'h0;
  assign _EVAL_420 = _EVAL_12 ^ 32'h1800000;
  assign _EVAL_620 = {1'b0,$signed(_EVAL_420)};
  assign _EVAL_135 = $signed(_EVAL_620) & $signed(-33'sh8000);
  assign _EVAL_566 = _EVAL_4 ^ 32'h20000000;
  assign _EVAL_616 = {1'b0,$signed(_EVAL_566)};
  assign _EVAL_258 = $signed(_EVAL_616) & $signed(-33'sh2000);
  assign _EVAL_593 = _EVAL_187 | _EVAL_0;
  assign _EVAL_114 = _EVAL_593 == 1'h0;
  assign _EVAL_72 = $signed(_EVAL_501) & $signed(-33'sh1000);
  assign _EVAL_352 = $signed(_EVAL_72);
  assign _EVAL_261 = $signed(_EVAL_352) == $signed(33'sh0);
  assign _EVAL_436 = _EVAL_27 ^ 32'hc000000;
  assign _EVAL_353 = {1'b0,$signed(_EVAL_436)};
  assign _EVAL_608 = $signed(_EVAL_353) & $signed(-33'sh4000000);
  assign _EVAL_390 = $signed(_EVAL_608);
  assign _EVAL_670 = $signed(_EVAL_390) == $signed(33'sh0);
  assign _EVAL_348 = _EVAL_261 | _EVAL_670;
  assign _EVAL_571 = _EVAL_27 ^ 32'h2000000;
  assign _EVAL_58 = {1'b0,$signed(_EVAL_571)};
  assign _EVAL_236 = $signed(_EVAL_58) & $signed(-33'sh10000);
  assign _EVAL_77 = $signed(_EVAL_236);
  assign _EVAL_525 = $signed(_EVAL_77) == $signed(33'sh0);
  assign _EVAL_169 = _EVAL_348 | _EVAL_525;
  assign _EVAL_585 = {1'b0,$signed(_EVAL_27)};
  assign _EVAL_277 = $signed(_EVAL_585) & $signed(-33'sh5000);
  assign _EVAL_611 = $signed(_EVAL_277);
  assign _EVAL_440 = $signed(_EVAL_611) == $signed(33'sh0);
  assign _EVAL_465 = _EVAL_169 | _EVAL_440;
  assign _EVAL_428 = _EVAL_27 ^ 32'h1800000;
  assign _EVAL_533 = {1'b0,$signed(_EVAL_428)};
  assign _EVAL_122 = $signed(_EVAL_533) & $signed(-33'sh8000);
  assign _EVAL_198 = $signed(_EVAL_122);
  assign _EVAL_598 = $signed(_EVAL_198) == $signed(33'sh0);
  assign _EVAL_232 = _EVAL_465 | _EVAL_598;
  assign _EVAL_85 = _EVAL_27 ^ 32'h1900000;
  assign _EVAL_205 = {1'b0,$signed(_EVAL_85)};
  assign _EVAL_438 = $signed(_EVAL_205) & $signed(-33'sh2000);
  assign _EVAL_263 = $signed(_EVAL_438);
  assign _EVAL_504 = $signed(_EVAL_263) == $signed(33'sh0);
  assign _EVAL_480 = _EVAL_232 | _EVAL_504;
  assign _EVAL_153 = _EVAL_4 ^ 32'h1900000;
  assign _EVAL_386 = {1'b0,$signed(_EVAL_153)};
  assign _EVAL_521 = $signed(_EVAL_386) & $signed(-33'sh2000);
  assign _EVAL_346 = $signed(_EVAL_521);
  assign _EVAL_409 = $signed(_EVAL_346) == $signed(33'sh0);
  assign _EVAL_242 = _EVAL_27 ^ 32'h40000000;
  assign _EVAL_38 = {1'b0,$signed(_EVAL_242)};
  assign _EVAL_381 = $signed(_EVAL_38) & $signed(-33'sh2000);
  assign _EVAL_513 = $signed(_EVAL_381);
  assign _EVAL_619 = $signed(_EVAL_513) == $signed(33'sh0);
  assign _EVAL_208 = _EVAL_619 | _EVAL_156;
  assign _EVAL_642 = _EVAL_208 | _EVAL_670;
  assign _EVAL_319 = _EVAL_642 | _EVAL_525;
  assign _EVAL_90 = _EVAL_319 | _EVAL_440;
  assign _EVAL_345 = _EVAL_90 | _EVAL_598;
  assign _EVAL_128 = _EVAL_345 | _EVAL_504;
  assign _EVAL_254 = _EVAL_27 ^ 32'h20000000;
  assign _EVAL_536 = {1'b0,$signed(_EVAL_254)};
  assign _EVAL_520 = $signed(_EVAL_536) & $signed(-33'sh2000);
  assign _EVAL_298 = $signed(_EVAL_520);
  assign _EVAL_527 = $signed(_EVAL_298) == $signed(33'sh0);
  assign _EVAL_229 = _EVAL_128 | _EVAL_527;
  assign _EVAL_638 = _EVAL_23 & _EVAL_9;
  assign _EVAL_147 = _EVAL_356 == 5'h0;
  assign _EVAL_237 = _EVAL_638 & _EVAL_147;
  assign _EVAL_288 = _EVAL_237 ? _EVAL_310 : 16'h0;
  assign _EVAL_481 = _EVAL_288[8:0];
  assign _EVAL_524 = _EVAL_481 | _EVAL_100;
  assign _EVAL_212 = _EVAL_524 >> _EVAL_2;
  assign _EVAL_247 = _EVAL_212[0];
  assign _EVAL_383 = _EVAL_247 | _EVAL_0;
  assign _EVAL_558 = _EVAL_383 == 1'h0;
  assign _EVAL_333 = _EVAL_182 & _EVAL_328;
  assign _EVAL_582 = _EVAL_464 & _EVAL_333;
  assign _EVAL_493 = _EVAL_315 | _EVAL_582;
  assign _EVAL_450 = _EVAL_590 == 1'h0;
  assign _EVAL_63 = _EVAL_333 & _EVAL_450;
  assign _EVAL_245 = _EVAL_55 & _EVAL_63;
  assign _EVAL_656 = _EVAL_493 | _EVAL_245;
  assign _EVAL_324 = _EVAL_2 == _EVAL_252;
  assign _EVAL_549 = _EVAL_324 | _EVAL_0;
  assign _EVAL_53 = _EVAL_447 == 5'h0;
  assign _EVAL_165 = _EVAL_641 & _EVAL_194;
  assign _EVAL_334 = _EVAL_61 | _EVAL_165;
  assign _EVAL_296 = _EVAL_194 & _EVAL_328;
  assign _EVAL_217 = _EVAL_464 & _EVAL_296;
  assign _EVAL_375 = _EVAL_334 | _EVAL_217;
  assign _EVAL_256 = _EVAL_296 & _EVAL_590;
  assign _EVAL_484 = _EVAL_55 & _EVAL_256;
  assign _EVAL_35 = _EVAL_375 | _EVAL_484;
  assign _EVAL_98 = _EVAL_296 & _EVAL_450;
  assign _EVAL_290 = _EVAL_55 & _EVAL_98;
  assign _EVAL_88 = _EVAL_375 | _EVAL_290;
  assign _EVAL_209 = _EVAL_464 & _EVAL_142;
  assign _EVAL_363 = _EVAL_334 | _EVAL_209;
  assign _EVAL_93 = _EVAL_55 & _EVAL_518;
  assign _EVAL_284 = _EVAL_363 | _EVAL_93;
  assign _EVAL_60 = _EVAL_142 & _EVAL_450;
  assign _EVAL_609 = _EVAL_55 & _EVAL_60;
  assign _EVAL_160 = _EVAL_363 | _EVAL_609;
  assign _EVAL_583 = _EVAL_333 & _EVAL_590;
  assign _EVAL_397 = _EVAL_55 & _EVAL_583;
  assign _EVAL_422 = _EVAL_493 | _EVAL_397;
  assign _EVAL_577 = _EVAL_591 & _EVAL_450;
  assign _EVAL_535 = _EVAL_55 & _EVAL_577;
  assign _EVAL_228 = _EVAL_176 | _EVAL_535;
  assign _EVAL_216 = {_EVAL_35,_EVAL_88,_EVAL_284,_EVAL_160,_EVAL_422,_EVAL_656,_EVAL_222,_EVAL_228};
  assign _EVAL_486 = _EVAL_1 == _EVAL_216;
  assign _EVAL_652 = _EVAL_12 ^ 32'h40000000;
  assign _EVAL_42 = {1'b0,$signed(_EVAL_652)};
  assign _EVAL_574 = $signed(_EVAL_42) & $signed(-33'sh2000);
  assign _EVAL_335 = $signed(_EVAL_574);
  assign _EVAL_91 = $signed(_EVAL_335) == $signed(33'sh0);
  assign _EVAL_151 = _EVAL_12 ^ 32'h80000000;
  assign _EVAL_271 = {1'b0,$signed(_EVAL_151)};
  assign _EVAL_597 = $signed(_EVAL_271) & $signed(-33'sh20000);
  assign _EVAL_378 = $signed(_EVAL_597);
  assign _EVAL_601 = $signed(_EVAL_378) == $signed(33'sh0);
  assign _EVAL_538 = _EVAL_91 | _EVAL_601;
  assign _EVAL_99 = _EVAL_12 ^ 32'h3000;
  assign _EVAL_241 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_139 = $signed(_EVAL_241) & $signed(-33'sh1000);
  assign _EVAL_512 = $signed(_EVAL_139);
  assign _EVAL_530 = $signed(_EVAL_512) == $signed(33'sh0);
  assign _EVAL_529 = _EVAL_538 | _EVAL_530;
  assign _EVAL_624 = _EVAL_12 ^ 32'hc000000;
  assign _EVAL_305 = {1'b0,$signed(_EVAL_624)};
  assign _EVAL_651 = $signed(_EVAL_305) & $signed(-33'sh4000000);
  assign _EVAL_410 = $signed(_EVAL_651);
  assign _EVAL_371 = $signed(_EVAL_410) == $signed(33'sh0);
  assign _EVAL_78 = _EVAL_529 | _EVAL_371;
  assign _EVAL_650 = _EVAL_78 | _EVAL_112;
  assign _EVAL_192 = $signed(_EVAL_330) & $signed(-33'sh1000);
  assign _EVAL_131 = $signed(_EVAL_192);
  assign _EVAL_373 = $signed(_EVAL_131) == $signed(33'sh0);
  assign _EVAL_400 = _EVAL_650 | _EVAL_373;
  assign _EVAL_565 = $signed(_EVAL_135);
  assign _EVAL_623 = $signed(_EVAL_565) == $signed(33'sh0);
  assign _EVAL_489 = _EVAL_400 | _EVAL_623;
  assign _EVAL_109 = _EVAL_12 ^ 32'h1900000;
  assign _EVAL_391 = {1'b0,$signed(_EVAL_109)};
  assign _EVAL_468 = $signed(_EVAL_391) & $signed(-33'sh2000);
  assign _EVAL_157 = $signed(_EVAL_468);
  assign _EVAL_562 = $signed(_EVAL_157) == $signed(33'sh0);
  assign _EVAL_202 = _EVAL_489 | _EVAL_562;
  assign _EVAL_528 = _EVAL_12 ^ 32'h4000;
  assign _EVAL_627 = {1'b0,$signed(_EVAL_528)};
  assign _EVAL_188 = $signed(_EVAL_627) & $signed(-33'sh1000);
  assign _EVAL_526 = $signed(_EVAL_188);
  assign _EVAL_259 = $signed(_EVAL_526) == $signed(33'sh0);
  assign _EVAL_637 = _EVAL_202 | _EVAL_259;
  assign _EVAL_64 = 23'hff << _EVAL_26;
  assign _EVAL_661 = _EVAL_64[7:0];
  assign _EVAL_654 = ~ _EVAL_661;
  assign _EVAL_49 = {{24'd0}, _EVAL_654};
  assign _EVAL_71 = _EVAL_30 <= 2'h2;
  assign _EVAL_276 = _EVAL_71 | _EVAL_0;
  assign _EVAL_369 = _EVAL_134 & _EVAL_261;
  assign _EVAL_411 = _EVAL_12 & _EVAL_49;
  assign _EVAL_441 = _EVAL_411 == 32'h0;
  assign _EVAL_226 = _EVAL_13[0];
  assign _EVAL_327 = _EVAL_654[7:3];
  assign _EVAL_653 = _EVAL_669 - 5'h1;
  assign _EVAL_546 = _EVAL_11 != 3'h0;
  assign _EVAL_515 = _EVAL_546 | _EVAL_0;
  assign _EVAL_569 = _EVAL_3 & _EVAL_6;
  assign _EVAL_201 = _EVAL_28[0];
  assign _EVAL_588 = 23'hff << _EVAL_22;
  assign _EVAL_482 = _EVAL_588[7:0];
  assign _EVAL_59 = ~ _EVAL_482;
  assign _EVAL_200 = _EVAL_59[7:3];
  assign _EVAL_451 = _EVAL_447 - 5'h1;
  assign _EVAL_382 = _EVAL_29 == 1'h0;
  assign _EVAL_349 = _EVAL_4 ^ 32'hc000000;
  assign _EVAL_459 = {1'b0,$signed(_EVAL_349)};
  assign _EVAL_97 = $signed(_EVAL_459) & $signed(-33'sh4000000);
  assign _EVAL_286 = $signed(_EVAL_97);
  assign _EVAL_523 = $signed(_EVAL_193);
  assign _EVAL_622 = $signed(_EVAL_230) == $signed(33'sh0);
  assign _EVAL_189 = {1'b0,$signed(_EVAL_168)};
  assign _EVAL_632 = $signed(_EVAL_189) & $signed(-33'sh20000);
  assign _EVAL_336 = $signed(_EVAL_632);
  assign _EVAL_243 = $signed(_EVAL_336) == $signed(33'sh0);
  assign _EVAL_266 = _EVAL_622 | _EVAL_243;
  assign _EVAL_467 = _EVAL_4 ^ 32'h3000;
  assign _EVAL_423 = {1'b0,$signed(_EVAL_467)};
  assign _EVAL_602 = $signed(_EVAL_423) & $signed(-33'sh1000);
  assign _EVAL_69 = $signed(_EVAL_602);
  assign _EVAL_268 = $signed(_EVAL_69) == $signed(33'sh0);
  assign _EVAL_476 = _EVAL_266 | _EVAL_268;
  assign _EVAL_444 = $signed(_EVAL_286) == $signed(33'sh0);
  assign _EVAL_488 = _EVAL_476 | _EVAL_444;
  assign _EVAL_248 = $signed(_EVAL_523) == $signed(33'sh0);
  assign _EVAL_607 = _EVAL_488 | _EVAL_248;
  assign _EVAL_70 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_446 = $signed(_EVAL_70) & $signed(-33'sh1000);
  assign _EVAL_351 = $signed(_EVAL_446);
  assign _EVAL_267 = $signed(_EVAL_351) == $signed(33'sh0);
  assign _EVAL_129 = _EVAL_607 | _EVAL_267;
  assign _EVAL_618 = $signed(_EVAL_398) & $signed(-33'sh8000);
  assign _EVAL_270 = $signed(_EVAL_618);
  assign _EVAL_119 = $signed(_EVAL_270) == $signed(33'sh0);
  assign _EVAL_197 = _EVAL_129 | _EVAL_119;
  assign _EVAL_394 = _EVAL_159 == 5'h0;
  assign _EVAL_218 = _EVAL_394 == 1'h0;
  assign _EVAL_347 = _EVAL_6 & _EVAL_218;
  assign _EVAL_615 = _EVAL_481 != 9'h0;
  assign _EVAL_257 = _EVAL_12 ^ 32'h20000000;
  assign _EVAL_195 = {1'b0,$signed(_EVAL_257)};
  assign _EVAL_463 = $signed(_EVAL_195) & $signed(-33'sh2000);
  assign _EVAL_174 = $signed(_EVAL_463);
  assign _EVAL_238 = $signed(_EVAL_174) == $signed(33'sh0);
  assign _EVAL_240 = _EVAL_637 | _EVAL_238;
  assign _EVAL_572 = _EVAL_240 | _EVAL_0;
  assign _EVAL_556 = _EVAL_572 == 1'h0;
  assign _EVAL_166 = _EVAL_100 >> _EVAL_25;
  assign _EVAL_121 = _EVAL_26 <= 4'h6;
  assign _EVAL_547 = _EVAL_19 <= 4'h6;
  assign _EVAL_399 = _EVAL_547 & _EVAL_229;
  assign _EVAL_517 = _EVAL_399 | _EVAL_369;
  assign _EVAL_393 = _EVAL_517 | _EVAL_0;
  assign _EVAL_339 = _EVAL_393 == 1'h0;
  assign _EVAL_502 = _EVAL_11 <= 3'h4;
  assign _EVAL_667 = _EVAL_149 + 32'h1;
  assign _EVAL_617 = _EVAL_25 == _EVAL_568;
  assign _EVAL_635 = _EVAL_617 | _EVAL_0;
  assign _EVAL_291 = _EVAL_635 == 1'h0;
  assign _EVAL_647 = _EVAL_120 == 5'h0;
  assign _EVAL_273 = _EVAL_569 & _EVAL_647;
  assign _EVAL_367 = _EVAL_28 == 3'h6;
  assign _EVAL_272 = _EVAL_367 == 1'h0;
  assign _EVAL_478 = _EVAL_273 & _EVAL_272;
  assign _EVAL_325 = 16'h1 << _EVAL_2;
  assign _EVAL_372 = _EVAL_478 ? _EVAL_325 : 16'h0;
  assign _EVAL_299 = _EVAL_372[8:0];
  assign _EVAL_265 = _EVAL_481 != _EVAL_299;
  assign _EVAL_289 = _EVAL_615 == 1'h0;
  assign _EVAL_111 = _EVAL_265 | _EVAL_289;
  assign _EVAL_460 = _EVAL_111 | _EVAL_0;
  assign _EVAL_323 = _EVAL_21 & _EVAL_7;
  assign _EVAL_595 = 2'h1 << _EVAL_24;
  assign _EVAL_673 = _EVAL_323 ? _EVAL_595 : 2'h0;
  assign _EVAL_457 = ~ _EVAL_673;
  assign _EVAL_124 = plusarg_reader_out == 32'h0;
  assign _EVAL_308 = _EVAL_28[1];
  assign _EVAL_433 = _EVAL_308 == 1'h0;
  assign _EVAL_118 = _EVAL_121 & _EVAL_601;
  assign _EVAL_340 = _EVAL_33 == 1'h0;
  assign _EVAL_81 = _EVAL_340 | _EVAL_0;
  assign _EVAL_303 = _EVAL_81 == 1'h0;
  assign _EVAL_606 = _EVAL_32 == _EVAL_219;
  assign _EVAL_552 = _EVAL_606 | _EVAL_0;
  assign _EVAL_662 = _EVAL_26 == _EVAL_113;
  assign _EVAL_152 = _EVAL_662 | _EVAL_0;
  assign _EVAL_294 = _EVAL_32 <= 3'h5;
  assign _EVAL_374 = _EVAL_294 | _EVAL_0;
  assign _EVAL_302 = _EVAL_374 == 1'h0;
  assign _EVAL_102 = _EVAL_10 == _EVAL_255;
  assign _EVAL_251 = _EVAL_102 | _EVAL_0;
  assign _EVAL_648 = _EVAL_251 == 1'h0;
  assign _EVAL_115 = _EVAL_10 == 3'h0;
  assign _EVAL_475 = _EVAL_9 & _EVAL_115;
  assign _EVAL_292 = _EVAL_10 == 3'h3;
  assign _EVAL_50 = _EVAL_9 & _EVAL_292;
  assign _EVAL_387 = _EVAL_547 & _EVAL_156;
  assign _EVAL_360 = _EVAL_387 | _EVAL_0;
  assign _EVAL_207 = _EVAL_360 == 1'h0;
  assign _EVAL_233 = _EVAL_14 == 1'h0;
  assign _EVAL_65 = _EVAL_280 >> _EVAL;
  assign _EVAL_39 = _EVAL_65[0];
  assign _EVAL_483 = _EVAL_39 == 1'h0;
  assign _EVAL_79 = _EVAL_483 | _EVAL_0;
  assign _EVAL_332 = _EVAL_79 == 1'h0;
  assign _EVAL_567 = _EVAL_28 == 3'h4;
  assign _EVAL_494 = ~ _EVAL_216;
  assign _EVAL_532 = _EVAL_1 & _EVAL_494;
  assign _EVAL_214 = _EVAL_120 - 5'h1;
  assign _EVAL_500 = _EVAL_32 == 3'h0;
  assign _EVAL_84 = _EVAL_500 | _EVAL_0;
  assign _EVAL_231 = _EVAL_84 == 1'h0;
  assign _EVAL_137 = _EVAL_369 | _EVAL_0;
  assign _EVAL_626 = 4'h6 == _EVAL_26;
  assign _EVAL_534 = _EVAL_11 == 3'h0;
  assign _EVAL_140 = _EVAL_534 | _EVAL_0;
  assign _EVAL_80 = _EVAL_140 == 1'h0;
  assign _EVAL_180 = _EVAL_13 == 3'h1;
  assign _EVAL_220 = _EVAL_358 == 5'h0;
  assign _EVAL_580 = _EVAL_220 == 1'h0;
  assign _EVAL_34 = 23'hff << _EVAL_19;
  assign _EVAL_264 = _EVAL_28 == 3'h1;
  assign _EVAL_495 = _EVAL_6 & _EVAL_264;
  assign _EVAL_223 = _EVAL_30 == _EVAL_540;
  assign _EVAL_430 = _EVAL_11 <= 3'h3;
  assign _EVAL_454 = _EVAL_430 | _EVAL_0;
  assign _EVAL_92 = _EVAL_454 == 1'h0;
  assign _EVAL_89 = 4'h6 == _EVAL_19;
  assign _EVAL_665 = _EVAL_123 ? _EVAL_89 : 1'h0;
  assign _EVAL_281 = _EVAL_665 | _EVAL_0;
  assign _EVAL_631 = _EVAL_34[7:0];
  assign _EVAL_664 = ~ _EVAL_631;
  assign _EVAL_603 = {{24'd0}, _EVAL_664};
  assign _EVAL_449 = _EVAL_27 & _EVAL_603;
  assign _EVAL_636 = _EVAL_449 == 32'h0;
  assign _EVAL_155 = _EVAL_10 == 3'h7;
  assign _EVAL_414 = _EVAL_13 == 3'h7;
  assign _EVAL_613 = _EVAL_16 & _EVAL_414;
  assign _EVAL_474 = _EVAL_10[2];
  assign _EVAL_235 = _EVAL_474 == 1'h0;
  assign _EVAL_301 = _EVAL_664[7:3];
  assign _EVAL_490 = _EVAL_197 | _EVAL_409;
  assign _EVAL_76 = $signed(_EVAL_491);
  assign _EVAL_196 = $signed(_EVAL_76) == $signed(33'sh0);
  assign _EVAL_573 = _EVAL_490 | _EVAL_196;
  assign _EVAL_341 = $signed(_EVAL_258);
  assign _EVAL_234 = $signed(_EVAL_341) == $signed(33'sh0);
  assign _EVAL_304 = _EVAL_573 | _EVAL_234;
  assign _EVAL_321 = _EVAL_304 | _EVAL_0;
  assign _EVAL_544 = _EVAL_321 == 1'h0;
  assign _EVAL_634 = _EVAL_569 & _EVAL_53;
  assign _EVAL_589 = _EVAL_28[2];
  assign _EVAL_621 = _EVAL_589 & _EVAL_433;
  assign _EVAL_594 = _EVAL_634 & _EVAL_621;
  assign _EVAL_519 = 2'h1 << _EVAL;
  assign _EVAL_659 = _EVAL_594 ? _EVAL_519 : 2'h0;
  assign _EVAL_396 = _EVAL_659 | _EVAL_280;
  assign _EVAL_107 = _EVAL_396 >> _EVAL_24;
  assign _EVAL_269 = _EVAL_107[0];
  assign _EVAL_511 = _EVAL_269 | _EVAL_0;
  assign _EVAL_470 = _EVAL_511 == 1'h0;
  assign _EVAL_110 = _EVAL_10 == 3'h6;
  assign _EVAL_178 = _EVAL_4 == _EVAL_82;
  assign _EVAL_437 = _EVAL_178 | _EVAL_0;
  assign _EVAL_311 = _EVAL_437 == 1'h0;
  assign _EVAL_542 = _EVAL_26 >= 4'h3;
  assign _EVAL_96 = _EVAL_13 == 3'h4;
  assign _EVAL_317 = _EVAL_492 | _EVAL_0;
  assign _EVAL_432 = _EVAL_233 | _EVAL_0;
  assign _EVAL_604 = _EVAL_19 <= 4'h2;
  assign _EVAL_408 = _EVAL_480 | _EVAL_527;
  assign _EVAL_473 = _EVAL_604 & _EVAL_408;
  assign _EVAL_625 = _EVAL_100 != 9'h0;
  assign _EVAL_599 = _EVAL_625 == 1'h0;
  assign _EVAL_581 = _EVAL_599 | _EVAL_124;
  assign _EVAL_145 = _EVAL_149 < plusarg_reader_out;
  assign _EVAL_507 = _EVAL_581 | _EVAL_145;
  assign _EVAL_162 = _EVAL_507 | _EVAL_0;
  assign _EVAL_388 = _EVAL_162 == 1'h0;
  assign _EVAL_366 = _EVAL_15 == _EVAL_417;
  assign _EVAL_350 = _EVAL_366 | _EVAL_0;
  assign _EVAL_541 = _EVAL_350 == 1'h0;
  assign _EVAL_56 = ~ _EVAL_299;
  assign _EVAL_314 = _EVAL_382 | _EVAL_0;
  assign _EVAL_282 = _EVAL_314 == 1'h0;
  assign _EVAL_283 = _EVAL_31 != 2'h2;
  assign _EVAL_40 = _EVAL_283 | _EVAL_0;
  assign _EVAL_586 = _EVAL_18 == _EVAL_150;
  assign _EVAL_164 = _EVAL_586 | _EVAL_0;
  assign _EVAL_179 = _EVAL_28 == _EVAL_138;
  assign _EVAL_41 = _EVAL_179 | _EVAL_0;
  assign _EVAL_297 = _EVAL_638 | _EVAL_569;
  assign _EVAL_359 = _EVAL_486 | _EVAL_0;
  assign _EVAL_668 = _EVAL_32 <= 3'h2;
  assign _EVAL_287 = _EVAL_668 | _EVAL_0;
  assign _EVAL_52 = _EVAL_287 == 1'h0;
  assign _EVAL_445 = _EVAL_19 == _EVAL_543;
  assign _EVAL_329 = _EVAL_445 | _EVAL_0;
  assign _EVAL_326 = _EVAL_28 <= 3'h6;
  assign _EVAL_37 = _EVAL_326 | _EVAL_0;
  assign _EVAL_628 = _EVAL_133 == 5'h0;
  assign _EVAL_357 = _EVAL_569 & _EVAL_394;
  assign _EVAL_561 = _EVAL_10 == 3'h1;
  assign _EVAL_225 = _EVAL_9 & _EVAL_561;
  assign _EVAL_62 = _EVAL_628 == 1'h0;
  assign _EVAL_285 = _EVAL_11 == _EVAL_424;
  assign _EVAL_657 = _EVAL_285 | _EVAL_0;
  assign _EVAL_362 = _EVAL_657 == 1'h0;
  assign _EVAL_579 = _EVAL_460 == 1'h0;
  assign _EVAL_54 = _EVAL_100 | _EVAL_481;
  assign _EVAL_338 = _EVAL_54 & _EVAL_56;
  assign _EVAL_469 = _EVAL_61 | _EVAL_0;
  assign _EVAL_439 = _EVAL_10 == 3'h2;
  assign _EVAL_537 = _EVAL_166[0];
  assign _EVAL_105 = _EVAL_31 <= 2'h2;
  assign _EVAL_630 = _EVAL_9 & _EVAL_62;
  assign _EVAL_610 = _EVAL_137 == 1'h0;
  assign _EVAL_74 = _EVAL_13 == 3'h5;
  assign _EVAL_215 = _EVAL_37 == 1'h0;
  assign _EVAL_514 = _EVAL_280 | _EVAL_659;
  assign _EVAL_600 = _EVAL_514 & _EVAL_457;
  assign _EVAL_204 = _EVAL_41 == 1'h0;
  assign _EVAL_307 = _EVAL_4 & 32'h3f;
  assign _EVAL_44 = _EVAL_307 == 32'h0;
  assign _EVAL_318 = _EVAL_636 | _EVAL_0;
  assign _EVAL_646 = _EVAL_9 & _EVAL_439;
  assign _EVAL_404 = _EVAL_6 & _EVAL_567;
  assign _EVAL_343 = _EVAL == _EVAL_425;
  assign _EVAL_419 = _EVAL_343 | _EVAL_0;
  assign _EVAL_45 = _EVAL_419 == 1'h0;
  assign _EVAL_175 = _EVAL_20 & _EVAL_580;
  assign _EVAL_503 = _EVAL_28 == 3'h0;
  assign _EVAL_392 = _EVAL_10 == 3'h4;
  assign _EVAL_101 = _EVAL_9 & _EVAL_392;
  assign _EVAL_418 = _EVAL_13 == 3'h0;
  assign _EVAL_413 = _EVAL_16 & _EVAL_418;
  assign _EVAL_106 = _EVAL_244 == 1'h0;
  assign _EVAL_427 = _EVAL_16 & _EVAL_106;
  assign _EVAL_184 = _EVAL_542 | _EVAL_0;
  assign _EVAL_86 = _EVAL_184 == 1'h0;
  assign _EVAL_354 = _EVAL_13 == 3'h2;
  assign _EVAL_564 = _EVAL_44 | _EVAL_0;
  assign _EVAL_434 = _EVAL_564 == 1'h0;
  assign _EVAL_672 = _EVAL_16 & _EVAL_354;
  assign _EVAL_278 = _EVAL_105 | _EVAL_0;
  assign _EVAL_148 = _EVAL_16 & _EVAL_180;
  assign _EVAL_163 = _EVAL_473 | _EVAL_0;
  assign _EVAL_555 = _EVAL_163 == 1'h0;
  assign _EVAL_385 = _EVAL_223 | _EVAL_0;
  assign _EVAL_553 = _EVAL_13 == _EVAL_415;
  assign _EVAL_104 = _EVAL_553 | _EVAL_0;
  assign _EVAL_344 = _EVAL_441 | _EVAL_0;
  assign _EVAL_36 = _EVAL_344 == 1'h0;
  assign _EVAL_510 = _EVAL_281 == 1'h0;
  assign _EVAL_246 = _EVAL_276 == 1'h0;
  assign _EVAL_563 = _EVAL_532 == 8'h0;
  assign _EVAL_506 = _EVAL_563 | _EVAL_0;
  assign _EVAL_260 = _EVAL_506 == 1'h0;
  assign _EVAL_253 = _EVAL_502 | _EVAL_0;
  assign _EVAL_361 = _EVAL_253 == 1'h0;
  assign _EVAL_87 = _EVAL_9 & _EVAL_110;
  assign _EVAL_472 = _EVAL_95 | _EVAL_0;
  assign _EVAL_125 = _EVAL_472 == 1'h0;
  assign _EVAL_126 = _EVAL_27 == _EVAL_407;
  assign _EVAL_43 = _EVAL_515 == 1'h0;
  assign _EVAL_640 = _EVAL_11 <= 3'h2;
  assign _EVAL_570 = _EVAL_640 | _EVAL_0;
  assign _EVAL_479 = _EVAL_570 == 1'h0;
  assign _EVAL_275 = _EVAL_28 == 3'h5;
  assign _EVAL_57 = _EVAL_278 == 1'h0;
  assign _EVAL_639 = _EVAL_9 & _EVAL_155;
  assign _EVAL_127 = _EVAL_104 == 1'h0;
  assign _EVAL_575 = _EVAL_16 & _EVAL_96;
  assign _EVAL_584 = _EVAL_6 & _EVAL_367;
  assign _EVAL_587 = _EVAL_16 & _EVAL_505;
  assign _EVAL_456 = _EVAL_164 == 1'h0;
  assign _EVAL_509 = _EVAL_17 & _EVAL_20;
  assign _EVAL_380 = _EVAL_509 & _EVAL_220;
  assign _EVAL_402 = _EVAL_552 == 1'h0;
  assign _EVAL_578 = _EVAL_359 == 1'h0;
  assign _EVAL_370 = _EVAL_16 & _EVAL_74;
  assign _EVAL_487 = _EVAL_469 == 1'h0;
  assign _EVAL_629 = _EVAL_22 == _EVAL_499;
  assign _EVAL_458 = _EVAL_118 | _EVAL_0;
  assign _EVAL_199 = _EVAL_68 | _EVAL_0;
  assign _EVAL_462 = _EVAL_199 == 1'h0;
  assign _EVAL_108 = _EVAL_537 == 1'h0;
  assign _EVAL_322 = _EVAL_108 | _EVAL_0;
  assign _EVAL_144 = _EVAL_31 == _EVAL_548;
  assign _EVAL_443 = _EVAL_6 & _EVAL_503;
  assign _EVAL_274 = _EVAL_10 == 3'h5;
  assign _EVAL_181 = _EVAL_133 - 5'h1;
  assign _EVAL_376 = _EVAL_638 & _EVAL_628;
  assign _EVAL_185 = _EVAL_322 == 1'h0;
  assign _EVAL_658 = _EVAL_329 == 1'h0;
  assign _EVAL_94 = _EVAL_293 ? _EVAL_626 : 1'h0;
  assign _EVAL_206 = _EVAL_94 | _EVAL_0;
  assign _EVAL_83 = _EVAL_9 & _EVAL_274;
  assign _EVAL_337 = _EVAL_629 | _EVAL_0;
  assign _EVAL_633 = _EVAL_337 == 1'h0;
  assign _EVAL_158 = _EVAL_6 & _EVAL_275;
  assign _EVAL_213 = _EVAL_458 == 1'h0;
  assign _EVAL_130 = _EVAL_40 == 1'h0;
  assign _EVAL_435 = _EVAL_152 == 1'h0;
  assign _EVAL_485 = _EVAL_432 == 1'h0;
  assign _EVAL_421 = _EVAL_144 | _EVAL_0;
  assign _EVAL_442 = _EVAL_421 == 1'h0;
  assign _EVAL_666 = _EVAL_206 == 1'h0;
  assign _EVAL_431 = _EVAL_549 == 1'h0;
  assign _EVAL_73 = _EVAL_318 == 1'h0;
  assign _EVAL_516 = _EVAL_6 & _EVAL_429;
  assign _EVAL_141 = _EVAL_126 | _EVAL_0;
  assign _EVAL_455 = _EVAL_385 == 1'h0;
  assign _EVAL_183 = _EVAL_317 == 1'h0;
  assign _EVAL_550 = _EVAL_141 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_82 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_100 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_113 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_120 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_133 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_138 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_149 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_150 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_159 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_219 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_252 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_255 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_280 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_356 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_358 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_407 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_415 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_417 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_424 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_425 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_447 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_499 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_540 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_543 = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_548 = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_559 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_568 = _RAND_26[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_669 = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_5) begin
    if (_EVAL_380) begin
      _EVAL_82 <= _EVAL_4;
    end
    if (_EVAL_0) begin
      _EVAL_100 <= 9'h0;
    end else begin
      _EVAL_100 <= _EVAL_338;
    end
    if (_EVAL_384) begin
      _EVAL_113 <= _EVAL_26;
    end
    if (_EVAL_0) begin
      _EVAL_120 <= 5'h0;
    end else begin
      if (_EVAL_569) begin
        if (_EVAL_647) begin
          if (_EVAL_201) begin
            _EVAL_120 <= _EVAL_200;
          end else begin
            _EVAL_120 <= 5'h0;
          end
        end else begin
          _EVAL_120 <= _EVAL_214;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_133 <= 5'h0;
    end else begin
      if (_EVAL_638) begin
        if (_EVAL_628) begin
          if (_EVAL_235) begin
            _EVAL_133 <= _EVAL_301;
          end else begin
            _EVAL_133 <= 5'h0;
          end
        end else begin
          _EVAL_133 <= _EVAL_181;
        end
      end
    end
    if (_EVAL_357) begin
      _EVAL_138 <= _EVAL_28;
    end
    if (_EVAL_0) begin
      _EVAL_149 <= 32'h0;
    end else begin
      if (_EVAL_297) begin
        _EVAL_149 <= 32'h0;
      end else begin
        _EVAL_149 <= _EVAL_667;
      end
    end
    if (_EVAL_357) begin
      _EVAL_150 <= _EVAL_18;
    end
    if (_EVAL_0) begin
      _EVAL_159 <= 5'h0;
    end else begin
      if (_EVAL_569) begin
        if (_EVAL_394) begin
          if (_EVAL_201) begin
            _EVAL_159 <= _EVAL_200;
          end else begin
            _EVAL_159 <= 5'h0;
          end
        end else begin
          _EVAL_159 <= _EVAL_497;
        end
      end
    end
    if (_EVAL_384) begin
      _EVAL_219 <= _EVAL_32;
    end
    if (_EVAL_357) begin
      _EVAL_252 <= _EVAL_2;
    end
    if (_EVAL_376) begin
      _EVAL_255 <= _EVAL_10;
    end
    if (_EVAL_0) begin
      _EVAL_280 <= 2'h0;
    end else begin
      _EVAL_280 <= _EVAL_600;
    end
    if (_EVAL_0) begin
      _EVAL_356 <= 5'h0;
    end else begin
      if (_EVAL_638) begin
        if (_EVAL_147) begin
          if (_EVAL_235) begin
            _EVAL_356 <= _EVAL_301;
          end else begin
            _EVAL_356 <= 5'h0;
          end
        end else begin
          _EVAL_356 <= _EVAL_365;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_358 <= 5'h0;
    end else begin
      if (_EVAL_509) begin
        if (_EVAL_220) begin
          _EVAL_358 <= 5'h0;
        end else begin
          _EVAL_358 <= _EVAL_171;
        end
      end
    end
    if (_EVAL_376) begin
      _EVAL_407 <= _EVAL_27;
    end
    if (_EVAL_384) begin
      _EVAL_415 <= _EVAL_13;
    end
    if (_EVAL_384) begin
      _EVAL_417 <= _EVAL_15;
    end
    if (_EVAL_376) begin
      _EVAL_424 <= _EVAL_11;
    end
    if (_EVAL_357) begin
      _EVAL_425 <= _EVAL;
    end
    if (_EVAL_0) begin
      _EVAL_447 <= 5'h0;
    end else begin
      if (_EVAL_569) begin
        if (_EVAL_53) begin
          if (_EVAL_201) begin
            _EVAL_447 <= _EVAL_200;
          end else begin
            _EVAL_447 <= 5'h0;
          end
        end else begin
          _EVAL_447 <= _EVAL_451;
        end
      end
    end
    if (_EVAL_357) begin
      _EVAL_499 <= _EVAL_22;
    end
    if (_EVAL_380) begin
      _EVAL_540 <= _EVAL_30;
    end
    if (_EVAL_376) begin
      _EVAL_543 <= _EVAL_19;
    end
    if (_EVAL_357) begin
      _EVAL_548 <= _EVAL_31;
    end
    if (_EVAL_384) begin
      _EVAL_559 <= _EVAL_12;
    end
    if (_EVAL_376) begin
      _EVAL_568 <= _EVAL_25;
    end
    if (_EVAL_0) begin
      _EVAL_669 <= 5'h0;
    end else begin
      if (_EVAL_403) begin
        if (_EVAL_244) begin
          if (_EVAL_226) begin
            _EVAL_669 <= _EVAL_327;
          end else begin
            _EVAL_669 <= 5'h0;
          end
        end else begin
          _EVAL_669 <= _EVAL_653;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_339) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24fe7ed9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_362) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(444051bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac61cc6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_478 & _EVAL_558) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_442) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2e9c7c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_339) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e834f2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(405e6fb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_402) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbccbc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(195b7ac2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_455) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(146ba626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ced1fa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_658) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_339) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928d024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a15a80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_578) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48d7420a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b9c5f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_479) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e02c24bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_435) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aedddd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_578) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a81fefb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_361) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_658) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e96267a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1adbf9de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcfd84c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea8fab60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_556) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c72ee8b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28fe7378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_479) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7beeaa5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(680cb602)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dc5495e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(921c1a16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75ee1b5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(213b834)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ed2bec5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a152b2c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34612e40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a7f4e00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf1bfb86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4663c30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6584e4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_442) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_434) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_556) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(939d64a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(955b0f2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(808746ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99f6a1c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f634ed72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13fa2aa8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854b5891)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1efbcb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55215411)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_556) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35ce3af6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_578) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2791f49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_362) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f1044b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cffcb94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f183ef82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89f2e6ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_633) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e3c617)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_388) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_541) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_339) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_435) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b5c82bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_579) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8734fbf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_578) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f5cb9f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_479) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c32862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd95fa21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cb8d297)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_510) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7748964)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3541aec6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_578) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_456) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1908618e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_648) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffbdc7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ebfd396)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36298647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_578) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3265bb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87427352)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff901680)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14e42990)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2336159b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_648) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f4992c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72d6e09a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b72a609)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(597f93ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ab6c6dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_578) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_470) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3aa3140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5827064a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(786276a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_594 & _EVAL_332) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(134998f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_339) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_579) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddcb1875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_510) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ceb482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11763208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_555) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e63b8f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_544) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4396d765)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70fae002)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caac4887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_434) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c959823)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_666) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cb63e31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_610) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7221690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_402) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_431) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9aee1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_541) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a9816bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f2f14e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5d0536e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c13124d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_556) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_412) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d1429)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_479) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_594 & _EVAL_332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(437d1942)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62f2a2a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_633) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_578) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33ee2561)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_555) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4bd3515)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_388) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c7da787)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_550) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eded9b56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bed3cc09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_555) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbb7436a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_666) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ef4a27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39c9b7dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f18aa5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_556) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(135f2920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb0e1834)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e63b2749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db474912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_578) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d75903e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ddd91e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc7a9af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_487) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ac1fc45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_544) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d01e617d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_556) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9a53be8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_361) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4c1d025)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7743c8cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35334d6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89a7ad9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29b65a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a6a9692)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_487) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb7ee4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c47485f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a740b84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cc2d6a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b67c6469)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_478 & _EVAL_558) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d804c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_555) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e30a9f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51904667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_455) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2cd9b46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(478c34e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bcc4b8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_431) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_339) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7480f1b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_578) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37bb0e72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397ba601)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_610) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(242fc5c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_645) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b44c6d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_495 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_456) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854e1c0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_550) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_516 & _EVAL_412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
