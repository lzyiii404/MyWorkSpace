//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module AXI4Shuffler_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [30:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [30:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits;
  wire [31:0] plusarg_reader_out;
  wire  MaxPeriodFibonacciLFSR__EVAL;
  wire  MaxPeriodFibonacciLFSR__EVAL_0;
  wire  MaxPeriodFibonacciLFSR__EVAL_1;
  wire  MaxPeriodFibonacciLFSR__EVAL_2;
  wire  MaxPeriodFibonacciLFSR__EVAL_3;
  wire  MaxPeriodFibonacciLFSR__EVAL_4;
  wire  MaxPeriodFibonacciLFSR__EVAL_5;
  wire  MaxPeriodFibonacciLFSR__EVAL_6;
  wire  MaxPeriodFibonacciLFSR__EVAL_7;
  wire  MaxPeriodFibonacciLFSR__EVAL_8;
  wire  MaxPeriodFibonacciLFSR__EVAL_9;
  wire  MaxPeriodFibonacciLFSR__EVAL_10;
  wire  MaxPeriodFibonacciLFSR__EVAL_11;
  wire  MaxPeriodFibonacciLFSR__EVAL_12;
  wire  MaxPeriodFibonacciLFSR__EVAL_13;
  wire  MaxPeriodFibonacciLFSR__EVAL_14;
  wire  MaxPeriodFibonacciLFSR__EVAL_15;
  wire  MaxPeriodFibonacciLFSR__EVAL_16;
  wire  MaxPeriodFibonacciLFSR__EVAL_17;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [3:0] Queue_1_io_enq_bits_data_id;
  wire [30:0] Queue_1_io_enq_bits_data_addr;
  wire [7:0] Queue_1_io_enq_bits_data_len;
  wire [2:0] Queue_1_io_enq_bits_data_size;
  wire [1:0] Queue_1_io_enq_bits_data_burst;
  wire  Queue_1_io_enq_bits_data_lock;
  wire [3:0] Queue_1_io_enq_bits_data_cache;
  wire [2:0] Queue_1_io_enq_bits_data_prot;
  wire [3:0] Queue_1_io_enq_bits_data_qos;
  wire [31:0] Queue_1_io_enq_bits_timestamp;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [3:0] Queue_1_io_deq_bits_data_id;
  wire [30:0] Queue_1_io_deq_bits_data_addr;
  wire [7:0] Queue_1_io_deq_bits_data_len;
  wire [2:0] Queue_1_io_deq_bits_data_size;
  wire [1:0] Queue_1_io_deq_bits_data_burst;
  wire  Queue_1_io_deq_bits_data_lock;
  wire [3:0] Queue_1_io_deq_bits_data_cache;
  wire [2:0] Queue_1_io_deq_bits_data_prot;
  wire [3:0] Queue_1_io_deq_bits_data_qos;
  wire [31:0] Queue_1_io_deq_bits_timestamp;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_data_id;
  wire [30:0] Queue_2_io_enq_bits_data_addr;
  wire [7:0] Queue_2_io_enq_bits_data_len;
  wire [2:0] Queue_2_io_enq_bits_data_size;
  wire [1:0] Queue_2_io_enq_bits_data_burst;
  wire  Queue_2_io_enq_bits_data_lock;
  wire [3:0] Queue_2_io_enq_bits_data_cache;
  wire [2:0] Queue_2_io_enq_bits_data_prot;
  wire [3:0] Queue_2_io_enq_bits_data_qos;
  wire [31:0] Queue_2_io_enq_bits_timestamp;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_data_id;
  wire [30:0] Queue_2_io_deq_bits_data_addr;
  wire [7:0] Queue_2_io_deq_bits_data_len;
  wire [2:0] Queue_2_io_deq_bits_data_size;
  wire [1:0] Queue_2_io_deq_bits_data_burst;
  wire  Queue_2_io_deq_bits_data_lock;
  wire [3:0] Queue_2_io_deq_bits_data_cache;
  wire [2:0] Queue_2_io_deq_bits_data_prot;
  wire [3:0] Queue_2_io_deq_bits_data_qos;
  wire [31:0] Queue_2_io_deq_bits_timestamp;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_data_id;
  wire [30:0] Queue_3_io_enq_bits_data_addr;
  wire [7:0] Queue_3_io_enq_bits_data_len;
  wire [2:0] Queue_3_io_enq_bits_data_size;
  wire [1:0] Queue_3_io_enq_bits_data_burst;
  wire  Queue_3_io_enq_bits_data_lock;
  wire [3:0] Queue_3_io_enq_bits_data_cache;
  wire [2:0] Queue_3_io_enq_bits_data_prot;
  wire [3:0] Queue_3_io_enq_bits_data_qos;
  wire [31:0] Queue_3_io_enq_bits_timestamp;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_data_id;
  wire [30:0] Queue_3_io_deq_bits_data_addr;
  wire [7:0] Queue_3_io_deq_bits_data_len;
  wire [2:0] Queue_3_io_deq_bits_data_size;
  wire [1:0] Queue_3_io_deq_bits_data_burst;
  wire  Queue_3_io_deq_bits_data_lock;
  wire [3:0] Queue_3_io_deq_bits_data_cache;
  wire [2:0] Queue_3_io_deq_bits_data_prot;
  wire [3:0] Queue_3_io_deq_bits_data_qos;
  wire [31:0] Queue_3_io_deq_bits_timestamp;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_data_id;
  wire [30:0] Queue_4_io_enq_bits_data_addr;
  wire [7:0] Queue_4_io_enq_bits_data_len;
  wire [2:0] Queue_4_io_enq_bits_data_size;
  wire [1:0] Queue_4_io_enq_bits_data_burst;
  wire  Queue_4_io_enq_bits_data_lock;
  wire [3:0] Queue_4_io_enq_bits_data_cache;
  wire [2:0] Queue_4_io_enq_bits_data_prot;
  wire [3:0] Queue_4_io_enq_bits_data_qos;
  wire [31:0] Queue_4_io_enq_bits_timestamp;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_data_id;
  wire [30:0] Queue_4_io_deq_bits_data_addr;
  wire [7:0] Queue_4_io_deq_bits_data_len;
  wire [2:0] Queue_4_io_deq_bits_data_size;
  wire [1:0] Queue_4_io_deq_bits_data_burst;
  wire  Queue_4_io_deq_bits_data_lock;
  wire [3:0] Queue_4_io_deq_bits_data_cache;
  wire [2:0] Queue_4_io_deq_bits_data_prot;
  wire [3:0] Queue_4_io_deq_bits_data_qos;
  wire [31:0] Queue_4_io_deq_bits_timestamp;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire [3:0] Queue_5_io_enq_bits_data_id;
  wire [30:0] Queue_5_io_enq_bits_data_addr;
  wire [7:0] Queue_5_io_enq_bits_data_len;
  wire [2:0] Queue_5_io_enq_bits_data_size;
  wire [1:0] Queue_5_io_enq_bits_data_burst;
  wire  Queue_5_io_enq_bits_data_lock;
  wire [3:0] Queue_5_io_enq_bits_data_cache;
  wire [2:0] Queue_5_io_enq_bits_data_prot;
  wire [3:0] Queue_5_io_enq_bits_data_qos;
  wire [31:0] Queue_5_io_enq_bits_timestamp;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire [3:0] Queue_5_io_deq_bits_data_id;
  wire [30:0] Queue_5_io_deq_bits_data_addr;
  wire [7:0] Queue_5_io_deq_bits_data_len;
  wire [2:0] Queue_5_io_deq_bits_data_size;
  wire [1:0] Queue_5_io_deq_bits_data_burst;
  wire  Queue_5_io_deq_bits_data_lock;
  wire [3:0] Queue_5_io_deq_bits_data_cache;
  wire [2:0] Queue_5_io_deq_bits_data_prot;
  wire [3:0] Queue_5_io_deq_bits_data_qos;
  wire [31:0] Queue_5_io_deq_bits_timestamp;
  wire  Queue_6_clock;
  wire  Queue_6_reset;
  wire  Queue_6_io_enq_ready;
  wire  Queue_6_io_enq_valid;
  wire [3:0] Queue_6_io_enq_bits_data_id;
  wire [30:0] Queue_6_io_enq_bits_data_addr;
  wire [7:0] Queue_6_io_enq_bits_data_len;
  wire [2:0] Queue_6_io_enq_bits_data_size;
  wire [1:0] Queue_6_io_enq_bits_data_burst;
  wire  Queue_6_io_enq_bits_data_lock;
  wire [3:0] Queue_6_io_enq_bits_data_cache;
  wire [2:0] Queue_6_io_enq_bits_data_prot;
  wire [3:0] Queue_6_io_enq_bits_data_qos;
  wire [31:0] Queue_6_io_enq_bits_timestamp;
  wire  Queue_6_io_deq_ready;
  wire  Queue_6_io_deq_valid;
  wire [3:0] Queue_6_io_deq_bits_data_id;
  wire [30:0] Queue_6_io_deq_bits_data_addr;
  wire [7:0] Queue_6_io_deq_bits_data_len;
  wire [2:0] Queue_6_io_deq_bits_data_size;
  wire [1:0] Queue_6_io_deq_bits_data_burst;
  wire  Queue_6_io_deq_bits_data_lock;
  wire [3:0] Queue_6_io_deq_bits_data_cache;
  wire [2:0] Queue_6_io_deq_bits_data_prot;
  wire [3:0] Queue_6_io_deq_bits_data_qos;
  wire [31:0] Queue_6_io_deq_bits_timestamp;
  wire  Queue_7_clock;
  wire  Queue_7_reset;
  wire  Queue_7_io_enq_ready;
  wire  Queue_7_io_enq_valid;
  wire [3:0] Queue_7_io_enq_bits_data_id;
  wire [30:0] Queue_7_io_enq_bits_data_addr;
  wire [7:0] Queue_7_io_enq_bits_data_len;
  wire [2:0] Queue_7_io_enq_bits_data_size;
  wire [1:0] Queue_7_io_enq_bits_data_burst;
  wire  Queue_7_io_enq_bits_data_lock;
  wire [3:0] Queue_7_io_enq_bits_data_cache;
  wire [2:0] Queue_7_io_enq_bits_data_prot;
  wire [3:0] Queue_7_io_enq_bits_data_qos;
  wire [31:0] Queue_7_io_enq_bits_timestamp;
  wire  Queue_7_io_deq_ready;
  wire  Queue_7_io_deq_valid;
  wire [3:0] Queue_7_io_deq_bits_data_id;
  wire [30:0] Queue_7_io_deq_bits_data_addr;
  wire [7:0] Queue_7_io_deq_bits_data_len;
  wire [2:0] Queue_7_io_deq_bits_data_size;
  wire [1:0] Queue_7_io_deq_bits_data_burst;
  wire  Queue_7_io_deq_bits_data_lock;
  wire [3:0] Queue_7_io_deq_bits_data_cache;
  wire [2:0] Queue_7_io_deq_bits_data_prot;
  wire [3:0] Queue_7_io_deq_bits_data_qos;
  wire [31:0] Queue_7_io_deq_bits_timestamp;
  wire  Queue_8_clock;
  wire  Queue_8_reset;
  wire  Queue_8_io_enq_ready;
  wire  Queue_8_io_enq_valid;
  wire [3:0] Queue_8_io_enq_bits_data_id;
  wire [30:0] Queue_8_io_enq_bits_data_addr;
  wire [7:0] Queue_8_io_enq_bits_data_len;
  wire [2:0] Queue_8_io_enq_bits_data_size;
  wire [1:0] Queue_8_io_enq_bits_data_burst;
  wire  Queue_8_io_enq_bits_data_lock;
  wire [3:0] Queue_8_io_enq_bits_data_cache;
  wire [2:0] Queue_8_io_enq_bits_data_prot;
  wire [3:0] Queue_8_io_enq_bits_data_qos;
  wire [31:0] Queue_8_io_enq_bits_timestamp;
  wire  Queue_8_io_deq_ready;
  wire  Queue_8_io_deq_valid;
  wire [3:0] Queue_8_io_deq_bits_data_id;
  wire [30:0] Queue_8_io_deq_bits_data_addr;
  wire [7:0] Queue_8_io_deq_bits_data_len;
  wire [2:0] Queue_8_io_deq_bits_data_size;
  wire [1:0] Queue_8_io_deq_bits_data_burst;
  wire  Queue_8_io_deq_bits_data_lock;
  wire [3:0] Queue_8_io_deq_bits_data_cache;
  wire [2:0] Queue_8_io_deq_bits_data_prot;
  wire [3:0] Queue_8_io_deq_bits_data_qos;
  wire [31:0] Queue_8_io_deq_bits_timestamp;
  wire  Queue_9_clock;
  wire  Queue_9_reset;
  wire  Queue_9_io_enq_ready;
  wire  Queue_9_io_enq_valid;
  wire [3:0] Queue_9_io_enq_bits_id;
  wire [30:0] Queue_9_io_enq_bits_addr;
  wire [7:0] Queue_9_io_enq_bits_len;
  wire [2:0] Queue_9_io_enq_bits_size;
  wire [1:0] Queue_9_io_enq_bits_burst;
  wire  Queue_9_io_deq_ready;
  wire  Queue_9_io_deq_valid;
  wire [3:0] Queue_9_io_deq_bits_id;
  wire [30:0] Queue_9_io_deq_bits_addr;
  wire [7:0] Queue_9_io_deq_bits_len;
  wire [2:0] Queue_9_io_deq_bits_size;
  wire [1:0] Queue_9_io_deq_bits_burst;
  wire  Queue_10_clock;
  wire  Queue_10_reset;
  wire  Queue_10_io_enq_ready;
  wire  Queue_10_io_enq_valid;
  wire [2:0] Queue_10_io_enq_bits;
  wire  Queue_10_io_deq_ready;
  wire  Queue_10_io_deq_valid;
  wire [2:0] Queue_10_io_deq_bits;
  wire  Queue_11_clock;
  wire  Queue_11_reset;
  wire  Queue_11_io_enq_ready;
  wire  Queue_11_io_enq_valid;
  wire [3:0] Queue_11_io_enq_bits_id;
  wire [30:0] Queue_11_io_enq_bits_addr;
  wire [7:0] Queue_11_io_enq_bits_len;
  wire [2:0] Queue_11_io_enq_bits_size;
  wire [1:0] Queue_11_io_enq_bits_burst;
  wire  Queue_11_io_deq_ready;
  wire  Queue_11_io_deq_valid;
  wire [3:0] Queue_11_io_deq_bits_id;
  wire [30:0] Queue_11_io_deq_bits_addr;
  wire [7:0] Queue_11_io_deq_bits_len;
  wire [2:0] Queue_11_io_deq_bits_size;
  wire [1:0] Queue_11_io_deq_bits_burst;
  wire  Queue_12_clock;
  wire  Queue_12_reset;
  wire  Queue_12_io_enq_ready;
  wire  Queue_12_io_enq_valid;
  wire [31:0] Queue_12_io_enq_bits_data;
  wire [3:0] Queue_12_io_enq_bits_strb;
  wire  Queue_12_io_enq_bits_last;
  wire  Queue_12_io_deq_ready;
  wire  Queue_12_io_deq_valid;
  wire [31:0] Queue_12_io_deq_bits_data;
  wire [3:0] Queue_12_io_deq_bits_strb;
  wire  Queue_12_io_deq_bits_last;
  wire  Queue_13_clock;
  wire  Queue_13_reset;
  wire  Queue_13_io_enq_ready;
  wire  Queue_13_io_enq_valid;
  wire [31:0] Queue_13_io_enq_bits_data;
  wire [3:0] Queue_13_io_enq_bits_strb;
  wire  Queue_13_io_enq_bits_last;
  wire  Queue_13_io_deq_ready;
  wire  Queue_13_io_deq_valid;
  wire [31:0] Queue_13_io_deq_bits_data;
  wire [3:0] Queue_13_io_deq_bits_strb;
  wire  Queue_13_io_deq_bits_last;
  wire  Queue_14_clock;
  wire  Queue_14_reset;
  wire  Queue_14_io_enq_ready;
  wire  Queue_14_io_enq_valid;
  wire [31:0] Queue_14_io_enq_bits_data;
  wire [3:0] Queue_14_io_enq_bits_strb;
  wire  Queue_14_io_enq_bits_last;
  wire  Queue_14_io_deq_ready;
  wire  Queue_14_io_deq_valid;
  wire [31:0] Queue_14_io_deq_bits_data;
  wire [3:0] Queue_14_io_deq_bits_strb;
  wire  Queue_14_io_deq_bits_last;
  wire  Queue_15_clock;
  wire  Queue_15_reset;
  wire  Queue_15_io_enq_ready;
  wire  Queue_15_io_enq_valid;
  wire [31:0] Queue_15_io_enq_bits_data;
  wire [3:0] Queue_15_io_enq_bits_strb;
  wire  Queue_15_io_enq_bits_last;
  wire  Queue_15_io_deq_ready;
  wire  Queue_15_io_deq_valid;
  wire [31:0] Queue_15_io_deq_bits_data;
  wire [3:0] Queue_15_io_deq_bits_strb;
  wire  Queue_15_io_deq_bits_last;
  wire  Queue_16_clock;
  wire  Queue_16_reset;
  wire  Queue_16_io_enq_ready;
  wire  Queue_16_io_enq_valid;
  wire [31:0] Queue_16_io_enq_bits_data;
  wire [3:0] Queue_16_io_enq_bits_strb;
  wire  Queue_16_io_enq_bits_last;
  wire  Queue_16_io_deq_ready;
  wire  Queue_16_io_deq_valid;
  wire [31:0] Queue_16_io_deq_bits_data;
  wire [3:0] Queue_16_io_deq_bits_strb;
  wire  Queue_16_io_deq_bits_last;
  wire  Queue_17_clock;
  wire  Queue_17_reset;
  wire  Queue_17_io_enq_ready;
  wire  Queue_17_io_enq_valid;
  wire [31:0] Queue_17_io_enq_bits_data;
  wire [3:0] Queue_17_io_enq_bits_strb;
  wire  Queue_17_io_enq_bits_last;
  wire  Queue_17_io_deq_ready;
  wire  Queue_17_io_deq_valid;
  wire [31:0] Queue_17_io_deq_bits_data;
  wire [3:0] Queue_17_io_deq_bits_strb;
  wire  Queue_17_io_deq_bits_last;
  wire  Queue_18_clock;
  wire  Queue_18_reset;
  wire  Queue_18_io_enq_ready;
  wire  Queue_18_io_enq_valid;
  wire [31:0] Queue_18_io_enq_bits_data;
  wire [3:0] Queue_18_io_enq_bits_strb;
  wire  Queue_18_io_enq_bits_last;
  wire  Queue_18_io_deq_ready;
  wire  Queue_18_io_deq_valid;
  wire [31:0] Queue_18_io_deq_bits_data;
  wire [3:0] Queue_18_io_deq_bits_strb;
  wire  Queue_18_io_deq_bits_last;
  wire  Queue_19_clock;
  wire  Queue_19_reset;
  wire  Queue_19_io_enq_ready;
  wire  Queue_19_io_enq_valid;
  wire [31:0] Queue_19_io_enq_bits_data;
  wire [3:0] Queue_19_io_enq_bits_strb;
  wire  Queue_19_io_enq_bits_last;
  wire  Queue_19_io_deq_ready;
  wire  Queue_19_io_deq_valid;
  wire [31:0] Queue_19_io_deq_bits_data;
  wire [3:0] Queue_19_io_deq_bits_strb;
  wire  Queue_19_io_deq_bits_last;
  wire [31:0] plusarg_reader_1_out;
  wire  MaxPeriodFibonacciLFSR_1__EVAL;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_17;
  wire  Queue_20_clock;
  wire  Queue_20_reset;
  wire  Queue_20_io_enq_ready;
  wire  Queue_20_io_enq_valid;
  wire [3:0] Queue_20_io_enq_bits_data_id;
  wire [30:0] Queue_20_io_enq_bits_data_addr;
  wire [7:0] Queue_20_io_enq_bits_data_len;
  wire [2:0] Queue_20_io_enq_bits_data_size;
  wire [1:0] Queue_20_io_enq_bits_data_burst;
  wire  Queue_20_io_enq_bits_data_lock;
  wire [3:0] Queue_20_io_enq_bits_data_cache;
  wire [2:0] Queue_20_io_enq_bits_data_prot;
  wire [3:0] Queue_20_io_enq_bits_data_qos;
  wire [31:0] Queue_20_io_enq_bits_timestamp;
  wire  Queue_20_io_deq_ready;
  wire  Queue_20_io_deq_valid;
  wire [3:0] Queue_20_io_deq_bits_data_id;
  wire [30:0] Queue_20_io_deq_bits_data_addr;
  wire [7:0] Queue_20_io_deq_bits_data_len;
  wire [2:0] Queue_20_io_deq_bits_data_size;
  wire [1:0] Queue_20_io_deq_bits_data_burst;
  wire  Queue_20_io_deq_bits_data_lock;
  wire [3:0] Queue_20_io_deq_bits_data_cache;
  wire [2:0] Queue_20_io_deq_bits_data_prot;
  wire [3:0] Queue_20_io_deq_bits_data_qos;
  wire [31:0] Queue_20_io_deq_bits_timestamp;
  wire  Queue_21_clock;
  wire  Queue_21_reset;
  wire  Queue_21_io_enq_ready;
  wire  Queue_21_io_enq_valid;
  wire [3:0] Queue_21_io_enq_bits_data_id;
  wire [30:0] Queue_21_io_enq_bits_data_addr;
  wire [7:0] Queue_21_io_enq_bits_data_len;
  wire [2:0] Queue_21_io_enq_bits_data_size;
  wire [1:0] Queue_21_io_enq_bits_data_burst;
  wire  Queue_21_io_enq_bits_data_lock;
  wire [3:0] Queue_21_io_enq_bits_data_cache;
  wire [2:0] Queue_21_io_enq_bits_data_prot;
  wire [3:0] Queue_21_io_enq_bits_data_qos;
  wire [31:0] Queue_21_io_enq_bits_timestamp;
  wire  Queue_21_io_deq_ready;
  wire  Queue_21_io_deq_valid;
  wire [3:0] Queue_21_io_deq_bits_data_id;
  wire [30:0] Queue_21_io_deq_bits_data_addr;
  wire [7:0] Queue_21_io_deq_bits_data_len;
  wire [2:0] Queue_21_io_deq_bits_data_size;
  wire [1:0] Queue_21_io_deq_bits_data_burst;
  wire  Queue_21_io_deq_bits_data_lock;
  wire [3:0] Queue_21_io_deq_bits_data_cache;
  wire [2:0] Queue_21_io_deq_bits_data_prot;
  wire [3:0] Queue_21_io_deq_bits_data_qos;
  wire [31:0] Queue_21_io_deq_bits_timestamp;
  wire  Queue_22_clock;
  wire  Queue_22_reset;
  wire  Queue_22_io_enq_ready;
  wire  Queue_22_io_enq_valid;
  wire [3:0] Queue_22_io_enq_bits_data_id;
  wire [30:0] Queue_22_io_enq_bits_data_addr;
  wire [7:0] Queue_22_io_enq_bits_data_len;
  wire [2:0] Queue_22_io_enq_bits_data_size;
  wire [1:0] Queue_22_io_enq_bits_data_burst;
  wire  Queue_22_io_enq_bits_data_lock;
  wire [3:0] Queue_22_io_enq_bits_data_cache;
  wire [2:0] Queue_22_io_enq_bits_data_prot;
  wire [3:0] Queue_22_io_enq_bits_data_qos;
  wire [31:0] Queue_22_io_enq_bits_timestamp;
  wire  Queue_22_io_deq_ready;
  wire  Queue_22_io_deq_valid;
  wire [3:0] Queue_22_io_deq_bits_data_id;
  wire [30:0] Queue_22_io_deq_bits_data_addr;
  wire [7:0] Queue_22_io_deq_bits_data_len;
  wire [2:0] Queue_22_io_deq_bits_data_size;
  wire [1:0] Queue_22_io_deq_bits_data_burst;
  wire  Queue_22_io_deq_bits_data_lock;
  wire [3:0] Queue_22_io_deq_bits_data_cache;
  wire [2:0] Queue_22_io_deq_bits_data_prot;
  wire [3:0] Queue_22_io_deq_bits_data_qos;
  wire [31:0] Queue_22_io_deq_bits_timestamp;
  wire  Queue_23_clock;
  wire  Queue_23_reset;
  wire  Queue_23_io_enq_ready;
  wire  Queue_23_io_enq_valid;
  wire [3:0] Queue_23_io_enq_bits_data_id;
  wire [30:0] Queue_23_io_enq_bits_data_addr;
  wire [7:0] Queue_23_io_enq_bits_data_len;
  wire [2:0] Queue_23_io_enq_bits_data_size;
  wire [1:0] Queue_23_io_enq_bits_data_burst;
  wire  Queue_23_io_enq_bits_data_lock;
  wire [3:0] Queue_23_io_enq_bits_data_cache;
  wire [2:0] Queue_23_io_enq_bits_data_prot;
  wire [3:0] Queue_23_io_enq_bits_data_qos;
  wire [31:0] Queue_23_io_enq_bits_timestamp;
  wire  Queue_23_io_deq_ready;
  wire  Queue_23_io_deq_valid;
  wire [3:0] Queue_23_io_deq_bits_data_id;
  wire [30:0] Queue_23_io_deq_bits_data_addr;
  wire [7:0] Queue_23_io_deq_bits_data_len;
  wire [2:0] Queue_23_io_deq_bits_data_size;
  wire [1:0] Queue_23_io_deq_bits_data_burst;
  wire  Queue_23_io_deq_bits_data_lock;
  wire [3:0] Queue_23_io_deq_bits_data_cache;
  wire [2:0] Queue_23_io_deq_bits_data_prot;
  wire [3:0] Queue_23_io_deq_bits_data_qos;
  wire [31:0] Queue_23_io_deq_bits_timestamp;
  wire  Queue_24_clock;
  wire  Queue_24_reset;
  wire  Queue_24_io_enq_ready;
  wire  Queue_24_io_enq_valid;
  wire [3:0] Queue_24_io_enq_bits_data_id;
  wire [30:0] Queue_24_io_enq_bits_data_addr;
  wire [7:0] Queue_24_io_enq_bits_data_len;
  wire [2:0] Queue_24_io_enq_bits_data_size;
  wire [1:0] Queue_24_io_enq_bits_data_burst;
  wire  Queue_24_io_enq_bits_data_lock;
  wire [3:0] Queue_24_io_enq_bits_data_cache;
  wire [2:0] Queue_24_io_enq_bits_data_prot;
  wire [3:0] Queue_24_io_enq_bits_data_qos;
  wire [31:0] Queue_24_io_enq_bits_timestamp;
  wire  Queue_24_io_deq_ready;
  wire  Queue_24_io_deq_valid;
  wire [3:0] Queue_24_io_deq_bits_data_id;
  wire [30:0] Queue_24_io_deq_bits_data_addr;
  wire [7:0] Queue_24_io_deq_bits_data_len;
  wire [2:0] Queue_24_io_deq_bits_data_size;
  wire [1:0] Queue_24_io_deq_bits_data_burst;
  wire  Queue_24_io_deq_bits_data_lock;
  wire [3:0] Queue_24_io_deq_bits_data_cache;
  wire [2:0] Queue_24_io_deq_bits_data_prot;
  wire [3:0] Queue_24_io_deq_bits_data_qos;
  wire [31:0] Queue_24_io_deq_bits_timestamp;
  wire  Queue_25_clock;
  wire  Queue_25_reset;
  wire  Queue_25_io_enq_ready;
  wire  Queue_25_io_enq_valid;
  wire [3:0] Queue_25_io_enq_bits_data_id;
  wire [30:0] Queue_25_io_enq_bits_data_addr;
  wire [7:0] Queue_25_io_enq_bits_data_len;
  wire [2:0] Queue_25_io_enq_bits_data_size;
  wire [1:0] Queue_25_io_enq_bits_data_burst;
  wire  Queue_25_io_enq_bits_data_lock;
  wire [3:0] Queue_25_io_enq_bits_data_cache;
  wire [2:0] Queue_25_io_enq_bits_data_prot;
  wire [3:0] Queue_25_io_enq_bits_data_qos;
  wire [31:0] Queue_25_io_enq_bits_timestamp;
  wire  Queue_25_io_deq_ready;
  wire  Queue_25_io_deq_valid;
  wire [3:0] Queue_25_io_deq_bits_data_id;
  wire [30:0] Queue_25_io_deq_bits_data_addr;
  wire [7:0] Queue_25_io_deq_bits_data_len;
  wire [2:0] Queue_25_io_deq_bits_data_size;
  wire [1:0] Queue_25_io_deq_bits_data_burst;
  wire  Queue_25_io_deq_bits_data_lock;
  wire [3:0] Queue_25_io_deq_bits_data_cache;
  wire [2:0] Queue_25_io_deq_bits_data_prot;
  wire [3:0] Queue_25_io_deq_bits_data_qos;
  wire [31:0] Queue_25_io_deq_bits_timestamp;
  wire  Queue_26_clock;
  wire  Queue_26_reset;
  wire  Queue_26_io_enq_ready;
  wire  Queue_26_io_enq_valid;
  wire [3:0] Queue_26_io_enq_bits_data_id;
  wire [30:0] Queue_26_io_enq_bits_data_addr;
  wire [7:0] Queue_26_io_enq_bits_data_len;
  wire [2:0] Queue_26_io_enq_bits_data_size;
  wire [1:0] Queue_26_io_enq_bits_data_burst;
  wire  Queue_26_io_enq_bits_data_lock;
  wire [3:0] Queue_26_io_enq_bits_data_cache;
  wire [2:0] Queue_26_io_enq_bits_data_prot;
  wire [3:0] Queue_26_io_enq_bits_data_qos;
  wire [31:0] Queue_26_io_enq_bits_timestamp;
  wire  Queue_26_io_deq_ready;
  wire  Queue_26_io_deq_valid;
  wire [3:0] Queue_26_io_deq_bits_data_id;
  wire [30:0] Queue_26_io_deq_bits_data_addr;
  wire [7:0] Queue_26_io_deq_bits_data_len;
  wire [2:0] Queue_26_io_deq_bits_data_size;
  wire [1:0] Queue_26_io_deq_bits_data_burst;
  wire  Queue_26_io_deq_bits_data_lock;
  wire [3:0] Queue_26_io_deq_bits_data_cache;
  wire [2:0] Queue_26_io_deq_bits_data_prot;
  wire [3:0] Queue_26_io_deq_bits_data_qos;
  wire [31:0] Queue_26_io_deq_bits_timestamp;
  wire  Queue_27_clock;
  wire  Queue_27_reset;
  wire  Queue_27_io_enq_ready;
  wire  Queue_27_io_enq_valid;
  wire [3:0] Queue_27_io_enq_bits_data_id;
  wire [30:0] Queue_27_io_enq_bits_data_addr;
  wire [7:0] Queue_27_io_enq_bits_data_len;
  wire [2:0] Queue_27_io_enq_bits_data_size;
  wire [1:0] Queue_27_io_enq_bits_data_burst;
  wire  Queue_27_io_enq_bits_data_lock;
  wire [3:0] Queue_27_io_enq_bits_data_cache;
  wire [2:0] Queue_27_io_enq_bits_data_prot;
  wire [3:0] Queue_27_io_enq_bits_data_qos;
  wire [31:0] Queue_27_io_enq_bits_timestamp;
  wire  Queue_27_io_deq_ready;
  wire  Queue_27_io_deq_valid;
  wire [3:0] Queue_27_io_deq_bits_data_id;
  wire [30:0] Queue_27_io_deq_bits_data_addr;
  wire [7:0] Queue_27_io_deq_bits_data_len;
  wire [2:0] Queue_27_io_deq_bits_data_size;
  wire [1:0] Queue_27_io_deq_bits_data_burst;
  wire  Queue_27_io_deq_bits_data_lock;
  wire [3:0] Queue_27_io_deq_bits_data_cache;
  wire [2:0] Queue_27_io_deq_bits_data_prot;
  wire [3:0] Queue_27_io_deq_bits_data_qos;
  wire [31:0] Queue_27_io_deq_bits_timestamp;
  wire  Queue_28_clock;
  wire  Queue_28_reset;
  wire  Queue_28_io_enq_ready;
  wire  Queue_28_io_enq_valid;
  wire [3:0] Queue_28_io_enq_bits_id;
  wire [30:0] Queue_28_io_enq_bits_addr;
  wire [7:0] Queue_28_io_enq_bits_len;
  wire [2:0] Queue_28_io_enq_bits_size;
  wire [1:0] Queue_28_io_enq_bits_burst;
  wire  Queue_28_io_deq_ready;
  wire  Queue_28_io_deq_valid;
  wire [3:0] Queue_28_io_deq_bits_id;
  wire [30:0] Queue_28_io_deq_bits_addr;
  wire [7:0] Queue_28_io_deq_bits_len;
  wire [2:0] Queue_28_io_deq_bits_size;
  wire [1:0] Queue_28_io_deq_bits_burst;
  wire [31:0] plusarg_reader_2_out;
  wire  MaxPeriodFibonacciLFSR_2__EVAL;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_2__EVAL_17;
  wire  Queue_29_clock;
  wire  Queue_29_reset;
  wire  Queue_29_io_enq_ready;
  wire  Queue_29_io_enq_valid;
  wire [3:0] Queue_29_io_enq_bits_data_id;
  wire [1:0] Queue_29_io_enq_bits_data_resp;
  wire [31:0] Queue_29_io_enq_bits_timestamp;
  wire  Queue_29_io_deq_ready;
  wire  Queue_29_io_deq_valid;
  wire [3:0] Queue_29_io_deq_bits_data_id;
  wire [1:0] Queue_29_io_deq_bits_data_resp;
  wire [31:0] Queue_29_io_deq_bits_timestamp;
  wire  Queue_30_clock;
  wire  Queue_30_reset;
  wire  Queue_30_io_enq_ready;
  wire  Queue_30_io_enq_valid;
  wire [3:0] Queue_30_io_enq_bits_data_id;
  wire [1:0] Queue_30_io_enq_bits_data_resp;
  wire [31:0] Queue_30_io_enq_bits_timestamp;
  wire  Queue_30_io_deq_ready;
  wire  Queue_30_io_deq_valid;
  wire [3:0] Queue_30_io_deq_bits_data_id;
  wire [1:0] Queue_30_io_deq_bits_data_resp;
  wire [31:0] Queue_30_io_deq_bits_timestamp;
  wire  Queue_31_clock;
  wire  Queue_31_reset;
  wire  Queue_31_io_enq_ready;
  wire  Queue_31_io_enq_valid;
  wire [3:0] Queue_31_io_enq_bits_data_id;
  wire [1:0] Queue_31_io_enq_bits_data_resp;
  wire [31:0] Queue_31_io_enq_bits_timestamp;
  wire  Queue_31_io_deq_ready;
  wire  Queue_31_io_deq_valid;
  wire [3:0] Queue_31_io_deq_bits_data_id;
  wire [1:0] Queue_31_io_deq_bits_data_resp;
  wire [31:0] Queue_31_io_deq_bits_timestamp;
  wire  Queue_32_clock;
  wire  Queue_32_reset;
  wire  Queue_32_io_enq_ready;
  wire  Queue_32_io_enq_valid;
  wire [3:0] Queue_32_io_enq_bits_data_id;
  wire [1:0] Queue_32_io_enq_bits_data_resp;
  wire [31:0] Queue_32_io_enq_bits_timestamp;
  wire  Queue_32_io_deq_ready;
  wire  Queue_32_io_deq_valid;
  wire [3:0] Queue_32_io_deq_bits_data_id;
  wire [1:0] Queue_32_io_deq_bits_data_resp;
  wire [31:0] Queue_32_io_deq_bits_timestamp;
  wire  Queue_33_clock;
  wire  Queue_33_reset;
  wire  Queue_33_io_enq_ready;
  wire  Queue_33_io_enq_valid;
  wire [3:0] Queue_33_io_enq_bits_data_id;
  wire [1:0] Queue_33_io_enq_bits_data_resp;
  wire [31:0] Queue_33_io_enq_bits_timestamp;
  wire  Queue_33_io_deq_ready;
  wire  Queue_33_io_deq_valid;
  wire [3:0] Queue_33_io_deq_bits_data_id;
  wire [1:0] Queue_33_io_deq_bits_data_resp;
  wire [31:0] Queue_33_io_deq_bits_timestamp;
  wire  Queue_34_clock;
  wire  Queue_34_reset;
  wire  Queue_34_io_enq_ready;
  wire  Queue_34_io_enq_valid;
  wire [3:0] Queue_34_io_enq_bits_data_id;
  wire [1:0] Queue_34_io_enq_bits_data_resp;
  wire [31:0] Queue_34_io_enq_bits_timestamp;
  wire  Queue_34_io_deq_ready;
  wire  Queue_34_io_deq_valid;
  wire [3:0] Queue_34_io_deq_bits_data_id;
  wire [1:0] Queue_34_io_deq_bits_data_resp;
  wire [31:0] Queue_34_io_deq_bits_timestamp;
  wire  Queue_35_clock;
  wire  Queue_35_reset;
  wire  Queue_35_io_enq_ready;
  wire  Queue_35_io_enq_valid;
  wire [3:0] Queue_35_io_enq_bits_data_id;
  wire [1:0] Queue_35_io_enq_bits_data_resp;
  wire [31:0] Queue_35_io_enq_bits_timestamp;
  wire  Queue_35_io_deq_ready;
  wire  Queue_35_io_deq_valid;
  wire [3:0] Queue_35_io_deq_bits_data_id;
  wire [1:0] Queue_35_io_deq_bits_data_resp;
  wire [31:0] Queue_35_io_deq_bits_timestamp;
  wire  Queue_36_clock;
  wire  Queue_36_reset;
  wire  Queue_36_io_enq_ready;
  wire  Queue_36_io_enq_valid;
  wire [3:0] Queue_36_io_enq_bits_data_id;
  wire [1:0] Queue_36_io_enq_bits_data_resp;
  wire [31:0] Queue_36_io_enq_bits_timestamp;
  wire  Queue_36_io_deq_ready;
  wire  Queue_36_io_deq_valid;
  wire [3:0] Queue_36_io_deq_bits_data_id;
  wire [1:0] Queue_36_io_deq_bits_data_resp;
  wire [31:0] Queue_36_io_deq_bits_timestamp;
  wire  Queue_37_clock;
  wire  Queue_37_reset;
  wire  Queue_37_io_enq_ready;
  wire  Queue_37_io_enq_valid;
  wire [3:0] Queue_37_io_enq_bits_id;
  wire [1:0] Queue_37_io_enq_bits_resp;
  wire  Queue_37_io_deq_ready;
  wire  Queue_37_io_deq_valid;
  wire [3:0] Queue_37_io_deq_bits_id;
  wire [1:0] Queue_37_io_deq_bits_resp;
  wire [31:0] plusarg_reader_3_out;
  wire  MaxPeriodFibonacciLFSR_3__EVAL;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_3__EVAL_17;
  wire  Queue_38_clock;
  wire  Queue_38_reset;
  wire  Queue_38_io_enq_ready;
  wire  Queue_38_io_enq_valid;
  wire [3:0] Queue_38_io_enq_bits_data_id;
  wire [31:0] Queue_38_io_enq_bits_data_data;
  wire [1:0] Queue_38_io_enq_bits_data_resp;
  wire  Queue_38_io_enq_bits_data_last;
  wire [31:0] Queue_38_io_enq_bits_timestamp;
  wire  Queue_38_io_deq_ready;
  wire  Queue_38_io_deq_valid;
  wire [3:0] Queue_38_io_deq_bits_data_id;
  wire [31:0] Queue_38_io_deq_bits_data_data;
  wire [1:0] Queue_38_io_deq_bits_data_resp;
  wire  Queue_38_io_deq_bits_data_last;
  wire [31:0] Queue_38_io_deq_bits_timestamp;
  wire  Queue_39_clock;
  wire  Queue_39_reset;
  wire  Queue_39_io_enq_ready;
  wire  Queue_39_io_enq_valid;
  wire [3:0] Queue_39_io_enq_bits_data_id;
  wire [31:0] Queue_39_io_enq_bits_data_data;
  wire [1:0] Queue_39_io_enq_bits_data_resp;
  wire  Queue_39_io_enq_bits_data_last;
  wire [31:0] Queue_39_io_enq_bits_timestamp;
  wire  Queue_39_io_deq_ready;
  wire  Queue_39_io_deq_valid;
  wire [3:0] Queue_39_io_deq_bits_data_id;
  wire [31:0] Queue_39_io_deq_bits_data_data;
  wire [1:0] Queue_39_io_deq_bits_data_resp;
  wire  Queue_39_io_deq_bits_data_last;
  wire [31:0] Queue_39_io_deq_bits_timestamp;
  wire  Queue_40_clock;
  wire  Queue_40_reset;
  wire  Queue_40_io_enq_ready;
  wire  Queue_40_io_enq_valid;
  wire [3:0] Queue_40_io_enq_bits_data_id;
  wire [31:0] Queue_40_io_enq_bits_data_data;
  wire [1:0] Queue_40_io_enq_bits_data_resp;
  wire  Queue_40_io_enq_bits_data_last;
  wire [31:0] Queue_40_io_enq_bits_timestamp;
  wire  Queue_40_io_deq_ready;
  wire  Queue_40_io_deq_valid;
  wire [3:0] Queue_40_io_deq_bits_data_id;
  wire [31:0] Queue_40_io_deq_bits_data_data;
  wire [1:0] Queue_40_io_deq_bits_data_resp;
  wire  Queue_40_io_deq_bits_data_last;
  wire [31:0] Queue_40_io_deq_bits_timestamp;
  wire  Queue_41_clock;
  wire  Queue_41_reset;
  wire  Queue_41_io_enq_ready;
  wire  Queue_41_io_enq_valid;
  wire [3:0] Queue_41_io_enq_bits_data_id;
  wire [31:0] Queue_41_io_enq_bits_data_data;
  wire [1:0] Queue_41_io_enq_bits_data_resp;
  wire  Queue_41_io_enq_bits_data_last;
  wire [31:0] Queue_41_io_enq_bits_timestamp;
  wire  Queue_41_io_deq_ready;
  wire  Queue_41_io_deq_valid;
  wire [3:0] Queue_41_io_deq_bits_data_id;
  wire [31:0] Queue_41_io_deq_bits_data_data;
  wire [1:0] Queue_41_io_deq_bits_data_resp;
  wire  Queue_41_io_deq_bits_data_last;
  wire [31:0] Queue_41_io_deq_bits_timestamp;
  wire  Queue_42_clock;
  wire  Queue_42_reset;
  wire  Queue_42_io_enq_ready;
  wire  Queue_42_io_enq_valid;
  wire [3:0] Queue_42_io_enq_bits_data_id;
  wire [31:0] Queue_42_io_enq_bits_data_data;
  wire [1:0] Queue_42_io_enq_bits_data_resp;
  wire  Queue_42_io_enq_bits_data_last;
  wire [31:0] Queue_42_io_enq_bits_timestamp;
  wire  Queue_42_io_deq_ready;
  wire  Queue_42_io_deq_valid;
  wire [3:0] Queue_42_io_deq_bits_data_id;
  wire [31:0] Queue_42_io_deq_bits_data_data;
  wire [1:0] Queue_42_io_deq_bits_data_resp;
  wire  Queue_42_io_deq_bits_data_last;
  wire [31:0] Queue_42_io_deq_bits_timestamp;
  wire  Queue_43_clock;
  wire  Queue_43_reset;
  wire  Queue_43_io_enq_ready;
  wire  Queue_43_io_enq_valid;
  wire [3:0] Queue_43_io_enq_bits_data_id;
  wire [31:0] Queue_43_io_enq_bits_data_data;
  wire [1:0] Queue_43_io_enq_bits_data_resp;
  wire  Queue_43_io_enq_bits_data_last;
  wire [31:0] Queue_43_io_enq_bits_timestamp;
  wire  Queue_43_io_deq_ready;
  wire  Queue_43_io_deq_valid;
  wire [3:0] Queue_43_io_deq_bits_data_id;
  wire [31:0] Queue_43_io_deq_bits_data_data;
  wire [1:0] Queue_43_io_deq_bits_data_resp;
  wire  Queue_43_io_deq_bits_data_last;
  wire [31:0] Queue_43_io_deq_bits_timestamp;
  wire  Queue_44_clock;
  wire  Queue_44_reset;
  wire  Queue_44_io_enq_ready;
  wire  Queue_44_io_enq_valid;
  wire [3:0] Queue_44_io_enq_bits_data_id;
  wire [31:0] Queue_44_io_enq_bits_data_data;
  wire [1:0] Queue_44_io_enq_bits_data_resp;
  wire  Queue_44_io_enq_bits_data_last;
  wire [31:0] Queue_44_io_enq_bits_timestamp;
  wire  Queue_44_io_deq_ready;
  wire  Queue_44_io_deq_valid;
  wire [3:0] Queue_44_io_deq_bits_data_id;
  wire [31:0] Queue_44_io_deq_bits_data_data;
  wire [1:0] Queue_44_io_deq_bits_data_resp;
  wire  Queue_44_io_deq_bits_data_last;
  wire [31:0] Queue_44_io_deq_bits_timestamp;
  wire  Queue_45_clock;
  wire  Queue_45_reset;
  wire  Queue_45_io_enq_ready;
  wire  Queue_45_io_enq_valid;
  wire [3:0] Queue_45_io_enq_bits_data_id;
  wire [31:0] Queue_45_io_enq_bits_data_data;
  wire [1:0] Queue_45_io_enq_bits_data_resp;
  wire  Queue_45_io_enq_bits_data_last;
  wire [31:0] Queue_45_io_enq_bits_timestamp;
  wire  Queue_45_io_deq_ready;
  wire  Queue_45_io_deq_valid;
  wire [3:0] Queue_45_io_deq_bits_data_id;
  wire [31:0] Queue_45_io_deq_bits_data_data;
  wire [1:0] Queue_45_io_deq_bits_data_resp;
  wire  Queue_45_io_deq_bits_data_last;
  wire [31:0] Queue_45_io_deq_bits_timestamp;
  wire  Queue_46_clock;
  wire  Queue_46_reset;
  wire  Queue_46_io_enq_ready;
  wire  Queue_46_io_enq_valid;
  wire [3:0] Queue_46_io_enq_bits_id;
  wire [31:0] Queue_46_io_enq_bits_data;
  wire [1:0] Queue_46_io_enq_bits_resp;
  wire  Queue_46_io_enq_bits_last;
  wire  Queue_46_io_deq_ready;
  wire  Queue_46_io_deq_valid;
  wire [3:0] Queue_46_io_deq_bits_id;
  wire [31:0] Queue_46_io_deq_bits_data;
  wire [1:0] Queue_46_io_deq_bits_resp;
  wire  Queue_46_io_deq_bits_last;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_2;
  wire [2:0] _GEN_3;
  wire [2:0] _GEN_4;
  wire [2:0] _GEN_5;
  wire [2:0] _GEN_6;
  wire [2:0] _GEN_7;
  wire [2:0] _GEN_8;
  wire [2:0] _GEN_9;
  wire [2:0] _GEN_10;
  wire [2:0] _GEN_11;
  wire [2:0] _GEN_12;
  wire [2:0] _GEN_13;
  wire [2:0] _GEN_14;
  wire [2:0] _GEN_15;
  wire  _T_71_7;
  wire  _T_71_6;
  wire  _T_71_5;
  wire  _T_71_4;
  wire  _T_71_3;
  wire  _T_71_2;
  wire  _T_71_1;
  wire  _T_71_0;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire [7:0] _T_19;
  wire [15:0] _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_39;
  wire  _T_40;
  wire  _T_41;
  wire  _T_42;
  wire  _T_43;
  wire [7:0] _T_51;
  wire [15:0] _T_59;
  wire  _T_60;
  wire  _T_9;
  wire  _T_64;
  wire  _T_65;
  wire  _T_6;
  reg [31:0] _T_10;
  reg [31:0] _RAND_0;
  wire [31:0] _T_12;
  wire  _T_63;
  wire [31:0] _T_67;
  wire [1:0] _T_68;
  wire [31:0] _GEN_156;
  wire [7:0] _T_73;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  _T_80;
  wire  _T_81;
  wire  _T_82;
  wire  _T_93;
  wire  _T_94;
  wire  _T_95;
  wire  _T_91_ready;
  reg  _T_140;
  reg [31:0] _RAND_1;
  wire  _T_141;
  wire  _T_135;
  wire  _T_136;
  wire  _T_137;
  wire  _T_129;
  wire  _T_130;
  wire  _T_131;
  wire  _T_123;
  wire  _T_124;
  wire  _T_125;
  wire  _T_117;
  wire  _T_118;
  wire  _T_119;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  _T_99;
  wire  _T_100;
  wire  _T_101;
  wire [7:0] _T_149;
  reg [7:0] _T_156;
  reg [31:0] _RAND_2;
  wire [7:0] _T_157;
  wire [7:0] _T_158;
  wire [15:0] _T_159;
  wire [14:0] _T_160;
  wire [15:0] _GEN_157;
  wire [15:0] _T_161;
  wire [13:0] _T_162;
  wire [15:0] _GEN_158;
  wire [15:0] _T_163;
  wire [11:0] _T_164;
  wire [15:0] _GEN_159;
  wire [15:0] _T_165;
  wire [14:0] _T_167;
  wire [15:0] _T_168;
  wire [15:0] _GEN_160;
  wire [15:0] _T_169;
  wire [7:0] _T_170;
  wire [7:0] _T_171;
  wire [7:0] _T_172;
  wire [7:0] _T_173;
  wire  _T_188;
  reg  _T_287_0;
  reg [31:0] _RAND_3;
  wire  _T_289_0;
  wire  _T_290;
  wire  _T_189;
  reg  _T_287_1;
  reg [31:0] _RAND_4;
  wire  _T_289_1;
  wire  _T_291;
  wire  _T_190;
  reg  _T_287_2;
  reg [31:0] _RAND_5;
  wire  _T_289_2;
  wire  _T_292;
  wire  _T_191;
  reg  _T_287_3;
  reg [31:0] _RAND_6;
  wire  _T_289_3;
  wire  _T_293;
  wire  _T_192;
  reg  _T_287_4;
  reg [31:0] _RAND_7;
  wire  _T_289_4;
  wire  _T_294;
  wire  _T_193;
  reg  _T_287_5;
  reg [31:0] _RAND_8;
  wire  _T_289_5;
  wire  _T_295;
  wire  _T_194;
  reg  _T_287_6;
  reg [31:0] _RAND_9;
  wire  _T_289_6;
  wire  _T_296;
  wire  _T_195;
  reg  _T_287_7;
  reg [31:0] _RAND_10;
  wire  _T_289_7;
  wire  _T_297;
  wire  _T_142;
  wire  _T_151;
  wire  _T_153;
  wire  _T_154;
  wire  _T_174;
  wire  _T_175;
  wire [7:0] _T_176;
  wire [8:0] _T_177;
  wire [7:0] _T_178;
  wire [7:0] _T_179;
  wire [9:0] _T_180;
  wire [7:0] _T_181;
  wire [7:0] _T_182;
  wire [11:0] _T_183;
  wire [7:0] _T_184;
  wire [7:0] _T_185;
  wire  _T_197;
  wire  _T_198;
  wire  _T_199;
  wire  _T_200;
  wire  _T_201;
  wire  _T_202;
  wire  _T_203;
  wire  _T_204;
  wire  _T_207;
  wire  _T_208;
  wire  _T_209;
  wire  _T_210;
  wire  _T_211;
  wire  _T_212;
  wire  _T_213;
  wire  _T_215;
  wire  _T_218;
  wire  _T_219;
  wire  _T_220;
  wire  _T_221;
  wire  _T_222;
  wire  _T_223;
  wire  _T_224;
  wire  _T_225;
  wire  _T_226;
  wire  _T_227;
  wire  _T_228;
  wire  _T_229;
  wire  _T_230;
  wire  _T_231;
  wire  _T_232;
  wire  _T_233;
  wire  _T_234;
  wire  _T_235;
  wire  _T_236;
  wire  _T_237;
  wire  _T_239;
  wire  _T_240;
  wire  _T_241;
  wire  _T_242;
  wire  _T_243;
  wire  _T_244;
  wire  _T_246;
  wire  _T_247;
  wire  _T_248;
  wire  _T_249;
  wire  _T_250;
  wire  _T_251;
  wire  _T_252;
  wire  _T_253;
  wire  _T_254;
  wire  _T_255;
  wire  _T_263;
  wire  _T_265;
  wire  _T_266;
  wire  _T_305;
  wire  _T_306;
  wire  _T_313;
  wire  _T_307;
  wire  _T_314;
  wire  _T_308;
  wire  _T_315;
  wire  _T_309;
  wire  _T_316;
  wire  _T_310;
  wire  _T_317;
  wire  _T_311;
  wire  _T_318;
  wire  _T_312;
  wire  _T_319;
  wire  _T_321;
  wire  _T_282;
  wire  _T_284;
  wire  _T_288_0;
  wire  _T_288_1;
  wire  _T_288_2;
  wire  _T_288_3;
  wire  _T_288_4;
  wire  _T_288_5;
  wire  _T_288_6;
  wire  _T_288_7;
  wire [2:0] _T_92_bits_prot;
  wire [3:0] _T_92_bits_qos;
  wire  _T_92_bits_lock;
  wire [3:0] _T_92_bits_cache;
  wire [2:0] _T_92_bits_size;
  wire [1:0] _T_92_bits_burst;
  wire [3:0] _T_92_bits_id;
  wire [30:0] _T_92_bits_addr;
  wire [7:0] _T_92_bits_len;
  wire [59:0] _T_329;
  wire [59:0] _T_330;
  wire [2:0] _T_98_bits_prot;
  wire [3:0] _T_98_bits_qos;
  wire  _T_98_bits_lock;
  wire [3:0] _T_98_bits_cache;
  wire [2:0] _T_98_bits_size;
  wire [1:0] _T_98_bits_burst;
  wire [3:0] _T_98_bits_id;
  wire [30:0] _T_98_bits_addr;
  wire [7:0] _T_98_bits_len;
  wire [59:0] _T_338;
  wire [59:0] _T_339;
  wire [2:0] _T_104_bits_prot;
  wire [3:0] _T_104_bits_qos;
  wire  _T_104_bits_lock;
  wire [3:0] _T_104_bits_cache;
  wire [2:0] _T_104_bits_size;
  wire [1:0] _T_104_bits_burst;
  wire [3:0] _T_104_bits_id;
  wire [30:0] _T_104_bits_addr;
  wire [7:0] _T_104_bits_len;
  wire [59:0] _T_347;
  wire [59:0] _T_348;
  wire [2:0] _T_110_bits_prot;
  wire [3:0] _T_110_bits_qos;
  wire  _T_110_bits_lock;
  wire [3:0] _T_110_bits_cache;
  wire [2:0] _T_110_bits_size;
  wire [1:0] _T_110_bits_burst;
  wire [3:0] _T_110_bits_id;
  wire [30:0] _T_110_bits_addr;
  wire [7:0] _T_110_bits_len;
  wire [59:0] _T_356;
  wire [59:0] _T_357;
  wire [2:0] _T_116_bits_prot;
  wire [3:0] _T_116_bits_qos;
  wire  _T_116_bits_lock;
  wire [3:0] _T_116_bits_cache;
  wire [2:0] _T_116_bits_size;
  wire [1:0] _T_116_bits_burst;
  wire [3:0] _T_116_bits_id;
  wire [30:0] _T_116_bits_addr;
  wire [7:0] _T_116_bits_len;
  wire [59:0] _T_365;
  wire [59:0] _T_366;
  wire [2:0] _T_122_bits_prot;
  wire [3:0] _T_122_bits_qos;
  wire  _T_122_bits_lock;
  wire [3:0] _T_122_bits_cache;
  wire [2:0] _T_122_bits_size;
  wire [1:0] _T_122_bits_burst;
  wire [3:0] _T_122_bits_id;
  wire [30:0] _T_122_bits_addr;
  wire [7:0] _T_122_bits_len;
  wire [59:0] _T_374;
  wire [59:0] _T_375;
  wire [2:0] _T_128_bits_prot;
  wire [3:0] _T_128_bits_qos;
  wire  _T_128_bits_lock;
  wire [3:0] _T_128_bits_cache;
  wire [2:0] _T_128_bits_size;
  wire [1:0] _T_128_bits_burst;
  wire [3:0] _T_128_bits_id;
  wire [30:0] _T_128_bits_addr;
  wire [7:0] _T_128_bits_len;
  wire [59:0] _T_383;
  wire [59:0] _T_384;
  wire [2:0] _T_134_bits_prot;
  wire [3:0] _T_134_bits_qos;
  wire  _T_134_bits_lock;
  wire [3:0] _T_134_bits_cache;
  wire [2:0] _T_134_bits_size;
  wire [1:0] _T_134_bits_burst;
  wire [3:0] _T_134_bits_id;
  wire [30:0] _T_134_bits_addr;
  wire [7:0] _T_134_bits_len;
  wire [59:0] _T_392;
  wire [59:0] _T_393;
  wire [59:0] _T_394;
  wire [59:0] _T_395;
  wire [59:0] _T_396;
  wire [59:0] _T_397;
  wire [59:0] _T_398;
  wire [59:0] _T_399;
  wire [59:0] _T_400;
  wire  _T_413_ready;
  wire  _T_412_valid;
  wire [3:0] _T_412_bits_id;
  wire [2:0] _GEN_26;
  wire [2:0] _GEN_27;
  wire [2:0] _GEN_28;
  wire [2:0] _GEN_29;
  wire [2:0] _GEN_30;
  wire [2:0] _GEN_31;
  wire [2:0] _GEN_32;
  wire [2:0] _GEN_33;
  wire [2:0] _GEN_34;
  wire [2:0] _GEN_35;
  wire [2:0] _GEN_36;
  wire [2:0] _GEN_37;
  wire [2:0] _GEN_38;
  wire [2:0] _GEN_39;
  wire [2:0] _T_4_bits;
  wire  _T_418_0;
  wire  _T_418_1;
  wire  _GEN_42;
  wire  _T_418_2;
  wire  _GEN_43;
  wire  _T_418_3;
  wire  _GEN_44;
  wire  _T_418_4;
  wire  _GEN_45;
  wire  _T_418_5;
  wire  _GEN_46;
  wire  _T_418_6;
  wire  _GEN_47;
  wire  _T_418_7;
  wire  _GEN_48;
  wire  _T_419;
  wire  _T_4_valid;
  wire [7:0] _T_423;
  wire  _T_425;
  wire  _T_426;
  wire  _T_427;
  wire  _T_428;
  wire  _T_429;
  wire  _T_430;
  wire  _T_431;
  wire  _T_432;
  wire  _T_433;
  wire [2:0] _T_414_bits;
  wire [31:0] _T_451_0_data;
  wire [3:0] _T_451_0_strb;
  wire  _T_451_0_last;
  wire [31:0] _T_451_1_data;
  wire [31:0] _GEN_52;
  wire [3:0] _T_451_1_strb;
  wire [3:0] _GEN_53;
  wire  _T_451_1_last;
  wire  _GEN_54;
  wire [31:0] _T_451_2_data;
  wire [31:0] _GEN_55;
  wire [3:0] _T_451_2_strb;
  wire [3:0] _GEN_56;
  wire  _T_451_2_last;
  wire  _GEN_57;
  wire [31:0] _T_451_3_data;
  wire [31:0] _GEN_58;
  wire [3:0] _T_451_3_strb;
  wire [3:0] _GEN_59;
  wire  _T_451_3_last;
  wire  _GEN_60;
  wire [31:0] _T_451_4_data;
  wire [31:0] _GEN_61;
  wire [3:0] _T_451_4_strb;
  wire [3:0] _GEN_62;
  wire  _T_451_4_last;
  wire  _GEN_63;
  wire [31:0] _T_451_5_data;
  wire [31:0] _GEN_64;
  wire [3:0] _T_451_5_strb;
  wire [3:0] _GEN_65;
  wire  _T_451_5_last;
  wire  _GEN_66;
  wire [31:0] _T_451_6_data;
  wire [31:0] _GEN_67;
  wire [3:0] _T_451_6_strb;
  wire [3:0] _GEN_68;
  wire  _T_451_6_last;
  wire  _GEN_69;
  wire [31:0] _T_451_7_data;
  wire [3:0] _T_451_7_strb;
  wire  _T_451_7_last;
  wire  _GEN_72;
  wire  _T_450_0;
  wire  _T_450_1;
  wire  _GEN_74;
  wire  _T_450_2;
  wire  _GEN_75;
  wire  _T_450_3;
  wire  _GEN_76;
  wire  _T_450_4;
  wire  _GEN_77;
  wire  _T_450_5;
  wire  _GEN_78;
  wire  _T_450_6;
  wire  _GEN_79;
  wire  _T_450_7;
  wire  _GEN_80;
  wire  _T_452;
  wire  _T_414_valid;
  wire [7:0] _T_456;
  wire  _T_458;
  wire  _T_459;
  wire  _T_460;
  wire  _T_461;
  wire  _T_462;
  wire  _T_463;
  wire  _T_464;
  wire  _T_465;
  wire  _T_466;
  wire  _T_483;
  reg [31:0] _T_484;
  reg [31:0] _RAND_11;
  wire [31:0] _T_486;
  wire [7:0] _T_493;
  wire [15:0] _T_501;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_506;
  wire  _T_507;
  wire  _T_508;
  wire  _T_509;
  wire  _T_510;
  wire  _T_511;
  wire  _T_512;
  wire  _T_513;
  wire  _T_514;
  wire  _T_515;
  wire  _T_516;
  wire  _T_517;
  wire [7:0] _T_525;
  wire [15:0] _T_533;
  wire  _T_534;
  wire  _T_536;
  wire  _T_537;
  wire [2:0] _GEN_82;
  wire [2:0] _GEN_83;
  wire [2:0] _GEN_84;
  wire [2:0] _GEN_85;
  wire [2:0] _GEN_86;
  wire [2:0] _GEN_87;
  wire [2:0] _GEN_88;
  wire [2:0] _GEN_89;
  wire [2:0] _GEN_90;
  wire [2:0] _GEN_91;
  wire [2:0] _GEN_92;
  wire [2:0] _GEN_93;
  wire [2:0] _GEN_94;
  wire [2:0] _GEN_95;
  wire [2:0] _GEN_96;
  wire  _T_545_7;
  wire  _T_545_6;
  wire  _T_545_5;
  wire  _T_545_4;
  wire  _T_545_3;
  wire  _T_545_2;
  wire  _T_545_1;
  wire  _T_545_0;
  wire  _GEN_98;
  wire  _GEN_99;
  wire  _GEN_100;
  wire  _GEN_101;
  wire  _GEN_102;
  wire  _GEN_103;
  wire  _GEN_104;
  wire [31:0] _T_541;
  wire [1:0] _T_542;
  wire [31:0] _GEN_161;
  wire [7:0] _T_547;
  wire  _T_549;
  wire  _T_550;
  wire  _T_551;
  wire  _T_552;
  wire  _T_553;
  wire  _T_554;
  wire  _T_555;
  wire  _T_556;
  wire  _T_567;
  wire  _T_568;
  wire  _T_569;
  wire  _T_565_ready;
  reg  _T_614;
  reg [31:0] _RAND_12;
  wire  _T_615;
  wire  _T_609;
  wire  _T_610;
  wire  _T_611;
  wire  _T_603;
  wire  _T_604;
  wire  _T_605;
  wire  _T_597;
  wire  _T_598;
  wire  _T_599;
  wire  _T_591;
  wire  _T_592;
  wire  _T_593;
  wire  _T_585;
  wire  _T_586;
  wire  _T_587;
  wire  _T_579;
  wire  _T_580;
  wire  _T_581;
  wire  _T_573;
  wire  _T_574;
  wire  _T_575;
  wire [7:0] _T_623;
  reg [7:0] _T_630;
  reg [31:0] _RAND_13;
  wire [7:0] _T_631;
  wire [7:0] _T_632;
  wire [15:0] _T_633;
  wire [14:0] _T_634;
  wire [15:0] _GEN_162;
  wire [15:0] _T_635;
  wire [13:0] _T_636;
  wire [15:0] _GEN_163;
  wire [15:0] _T_637;
  wire [11:0] _T_638;
  wire [15:0] _GEN_164;
  wire [15:0] _T_639;
  wire [14:0] _T_641;
  wire [15:0] _T_642;
  wire [15:0] _GEN_165;
  wire [15:0] _T_643;
  wire [7:0] _T_644;
  wire [7:0] _T_645;
  wire [7:0] _T_646;
  wire [7:0] _T_647;
  wire  _T_662;
  reg  _T_761_0;
  reg [31:0] _RAND_14;
  wire  _T_763_0;
  wire  _T_764;
  wire  _T_663;
  reg  _T_761_1;
  reg [31:0] _RAND_15;
  wire  _T_763_1;
  wire  _T_765;
  wire  _T_664;
  reg  _T_761_2;
  reg [31:0] _RAND_16;
  wire  _T_763_2;
  wire  _T_766;
  wire  _T_665;
  reg  _T_761_3;
  reg [31:0] _RAND_17;
  wire  _T_763_3;
  wire  _T_767;
  wire  _T_666;
  reg  _T_761_4;
  reg [31:0] _RAND_18;
  wire  _T_763_4;
  wire  _T_768;
  wire  _T_667;
  reg  _T_761_5;
  reg [31:0] _RAND_19;
  wire  _T_763_5;
  wire  _T_769;
  wire  _T_668;
  reg  _T_761_6;
  reg [31:0] _RAND_20;
  wire  _T_763_6;
  wire  _T_770;
  wire  _T_669;
  reg  _T_761_7;
  reg [31:0] _RAND_21;
  wire  _T_763_7;
  wire  _T_771;
  wire  _T_616;
  wire  _T_625;
  wire  _T_627;
  wire  _T_628;
  wire  _T_648;
  wire  _T_649;
  wire [7:0] _T_650;
  wire [8:0] _T_651;
  wire [7:0] _T_652;
  wire [7:0] _T_653;
  wire [9:0] _T_654;
  wire [7:0] _T_655;
  wire [7:0] _T_656;
  wire [11:0] _T_657;
  wire [7:0] _T_658;
  wire [7:0] _T_659;
  wire  _T_671;
  wire  _T_672;
  wire  _T_673;
  wire  _T_674;
  wire  _T_675;
  wire  _T_676;
  wire  _T_677;
  wire  _T_678;
  wire  _T_681;
  wire  _T_682;
  wire  _T_683;
  wire  _T_684;
  wire  _T_685;
  wire  _T_686;
  wire  _T_687;
  wire  _T_689;
  wire  _T_692;
  wire  _T_693;
  wire  _T_694;
  wire  _T_695;
  wire  _T_696;
  wire  _T_697;
  wire  _T_698;
  wire  _T_699;
  wire  _T_700;
  wire  _T_701;
  wire  _T_702;
  wire  _T_703;
  wire  _T_704;
  wire  _T_705;
  wire  _T_706;
  wire  _T_707;
  wire  _T_708;
  wire  _T_709;
  wire  _T_710;
  wire  _T_711;
  wire  _T_713;
  wire  _T_714;
  wire  _T_715;
  wire  _T_716;
  wire  _T_717;
  wire  _T_718;
  wire  _T_720;
  wire  _T_721;
  wire  _T_722;
  wire  _T_723;
  wire  _T_724;
  wire  _T_725;
  wire  _T_726;
  wire  _T_727;
  wire  _T_728;
  wire  _T_729;
  wire  _T_737;
  wire  _T_739;
  wire  _T_740;
  wire  _T_779;
  wire  _T_780;
  wire  _T_787;
  wire  _T_781;
  wire  _T_788;
  wire  _T_782;
  wire  _T_789;
  wire  _T_783;
  wire  _T_790;
  wire  _T_784;
  wire  _T_791;
  wire  _T_785;
  wire  _T_792;
  wire  _T_786;
  wire  _T_793;
  wire  _T_795;
  wire  _T_756;
  wire  _T_758;
  wire  _T_762_0;
  wire  _T_762_1;
  wire  _T_762_2;
  wire  _T_762_3;
  wire  _T_762_4;
  wire  _T_762_5;
  wire  _T_762_6;
  wire  _T_762_7;
  wire [2:0] _T_566_bits_prot;
  wire [3:0] _T_566_bits_qos;
  wire  _T_566_bits_lock;
  wire [3:0] _T_566_bits_cache;
  wire [2:0] _T_566_bits_size;
  wire [1:0] _T_566_bits_burst;
  wire [3:0] _T_566_bits_id;
  wire [30:0] _T_566_bits_addr;
  wire [7:0] _T_566_bits_len;
  wire [59:0] _T_803;
  wire [59:0] _T_804;
  wire [2:0] _T_572_bits_prot;
  wire [3:0] _T_572_bits_qos;
  wire  _T_572_bits_lock;
  wire [3:0] _T_572_bits_cache;
  wire [2:0] _T_572_bits_size;
  wire [1:0] _T_572_bits_burst;
  wire [3:0] _T_572_bits_id;
  wire [30:0] _T_572_bits_addr;
  wire [7:0] _T_572_bits_len;
  wire [59:0] _T_812;
  wire [59:0] _T_813;
  wire [2:0] _T_578_bits_prot;
  wire [3:0] _T_578_bits_qos;
  wire  _T_578_bits_lock;
  wire [3:0] _T_578_bits_cache;
  wire [2:0] _T_578_bits_size;
  wire [1:0] _T_578_bits_burst;
  wire [3:0] _T_578_bits_id;
  wire [30:0] _T_578_bits_addr;
  wire [7:0] _T_578_bits_len;
  wire [59:0] _T_821;
  wire [59:0] _T_822;
  wire [2:0] _T_584_bits_prot;
  wire [3:0] _T_584_bits_qos;
  wire  _T_584_bits_lock;
  wire [3:0] _T_584_bits_cache;
  wire [2:0] _T_584_bits_size;
  wire [1:0] _T_584_bits_burst;
  wire [3:0] _T_584_bits_id;
  wire [30:0] _T_584_bits_addr;
  wire [7:0] _T_584_bits_len;
  wire [59:0] _T_830;
  wire [59:0] _T_831;
  wire [2:0] _T_590_bits_prot;
  wire [3:0] _T_590_bits_qos;
  wire  _T_590_bits_lock;
  wire [3:0] _T_590_bits_cache;
  wire [2:0] _T_590_bits_size;
  wire [1:0] _T_590_bits_burst;
  wire [3:0] _T_590_bits_id;
  wire [30:0] _T_590_bits_addr;
  wire [7:0] _T_590_bits_len;
  wire [59:0] _T_839;
  wire [59:0] _T_840;
  wire [2:0] _T_596_bits_prot;
  wire [3:0] _T_596_bits_qos;
  wire  _T_596_bits_lock;
  wire [3:0] _T_596_bits_cache;
  wire [2:0] _T_596_bits_size;
  wire [1:0] _T_596_bits_burst;
  wire [3:0] _T_596_bits_id;
  wire [30:0] _T_596_bits_addr;
  wire [7:0] _T_596_bits_len;
  wire [59:0] _T_848;
  wire [59:0] _T_849;
  wire [2:0] _T_602_bits_prot;
  wire [3:0] _T_602_bits_qos;
  wire  _T_602_bits_lock;
  wire [3:0] _T_602_bits_cache;
  wire [2:0] _T_602_bits_size;
  wire [1:0] _T_602_bits_burst;
  wire [3:0] _T_602_bits_id;
  wire [30:0] _T_602_bits_addr;
  wire [7:0] _T_602_bits_len;
  wire [59:0] _T_857;
  wire [59:0] _T_858;
  wire [2:0] _T_608_bits_prot;
  wire [3:0] _T_608_bits_qos;
  wire  _T_608_bits_lock;
  wire [3:0] _T_608_bits_cache;
  wire [2:0] _T_608_bits_size;
  wire [1:0] _T_608_bits_burst;
  wire [3:0] _T_608_bits_id;
  wire [30:0] _T_608_bits_addr;
  wire [7:0] _T_608_bits_len;
  wire [59:0] _T_866;
  wire [59:0] _T_867;
  wire [59:0] _T_868;
  wire [59:0] _T_869;
  wire [59:0] _T_870;
  wire [59:0] _T_871;
  wire [59:0] _T_872;
  wire [59:0] _T_873;
  wire [59:0] _T_874;
  wire  _T_888;
  reg [31:0] _T_889;
  reg [31:0] _RAND_22;
  wire [31:0] _T_891;
  wire [7:0] _T_898;
  wire [15:0] _T_906;
  wire  _T_907;
  wire  _T_908;
  wire  _T_909;
  wire  _T_910;
  wire  _T_911;
  wire  _T_912;
  wire  _T_913;
  wire  _T_914;
  wire  _T_915;
  wire  _T_916;
  wire  _T_917;
  wire  _T_918;
  wire  _T_919;
  wire  _T_920;
  wire  _T_921;
  wire  _T_922;
  wire [7:0] _T_930;
  wire [15:0] _T_938;
  wire [2:0] _GEN_107;
  wire [2:0] _GEN_108;
  wire [2:0] _GEN_109;
  wire [2:0] _GEN_110;
  wire [2:0] _GEN_111;
  wire [2:0] _GEN_112;
  wire [2:0] _GEN_113;
  wire [2:0] _GEN_114;
  wire [2:0] _GEN_115;
  wire [2:0] _GEN_116;
  wire [2:0] _GEN_117;
  wire [2:0] _GEN_118;
  wire [2:0] _GEN_119;
  wire [2:0] _GEN_120;
  wire [2:0] _GEN_121;
  wire  _T_950_7;
  wire  _T_950_6;
  wire  _T_950_5;
  wire  _T_950_4;
  wire  _T_950_3;
  wire  _T_950_2;
  wire  _T_950_1;
  wire  _T_950_0;
  wire  _GEN_123;
  wire  _GEN_124;
  wire  _GEN_125;
  wire  _GEN_126;
  wire  _GEN_127;
  wire  _GEN_128;
  wire [31:0] _T_946;
  wire [1:0] _T_947;
  wire [31:0] _GEN_166;
  wire [7:0] _T_952;
  wire  _T_954;
  wire  _T_955;
  wire  _T_956;
  wire  _T_957;
  wire  _T_958;
  wire  _T_959;
  wire  _T_960;
  wire  _T_961;
  wire  _T_972;
  wire  _T_973;
  wire  _T_974;
  wire  _T_970_ready;
  reg  _T_1019;
  reg [31:0] _RAND_23;
  wire  _T_1020;
  wire  _T_1014;
  wire  _T_1015;
  wire  _T_1016;
  wire  _T_1008;
  wire  _T_1009;
  wire  _T_1010;
  wire  _T_1002;
  wire  _T_1003;
  wire  _T_1004;
  wire  _T_996;
  wire  _T_997;
  wire  _T_998;
  wire  _T_990;
  wire  _T_991;
  wire  _T_992;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire  _T_978;
  wire  _T_979;
  wire  _T_980;
  wire [7:0] _T_1028;
  reg [7:0] _T_1035;
  reg [31:0] _RAND_24;
  wire [7:0] _T_1036;
  wire [7:0] _T_1037;
  wire [15:0] _T_1038;
  wire [14:0] _T_1039;
  wire [15:0] _GEN_167;
  wire [15:0] _T_1040;
  wire [13:0] _T_1041;
  wire [15:0] _GEN_168;
  wire [15:0] _T_1042;
  wire [11:0] _T_1043;
  wire [15:0] _GEN_169;
  wire [15:0] _T_1044;
  wire [14:0] _T_1046;
  wire [15:0] _T_1047;
  wire [15:0] _GEN_170;
  wire [15:0] _T_1048;
  wire [7:0] _T_1049;
  wire [7:0] _T_1050;
  wire [7:0] _T_1051;
  wire [7:0] _T_1052;
  wire  _T_1067;
  reg  _T_1166_0;
  reg [31:0] _RAND_25;
  wire  _T_1168_0;
  wire  _T_1169;
  wire  _T_1068;
  reg  _T_1166_1;
  reg [31:0] _RAND_26;
  wire  _T_1168_1;
  wire  _T_1170;
  wire  _T_1069;
  reg  _T_1166_2;
  reg [31:0] _RAND_27;
  wire  _T_1168_2;
  wire  _T_1171;
  wire  _T_1070;
  reg  _T_1166_3;
  reg [31:0] _RAND_28;
  wire  _T_1168_3;
  wire  _T_1172;
  wire  _T_1071;
  reg  _T_1166_4;
  reg [31:0] _RAND_29;
  wire  _T_1168_4;
  wire  _T_1173;
  wire  _T_1072;
  reg  _T_1166_5;
  reg [31:0] _RAND_30;
  wire  _T_1168_5;
  wire  _T_1174;
  wire  _T_1073;
  reg  _T_1166_6;
  reg [31:0] _RAND_31;
  wire  _T_1168_6;
  wire  _T_1175;
  wire  _T_1074;
  reg  _T_1166_7;
  reg [31:0] _RAND_32;
  wire  _T_1168_7;
  wire  _T_1176;
  wire  _T_1021;
  wire  _T_1030;
  wire  _T_1032;
  wire  _T_1033;
  wire  _T_1053;
  wire  _T_1054;
  wire [7:0] _T_1055;
  wire [8:0] _T_1056;
  wire [7:0] _T_1057;
  wire [7:0] _T_1058;
  wire [9:0] _T_1059;
  wire [7:0] _T_1060;
  wire [7:0] _T_1061;
  wire [11:0] _T_1062;
  wire [7:0] _T_1063;
  wire [7:0] _T_1064;
  wire  _T_1076;
  wire  _T_1077;
  wire  _T_1078;
  wire  _T_1079;
  wire  _T_1080;
  wire  _T_1081;
  wire  _T_1082;
  wire  _T_1083;
  wire  _T_1086;
  wire  _T_1087;
  wire  _T_1088;
  wire  _T_1089;
  wire  _T_1090;
  wire  _T_1091;
  wire  _T_1092;
  wire  _T_1094;
  wire  _T_1097;
  wire  _T_1098;
  wire  _T_1099;
  wire  _T_1100;
  wire  _T_1101;
  wire  _T_1102;
  wire  _T_1103;
  wire  _T_1104;
  wire  _T_1105;
  wire  _T_1106;
  wire  _T_1107;
  wire  _T_1108;
  wire  _T_1109;
  wire  _T_1110;
  wire  _T_1111;
  wire  _T_1112;
  wire  _T_1113;
  wire  _T_1114;
  wire  _T_1115;
  wire  _T_1116;
  wire  _T_1118;
  wire  _T_1119;
  wire  _T_1120;
  wire  _T_1121;
  wire  _T_1122;
  wire  _T_1123;
  wire  _T_1125;
  wire  _T_1126;
  wire  _T_1127;
  wire  _T_1128;
  wire  _T_1129;
  wire  _T_1130;
  wire  _T_1131;
  wire  _T_1132;
  wire  _T_1133;
  wire  _T_1134;
  wire  _T_1142;
  wire  _T_1144;
  wire  _T_1145;
  wire  _T_1184;
  wire  _T_1185;
  wire  _T_1192;
  wire  _T_1186;
  wire  _T_1193;
  wire  _T_1187;
  wire  _T_1194;
  wire  _T_1188;
  wire  _T_1195;
  wire  _T_1189;
  wire  _T_1196;
  wire  _T_1190;
  wire  _T_1197;
  wire  _T_1191;
  wire  _T_1198;
  wire  _T_1200;
  wire  _T_1161;
  wire  _T_1163;
  wire  _T_1167_0;
  wire  _T_1167_1;
  wire  _T_1167_2;
  wire  _T_1167_3;
  wire  _T_1167_4;
  wire  _T_1167_5;
  wire  _T_1167_6;
  wire  _T_1167_7;
  wire [3:0] _T_971_bits_id;
  wire [1:0] _T_971_bits_resp;
  wire [5:0] _T_1201;
  wire [5:0] _T_1202;
  wire [3:0] _T_977_bits_id;
  wire [1:0] _T_977_bits_resp;
  wire [5:0] _T_1203;
  wire [5:0] _T_1204;
  wire [3:0] _T_983_bits_id;
  wire [1:0] _T_983_bits_resp;
  wire [5:0] _T_1205;
  wire [5:0] _T_1206;
  wire [3:0] _T_989_bits_id;
  wire [1:0] _T_989_bits_resp;
  wire [5:0] _T_1207;
  wire [5:0] _T_1208;
  wire [3:0] _T_995_bits_id;
  wire [1:0] _T_995_bits_resp;
  wire [5:0] _T_1209;
  wire [5:0] _T_1210;
  wire [3:0] _T_1001_bits_id;
  wire [1:0] _T_1001_bits_resp;
  wire [5:0] _T_1211;
  wire [5:0] _T_1212;
  wire [3:0] _T_1007_bits_id;
  wire [1:0] _T_1007_bits_resp;
  wire [5:0] _T_1213;
  wire [5:0] _T_1214;
  wire [3:0] _T_1013_bits_id;
  wire [1:0] _T_1013_bits_resp;
  wire [5:0] _T_1215;
  wire [5:0] _T_1216;
  wire [5:0] _T_1217;
  wire [5:0] _T_1218;
  wire [5:0] _T_1219;
  wire [5:0] _T_1220;
  wire [5:0] _T_1221;
  wire [5:0] _T_1222;
  wire [5:0] _T_1223;
  wire  _T_1230;
  reg [31:0] _T_1231;
  reg [31:0] _RAND_33;
  wire [31:0] _T_1233;
  wire [7:0] _T_1240;
  wire [15:0] _T_1248;
  wire  _T_1249;
  wire  _T_1250;
  wire  _T_1251;
  wire  _T_1252;
  wire  _T_1253;
  wire  _T_1254;
  wire  _T_1255;
  wire  _T_1256;
  wire  _T_1257;
  wire  _T_1258;
  wire  _T_1259;
  wire  _T_1260;
  wire  _T_1261;
  wire  _T_1262;
  wire  _T_1263;
  wire  _T_1264;
  wire [7:0] _T_1272;
  wire [15:0] _T_1280;
  wire [2:0] _GEN_132;
  wire [2:0] _GEN_133;
  wire [2:0] _GEN_134;
  wire [2:0] _GEN_135;
  wire [2:0] _GEN_136;
  wire [2:0] _GEN_137;
  wire [2:0] _GEN_138;
  wire [2:0] _GEN_139;
  wire [2:0] _GEN_140;
  wire [2:0] _GEN_141;
  wire [2:0] _GEN_142;
  wire [2:0] _GEN_143;
  wire [2:0] _GEN_144;
  wire [2:0] _GEN_145;
  wire [2:0] _GEN_146;
  wire  _T_1292_7;
  wire  _T_1292_6;
  wire  _T_1292_5;
  wire  _T_1292_4;
  wire  _T_1292_3;
  wire  _T_1292_2;
  wire  _T_1292_1;
  wire  _T_1292_0;
  wire  _GEN_148;
  wire  _GEN_149;
  wire  _GEN_150;
  wire  _GEN_151;
  wire  _GEN_152;
  wire  _GEN_153;
  wire [31:0] _T_1288;
  wire [1:0] _T_1289;
  wire [31:0] _GEN_171;
  wire [7:0] _T_1294;
  wire  _T_1296;
  wire  _T_1297;
  wire  _T_1298;
  wire  _T_1299;
  wire  _T_1300;
  wire  _T_1301;
  wire  _T_1302;
  wire  _T_1303;
  wire  _T_1314;
  wire  _T_1315;
  wire  _T_1316;
  wire  _T_1312_ready;
  reg  _T_1361;
  reg [31:0] _RAND_34;
  wire  _T_1362;
  wire  _T_1356;
  wire  _T_1357;
  wire  _T_1358;
  wire  _T_1350;
  wire  _T_1351;
  wire  _T_1352;
  wire  _T_1344;
  wire  _T_1345;
  wire  _T_1346;
  wire  _T_1338;
  wire  _T_1339;
  wire  _T_1340;
  wire  _T_1332;
  wire  _T_1333;
  wire  _T_1334;
  wire  _T_1326;
  wire  _T_1327;
  wire  _T_1328;
  wire  _T_1320;
  wire  _T_1321;
  wire  _T_1322;
  wire [7:0] _T_1370;
  reg [7:0] _T_1377;
  reg [31:0] _RAND_35;
  wire [7:0] _T_1378;
  wire [7:0] _T_1379;
  wire [15:0] _T_1380;
  wire [14:0] _T_1381;
  wire [15:0] _GEN_172;
  wire [15:0] _T_1382;
  wire [13:0] _T_1383;
  wire [15:0] _GEN_173;
  wire [15:0] _T_1384;
  wire [11:0] _T_1385;
  wire [15:0] _GEN_174;
  wire [15:0] _T_1386;
  wire [14:0] _T_1388;
  wire [15:0] _T_1389;
  wire [15:0] _GEN_175;
  wire [15:0] _T_1390;
  wire [7:0] _T_1391;
  wire [7:0] _T_1392;
  wire [7:0] _T_1393;
  wire [7:0] _T_1394;
  wire  _T_1409;
  reg  _T_1508_0;
  reg [31:0] _RAND_36;
  wire  _T_1510_0;
  wire  _T_1511;
  wire  _T_1410;
  reg  _T_1508_1;
  reg [31:0] _RAND_37;
  wire  _T_1510_1;
  wire  _T_1512;
  wire  _T_1411;
  reg  _T_1508_2;
  reg [31:0] _RAND_38;
  wire  _T_1510_2;
  wire  _T_1513;
  wire  _T_1412;
  reg  _T_1508_3;
  reg [31:0] _RAND_39;
  wire  _T_1510_3;
  wire  _T_1514;
  wire  _T_1413;
  reg  _T_1508_4;
  reg [31:0] _RAND_40;
  wire  _T_1510_4;
  wire  _T_1515;
  wire  _T_1414;
  reg  _T_1508_5;
  reg [31:0] _RAND_41;
  wire  _T_1510_5;
  wire  _T_1516;
  wire  _T_1415;
  reg  _T_1508_6;
  reg [31:0] _RAND_42;
  wire  _T_1510_6;
  wire  _T_1517;
  wire  _T_1416;
  reg  _T_1508_7;
  reg [31:0] _RAND_43;
  wire  _T_1510_7;
  wire  _T_1518;
  wire  _T_1363;
  wire  _T_1372;
  wire  _T_1374;
  wire  _T_1375;
  wire  _T_1395;
  wire  _T_1396;
  wire [7:0] _T_1397;
  wire [8:0] _T_1398;
  wire [7:0] _T_1399;
  wire [7:0] _T_1400;
  wire [9:0] _T_1401;
  wire [7:0] _T_1402;
  wire [7:0] _T_1403;
  wire [11:0] _T_1404;
  wire [7:0] _T_1405;
  wire [7:0] _T_1406;
  wire  _T_1418;
  wire  _T_1419;
  wire  _T_1420;
  wire  _T_1421;
  wire  _T_1422;
  wire  _T_1423;
  wire  _T_1424;
  wire  _T_1425;
  wire  _T_1428;
  wire  _T_1429;
  wire  _T_1430;
  wire  _T_1431;
  wire  _T_1432;
  wire  _T_1433;
  wire  _T_1434;
  wire  _T_1436;
  wire  _T_1439;
  wire  _T_1440;
  wire  _T_1441;
  wire  _T_1442;
  wire  _T_1443;
  wire  _T_1444;
  wire  _T_1445;
  wire  _T_1446;
  wire  _T_1447;
  wire  _T_1448;
  wire  _T_1449;
  wire  _T_1450;
  wire  _T_1451;
  wire  _T_1452;
  wire  _T_1453;
  wire  _T_1454;
  wire  _T_1455;
  wire  _T_1456;
  wire  _T_1457;
  wire  _T_1458;
  wire  _T_1460;
  wire  _T_1461;
  wire  _T_1462;
  wire  _T_1463;
  wire  _T_1464;
  wire  _T_1465;
  wire  _T_1467;
  wire  _T_1468;
  wire  _T_1469;
  wire  _T_1470;
  wire  _T_1471;
  wire  _T_1472;
  wire  _T_1473;
  wire  _T_1474;
  wire  _T_1475;
  wire  _T_1476;
  wire  _T_1484;
  wire  _T_1486;
  wire  _T_1487;
  wire  _T_1526;
  wire  _T_1527;
  wire  _T_1534;
  wire  _T_1528;
  wire  _T_1535;
  wire  _T_1529;
  wire  _T_1536;
  wire  _T_1530;
  wire  _T_1537;
  wire  _T_1531;
  wire  _T_1538;
  wire  _T_1532;
  wire  _T_1539;
  wire  _T_1533;
  wire  _T_1540;
  wire  _T_1542;
  wire  _T_1503;
  wire  _T_1505;
  wire  _T_1509_0;
  wire  _T_1509_1;
  wire  _T_1509_2;
  wire  _T_1509_3;
  wire  _T_1509_4;
  wire  _T_1509_5;
  wire  _T_1509_6;
  wire  _T_1509_7;
  wire [1:0] _T_1313_bits_resp;
  wire  _T_1313_bits_last;
  wire [3:0] _T_1313_bits_id;
  wire [31:0] _T_1313_bits_data;
  wire [38:0] _T_1545;
  wire [38:0] _T_1546;
  wire [1:0] _T_1319_bits_resp;
  wire  _T_1319_bits_last;
  wire [3:0] _T_1319_bits_id;
  wire [31:0] _T_1319_bits_data;
  wire [38:0] _T_1549;
  wire [38:0] _T_1550;
  wire [1:0] _T_1325_bits_resp;
  wire  _T_1325_bits_last;
  wire [3:0] _T_1325_bits_id;
  wire [31:0] _T_1325_bits_data;
  wire [38:0] _T_1553;
  wire [38:0] _T_1554;
  wire [1:0] _T_1331_bits_resp;
  wire  _T_1331_bits_last;
  wire [3:0] _T_1331_bits_id;
  wire [31:0] _T_1331_bits_data;
  wire [38:0] _T_1557;
  wire [38:0] _T_1558;
  wire [1:0] _T_1337_bits_resp;
  wire  _T_1337_bits_last;
  wire [3:0] _T_1337_bits_id;
  wire [31:0] _T_1337_bits_data;
  wire [38:0] _T_1561;
  wire [38:0] _T_1562;
  wire [1:0] _T_1343_bits_resp;
  wire  _T_1343_bits_last;
  wire [3:0] _T_1343_bits_id;
  wire [31:0] _T_1343_bits_data;
  wire [38:0] _T_1565;
  wire [38:0] _T_1566;
  wire [1:0] _T_1349_bits_resp;
  wire  _T_1349_bits_last;
  wire [3:0] _T_1349_bits_id;
  wire [31:0] _T_1349_bits_data;
  wire [38:0] _T_1569;
  wire [38:0] _T_1570;
  wire [1:0] _T_1355_bits_resp;
  wire  _T_1355_bits_last;
  wire [3:0] _T_1355_bits_id;
  wire [31:0] _T_1355_bits_data;
  wire [38:0] _T_1573;
  wire [38:0] _T_1574;
  wire [38:0] _T_1575;
  wire [38:0] _T_1576;
  wire [38:0] _T_1577;
  wire [38:0] _T_1578;
  wire [38:0] _T_1579;
  wire [38:0] _T_1580;
  wire [38:0] _T_1581;
  Queue_107 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR (
    ._EVAL(MaxPeriodFibonacciLFSR__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR__EVAL_17)
  );
  Queue_108 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data_id(Queue_1_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_1_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_1_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_1_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_1_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_1_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_1_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_1_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_1_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_1_io_enq_bits_timestamp),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data_id(Queue_1_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_1_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_1_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_1_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_1_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_1_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_1_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_1_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_1_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_1_io_deq_bits_timestamp)
  );
  Queue_108 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data_id(Queue_2_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_2_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_2_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_2_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_2_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_2_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_2_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_2_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_2_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_2_io_enq_bits_timestamp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data_id(Queue_2_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_2_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_2_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_2_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_2_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_2_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_2_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_2_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_2_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_2_io_deq_bits_timestamp)
  );
  Queue_108 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_data_id(Queue_3_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_3_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_3_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_3_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_3_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_3_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_3_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_3_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_3_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_3_io_enq_bits_timestamp),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_data_id(Queue_3_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_3_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_3_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_3_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_3_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_3_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_3_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_3_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_3_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_3_io_deq_bits_timestamp)
  );
  Queue_108 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_data_id(Queue_4_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_4_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_4_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_4_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_4_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_4_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_4_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_4_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_4_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_4_io_enq_bits_timestamp),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_data_id(Queue_4_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_4_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_4_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_4_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_4_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_4_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_4_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_4_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_4_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_4_io_deq_bits_timestamp)
  );
  Queue_108 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_data_id(Queue_5_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_5_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_5_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_5_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_5_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_5_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_5_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_5_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_5_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_5_io_enq_bits_timestamp),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_data_id(Queue_5_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_5_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_5_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_5_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_5_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_5_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_5_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_5_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_5_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_5_io_deq_bits_timestamp)
  );
  Queue_108 Queue_6 (
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits_data_id(Queue_6_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_6_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_6_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_6_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_6_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_6_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_6_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_6_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_6_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_6_io_enq_bits_timestamp),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits_data_id(Queue_6_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_6_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_6_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_6_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_6_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_6_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_6_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_6_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_6_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_6_io_deq_bits_timestamp)
  );
  Queue_108 Queue_7 (
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits_data_id(Queue_7_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_7_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_7_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_7_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_7_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_7_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_7_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_7_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_7_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_7_io_enq_bits_timestamp),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits_data_id(Queue_7_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_7_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_7_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_7_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_7_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_7_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_7_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_7_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_7_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_7_io_deq_bits_timestamp)
  );
  Queue_108 Queue_8 (
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits_data_id(Queue_8_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_8_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_8_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_8_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_8_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_8_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_8_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_8_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_8_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_8_io_enq_bits_timestamp),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits_data_id(Queue_8_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_8_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_8_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_8_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_8_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_8_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_8_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_8_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_8_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_8_io_deq_bits_timestamp)
  );
  Queue_116 Queue_9 (
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits_id(Queue_9_io_enq_bits_id),
    .io_enq_bits_addr(Queue_9_io_enq_bits_addr),
    .io_enq_bits_len(Queue_9_io_enq_bits_len),
    .io_enq_bits_size(Queue_9_io_enq_bits_size),
    .io_enq_bits_burst(Queue_9_io_enq_bits_burst),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits_id(Queue_9_io_deq_bits_id),
    .io_deq_bits_addr(Queue_9_io_deq_bits_addr),
    .io_deq_bits_len(Queue_9_io_deq_bits_len),
    .io_deq_bits_size(Queue_9_io_deq_bits_size),
    .io_deq_bits_burst(Queue_9_io_deq_bits_burst)
  );
  Queue_107 Queue_10 (
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits(Queue_10_io_enq_bits),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits(Queue_10_io_deq_bits)
  );
  Queue_116 Queue_11 (
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits_id(Queue_11_io_enq_bits_id),
    .io_enq_bits_addr(Queue_11_io_enq_bits_addr),
    .io_enq_bits_len(Queue_11_io_enq_bits_len),
    .io_enq_bits_size(Queue_11_io_enq_bits_size),
    .io_enq_bits_burst(Queue_11_io_enq_bits_burst),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits_id(Queue_11_io_deq_bits_id),
    .io_deq_bits_addr(Queue_11_io_deq_bits_addr),
    .io_deq_bits_len(Queue_11_io_deq_bits_len),
    .io_deq_bits_size(Queue_11_io_deq_bits_size),
    .io_deq_bits_burst(Queue_11_io_deq_bits_burst)
  );
  Queue_119 Queue_12 (
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits_data(Queue_12_io_enq_bits_data),
    .io_enq_bits_strb(Queue_12_io_enq_bits_strb),
    .io_enq_bits_last(Queue_12_io_enq_bits_last),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits_data(Queue_12_io_deq_bits_data),
    .io_deq_bits_strb(Queue_12_io_deq_bits_strb),
    .io_deq_bits_last(Queue_12_io_deq_bits_last)
  );
  Queue_119 Queue_13 (
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits_data(Queue_13_io_enq_bits_data),
    .io_enq_bits_strb(Queue_13_io_enq_bits_strb),
    .io_enq_bits_last(Queue_13_io_enq_bits_last),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits_data(Queue_13_io_deq_bits_data),
    .io_deq_bits_strb(Queue_13_io_deq_bits_strb),
    .io_deq_bits_last(Queue_13_io_deq_bits_last)
  );
  Queue_119 Queue_14 (
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits_data(Queue_14_io_enq_bits_data),
    .io_enq_bits_strb(Queue_14_io_enq_bits_strb),
    .io_enq_bits_last(Queue_14_io_enq_bits_last),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits_data(Queue_14_io_deq_bits_data),
    .io_deq_bits_strb(Queue_14_io_deq_bits_strb),
    .io_deq_bits_last(Queue_14_io_deq_bits_last)
  );
  Queue_119 Queue_15 (
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits_data(Queue_15_io_enq_bits_data),
    .io_enq_bits_strb(Queue_15_io_enq_bits_strb),
    .io_enq_bits_last(Queue_15_io_enq_bits_last),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits_data(Queue_15_io_deq_bits_data),
    .io_deq_bits_strb(Queue_15_io_deq_bits_strb),
    .io_deq_bits_last(Queue_15_io_deq_bits_last)
  );
  Queue_119 Queue_16 (
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits_data(Queue_16_io_enq_bits_data),
    .io_enq_bits_strb(Queue_16_io_enq_bits_strb),
    .io_enq_bits_last(Queue_16_io_enq_bits_last),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits_data(Queue_16_io_deq_bits_data),
    .io_deq_bits_strb(Queue_16_io_deq_bits_strb),
    .io_deq_bits_last(Queue_16_io_deq_bits_last)
  );
  Queue_119 Queue_17 (
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits_data(Queue_17_io_enq_bits_data),
    .io_enq_bits_strb(Queue_17_io_enq_bits_strb),
    .io_enq_bits_last(Queue_17_io_enq_bits_last),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits_data(Queue_17_io_deq_bits_data),
    .io_deq_bits_strb(Queue_17_io_deq_bits_strb),
    .io_deq_bits_last(Queue_17_io_deq_bits_last)
  );
  Queue_119 Queue_18 (
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits_data(Queue_18_io_enq_bits_data),
    .io_enq_bits_strb(Queue_18_io_enq_bits_strb),
    .io_enq_bits_last(Queue_18_io_enq_bits_last),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits_data(Queue_18_io_deq_bits_data),
    .io_deq_bits_strb(Queue_18_io_deq_bits_strb),
    .io_deq_bits_last(Queue_18_io_deq_bits_last)
  );
  Queue_119 Queue_19 (
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits_data(Queue_19_io_enq_bits_data),
    .io_enq_bits_strb(Queue_19_io_enq_bits_strb),
    .io_enq_bits_last(Queue_19_io_enq_bits_last),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits_data(Queue_19_io_deq_bits_data),
    .io_deq_bits_strb(Queue_19_io_deq_bits_strb),
    .io_deq_bits_last(Queue_19_io_deq_bits_last)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 (
    .out(plusarg_reader_1_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_1 (
    ._EVAL(MaxPeriodFibonacciLFSR_1__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_1__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_1__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_1__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_1__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_1__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_1__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_1__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_1__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_1__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_1__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_1__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_1__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_1__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_1__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_1__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_1__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_1__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_1__EVAL_17)
  );
  Queue_108 Queue_20 (
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits_data_id(Queue_20_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_20_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_20_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_20_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_20_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_20_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_20_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_20_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_20_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_20_io_enq_bits_timestamp),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits_data_id(Queue_20_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_20_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_20_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_20_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_20_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_20_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_20_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_20_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_20_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_20_io_deq_bits_timestamp)
  );
  Queue_108 Queue_21 (
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits_data_id(Queue_21_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_21_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_21_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_21_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_21_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_21_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_21_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_21_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_21_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_21_io_enq_bits_timestamp),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits_data_id(Queue_21_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_21_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_21_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_21_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_21_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_21_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_21_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_21_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_21_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_21_io_deq_bits_timestamp)
  );
  Queue_108 Queue_22 (
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits_data_id(Queue_22_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_22_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_22_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_22_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_22_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_22_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_22_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_22_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_22_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_22_io_enq_bits_timestamp),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits_data_id(Queue_22_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_22_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_22_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_22_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_22_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_22_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_22_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_22_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_22_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_22_io_deq_bits_timestamp)
  );
  Queue_108 Queue_23 (
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits_data_id(Queue_23_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_23_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_23_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_23_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_23_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_23_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_23_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_23_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_23_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_23_io_enq_bits_timestamp),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits_data_id(Queue_23_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_23_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_23_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_23_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_23_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_23_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_23_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_23_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_23_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_23_io_deq_bits_timestamp)
  );
  Queue_108 Queue_24 (
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits_data_id(Queue_24_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_24_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_24_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_24_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_24_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_24_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_24_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_24_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_24_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_24_io_enq_bits_timestamp),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits_data_id(Queue_24_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_24_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_24_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_24_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_24_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_24_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_24_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_24_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_24_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_24_io_deq_bits_timestamp)
  );
  Queue_108 Queue_25 (
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits_data_id(Queue_25_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_25_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_25_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_25_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_25_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_25_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_25_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_25_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_25_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_25_io_enq_bits_timestamp),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits_data_id(Queue_25_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_25_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_25_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_25_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_25_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_25_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_25_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_25_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_25_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_25_io_deq_bits_timestamp)
  );
  Queue_108 Queue_26 (
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits_data_id(Queue_26_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_26_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_26_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_26_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_26_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_26_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_26_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_26_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_26_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_26_io_enq_bits_timestamp),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits_data_id(Queue_26_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_26_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_26_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_26_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_26_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_26_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_26_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_26_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_26_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_26_io_deq_bits_timestamp)
  );
  Queue_108 Queue_27 (
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits_data_id(Queue_27_io_enq_bits_data_id),
    .io_enq_bits_data_addr(Queue_27_io_enq_bits_data_addr),
    .io_enq_bits_data_len(Queue_27_io_enq_bits_data_len),
    .io_enq_bits_data_size(Queue_27_io_enq_bits_data_size),
    .io_enq_bits_data_burst(Queue_27_io_enq_bits_data_burst),
    .io_enq_bits_data_lock(Queue_27_io_enq_bits_data_lock),
    .io_enq_bits_data_cache(Queue_27_io_enq_bits_data_cache),
    .io_enq_bits_data_prot(Queue_27_io_enq_bits_data_prot),
    .io_enq_bits_data_qos(Queue_27_io_enq_bits_data_qos),
    .io_enq_bits_timestamp(Queue_27_io_enq_bits_timestamp),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits_data_id(Queue_27_io_deq_bits_data_id),
    .io_deq_bits_data_addr(Queue_27_io_deq_bits_data_addr),
    .io_deq_bits_data_len(Queue_27_io_deq_bits_data_len),
    .io_deq_bits_data_size(Queue_27_io_deq_bits_data_size),
    .io_deq_bits_data_burst(Queue_27_io_deq_bits_data_burst),
    .io_deq_bits_data_lock(Queue_27_io_deq_bits_data_lock),
    .io_deq_bits_data_cache(Queue_27_io_deq_bits_data_cache),
    .io_deq_bits_data_prot(Queue_27_io_deq_bits_data_prot),
    .io_deq_bits_data_qos(Queue_27_io_deq_bits_data_qos),
    .io_deq_bits_timestamp(Queue_27_io_deq_bits_timestamp)
  );
  Queue_116 Queue_28 (
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits_id(Queue_28_io_enq_bits_id),
    .io_enq_bits_addr(Queue_28_io_enq_bits_addr),
    .io_enq_bits_len(Queue_28_io_enq_bits_len),
    .io_enq_bits_size(Queue_28_io_enq_bits_size),
    .io_enq_bits_burst(Queue_28_io_enq_bits_burst),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits_id(Queue_28_io_deq_bits_id),
    .io_deq_bits_addr(Queue_28_io_deq_bits_addr),
    .io_deq_bits_len(Queue_28_io_deq_bits_len),
    .io_deq_bits_size(Queue_28_io_deq_bits_size),
    .io_deq_bits_burst(Queue_28_io_deq_bits_burst)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_2 (
    .out(plusarg_reader_2_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_2 (
    ._EVAL(MaxPeriodFibonacciLFSR_2__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_2__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_2__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_2__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_2__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_2__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_2__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_2__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_2__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_2__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_2__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_2__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_2__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_2__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_2__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_2__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_2__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_2__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_2__EVAL_17)
  );
  Queue_136 Queue_29 (
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits_data_id(Queue_29_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_29_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_29_io_enq_bits_timestamp),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits_data_id(Queue_29_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_29_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_29_io_deq_bits_timestamp)
  );
  Queue_136 Queue_30 (
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits_data_id(Queue_30_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_30_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_30_io_enq_bits_timestamp),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits_data_id(Queue_30_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_30_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_30_io_deq_bits_timestamp)
  );
  Queue_136 Queue_31 (
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits_data_id(Queue_31_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_31_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_31_io_enq_bits_timestamp),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits_data_id(Queue_31_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_31_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_31_io_deq_bits_timestamp)
  );
  Queue_136 Queue_32 (
    .clock(Queue_32_clock),
    .reset(Queue_32_reset),
    .io_enq_ready(Queue_32_io_enq_ready),
    .io_enq_valid(Queue_32_io_enq_valid),
    .io_enq_bits_data_id(Queue_32_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_32_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_32_io_enq_bits_timestamp),
    .io_deq_ready(Queue_32_io_deq_ready),
    .io_deq_valid(Queue_32_io_deq_valid),
    .io_deq_bits_data_id(Queue_32_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_32_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_32_io_deq_bits_timestamp)
  );
  Queue_136 Queue_33 (
    .clock(Queue_33_clock),
    .reset(Queue_33_reset),
    .io_enq_ready(Queue_33_io_enq_ready),
    .io_enq_valid(Queue_33_io_enq_valid),
    .io_enq_bits_data_id(Queue_33_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_33_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_33_io_enq_bits_timestamp),
    .io_deq_ready(Queue_33_io_deq_ready),
    .io_deq_valid(Queue_33_io_deq_valid),
    .io_deq_bits_data_id(Queue_33_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_33_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_33_io_deq_bits_timestamp)
  );
  Queue_136 Queue_34 (
    .clock(Queue_34_clock),
    .reset(Queue_34_reset),
    .io_enq_ready(Queue_34_io_enq_ready),
    .io_enq_valid(Queue_34_io_enq_valid),
    .io_enq_bits_data_id(Queue_34_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_34_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_34_io_enq_bits_timestamp),
    .io_deq_ready(Queue_34_io_deq_ready),
    .io_deq_valid(Queue_34_io_deq_valid),
    .io_deq_bits_data_id(Queue_34_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_34_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_34_io_deq_bits_timestamp)
  );
  Queue_136 Queue_35 (
    .clock(Queue_35_clock),
    .reset(Queue_35_reset),
    .io_enq_ready(Queue_35_io_enq_ready),
    .io_enq_valid(Queue_35_io_enq_valid),
    .io_enq_bits_data_id(Queue_35_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_35_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_35_io_enq_bits_timestamp),
    .io_deq_ready(Queue_35_io_deq_ready),
    .io_deq_valid(Queue_35_io_deq_valid),
    .io_deq_bits_data_id(Queue_35_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_35_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_35_io_deq_bits_timestamp)
  );
  Queue_136 Queue_36 (
    .clock(Queue_36_clock),
    .reset(Queue_36_reset),
    .io_enq_ready(Queue_36_io_enq_ready),
    .io_enq_valid(Queue_36_io_enq_valid),
    .io_enq_bits_data_id(Queue_36_io_enq_bits_data_id),
    .io_enq_bits_data_resp(Queue_36_io_enq_bits_data_resp),
    .io_enq_bits_timestamp(Queue_36_io_enq_bits_timestamp),
    .io_deq_ready(Queue_36_io_deq_ready),
    .io_deq_valid(Queue_36_io_deq_valid),
    .io_deq_bits_data_id(Queue_36_io_deq_bits_data_id),
    .io_deq_bits_data_resp(Queue_36_io_deq_bits_data_resp),
    .io_deq_bits_timestamp(Queue_36_io_deq_bits_timestamp)
  );
  Queue_144 Queue_37 (
    .clock(Queue_37_clock),
    .reset(Queue_37_reset),
    .io_enq_ready(Queue_37_io_enq_ready),
    .io_enq_valid(Queue_37_io_enq_valid),
    .io_enq_bits_id(Queue_37_io_enq_bits_id),
    .io_enq_bits_resp(Queue_37_io_enq_bits_resp),
    .io_deq_ready(Queue_37_io_deq_ready),
    .io_deq_valid(Queue_37_io_deq_valid),
    .io_deq_bits_id(Queue_37_io_deq_bits_id),
    .io_deq_bits_resp(Queue_37_io_deq_bits_resp)
  );
  plusarg_reader #(.FORMAT("disable_axi4_shuffling=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_3 (
    .out(plusarg_reader_3_out)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_3 (
    ._EVAL(MaxPeriodFibonacciLFSR_3__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_3__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_3__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_3__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_3__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_3__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_3__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_3__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_3__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_3__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_3__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_3__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_3__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_3__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_3__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_3__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_3__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_3__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_3__EVAL_17)
  );
  Queue_145 Queue_38 (
    .clock(Queue_38_clock),
    .reset(Queue_38_reset),
    .io_enq_ready(Queue_38_io_enq_ready),
    .io_enq_valid(Queue_38_io_enq_valid),
    .io_enq_bits_data_id(Queue_38_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_38_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_38_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_38_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_38_io_enq_bits_timestamp),
    .io_deq_ready(Queue_38_io_deq_ready),
    .io_deq_valid(Queue_38_io_deq_valid),
    .io_deq_bits_data_id(Queue_38_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_38_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_38_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_38_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_38_io_deq_bits_timestamp)
  );
  Queue_145 Queue_39 (
    .clock(Queue_39_clock),
    .reset(Queue_39_reset),
    .io_enq_ready(Queue_39_io_enq_ready),
    .io_enq_valid(Queue_39_io_enq_valid),
    .io_enq_bits_data_id(Queue_39_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_39_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_39_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_39_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_39_io_enq_bits_timestamp),
    .io_deq_ready(Queue_39_io_deq_ready),
    .io_deq_valid(Queue_39_io_deq_valid),
    .io_deq_bits_data_id(Queue_39_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_39_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_39_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_39_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_39_io_deq_bits_timestamp)
  );
  Queue_145 Queue_40 (
    .clock(Queue_40_clock),
    .reset(Queue_40_reset),
    .io_enq_ready(Queue_40_io_enq_ready),
    .io_enq_valid(Queue_40_io_enq_valid),
    .io_enq_bits_data_id(Queue_40_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_40_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_40_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_40_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_40_io_enq_bits_timestamp),
    .io_deq_ready(Queue_40_io_deq_ready),
    .io_deq_valid(Queue_40_io_deq_valid),
    .io_deq_bits_data_id(Queue_40_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_40_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_40_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_40_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_40_io_deq_bits_timestamp)
  );
  Queue_145 Queue_41 (
    .clock(Queue_41_clock),
    .reset(Queue_41_reset),
    .io_enq_ready(Queue_41_io_enq_ready),
    .io_enq_valid(Queue_41_io_enq_valid),
    .io_enq_bits_data_id(Queue_41_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_41_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_41_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_41_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_41_io_enq_bits_timestamp),
    .io_deq_ready(Queue_41_io_deq_ready),
    .io_deq_valid(Queue_41_io_deq_valid),
    .io_deq_bits_data_id(Queue_41_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_41_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_41_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_41_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_41_io_deq_bits_timestamp)
  );
  Queue_145 Queue_42 (
    .clock(Queue_42_clock),
    .reset(Queue_42_reset),
    .io_enq_ready(Queue_42_io_enq_ready),
    .io_enq_valid(Queue_42_io_enq_valid),
    .io_enq_bits_data_id(Queue_42_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_42_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_42_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_42_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_42_io_enq_bits_timestamp),
    .io_deq_ready(Queue_42_io_deq_ready),
    .io_deq_valid(Queue_42_io_deq_valid),
    .io_deq_bits_data_id(Queue_42_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_42_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_42_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_42_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_42_io_deq_bits_timestamp)
  );
  Queue_145 Queue_43 (
    .clock(Queue_43_clock),
    .reset(Queue_43_reset),
    .io_enq_ready(Queue_43_io_enq_ready),
    .io_enq_valid(Queue_43_io_enq_valid),
    .io_enq_bits_data_id(Queue_43_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_43_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_43_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_43_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_43_io_enq_bits_timestamp),
    .io_deq_ready(Queue_43_io_deq_ready),
    .io_deq_valid(Queue_43_io_deq_valid),
    .io_deq_bits_data_id(Queue_43_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_43_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_43_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_43_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_43_io_deq_bits_timestamp)
  );
  Queue_145 Queue_44 (
    .clock(Queue_44_clock),
    .reset(Queue_44_reset),
    .io_enq_ready(Queue_44_io_enq_ready),
    .io_enq_valid(Queue_44_io_enq_valid),
    .io_enq_bits_data_id(Queue_44_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_44_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_44_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_44_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_44_io_enq_bits_timestamp),
    .io_deq_ready(Queue_44_io_deq_ready),
    .io_deq_valid(Queue_44_io_deq_valid),
    .io_deq_bits_data_id(Queue_44_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_44_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_44_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_44_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_44_io_deq_bits_timestamp)
  );
  Queue_145 Queue_45 (
    .clock(Queue_45_clock),
    .reset(Queue_45_reset),
    .io_enq_ready(Queue_45_io_enq_ready),
    .io_enq_valid(Queue_45_io_enq_valid),
    .io_enq_bits_data_id(Queue_45_io_enq_bits_data_id),
    .io_enq_bits_data_data(Queue_45_io_enq_bits_data_data),
    .io_enq_bits_data_resp(Queue_45_io_enq_bits_data_resp),
    .io_enq_bits_data_last(Queue_45_io_enq_bits_data_last),
    .io_enq_bits_timestamp(Queue_45_io_enq_bits_timestamp),
    .io_deq_ready(Queue_45_io_deq_ready),
    .io_deq_valid(Queue_45_io_deq_valid),
    .io_deq_bits_data_id(Queue_45_io_deq_bits_data_id),
    .io_deq_bits_data_data(Queue_45_io_deq_bits_data_data),
    .io_deq_bits_data_resp(Queue_45_io_deq_bits_data_resp),
    .io_deq_bits_data_last(Queue_45_io_deq_bits_data_last),
    .io_deq_bits_timestamp(Queue_45_io_deq_bits_timestamp)
  );
  Queue_153 Queue_46 (
    .clock(Queue_46_clock),
    .reset(Queue_46_reset),
    .io_enq_ready(Queue_46_io_enq_ready),
    .io_enq_valid(Queue_46_io_enq_valid),
    .io_enq_bits_id(Queue_46_io_enq_bits_id),
    .io_enq_bits_data(Queue_46_io_enq_bits_data),
    .io_enq_bits_resp(Queue_46_io_enq_bits_resp),
    .io_enq_bits_last(Queue_46_io_enq_bits_last),
    .io_deq_ready(Queue_46_io_deq_ready),
    .io_deq_valid(Queue_46_io_deq_valid),
    .io_deq_bits_id(Queue_46_io_deq_bits_id),
    .io_deq_bits_data(Queue_46_io_deq_bits_data),
    .io_deq_bits_resp(Queue_46_io_deq_bits_resp),
    .io_deq_bits_last(Queue_46_io_deq_bits_last)
  );
  assign _GEN_1 = 4'h1 == auto_in_aw_bits_id ? 3'h0 : 3'h5;
  assign _GEN_2 = 4'h2 == auto_in_aw_bits_id ? 3'h5 : _GEN_1;
  assign _GEN_3 = 4'h3 == auto_in_aw_bits_id ? 3'h0 : _GEN_2;
  assign _GEN_4 = 4'h4 == auto_in_aw_bits_id ? 3'h2 : _GEN_3;
  assign _GEN_5 = 4'h5 == auto_in_aw_bits_id ? 3'h7 : _GEN_4;
  assign _GEN_6 = 4'h6 == auto_in_aw_bits_id ? 3'h2 : _GEN_5;
  assign _GEN_7 = 4'h7 == auto_in_aw_bits_id ? 3'h5 : _GEN_6;
  assign _GEN_8 = 4'h8 == auto_in_aw_bits_id ? 3'h5 : _GEN_7;
  assign _GEN_9 = 4'h9 == auto_in_aw_bits_id ? 3'h0 : _GEN_8;
  assign _GEN_10 = 4'ha == auto_in_aw_bits_id ? 3'h7 : _GEN_9;
  assign _GEN_11 = 4'hb == auto_in_aw_bits_id ? 3'h3 : _GEN_10;
  assign _GEN_12 = 4'hc == auto_in_aw_bits_id ? 3'h2 : _GEN_11;
  assign _GEN_13 = 4'hd == auto_in_aw_bits_id ? 3'h3 : _GEN_12;
  assign _GEN_14 = 4'he == auto_in_aw_bits_id ? 3'h2 : _GEN_13;
  assign _GEN_15 = 4'hf == auto_in_aw_bits_id ? 3'h5 : _GEN_14;
  assign _T_71_7 = Queue_8_io_enq_ready;
  assign _T_71_6 = Queue_7_io_enq_ready;
  assign _T_71_5 = Queue_6_io_enq_ready;
  assign _T_71_4 = Queue_5_io_enq_ready;
  assign _T_71_3 = Queue_4_io_enq_ready;
  assign _T_71_2 = Queue_3_io_enq_ready;
  assign _T_71_1 = Queue_2_io_enq_ready;
  assign _T_71_0 = Queue_1_io_enq_ready;
  assign _GEN_17 = 3'h1 == _GEN_15 ? _T_71_1 : _T_71_0;
  assign _GEN_18 = 3'h2 == _GEN_15 ? _T_71_2 : _GEN_17;
  assign _GEN_19 = 3'h3 == _GEN_15 ? _T_71_3 : _GEN_18;
  assign _GEN_20 = 3'h4 == _GEN_15 ? _T_71_4 : _GEN_19;
  assign _GEN_21 = 3'h5 == _GEN_15 ? _T_71_5 : _GEN_20;
  assign _GEN_22 = 3'h6 == _GEN_15 ? _T_71_6 : _GEN_21;
  assign _GEN_23 = 3'h7 == _GEN_15 ? _T_71_7 : _GEN_22;
  assign _T_19 = {MaxPeriodFibonacciLFSR__EVAL_12,MaxPeriodFibonacciLFSR__EVAL_11,MaxPeriodFibonacciLFSR__EVAL_3,MaxPeriodFibonacciLFSR__EVAL_16,MaxPeriodFibonacciLFSR__EVAL_8,MaxPeriodFibonacciLFSR__EVAL_10,MaxPeriodFibonacciLFSR__EVAL_14,MaxPeriodFibonacciLFSR__EVAL_7};
  assign _T_27 = {MaxPeriodFibonacciLFSR__EVAL_0,MaxPeriodFibonacciLFSR__EVAL_17,MaxPeriodFibonacciLFSR__EVAL_1,MaxPeriodFibonacciLFSR__EVAL,MaxPeriodFibonacciLFSR__EVAL_5,MaxPeriodFibonacciLFSR__EVAL_4,MaxPeriodFibonacciLFSR__EVAL_6,MaxPeriodFibonacciLFSR__EVAL_2,_T_19};
  assign _T_28 = _T_27[0];
  assign _T_29 = _T_27[1];
  assign _T_30 = _T_27[2];
  assign _T_31 = _T_27[3];
  assign _T_32 = _T_27[4];
  assign _T_33 = _T_27[5];
  assign _T_34 = _T_27[6];
  assign _T_35 = _T_27[7];
  assign _T_36 = _T_27[8];
  assign _T_37 = _T_27[9];
  assign _T_38 = _T_27[10];
  assign _T_39 = _T_27[11];
  assign _T_40 = _T_27[12];
  assign _T_41 = _T_27[13];
  assign _T_42 = _T_27[14];
  assign _T_43 = _T_27[15];
  assign _T_51 = {_T_36,_T_37,_T_38,_T_39,_T_40,_T_41,_T_42,_T_43};
  assign _T_59 = {_T_28,_T_29,_T_30,_T_31,_T_32,_T_33,_T_34,_T_35,_T_51};
  assign _T_60 = 16'h7fff <= _T_59;
  assign _T_9 = plusarg_reader_out[0];
  assign _T_64 = _T_60 | _T_9;
  assign _T_65 = _GEN_23 & _T_64;
  assign _T_6 = auto_in_aw_valid & Queue_io_enq_ready;
  assign _T_12 = _T_10 + 32'h1;
  assign _T_63 = _T_6 & _T_64;
  assign _T_67 = _T_10 + 32'h2;
  assign _T_68 = _T_59[1:0];
  assign _GEN_156 = {{30'd0}, _T_68};
  assign _T_73 = 8'h1 << _GEN_15;
  assign _T_75 = _T_73[0];
  assign _T_76 = _T_73[1];
  assign _T_77 = _T_73[2];
  assign _T_78 = _T_73[3];
  assign _T_79 = _T_73[4];
  assign _T_80 = _T_73[5];
  assign _T_81 = _T_73[6];
  assign _T_82 = _T_73[7];
  assign _T_93 = Queue_1_io_deq_bits_timestamp <= _T_10;
  assign _T_94 = _T_93 | _T_9;
  assign _T_95 = Queue_1_io_deq_valid & _T_94;
  assign _T_91_ready = Queue_9_io_enq_ready;
  assign _T_141 = _T_140 == 1'h0;
  assign _T_135 = Queue_8_io_deq_bits_timestamp <= _T_10;
  assign _T_136 = _T_135 | _T_9;
  assign _T_137 = Queue_8_io_deq_valid & _T_136;
  assign _T_129 = Queue_7_io_deq_bits_timestamp <= _T_10;
  assign _T_130 = _T_129 | _T_9;
  assign _T_131 = Queue_7_io_deq_valid & _T_130;
  assign _T_123 = Queue_6_io_deq_bits_timestamp <= _T_10;
  assign _T_124 = _T_123 | _T_9;
  assign _T_125 = Queue_6_io_deq_valid & _T_124;
  assign _T_117 = Queue_5_io_deq_bits_timestamp <= _T_10;
  assign _T_118 = _T_117 | _T_9;
  assign _T_119 = Queue_5_io_deq_valid & _T_118;
  assign _T_111 = Queue_4_io_deq_bits_timestamp <= _T_10;
  assign _T_112 = _T_111 | _T_9;
  assign _T_113 = Queue_4_io_deq_valid & _T_112;
  assign _T_105 = Queue_3_io_deq_bits_timestamp <= _T_10;
  assign _T_106 = _T_105 | _T_9;
  assign _T_107 = Queue_3_io_deq_valid & _T_106;
  assign _T_99 = Queue_2_io_deq_bits_timestamp <= _T_10;
  assign _T_100 = _T_99 | _T_9;
  assign _T_101 = Queue_2_io_deq_valid & _T_100;
  assign _T_149 = {_T_137,_T_131,_T_125,_T_119,_T_113,_T_107,_T_101,_T_95};
  assign _T_157 = ~ _T_156;
  assign _T_158 = _T_149 & _T_157;
  assign _T_159 = {_T_158,_T_137,_T_131,_T_125,_T_119,_T_113,_T_107,_T_101,_T_95};
  assign _T_160 = _T_159[15:1];
  assign _GEN_157 = {{1'd0}, _T_160};
  assign _T_161 = _T_159 | _GEN_157;
  assign _T_162 = _T_161[15:2];
  assign _GEN_158 = {{2'd0}, _T_162};
  assign _T_163 = _T_161 | _GEN_158;
  assign _T_164 = _T_163[15:4];
  assign _GEN_159 = {{4'd0}, _T_164};
  assign _T_165 = _T_163 | _GEN_159;
  assign _T_167 = _T_165[15:1];
  assign _T_168 = {_T_156, 8'h0};
  assign _GEN_160 = {{1'd0}, _T_167};
  assign _T_169 = _GEN_160 | _T_168;
  assign _T_170 = _T_169[15:8];
  assign _T_171 = _T_169[7:0];
  assign _T_172 = _T_170 & _T_171;
  assign _T_173 = ~ _T_172;
  assign _T_188 = _T_173[0];
  assign _T_289_0 = _T_141 ? _T_188 : _T_287_0;
  assign _T_290 = _T_91_ready & _T_289_0;
  assign _T_189 = _T_173[1];
  assign _T_289_1 = _T_141 ? _T_189 : _T_287_1;
  assign _T_291 = _T_91_ready & _T_289_1;
  assign _T_190 = _T_173[2];
  assign _T_289_2 = _T_141 ? _T_190 : _T_287_2;
  assign _T_292 = _T_91_ready & _T_289_2;
  assign _T_191 = _T_173[3];
  assign _T_289_3 = _T_141 ? _T_191 : _T_287_3;
  assign _T_293 = _T_91_ready & _T_289_3;
  assign _T_192 = _T_173[4];
  assign _T_289_4 = _T_141 ? _T_192 : _T_287_4;
  assign _T_294 = _T_91_ready & _T_289_4;
  assign _T_193 = _T_173[5];
  assign _T_289_5 = _T_141 ? _T_193 : _T_287_5;
  assign _T_295 = _T_91_ready & _T_289_5;
  assign _T_194 = _T_173[6];
  assign _T_289_6 = _T_141 ? _T_194 : _T_287_6;
  assign _T_296 = _T_91_ready & _T_289_6;
  assign _T_195 = _T_173[7];
  assign _T_289_7 = _T_141 ? _T_195 : _T_287_7;
  assign _T_297 = _T_91_ready & _T_289_7;
  assign _T_142 = _T_141 & _T_91_ready;
  assign _T_151 = _T_149 == _T_149;
  assign _T_153 = _T_151 | reset;
  assign _T_154 = _T_153 == 1'h0;
  assign _T_174 = _T_149 != 8'h0;
  assign _T_175 = _T_142 & _T_174;
  assign _T_176 = _T_173 & _T_149;
  assign _T_177 = {_T_176, 1'h0};
  assign _T_178 = _T_177[7:0];
  assign _T_179 = _T_176 | _T_178;
  assign _T_180 = {_T_179, 2'h0};
  assign _T_181 = _T_180[7:0];
  assign _T_182 = _T_179 | _T_181;
  assign _T_183 = {_T_182, 4'h0};
  assign _T_184 = _T_183[7:0];
  assign _T_185 = _T_182 | _T_184;
  assign _T_197 = _T_188 & _T_95;
  assign _T_198 = _T_189 & _T_101;
  assign _T_199 = _T_190 & _T_107;
  assign _T_200 = _T_191 & _T_113;
  assign _T_201 = _T_192 & _T_119;
  assign _T_202 = _T_193 & _T_125;
  assign _T_203 = _T_194 & _T_131;
  assign _T_204 = _T_195 & _T_137;
  assign _T_207 = _T_197 | _T_198;
  assign _T_208 = _T_207 | _T_199;
  assign _T_209 = _T_208 | _T_200;
  assign _T_210 = _T_209 | _T_201;
  assign _T_211 = _T_210 | _T_202;
  assign _T_212 = _T_211 | _T_203;
  assign _T_213 = _T_212 | _T_204;
  assign _T_215 = _T_197 == 1'h0;
  assign _T_218 = _T_198 == 1'h0;
  assign _T_219 = _T_215 | _T_218;
  assign _T_220 = _T_207 == 1'h0;
  assign _T_221 = _T_199 == 1'h0;
  assign _T_222 = _T_220 | _T_221;
  assign _T_223 = _T_208 == 1'h0;
  assign _T_224 = _T_200 == 1'h0;
  assign _T_225 = _T_223 | _T_224;
  assign _T_226 = _T_209 == 1'h0;
  assign _T_227 = _T_201 == 1'h0;
  assign _T_228 = _T_226 | _T_227;
  assign _T_229 = _T_210 == 1'h0;
  assign _T_230 = _T_202 == 1'h0;
  assign _T_231 = _T_229 | _T_230;
  assign _T_232 = _T_211 == 1'h0;
  assign _T_233 = _T_203 == 1'h0;
  assign _T_234 = _T_232 | _T_233;
  assign _T_235 = _T_212 == 1'h0;
  assign _T_236 = _T_204 == 1'h0;
  assign _T_237 = _T_235 | _T_236;
  assign _T_239 = _T_219 & _T_222;
  assign _T_240 = _T_239 & _T_225;
  assign _T_241 = _T_240 & _T_228;
  assign _T_242 = _T_241 & _T_231;
  assign _T_243 = _T_242 & _T_234;
  assign _T_244 = _T_243 & _T_237;
  assign _T_246 = _T_244 | reset;
  assign _T_247 = _T_246 == 1'h0;
  assign _T_248 = _T_95 | _T_101;
  assign _T_249 = _T_248 | _T_107;
  assign _T_250 = _T_249 | _T_113;
  assign _T_251 = _T_250 | _T_119;
  assign _T_252 = _T_251 | _T_125;
  assign _T_253 = _T_252 | _T_131;
  assign _T_254 = _T_253 | _T_137;
  assign _T_255 = _T_254 == 1'h0;
  assign _T_263 = _T_255 | _T_213;
  assign _T_265 = _T_263 | reset;
  assign _T_266 = _T_265 == 1'h0;
  assign _T_305 = _T_287_0 ? _T_95 : 1'h0;
  assign _T_306 = _T_287_1 ? _T_101 : 1'h0;
  assign _T_313 = _T_305 | _T_306;
  assign _T_307 = _T_287_2 ? _T_107 : 1'h0;
  assign _T_314 = _T_313 | _T_307;
  assign _T_308 = _T_287_3 ? _T_113 : 1'h0;
  assign _T_315 = _T_314 | _T_308;
  assign _T_309 = _T_287_4 ? _T_119 : 1'h0;
  assign _T_316 = _T_315 | _T_309;
  assign _T_310 = _T_287_5 ? _T_125 : 1'h0;
  assign _T_317 = _T_316 | _T_310;
  assign _T_311 = _T_287_6 ? _T_131 : 1'h0;
  assign _T_318 = _T_317 | _T_311;
  assign _T_312 = _T_287_7 ? _T_137 : 1'h0;
  assign _T_319 = _T_318 | _T_312;
  assign _T_321 = _T_141 ? _T_254 : _T_319;
  assign _T_282 = _T_91_ready & _T_321;
  assign _T_284 = _T_140 - _T_282;
  assign _T_288_0 = _T_141 ? _T_197 : _T_287_0;
  assign _T_288_1 = _T_141 ? _T_198 : _T_287_1;
  assign _T_288_2 = _T_141 ? _T_199 : _T_287_2;
  assign _T_288_3 = _T_141 ? _T_200 : _T_287_3;
  assign _T_288_4 = _T_141 ? _T_201 : _T_287_4;
  assign _T_288_5 = _T_141 ? _T_202 : _T_287_5;
  assign _T_288_6 = _T_141 ? _T_203 : _T_287_6;
  assign _T_288_7 = _T_141 ? _T_204 : _T_287_7;
  assign _T_92_bits_prot = Queue_1_io_deq_bits_data_prot;
  assign _T_92_bits_qos = Queue_1_io_deq_bits_data_qos;
  assign _T_92_bits_lock = Queue_1_io_deq_bits_data_lock;
  assign _T_92_bits_cache = Queue_1_io_deq_bits_data_cache;
  assign _T_92_bits_size = Queue_1_io_deq_bits_data_size;
  assign _T_92_bits_burst = Queue_1_io_deq_bits_data_burst;
  assign _T_92_bits_id = Queue_1_io_deq_bits_data_id;
  assign _T_92_bits_addr = Queue_1_io_deq_bits_data_addr;
  assign _T_92_bits_len = Queue_1_io_deq_bits_data_len;
  assign _T_329 = {_T_92_bits_id,_T_92_bits_addr,_T_92_bits_len,_T_92_bits_size,_T_92_bits_burst,_T_92_bits_lock,_T_92_bits_cache,_T_92_bits_prot,_T_92_bits_qos};
  assign _T_330 = _T_288_0 ? _T_329 : 60'h0;
  assign _T_98_bits_prot = Queue_2_io_deq_bits_data_prot;
  assign _T_98_bits_qos = Queue_2_io_deq_bits_data_qos;
  assign _T_98_bits_lock = Queue_2_io_deq_bits_data_lock;
  assign _T_98_bits_cache = Queue_2_io_deq_bits_data_cache;
  assign _T_98_bits_size = Queue_2_io_deq_bits_data_size;
  assign _T_98_bits_burst = Queue_2_io_deq_bits_data_burst;
  assign _T_98_bits_id = Queue_2_io_deq_bits_data_id;
  assign _T_98_bits_addr = Queue_2_io_deq_bits_data_addr;
  assign _T_98_bits_len = Queue_2_io_deq_bits_data_len;
  assign _T_338 = {_T_98_bits_id,_T_98_bits_addr,_T_98_bits_len,_T_98_bits_size,_T_98_bits_burst,_T_98_bits_lock,_T_98_bits_cache,_T_98_bits_prot,_T_98_bits_qos};
  assign _T_339 = _T_288_1 ? _T_338 : 60'h0;
  assign _T_104_bits_prot = Queue_3_io_deq_bits_data_prot;
  assign _T_104_bits_qos = Queue_3_io_deq_bits_data_qos;
  assign _T_104_bits_lock = Queue_3_io_deq_bits_data_lock;
  assign _T_104_bits_cache = Queue_3_io_deq_bits_data_cache;
  assign _T_104_bits_size = Queue_3_io_deq_bits_data_size;
  assign _T_104_bits_burst = Queue_3_io_deq_bits_data_burst;
  assign _T_104_bits_id = Queue_3_io_deq_bits_data_id;
  assign _T_104_bits_addr = Queue_3_io_deq_bits_data_addr;
  assign _T_104_bits_len = Queue_3_io_deq_bits_data_len;
  assign _T_347 = {_T_104_bits_id,_T_104_bits_addr,_T_104_bits_len,_T_104_bits_size,_T_104_bits_burst,_T_104_bits_lock,_T_104_bits_cache,_T_104_bits_prot,_T_104_bits_qos};
  assign _T_348 = _T_288_2 ? _T_347 : 60'h0;
  assign _T_110_bits_prot = Queue_4_io_deq_bits_data_prot;
  assign _T_110_bits_qos = Queue_4_io_deq_bits_data_qos;
  assign _T_110_bits_lock = Queue_4_io_deq_bits_data_lock;
  assign _T_110_bits_cache = Queue_4_io_deq_bits_data_cache;
  assign _T_110_bits_size = Queue_4_io_deq_bits_data_size;
  assign _T_110_bits_burst = Queue_4_io_deq_bits_data_burst;
  assign _T_110_bits_id = Queue_4_io_deq_bits_data_id;
  assign _T_110_bits_addr = Queue_4_io_deq_bits_data_addr;
  assign _T_110_bits_len = Queue_4_io_deq_bits_data_len;
  assign _T_356 = {_T_110_bits_id,_T_110_bits_addr,_T_110_bits_len,_T_110_bits_size,_T_110_bits_burst,_T_110_bits_lock,_T_110_bits_cache,_T_110_bits_prot,_T_110_bits_qos};
  assign _T_357 = _T_288_3 ? _T_356 : 60'h0;
  assign _T_116_bits_prot = Queue_5_io_deq_bits_data_prot;
  assign _T_116_bits_qos = Queue_5_io_deq_bits_data_qos;
  assign _T_116_bits_lock = Queue_5_io_deq_bits_data_lock;
  assign _T_116_bits_cache = Queue_5_io_deq_bits_data_cache;
  assign _T_116_bits_size = Queue_5_io_deq_bits_data_size;
  assign _T_116_bits_burst = Queue_5_io_deq_bits_data_burst;
  assign _T_116_bits_id = Queue_5_io_deq_bits_data_id;
  assign _T_116_bits_addr = Queue_5_io_deq_bits_data_addr;
  assign _T_116_bits_len = Queue_5_io_deq_bits_data_len;
  assign _T_365 = {_T_116_bits_id,_T_116_bits_addr,_T_116_bits_len,_T_116_bits_size,_T_116_bits_burst,_T_116_bits_lock,_T_116_bits_cache,_T_116_bits_prot,_T_116_bits_qos};
  assign _T_366 = _T_288_4 ? _T_365 : 60'h0;
  assign _T_122_bits_prot = Queue_6_io_deq_bits_data_prot;
  assign _T_122_bits_qos = Queue_6_io_deq_bits_data_qos;
  assign _T_122_bits_lock = Queue_6_io_deq_bits_data_lock;
  assign _T_122_bits_cache = Queue_6_io_deq_bits_data_cache;
  assign _T_122_bits_size = Queue_6_io_deq_bits_data_size;
  assign _T_122_bits_burst = Queue_6_io_deq_bits_data_burst;
  assign _T_122_bits_id = Queue_6_io_deq_bits_data_id;
  assign _T_122_bits_addr = Queue_6_io_deq_bits_data_addr;
  assign _T_122_bits_len = Queue_6_io_deq_bits_data_len;
  assign _T_374 = {_T_122_bits_id,_T_122_bits_addr,_T_122_bits_len,_T_122_bits_size,_T_122_bits_burst,_T_122_bits_lock,_T_122_bits_cache,_T_122_bits_prot,_T_122_bits_qos};
  assign _T_375 = _T_288_5 ? _T_374 : 60'h0;
  assign _T_128_bits_prot = Queue_7_io_deq_bits_data_prot;
  assign _T_128_bits_qos = Queue_7_io_deq_bits_data_qos;
  assign _T_128_bits_lock = Queue_7_io_deq_bits_data_lock;
  assign _T_128_bits_cache = Queue_7_io_deq_bits_data_cache;
  assign _T_128_bits_size = Queue_7_io_deq_bits_data_size;
  assign _T_128_bits_burst = Queue_7_io_deq_bits_data_burst;
  assign _T_128_bits_id = Queue_7_io_deq_bits_data_id;
  assign _T_128_bits_addr = Queue_7_io_deq_bits_data_addr;
  assign _T_128_bits_len = Queue_7_io_deq_bits_data_len;
  assign _T_383 = {_T_128_bits_id,_T_128_bits_addr,_T_128_bits_len,_T_128_bits_size,_T_128_bits_burst,_T_128_bits_lock,_T_128_bits_cache,_T_128_bits_prot,_T_128_bits_qos};
  assign _T_384 = _T_288_6 ? _T_383 : 60'h0;
  assign _T_134_bits_prot = Queue_8_io_deq_bits_data_prot;
  assign _T_134_bits_qos = Queue_8_io_deq_bits_data_qos;
  assign _T_134_bits_lock = Queue_8_io_deq_bits_data_lock;
  assign _T_134_bits_cache = Queue_8_io_deq_bits_data_cache;
  assign _T_134_bits_size = Queue_8_io_deq_bits_data_size;
  assign _T_134_bits_burst = Queue_8_io_deq_bits_data_burst;
  assign _T_134_bits_id = Queue_8_io_deq_bits_data_id;
  assign _T_134_bits_addr = Queue_8_io_deq_bits_data_addr;
  assign _T_134_bits_len = Queue_8_io_deq_bits_data_len;
  assign _T_392 = {_T_134_bits_id,_T_134_bits_addr,_T_134_bits_len,_T_134_bits_size,_T_134_bits_burst,_T_134_bits_lock,_T_134_bits_cache,_T_134_bits_prot,_T_134_bits_qos};
  assign _T_393 = _T_288_7 ? _T_392 : 60'h0;
  assign _T_394 = _T_330 | _T_339;
  assign _T_395 = _T_394 | _T_348;
  assign _T_396 = _T_395 | _T_357;
  assign _T_397 = _T_396 | _T_366;
  assign _T_398 = _T_397 | _T_375;
  assign _T_399 = _T_398 | _T_384;
  assign _T_400 = _T_399 | _T_393;
  assign _T_413_ready = Queue_11_io_enq_ready;
  assign _T_412_valid = Queue_9_io_deq_valid;
  assign _T_412_bits_id = Queue_9_io_deq_bits_id;
  assign _GEN_26 = 4'h1 == _T_412_bits_id ? 3'h0 : 3'h5;
  assign _GEN_27 = 4'h2 == _T_412_bits_id ? 3'h5 : _GEN_26;
  assign _GEN_28 = 4'h3 == _T_412_bits_id ? 3'h0 : _GEN_27;
  assign _GEN_29 = 4'h4 == _T_412_bits_id ? 3'h2 : _GEN_28;
  assign _GEN_30 = 4'h5 == _T_412_bits_id ? 3'h7 : _GEN_29;
  assign _GEN_31 = 4'h6 == _T_412_bits_id ? 3'h2 : _GEN_30;
  assign _GEN_32 = 4'h7 == _T_412_bits_id ? 3'h5 : _GEN_31;
  assign _GEN_33 = 4'h8 == _T_412_bits_id ? 3'h5 : _GEN_32;
  assign _GEN_34 = 4'h9 == _T_412_bits_id ? 3'h0 : _GEN_33;
  assign _GEN_35 = 4'ha == _T_412_bits_id ? 3'h7 : _GEN_34;
  assign _GEN_36 = 4'hb == _T_412_bits_id ? 3'h3 : _GEN_35;
  assign _GEN_37 = 4'hc == _T_412_bits_id ? 3'h2 : _GEN_36;
  assign _GEN_38 = 4'hd == _T_412_bits_id ? 3'h3 : _GEN_37;
  assign _GEN_39 = 4'he == _T_412_bits_id ? 3'h2 : _GEN_38;
  assign _T_4_bits = Queue_io_deq_bits;
  assign _T_418_0 = Queue_12_io_enq_ready;
  assign _T_418_1 = Queue_13_io_enq_ready;
  assign _GEN_42 = 3'h1 == _T_4_bits ? _T_418_1 : _T_418_0;
  assign _T_418_2 = Queue_14_io_enq_ready;
  assign _GEN_43 = 3'h2 == _T_4_bits ? _T_418_2 : _GEN_42;
  assign _T_418_3 = Queue_15_io_enq_ready;
  assign _GEN_44 = 3'h3 == _T_4_bits ? _T_418_3 : _GEN_43;
  assign _T_418_4 = Queue_16_io_enq_ready;
  assign _GEN_45 = 3'h4 == _T_4_bits ? _T_418_4 : _GEN_44;
  assign _T_418_5 = Queue_17_io_enq_ready;
  assign _GEN_46 = 3'h5 == _T_4_bits ? _T_418_5 : _GEN_45;
  assign _T_418_6 = Queue_18_io_enq_ready;
  assign _GEN_47 = 3'h6 == _T_4_bits ? _T_418_6 : _GEN_46;
  assign _T_418_7 = Queue_19_io_enq_ready;
  assign _GEN_48 = 3'h7 == _T_4_bits ? _T_418_7 : _GEN_47;
  assign _T_419 = auto_in_w_bits_last & _GEN_48;
  assign _T_4_valid = Queue_io_deq_valid;
  assign _T_423 = 8'h1 << _T_4_bits;
  assign _T_425 = _T_423[0];
  assign _T_426 = _T_423[1];
  assign _T_427 = _T_423[2];
  assign _T_428 = _T_423[3];
  assign _T_429 = _T_423[4];
  assign _T_430 = _T_423[5];
  assign _T_431 = _T_423[6];
  assign _T_432 = _T_423[7];
  assign _T_433 = _T_4_valid & auto_in_w_valid;
  assign _T_414_bits = Queue_10_io_deq_bits;
  assign _T_451_0_data = Queue_12_io_deq_bits_data;
  assign _T_451_0_strb = Queue_12_io_deq_bits_strb;
  assign _T_451_0_last = Queue_12_io_deq_bits_last;
  assign _T_451_1_data = Queue_13_io_deq_bits_data;
  assign _GEN_52 = 3'h1 == _T_414_bits ? _T_451_1_data : _T_451_0_data;
  assign _T_451_1_strb = Queue_13_io_deq_bits_strb;
  assign _GEN_53 = 3'h1 == _T_414_bits ? _T_451_1_strb : _T_451_0_strb;
  assign _T_451_1_last = Queue_13_io_deq_bits_last;
  assign _GEN_54 = 3'h1 == _T_414_bits ? _T_451_1_last : _T_451_0_last;
  assign _T_451_2_data = Queue_14_io_deq_bits_data;
  assign _GEN_55 = 3'h2 == _T_414_bits ? _T_451_2_data : _GEN_52;
  assign _T_451_2_strb = Queue_14_io_deq_bits_strb;
  assign _GEN_56 = 3'h2 == _T_414_bits ? _T_451_2_strb : _GEN_53;
  assign _T_451_2_last = Queue_14_io_deq_bits_last;
  assign _GEN_57 = 3'h2 == _T_414_bits ? _T_451_2_last : _GEN_54;
  assign _T_451_3_data = Queue_15_io_deq_bits_data;
  assign _GEN_58 = 3'h3 == _T_414_bits ? _T_451_3_data : _GEN_55;
  assign _T_451_3_strb = Queue_15_io_deq_bits_strb;
  assign _GEN_59 = 3'h3 == _T_414_bits ? _T_451_3_strb : _GEN_56;
  assign _T_451_3_last = Queue_15_io_deq_bits_last;
  assign _GEN_60 = 3'h3 == _T_414_bits ? _T_451_3_last : _GEN_57;
  assign _T_451_4_data = Queue_16_io_deq_bits_data;
  assign _GEN_61 = 3'h4 == _T_414_bits ? _T_451_4_data : _GEN_58;
  assign _T_451_4_strb = Queue_16_io_deq_bits_strb;
  assign _GEN_62 = 3'h4 == _T_414_bits ? _T_451_4_strb : _GEN_59;
  assign _T_451_4_last = Queue_16_io_deq_bits_last;
  assign _GEN_63 = 3'h4 == _T_414_bits ? _T_451_4_last : _GEN_60;
  assign _T_451_5_data = Queue_17_io_deq_bits_data;
  assign _GEN_64 = 3'h5 == _T_414_bits ? _T_451_5_data : _GEN_61;
  assign _T_451_5_strb = Queue_17_io_deq_bits_strb;
  assign _GEN_65 = 3'h5 == _T_414_bits ? _T_451_5_strb : _GEN_62;
  assign _T_451_5_last = Queue_17_io_deq_bits_last;
  assign _GEN_66 = 3'h5 == _T_414_bits ? _T_451_5_last : _GEN_63;
  assign _T_451_6_data = Queue_18_io_deq_bits_data;
  assign _GEN_67 = 3'h6 == _T_414_bits ? _T_451_6_data : _GEN_64;
  assign _T_451_6_strb = Queue_18_io_deq_bits_strb;
  assign _GEN_68 = 3'h6 == _T_414_bits ? _T_451_6_strb : _GEN_65;
  assign _T_451_6_last = Queue_18_io_deq_bits_last;
  assign _GEN_69 = 3'h6 == _T_414_bits ? _T_451_6_last : _GEN_66;
  assign _T_451_7_data = Queue_19_io_deq_bits_data;
  assign _T_451_7_strb = Queue_19_io_deq_bits_strb;
  assign _T_451_7_last = Queue_19_io_deq_bits_last;
  assign _GEN_72 = 3'h7 == _T_414_bits ? _T_451_7_last : _GEN_69;
  assign _T_450_0 = Queue_12_io_deq_valid;
  assign _T_450_1 = Queue_13_io_deq_valid;
  assign _GEN_74 = 3'h1 == _T_414_bits ? _T_450_1 : _T_450_0;
  assign _T_450_2 = Queue_14_io_deq_valid;
  assign _GEN_75 = 3'h2 == _T_414_bits ? _T_450_2 : _GEN_74;
  assign _T_450_3 = Queue_15_io_deq_valid;
  assign _GEN_76 = 3'h3 == _T_414_bits ? _T_450_3 : _GEN_75;
  assign _T_450_4 = Queue_16_io_deq_valid;
  assign _GEN_77 = 3'h4 == _T_414_bits ? _T_450_4 : _GEN_76;
  assign _T_450_5 = Queue_17_io_deq_valid;
  assign _GEN_78 = 3'h5 == _T_414_bits ? _T_450_5 : _GEN_77;
  assign _T_450_6 = Queue_18_io_deq_valid;
  assign _GEN_79 = 3'h6 == _T_414_bits ? _T_450_6 : _GEN_78;
  assign _T_450_7 = Queue_19_io_deq_valid;
  assign _GEN_80 = 3'h7 == _T_414_bits ? _T_450_7 : _GEN_79;
  assign _T_452 = _GEN_72 & _GEN_80;
  assign _T_414_valid = Queue_10_io_deq_valid;
  assign _T_456 = 8'h1 << _T_414_bits;
  assign _T_458 = _T_456[0];
  assign _T_459 = _T_456[1];
  assign _T_460 = _T_456[2];
  assign _T_461 = _T_456[3];
  assign _T_462 = _T_456[4];
  assign _T_463 = _T_456[5];
  assign _T_464 = _T_456[6];
  assign _T_465 = _T_456[7];
  assign _T_466 = _T_414_valid & auto_out_w_ready;
  assign _T_483 = plusarg_reader_1_out[0];
  assign _T_486 = _T_484 + 32'h1;
  assign _T_493 = {MaxPeriodFibonacciLFSR_1__EVAL_12,MaxPeriodFibonacciLFSR_1__EVAL_11,MaxPeriodFibonacciLFSR_1__EVAL_3,MaxPeriodFibonacciLFSR_1__EVAL_16,MaxPeriodFibonacciLFSR_1__EVAL_8,MaxPeriodFibonacciLFSR_1__EVAL_10,MaxPeriodFibonacciLFSR_1__EVAL_14,MaxPeriodFibonacciLFSR_1__EVAL_7};
  assign _T_501 = {MaxPeriodFibonacciLFSR_1__EVAL_0,MaxPeriodFibonacciLFSR_1__EVAL_17,MaxPeriodFibonacciLFSR_1__EVAL_1,MaxPeriodFibonacciLFSR_1__EVAL,MaxPeriodFibonacciLFSR_1__EVAL_5,MaxPeriodFibonacciLFSR_1__EVAL_4,MaxPeriodFibonacciLFSR_1__EVAL_6,MaxPeriodFibonacciLFSR_1__EVAL_2,_T_493};
  assign _T_502 = _T_501[0];
  assign _T_503 = _T_501[1];
  assign _T_504 = _T_501[2];
  assign _T_505 = _T_501[3];
  assign _T_506 = _T_501[4];
  assign _T_507 = _T_501[5];
  assign _T_508 = _T_501[6];
  assign _T_509 = _T_501[7];
  assign _T_510 = _T_501[8];
  assign _T_511 = _T_501[9];
  assign _T_512 = _T_501[10];
  assign _T_513 = _T_501[11];
  assign _T_514 = _T_501[12];
  assign _T_515 = _T_501[13];
  assign _T_516 = _T_501[14];
  assign _T_517 = _T_501[15];
  assign _T_525 = {_T_510,_T_511,_T_512,_T_513,_T_514,_T_515,_T_516,_T_517};
  assign _T_533 = {_T_502,_T_503,_T_504,_T_505,_T_506,_T_507,_T_508,_T_509,_T_525};
  assign _T_534 = 16'h7fff <= _T_533;
  assign _T_536 = _T_534 | _T_483;
  assign _T_537 = auto_in_ar_valid & _T_536;
  assign _GEN_82 = 4'h1 == auto_in_ar_bits_id ? 3'h0 : 3'h5;
  assign _GEN_83 = 4'h2 == auto_in_ar_bits_id ? 3'h5 : _GEN_82;
  assign _GEN_84 = 4'h3 == auto_in_ar_bits_id ? 3'h0 : _GEN_83;
  assign _GEN_85 = 4'h4 == auto_in_ar_bits_id ? 3'h2 : _GEN_84;
  assign _GEN_86 = 4'h5 == auto_in_ar_bits_id ? 3'h7 : _GEN_85;
  assign _GEN_87 = 4'h6 == auto_in_ar_bits_id ? 3'h2 : _GEN_86;
  assign _GEN_88 = 4'h7 == auto_in_ar_bits_id ? 3'h5 : _GEN_87;
  assign _GEN_89 = 4'h8 == auto_in_ar_bits_id ? 3'h5 : _GEN_88;
  assign _GEN_90 = 4'h9 == auto_in_ar_bits_id ? 3'h0 : _GEN_89;
  assign _GEN_91 = 4'ha == auto_in_ar_bits_id ? 3'h7 : _GEN_90;
  assign _GEN_92 = 4'hb == auto_in_ar_bits_id ? 3'h3 : _GEN_91;
  assign _GEN_93 = 4'hc == auto_in_ar_bits_id ? 3'h2 : _GEN_92;
  assign _GEN_94 = 4'hd == auto_in_ar_bits_id ? 3'h3 : _GEN_93;
  assign _GEN_95 = 4'he == auto_in_ar_bits_id ? 3'h2 : _GEN_94;
  assign _GEN_96 = 4'hf == auto_in_ar_bits_id ? 3'h5 : _GEN_95;
  assign _T_545_7 = Queue_27_io_enq_ready;
  assign _T_545_6 = Queue_26_io_enq_ready;
  assign _T_545_5 = Queue_25_io_enq_ready;
  assign _T_545_4 = Queue_24_io_enq_ready;
  assign _T_545_3 = Queue_23_io_enq_ready;
  assign _T_545_2 = Queue_22_io_enq_ready;
  assign _T_545_1 = Queue_21_io_enq_ready;
  assign _T_545_0 = Queue_20_io_enq_ready;
  assign _GEN_98 = 3'h1 == _GEN_96 ? _T_545_1 : _T_545_0;
  assign _GEN_99 = 3'h2 == _GEN_96 ? _T_545_2 : _GEN_98;
  assign _GEN_100 = 3'h3 == _GEN_96 ? _T_545_3 : _GEN_99;
  assign _GEN_101 = 3'h4 == _GEN_96 ? _T_545_4 : _GEN_100;
  assign _GEN_102 = 3'h5 == _GEN_96 ? _T_545_5 : _GEN_101;
  assign _GEN_103 = 3'h6 == _GEN_96 ? _T_545_6 : _GEN_102;
  assign _GEN_104 = 3'h7 == _GEN_96 ? _T_545_7 : _GEN_103;
  assign _T_541 = _T_484 + 32'h2;
  assign _T_542 = _T_533[1:0];
  assign _GEN_161 = {{30'd0}, _T_542};
  assign _T_547 = 8'h1 << _GEN_96;
  assign _T_549 = _T_547[0];
  assign _T_550 = _T_547[1];
  assign _T_551 = _T_547[2];
  assign _T_552 = _T_547[3];
  assign _T_553 = _T_547[4];
  assign _T_554 = _T_547[5];
  assign _T_555 = _T_547[6];
  assign _T_556 = _T_547[7];
  assign _T_567 = Queue_20_io_deq_bits_timestamp <= _T_484;
  assign _T_568 = _T_567 | _T_483;
  assign _T_569 = Queue_20_io_deq_valid & _T_568;
  assign _T_565_ready = Queue_28_io_enq_ready;
  assign _T_615 = _T_614 == 1'h0;
  assign _T_609 = Queue_27_io_deq_bits_timestamp <= _T_484;
  assign _T_610 = _T_609 | _T_483;
  assign _T_611 = Queue_27_io_deq_valid & _T_610;
  assign _T_603 = Queue_26_io_deq_bits_timestamp <= _T_484;
  assign _T_604 = _T_603 | _T_483;
  assign _T_605 = Queue_26_io_deq_valid & _T_604;
  assign _T_597 = Queue_25_io_deq_bits_timestamp <= _T_484;
  assign _T_598 = _T_597 | _T_483;
  assign _T_599 = Queue_25_io_deq_valid & _T_598;
  assign _T_591 = Queue_24_io_deq_bits_timestamp <= _T_484;
  assign _T_592 = _T_591 | _T_483;
  assign _T_593 = Queue_24_io_deq_valid & _T_592;
  assign _T_585 = Queue_23_io_deq_bits_timestamp <= _T_484;
  assign _T_586 = _T_585 | _T_483;
  assign _T_587 = Queue_23_io_deq_valid & _T_586;
  assign _T_579 = Queue_22_io_deq_bits_timestamp <= _T_484;
  assign _T_580 = _T_579 | _T_483;
  assign _T_581 = Queue_22_io_deq_valid & _T_580;
  assign _T_573 = Queue_21_io_deq_bits_timestamp <= _T_484;
  assign _T_574 = _T_573 | _T_483;
  assign _T_575 = Queue_21_io_deq_valid & _T_574;
  assign _T_623 = {_T_611,_T_605,_T_599,_T_593,_T_587,_T_581,_T_575,_T_569};
  assign _T_631 = ~ _T_630;
  assign _T_632 = _T_623 & _T_631;
  assign _T_633 = {_T_632,_T_611,_T_605,_T_599,_T_593,_T_587,_T_581,_T_575,_T_569};
  assign _T_634 = _T_633[15:1];
  assign _GEN_162 = {{1'd0}, _T_634};
  assign _T_635 = _T_633 | _GEN_162;
  assign _T_636 = _T_635[15:2];
  assign _GEN_163 = {{2'd0}, _T_636};
  assign _T_637 = _T_635 | _GEN_163;
  assign _T_638 = _T_637[15:4];
  assign _GEN_164 = {{4'd0}, _T_638};
  assign _T_639 = _T_637 | _GEN_164;
  assign _T_641 = _T_639[15:1];
  assign _T_642 = {_T_630, 8'h0};
  assign _GEN_165 = {{1'd0}, _T_641};
  assign _T_643 = _GEN_165 | _T_642;
  assign _T_644 = _T_643[15:8];
  assign _T_645 = _T_643[7:0];
  assign _T_646 = _T_644 & _T_645;
  assign _T_647 = ~ _T_646;
  assign _T_662 = _T_647[0];
  assign _T_763_0 = _T_615 ? _T_662 : _T_761_0;
  assign _T_764 = _T_565_ready & _T_763_0;
  assign _T_663 = _T_647[1];
  assign _T_763_1 = _T_615 ? _T_663 : _T_761_1;
  assign _T_765 = _T_565_ready & _T_763_1;
  assign _T_664 = _T_647[2];
  assign _T_763_2 = _T_615 ? _T_664 : _T_761_2;
  assign _T_766 = _T_565_ready & _T_763_2;
  assign _T_665 = _T_647[3];
  assign _T_763_3 = _T_615 ? _T_665 : _T_761_3;
  assign _T_767 = _T_565_ready & _T_763_3;
  assign _T_666 = _T_647[4];
  assign _T_763_4 = _T_615 ? _T_666 : _T_761_4;
  assign _T_768 = _T_565_ready & _T_763_4;
  assign _T_667 = _T_647[5];
  assign _T_763_5 = _T_615 ? _T_667 : _T_761_5;
  assign _T_769 = _T_565_ready & _T_763_5;
  assign _T_668 = _T_647[6];
  assign _T_763_6 = _T_615 ? _T_668 : _T_761_6;
  assign _T_770 = _T_565_ready & _T_763_6;
  assign _T_669 = _T_647[7];
  assign _T_763_7 = _T_615 ? _T_669 : _T_761_7;
  assign _T_771 = _T_565_ready & _T_763_7;
  assign _T_616 = _T_615 & _T_565_ready;
  assign _T_625 = _T_623 == _T_623;
  assign _T_627 = _T_625 | reset;
  assign _T_628 = _T_627 == 1'h0;
  assign _T_648 = _T_623 != 8'h0;
  assign _T_649 = _T_616 & _T_648;
  assign _T_650 = _T_647 & _T_623;
  assign _T_651 = {_T_650, 1'h0};
  assign _T_652 = _T_651[7:0];
  assign _T_653 = _T_650 | _T_652;
  assign _T_654 = {_T_653, 2'h0};
  assign _T_655 = _T_654[7:0];
  assign _T_656 = _T_653 | _T_655;
  assign _T_657 = {_T_656, 4'h0};
  assign _T_658 = _T_657[7:0];
  assign _T_659 = _T_656 | _T_658;
  assign _T_671 = _T_662 & _T_569;
  assign _T_672 = _T_663 & _T_575;
  assign _T_673 = _T_664 & _T_581;
  assign _T_674 = _T_665 & _T_587;
  assign _T_675 = _T_666 & _T_593;
  assign _T_676 = _T_667 & _T_599;
  assign _T_677 = _T_668 & _T_605;
  assign _T_678 = _T_669 & _T_611;
  assign _T_681 = _T_671 | _T_672;
  assign _T_682 = _T_681 | _T_673;
  assign _T_683 = _T_682 | _T_674;
  assign _T_684 = _T_683 | _T_675;
  assign _T_685 = _T_684 | _T_676;
  assign _T_686 = _T_685 | _T_677;
  assign _T_687 = _T_686 | _T_678;
  assign _T_689 = _T_671 == 1'h0;
  assign _T_692 = _T_672 == 1'h0;
  assign _T_693 = _T_689 | _T_692;
  assign _T_694 = _T_681 == 1'h0;
  assign _T_695 = _T_673 == 1'h0;
  assign _T_696 = _T_694 | _T_695;
  assign _T_697 = _T_682 == 1'h0;
  assign _T_698 = _T_674 == 1'h0;
  assign _T_699 = _T_697 | _T_698;
  assign _T_700 = _T_683 == 1'h0;
  assign _T_701 = _T_675 == 1'h0;
  assign _T_702 = _T_700 | _T_701;
  assign _T_703 = _T_684 == 1'h0;
  assign _T_704 = _T_676 == 1'h0;
  assign _T_705 = _T_703 | _T_704;
  assign _T_706 = _T_685 == 1'h0;
  assign _T_707 = _T_677 == 1'h0;
  assign _T_708 = _T_706 | _T_707;
  assign _T_709 = _T_686 == 1'h0;
  assign _T_710 = _T_678 == 1'h0;
  assign _T_711 = _T_709 | _T_710;
  assign _T_713 = _T_693 & _T_696;
  assign _T_714 = _T_713 & _T_699;
  assign _T_715 = _T_714 & _T_702;
  assign _T_716 = _T_715 & _T_705;
  assign _T_717 = _T_716 & _T_708;
  assign _T_718 = _T_717 & _T_711;
  assign _T_720 = _T_718 | reset;
  assign _T_721 = _T_720 == 1'h0;
  assign _T_722 = _T_569 | _T_575;
  assign _T_723 = _T_722 | _T_581;
  assign _T_724 = _T_723 | _T_587;
  assign _T_725 = _T_724 | _T_593;
  assign _T_726 = _T_725 | _T_599;
  assign _T_727 = _T_726 | _T_605;
  assign _T_728 = _T_727 | _T_611;
  assign _T_729 = _T_728 == 1'h0;
  assign _T_737 = _T_729 | _T_687;
  assign _T_739 = _T_737 | reset;
  assign _T_740 = _T_739 == 1'h0;
  assign _T_779 = _T_761_0 ? _T_569 : 1'h0;
  assign _T_780 = _T_761_1 ? _T_575 : 1'h0;
  assign _T_787 = _T_779 | _T_780;
  assign _T_781 = _T_761_2 ? _T_581 : 1'h0;
  assign _T_788 = _T_787 | _T_781;
  assign _T_782 = _T_761_3 ? _T_587 : 1'h0;
  assign _T_789 = _T_788 | _T_782;
  assign _T_783 = _T_761_4 ? _T_593 : 1'h0;
  assign _T_790 = _T_789 | _T_783;
  assign _T_784 = _T_761_5 ? _T_599 : 1'h0;
  assign _T_791 = _T_790 | _T_784;
  assign _T_785 = _T_761_6 ? _T_605 : 1'h0;
  assign _T_792 = _T_791 | _T_785;
  assign _T_786 = _T_761_7 ? _T_611 : 1'h0;
  assign _T_793 = _T_792 | _T_786;
  assign _T_795 = _T_615 ? _T_728 : _T_793;
  assign _T_756 = _T_565_ready & _T_795;
  assign _T_758 = _T_614 - _T_756;
  assign _T_762_0 = _T_615 ? _T_671 : _T_761_0;
  assign _T_762_1 = _T_615 ? _T_672 : _T_761_1;
  assign _T_762_2 = _T_615 ? _T_673 : _T_761_2;
  assign _T_762_3 = _T_615 ? _T_674 : _T_761_3;
  assign _T_762_4 = _T_615 ? _T_675 : _T_761_4;
  assign _T_762_5 = _T_615 ? _T_676 : _T_761_5;
  assign _T_762_6 = _T_615 ? _T_677 : _T_761_6;
  assign _T_762_7 = _T_615 ? _T_678 : _T_761_7;
  assign _T_566_bits_prot = Queue_20_io_deq_bits_data_prot;
  assign _T_566_bits_qos = Queue_20_io_deq_bits_data_qos;
  assign _T_566_bits_lock = Queue_20_io_deq_bits_data_lock;
  assign _T_566_bits_cache = Queue_20_io_deq_bits_data_cache;
  assign _T_566_bits_size = Queue_20_io_deq_bits_data_size;
  assign _T_566_bits_burst = Queue_20_io_deq_bits_data_burst;
  assign _T_566_bits_id = Queue_20_io_deq_bits_data_id;
  assign _T_566_bits_addr = Queue_20_io_deq_bits_data_addr;
  assign _T_566_bits_len = Queue_20_io_deq_bits_data_len;
  assign _T_803 = {_T_566_bits_id,_T_566_bits_addr,_T_566_bits_len,_T_566_bits_size,_T_566_bits_burst,_T_566_bits_lock,_T_566_bits_cache,_T_566_bits_prot,_T_566_bits_qos};
  assign _T_804 = _T_762_0 ? _T_803 : 60'h0;
  assign _T_572_bits_prot = Queue_21_io_deq_bits_data_prot;
  assign _T_572_bits_qos = Queue_21_io_deq_bits_data_qos;
  assign _T_572_bits_lock = Queue_21_io_deq_bits_data_lock;
  assign _T_572_bits_cache = Queue_21_io_deq_bits_data_cache;
  assign _T_572_bits_size = Queue_21_io_deq_bits_data_size;
  assign _T_572_bits_burst = Queue_21_io_deq_bits_data_burst;
  assign _T_572_bits_id = Queue_21_io_deq_bits_data_id;
  assign _T_572_bits_addr = Queue_21_io_deq_bits_data_addr;
  assign _T_572_bits_len = Queue_21_io_deq_bits_data_len;
  assign _T_812 = {_T_572_bits_id,_T_572_bits_addr,_T_572_bits_len,_T_572_bits_size,_T_572_bits_burst,_T_572_bits_lock,_T_572_bits_cache,_T_572_bits_prot,_T_572_bits_qos};
  assign _T_813 = _T_762_1 ? _T_812 : 60'h0;
  assign _T_578_bits_prot = Queue_22_io_deq_bits_data_prot;
  assign _T_578_bits_qos = Queue_22_io_deq_bits_data_qos;
  assign _T_578_bits_lock = Queue_22_io_deq_bits_data_lock;
  assign _T_578_bits_cache = Queue_22_io_deq_bits_data_cache;
  assign _T_578_bits_size = Queue_22_io_deq_bits_data_size;
  assign _T_578_bits_burst = Queue_22_io_deq_bits_data_burst;
  assign _T_578_bits_id = Queue_22_io_deq_bits_data_id;
  assign _T_578_bits_addr = Queue_22_io_deq_bits_data_addr;
  assign _T_578_bits_len = Queue_22_io_deq_bits_data_len;
  assign _T_821 = {_T_578_bits_id,_T_578_bits_addr,_T_578_bits_len,_T_578_bits_size,_T_578_bits_burst,_T_578_bits_lock,_T_578_bits_cache,_T_578_bits_prot,_T_578_bits_qos};
  assign _T_822 = _T_762_2 ? _T_821 : 60'h0;
  assign _T_584_bits_prot = Queue_23_io_deq_bits_data_prot;
  assign _T_584_bits_qos = Queue_23_io_deq_bits_data_qos;
  assign _T_584_bits_lock = Queue_23_io_deq_bits_data_lock;
  assign _T_584_bits_cache = Queue_23_io_deq_bits_data_cache;
  assign _T_584_bits_size = Queue_23_io_deq_bits_data_size;
  assign _T_584_bits_burst = Queue_23_io_deq_bits_data_burst;
  assign _T_584_bits_id = Queue_23_io_deq_bits_data_id;
  assign _T_584_bits_addr = Queue_23_io_deq_bits_data_addr;
  assign _T_584_bits_len = Queue_23_io_deq_bits_data_len;
  assign _T_830 = {_T_584_bits_id,_T_584_bits_addr,_T_584_bits_len,_T_584_bits_size,_T_584_bits_burst,_T_584_bits_lock,_T_584_bits_cache,_T_584_bits_prot,_T_584_bits_qos};
  assign _T_831 = _T_762_3 ? _T_830 : 60'h0;
  assign _T_590_bits_prot = Queue_24_io_deq_bits_data_prot;
  assign _T_590_bits_qos = Queue_24_io_deq_bits_data_qos;
  assign _T_590_bits_lock = Queue_24_io_deq_bits_data_lock;
  assign _T_590_bits_cache = Queue_24_io_deq_bits_data_cache;
  assign _T_590_bits_size = Queue_24_io_deq_bits_data_size;
  assign _T_590_bits_burst = Queue_24_io_deq_bits_data_burst;
  assign _T_590_bits_id = Queue_24_io_deq_bits_data_id;
  assign _T_590_bits_addr = Queue_24_io_deq_bits_data_addr;
  assign _T_590_bits_len = Queue_24_io_deq_bits_data_len;
  assign _T_839 = {_T_590_bits_id,_T_590_bits_addr,_T_590_bits_len,_T_590_bits_size,_T_590_bits_burst,_T_590_bits_lock,_T_590_bits_cache,_T_590_bits_prot,_T_590_bits_qos};
  assign _T_840 = _T_762_4 ? _T_839 : 60'h0;
  assign _T_596_bits_prot = Queue_25_io_deq_bits_data_prot;
  assign _T_596_bits_qos = Queue_25_io_deq_bits_data_qos;
  assign _T_596_bits_lock = Queue_25_io_deq_bits_data_lock;
  assign _T_596_bits_cache = Queue_25_io_deq_bits_data_cache;
  assign _T_596_bits_size = Queue_25_io_deq_bits_data_size;
  assign _T_596_bits_burst = Queue_25_io_deq_bits_data_burst;
  assign _T_596_bits_id = Queue_25_io_deq_bits_data_id;
  assign _T_596_bits_addr = Queue_25_io_deq_bits_data_addr;
  assign _T_596_bits_len = Queue_25_io_deq_bits_data_len;
  assign _T_848 = {_T_596_bits_id,_T_596_bits_addr,_T_596_bits_len,_T_596_bits_size,_T_596_bits_burst,_T_596_bits_lock,_T_596_bits_cache,_T_596_bits_prot,_T_596_bits_qos};
  assign _T_849 = _T_762_5 ? _T_848 : 60'h0;
  assign _T_602_bits_prot = Queue_26_io_deq_bits_data_prot;
  assign _T_602_bits_qos = Queue_26_io_deq_bits_data_qos;
  assign _T_602_bits_lock = Queue_26_io_deq_bits_data_lock;
  assign _T_602_bits_cache = Queue_26_io_deq_bits_data_cache;
  assign _T_602_bits_size = Queue_26_io_deq_bits_data_size;
  assign _T_602_bits_burst = Queue_26_io_deq_bits_data_burst;
  assign _T_602_bits_id = Queue_26_io_deq_bits_data_id;
  assign _T_602_bits_addr = Queue_26_io_deq_bits_data_addr;
  assign _T_602_bits_len = Queue_26_io_deq_bits_data_len;
  assign _T_857 = {_T_602_bits_id,_T_602_bits_addr,_T_602_bits_len,_T_602_bits_size,_T_602_bits_burst,_T_602_bits_lock,_T_602_bits_cache,_T_602_bits_prot,_T_602_bits_qos};
  assign _T_858 = _T_762_6 ? _T_857 : 60'h0;
  assign _T_608_bits_prot = Queue_27_io_deq_bits_data_prot;
  assign _T_608_bits_qos = Queue_27_io_deq_bits_data_qos;
  assign _T_608_bits_lock = Queue_27_io_deq_bits_data_lock;
  assign _T_608_bits_cache = Queue_27_io_deq_bits_data_cache;
  assign _T_608_bits_size = Queue_27_io_deq_bits_data_size;
  assign _T_608_bits_burst = Queue_27_io_deq_bits_data_burst;
  assign _T_608_bits_id = Queue_27_io_deq_bits_data_id;
  assign _T_608_bits_addr = Queue_27_io_deq_bits_data_addr;
  assign _T_608_bits_len = Queue_27_io_deq_bits_data_len;
  assign _T_866 = {_T_608_bits_id,_T_608_bits_addr,_T_608_bits_len,_T_608_bits_size,_T_608_bits_burst,_T_608_bits_lock,_T_608_bits_cache,_T_608_bits_prot,_T_608_bits_qos};
  assign _T_867 = _T_762_7 ? _T_866 : 60'h0;
  assign _T_868 = _T_804 | _T_813;
  assign _T_869 = _T_868 | _T_822;
  assign _T_870 = _T_869 | _T_831;
  assign _T_871 = _T_870 | _T_840;
  assign _T_872 = _T_871 | _T_849;
  assign _T_873 = _T_872 | _T_858;
  assign _T_874 = _T_873 | _T_867;
  assign _T_888 = plusarg_reader_2_out[0];
  assign _T_891 = _T_889 + 32'h1;
  assign _T_898 = {MaxPeriodFibonacciLFSR_2__EVAL_12,MaxPeriodFibonacciLFSR_2__EVAL_11,MaxPeriodFibonacciLFSR_2__EVAL_3,MaxPeriodFibonacciLFSR_2__EVAL_16,MaxPeriodFibonacciLFSR_2__EVAL_8,MaxPeriodFibonacciLFSR_2__EVAL_10,MaxPeriodFibonacciLFSR_2__EVAL_14,MaxPeriodFibonacciLFSR_2__EVAL_7};
  assign _T_906 = {MaxPeriodFibonacciLFSR_2__EVAL_0,MaxPeriodFibonacciLFSR_2__EVAL_17,MaxPeriodFibonacciLFSR_2__EVAL_1,MaxPeriodFibonacciLFSR_2__EVAL,MaxPeriodFibonacciLFSR_2__EVAL_5,MaxPeriodFibonacciLFSR_2__EVAL_4,MaxPeriodFibonacciLFSR_2__EVAL_6,MaxPeriodFibonacciLFSR_2__EVAL_2,_T_898};
  assign _T_907 = _T_906[0];
  assign _T_908 = _T_906[1];
  assign _T_909 = _T_906[2];
  assign _T_910 = _T_906[3];
  assign _T_911 = _T_906[4];
  assign _T_912 = _T_906[5];
  assign _T_913 = _T_906[6];
  assign _T_914 = _T_906[7];
  assign _T_915 = _T_906[8];
  assign _T_916 = _T_906[9];
  assign _T_917 = _T_906[10];
  assign _T_918 = _T_906[11];
  assign _T_919 = _T_906[12];
  assign _T_920 = _T_906[13];
  assign _T_921 = _T_906[14];
  assign _T_922 = _T_906[15];
  assign _T_930 = {_T_915,_T_916,_T_917,_T_918,_T_919,_T_920,_T_921,_T_922};
  assign _T_938 = {_T_907,_T_908,_T_909,_T_910,_T_911,_T_912,_T_913,_T_914,_T_930};
  assign _GEN_107 = 4'h1 == auto_out_b_bits_id ? 3'h0 : 3'h5;
  assign _GEN_108 = 4'h2 == auto_out_b_bits_id ? 3'h5 : _GEN_107;
  assign _GEN_109 = 4'h3 == auto_out_b_bits_id ? 3'h0 : _GEN_108;
  assign _GEN_110 = 4'h4 == auto_out_b_bits_id ? 3'h2 : _GEN_109;
  assign _GEN_111 = 4'h5 == auto_out_b_bits_id ? 3'h7 : _GEN_110;
  assign _GEN_112 = 4'h6 == auto_out_b_bits_id ? 3'h2 : _GEN_111;
  assign _GEN_113 = 4'h7 == auto_out_b_bits_id ? 3'h5 : _GEN_112;
  assign _GEN_114 = 4'h8 == auto_out_b_bits_id ? 3'h5 : _GEN_113;
  assign _GEN_115 = 4'h9 == auto_out_b_bits_id ? 3'h0 : _GEN_114;
  assign _GEN_116 = 4'ha == auto_out_b_bits_id ? 3'h7 : _GEN_115;
  assign _GEN_117 = 4'hb == auto_out_b_bits_id ? 3'h3 : _GEN_116;
  assign _GEN_118 = 4'hc == auto_out_b_bits_id ? 3'h2 : _GEN_117;
  assign _GEN_119 = 4'hd == auto_out_b_bits_id ? 3'h3 : _GEN_118;
  assign _GEN_120 = 4'he == auto_out_b_bits_id ? 3'h2 : _GEN_119;
  assign _GEN_121 = 4'hf == auto_out_b_bits_id ? 3'h5 : _GEN_120;
  assign _T_950_7 = Queue_36_io_enq_ready;
  assign _T_950_6 = Queue_35_io_enq_ready;
  assign _T_950_5 = Queue_34_io_enq_ready;
  assign _T_950_4 = Queue_33_io_enq_ready;
  assign _T_950_3 = Queue_32_io_enq_ready;
  assign _T_950_2 = Queue_31_io_enq_ready;
  assign _T_950_1 = Queue_30_io_enq_ready;
  assign _T_950_0 = Queue_29_io_enq_ready;
  assign _GEN_123 = 3'h1 == _GEN_121 ? _T_950_1 : _T_950_0;
  assign _GEN_124 = 3'h2 == _GEN_121 ? _T_950_2 : _GEN_123;
  assign _GEN_125 = 3'h3 == _GEN_121 ? _T_950_3 : _GEN_124;
  assign _GEN_126 = 3'h4 == _GEN_121 ? _T_950_4 : _GEN_125;
  assign _GEN_127 = 3'h5 == _GEN_121 ? _T_950_5 : _GEN_126;
  assign _GEN_128 = 3'h6 == _GEN_121 ? _T_950_6 : _GEN_127;
  assign _T_946 = _T_889 + 32'h2;
  assign _T_947 = _T_938[1:0];
  assign _GEN_166 = {{30'd0}, _T_947};
  assign _T_952 = 8'h1 << _GEN_121;
  assign _T_954 = _T_952[0];
  assign _T_955 = _T_952[1];
  assign _T_956 = _T_952[2];
  assign _T_957 = _T_952[3];
  assign _T_958 = _T_952[4];
  assign _T_959 = _T_952[5];
  assign _T_960 = _T_952[6];
  assign _T_961 = _T_952[7];
  assign _T_972 = Queue_29_io_deq_bits_timestamp <= _T_889;
  assign _T_973 = _T_972 | _T_888;
  assign _T_974 = Queue_29_io_deq_valid & _T_973;
  assign _T_970_ready = Queue_37_io_enq_ready;
  assign _T_1020 = _T_1019 == 1'h0;
  assign _T_1014 = Queue_36_io_deq_bits_timestamp <= _T_889;
  assign _T_1015 = _T_1014 | _T_888;
  assign _T_1016 = Queue_36_io_deq_valid & _T_1015;
  assign _T_1008 = Queue_35_io_deq_bits_timestamp <= _T_889;
  assign _T_1009 = _T_1008 | _T_888;
  assign _T_1010 = Queue_35_io_deq_valid & _T_1009;
  assign _T_1002 = Queue_34_io_deq_bits_timestamp <= _T_889;
  assign _T_1003 = _T_1002 | _T_888;
  assign _T_1004 = Queue_34_io_deq_valid & _T_1003;
  assign _T_996 = Queue_33_io_deq_bits_timestamp <= _T_889;
  assign _T_997 = _T_996 | _T_888;
  assign _T_998 = Queue_33_io_deq_valid & _T_997;
  assign _T_990 = Queue_32_io_deq_bits_timestamp <= _T_889;
  assign _T_991 = _T_990 | _T_888;
  assign _T_992 = Queue_32_io_deq_valid & _T_991;
  assign _T_984 = Queue_31_io_deq_bits_timestamp <= _T_889;
  assign _T_985 = _T_984 | _T_888;
  assign _T_986 = Queue_31_io_deq_valid & _T_985;
  assign _T_978 = Queue_30_io_deq_bits_timestamp <= _T_889;
  assign _T_979 = _T_978 | _T_888;
  assign _T_980 = Queue_30_io_deq_valid & _T_979;
  assign _T_1028 = {_T_1016,_T_1010,_T_1004,_T_998,_T_992,_T_986,_T_980,_T_974};
  assign _T_1036 = ~ _T_1035;
  assign _T_1037 = _T_1028 & _T_1036;
  assign _T_1038 = {_T_1037,_T_1016,_T_1010,_T_1004,_T_998,_T_992,_T_986,_T_980,_T_974};
  assign _T_1039 = _T_1038[15:1];
  assign _GEN_167 = {{1'd0}, _T_1039};
  assign _T_1040 = _T_1038 | _GEN_167;
  assign _T_1041 = _T_1040[15:2];
  assign _GEN_168 = {{2'd0}, _T_1041};
  assign _T_1042 = _T_1040 | _GEN_168;
  assign _T_1043 = _T_1042[15:4];
  assign _GEN_169 = {{4'd0}, _T_1043};
  assign _T_1044 = _T_1042 | _GEN_169;
  assign _T_1046 = _T_1044[15:1];
  assign _T_1047 = {_T_1035, 8'h0};
  assign _GEN_170 = {{1'd0}, _T_1046};
  assign _T_1048 = _GEN_170 | _T_1047;
  assign _T_1049 = _T_1048[15:8];
  assign _T_1050 = _T_1048[7:0];
  assign _T_1051 = _T_1049 & _T_1050;
  assign _T_1052 = ~ _T_1051;
  assign _T_1067 = _T_1052[0];
  assign _T_1168_0 = _T_1020 ? _T_1067 : _T_1166_0;
  assign _T_1169 = _T_970_ready & _T_1168_0;
  assign _T_1068 = _T_1052[1];
  assign _T_1168_1 = _T_1020 ? _T_1068 : _T_1166_1;
  assign _T_1170 = _T_970_ready & _T_1168_1;
  assign _T_1069 = _T_1052[2];
  assign _T_1168_2 = _T_1020 ? _T_1069 : _T_1166_2;
  assign _T_1171 = _T_970_ready & _T_1168_2;
  assign _T_1070 = _T_1052[3];
  assign _T_1168_3 = _T_1020 ? _T_1070 : _T_1166_3;
  assign _T_1172 = _T_970_ready & _T_1168_3;
  assign _T_1071 = _T_1052[4];
  assign _T_1168_4 = _T_1020 ? _T_1071 : _T_1166_4;
  assign _T_1173 = _T_970_ready & _T_1168_4;
  assign _T_1072 = _T_1052[5];
  assign _T_1168_5 = _T_1020 ? _T_1072 : _T_1166_5;
  assign _T_1174 = _T_970_ready & _T_1168_5;
  assign _T_1073 = _T_1052[6];
  assign _T_1168_6 = _T_1020 ? _T_1073 : _T_1166_6;
  assign _T_1175 = _T_970_ready & _T_1168_6;
  assign _T_1074 = _T_1052[7];
  assign _T_1168_7 = _T_1020 ? _T_1074 : _T_1166_7;
  assign _T_1176 = _T_970_ready & _T_1168_7;
  assign _T_1021 = _T_1020 & _T_970_ready;
  assign _T_1030 = _T_1028 == _T_1028;
  assign _T_1032 = _T_1030 | reset;
  assign _T_1033 = _T_1032 == 1'h0;
  assign _T_1053 = _T_1028 != 8'h0;
  assign _T_1054 = _T_1021 & _T_1053;
  assign _T_1055 = _T_1052 & _T_1028;
  assign _T_1056 = {_T_1055, 1'h0};
  assign _T_1057 = _T_1056[7:0];
  assign _T_1058 = _T_1055 | _T_1057;
  assign _T_1059 = {_T_1058, 2'h0};
  assign _T_1060 = _T_1059[7:0];
  assign _T_1061 = _T_1058 | _T_1060;
  assign _T_1062 = {_T_1061, 4'h0};
  assign _T_1063 = _T_1062[7:0];
  assign _T_1064 = _T_1061 | _T_1063;
  assign _T_1076 = _T_1067 & _T_974;
  assign _T_1077 = _T_1068 & _T_980;
  assign _T_1078 = _T_1069 & _T_986;
  assign _T_1079 = _T_1070 & _T_992;
  assign _T_1080 = _T_1071 & _T_998;
  assign _T_1081 = _T_1072 & _T_1004;
  assign _T_1082 = _T_1073 & _T_1010;
  assign _T_1083 = _T_1074 & _T_1016;
  assign _T_1086 = _T_1076 | _T_1077;
  assign _T_1087 = _T_1086 | _T_1078;
  assign _T_1088 = _T_1087 | _T_1079;
  assign _T_1089 = _T_1088 | _T_1080;
  assign _T_1090 = _T_1089 | _T_1081;
  assign _T_1091 = _T_1090 | _T_1082;
  assign _T_1092 = _T_1091 | _T_1083;
  assign _T_1094 = _T_1076 == 1'h0;
  assign _T_1097 = _T_1077 == 1'h0;
  assign _T_1098 = _T_1094 | _T_1097;
  assign _T_1099 = _T_1086 == 1'h0;
  assign _T_1100 = _T_1078 == 1'h0;
  assign _T_1101 = _T_1099 | _T_1100;
  assign _T_1102 = _T_1087 == 1'h0;
  assign _T_1103 = _T_1079 == 1'h0;
  assign _T_1104 = _T_1102 | _T_1103;
  assign _T_1105 = _T_1088 == 1'h0;
  assign _T_1106 = _T_1080 == 1'h0;
  assign _T_1107 = _T_1105 | _T_1106;
  assign _T_1108 = _T_1089 == 1'h0;
  assign _T_1109 = _T_1081 == 1'h0;
  assign _T_1110 = _T_1108 | _T_1109;
  assign _T_1111 = _T_1090 == 1'h0;
  assign _T_1112 = _T_1082 == 1'h0;
  assign _T_1113 = _T_1111 | _T_1112;
  assign _T_1114 = _T_1091 == 1'h0;
  assign _T_1115 = _T_1083 == 1'h0;
  assign _T_1116 = _T_1114 | _T_1115;
  assign _T_1118 = _T_1098 & _T_1101;
  assign _T_1119 = _T_1118 & _T_1104;
  assign _T_1120 = _T_1119 & _T_1107;
  assign _T_1121 = _T_1120 & _T_1110;
  assign _T_1122 = _T_1121 & _T_1113;
  assign _T_1123 = _T_1122 & _T_1116;
  assign _T_1125 = _T_1123 | reset;
  assign _T_1126 = _T_1125 == 1'h0;
  assign _T_1127 = _T_974 | _T_980;
  assign _T_1128 = _T_1127 | _T_986;
  assign _T_1129 = _T_1128 | _T_992;
  assign _T_1130 = _T_1129 | _T_998;
  assign _T_1131 = _T_1130 | _T_1004;
  assign _T_1132 = _T_1131 | _T_1010;
  assign _T_1133 = _T_1132 | _T_1016;
  assign _T_1134 = _T_1133 == 1'h0;
  assign _T_1142 = _T_1134 | _T_1092;
  assign _T_1144 = _T_1142 | reset;
  assign _T_1145 = _T_1144 == 1'h0;
  assign _T_1184 = _T_1166_0 ? _T_974 : 1'h0;
  assign _T_1185 = _T_1166_1 ? _T_980 : 1'h0;
  assign _T_1192 = _T_1184 | _T_1185;
  assign _T_1186 = _T_1166_2 ? _T_986 : 1'h0;
  assign _T_1193 = _T_1192 | _T_1186;
  assign _T_1187 = _T_1166_3 ? _T_992 : 1'h0;
  assign _T_1194 = _T_1193 | _T_1187;
  assign _T_1188 = _T_1166_4 ? _T_998 : 1'h0;
  assign _T_1195 = _T_1194 | _T_1188;
  assign _T_1189 = _T_1166_5 ? _T_1004 : 1'h0;
  assign _T_1196 = _T_1195 | _T_1189;
  assign _T_1190 = _T_1166_6 ? _T_1010 : 1'h0;
  assign _T_1197 = _T_1196 | _T_1190;
  assign _T_1191 = _T_1166_7 ? _T_1016 : 1'h0;
  assign _T_1198 = _T_1197 | _T_1191;
  assign _T_1200 = _T_1020 ? _T_1133 : _T_1198;
  assign _T_1161 = _T_970_ready & _T_1200;
  assign _T_1163 = _T_1019 - _T_1161;
  assign _T_1167_0 = _T_1020 ? _T_1076 : _T_1166_0;
  assign _T_1167_1 = _T_1020 ? _T_1077 : _T_1166_1;
  assign _T_1167_2 = _T_1020 ? _T_1078 : _T_1166_2;
  assign _T_1167_3 = _T_1020 ? _T_1079 : _T_1166_3;
  assign _T_1167_4 = _T_1020 ? _T_1080 : _T_1166_4;
  assign _T_1167_5 = _T_1020 ? _T_1081 : _T_1166_5;
  assign _T_1167_6 = _T_1020 ? _T_1082 : _T_1166_6;
  assign _T_1167_7 = _T_1020 ? _T_1083 : _T_1166_7;
  assign _T_971_bits_id = Queue_29_io_deq_bits_data_id;
  assign _T_971_bits_resp = Queue_29_io_deq_bits_data_resp;
  assign _T_1201 = {_T_971_bits_id,_T_971_bits_resp};
  assign _T_1202 = _T_1167_0 ? _T_1201 : 6'h0;
  assign _T_977_bits_id = Queue_30_io_deq_bits_data_id;
  assign _T_977_bits_resp = Queue_30_io_deq_bits_data_resp;
  assign _T_1203 = {_T_977_bits_id,_T_977_bits_resp};
  assign _T_1204 = _T_1167_1 ? _T_1203 : 6'h0;
  assign _T_983_bits_id = Queue_31_io_deq_bits_data_id;
  assign _T_983_bits_resp = Queue_31_io_deq_bits_data_resp;
  assign _T_1205 = {_T_983_bits_id,_T_983_bits_resp};
  assign _T_1206 = _T_1167_2 ? _T_1205 : 6'h0;
  assign _T_989_bits_id = Queue_32_io_deq_bits_data_id;
  assign _T_989_bits_resp = Queue_32_io_deq_bits_data_resp;
  assign _T_1207 = {_T_989_bits_id,_T_989_bits_resp};
  assign _T_1208 = _T_1167_3 ? _T_1207 : 6'h0;
  assign _T_995_bits_id = Queue_33_io_deq_bits_data_id;
  assign _T_995_bits_resp = Queue_33_io_deq_bits_data_resp;
  assign _T_1209 = {_T_995_bits_id,_T_995_bits_resp};
  assign _T_1210 = _T_1167_4 ? _T_1209 : 6'h0;
  assign _T_1001_bits_id = Queue_34_io_deq_bits_data_id;
  assign _T_1001_bits_resp = Queue_34_io_deq_bits_data_resp;
  assign _T_1211 = {_T_1001_bits_id,_T_1001_bits_resp};
  assign _T_1212 = _T_1167_5 ? _T_1211 : 6'h0;
  assign _T_1007_bits_id = Queue_35_io_deq_bits_data_id;
  assign _T_1007_bits_resp = Queue_35_io_deq_bits_data_resp;
  assign _T_1213 = {_T_1007_bits_id,_T_1007_bits_resp};
  assign _T_1214 = _T_1167_6 ? _T_1213 : 6'h0;
  assign _T_1013_bits_id = Queue_36_io_deq_bits_data_id;
  assign _T_1013_bits_resp = Queue_36_io_deq_bits_data_resp;
  assign _T_1215 = {_T_1013_bits_id,_T_1013_bits_resp};
  assign _T_1216 = _T_1167_7 ? _T_1215 : 6'h0;
  assign _T_1217 = _T_1202 | _T_1204;
  assign _T_1218 = _T_1217 | _T_1206;
  assign _T_1219 = _T_1218 | _T_1208;
  assign _T_1220 = _T_1219 | _T_1210;
  assign _T_1221 = _T_1220 | _T_1212;
  assign _T_1222 = _T_1221 | _T_1214;
  assign _T_1223 = _T_1222 | _T_1216;
  assign _T_1230 = plusarg_reader_3_out[0];
  assign _T_1233 = _T_1231 + 32'h1;
  assign _T_1240 = {MaxPeriodFibonacciLFSR_3__EVAL_12,MaxPeriodFibonacciLFSR_3__EVAL_11,MaxPeriodFibonacciLFSR_3__EVAL_3,MaxPeriodFibonacciLFSR_3__EVAL_16,MaxPeriodFibonacciLFSR_3__EVAL_8,MaxPeriodFibonacciLFSR_3__EVAL_10,MaxPeriodFibonacciLFSR_3__EVAL_14,MaxPeriodFibonacciLFSR_3__EVAL_7};
  assign _T_1248 = {MaxPeriodFibonacciLFSR_3__EVAL_0,MaxPeriodFibonacciLFSR_3__EVAL_17,MaxPeriodFibonacciLFSR_3__EVAL_1,MaxPeriodFibonacciLFSR_3__EVAL,MaxPeriodFibonacciLFSR_3__EVAL_5,MaxPeriodFibonacciLFSR_3__EVAL_4,MaxPeriodFibonacciLFSR_3__EVAL_6,MaxPeriodFibonacciLFSR_3__EVAL_2,_T_1240};
  assign _T_1249 = _T_1248[0];
  assign _T_1250 = _T_1248[1];
  assign _T_1251 = _T_1248[2];
  assign _T_1252 = _T_1248[3];
  assign _T_1253 = _T_1248[4];
  assign _T_1254 = _T_1248[5];
  assign _T_1255 = _T_1248[6];
  assign _T_1256 = _T_1248[7];
  assign _T_1257 = _T_1248[8];
  assign _T_1258 = _T_1248[9];
  assign _T_1259 = _T_1248[10];
  assign _T_1260 = _T_1248[11];
  assign _T_1261 = _T_1248[12];
  assign _T_1262 = _T_1248[13];
  assign _T_1263 = _T_1248[14];
  assign _T_1264 = _T_1248[15];
  assign _T_1272 = {_T_1257,_T_1258,_T_1259,_T_1260,_T_1261,_T_1262,_T_1263,_T_1264};
  assign _T_1280 = {_T_1249,_T_1250,_T_1251,_T_1252,_T_1253,_T_1254,_T_1255,_T_1256,_T_1272};
  assign _GEN_132 = 4'h1 == auto_out_r_bits_id ? 3'h0 : 3'h5;
  assign _GEN_133 = 4'h2 == auto_out_r_bits_id ? 3'h5 : _GEN_132;
  assign _GEN_134 = 4'h3 == auto_out_r_bits_id ? 3'h0 : _GEN_133;
  assign _GEN_135 = 4'h4 == auto_out_r_bits_id ? 3'h2 : _GEN_134;
  assign _GEN_136 = 4'h5 == auto_out_r_bits_id ? 3'h7 : _GEN_135;
  assign _GEN_137 = 4'h6 == auto_out_r_bits_id ? 3'h2 : _GEN_136;
  assign _GEN_138 = 4'h7 == auto_out_r_bits_id ? 3'h5 : _GEN_137;
  assign _GEN_139 = 4'h8 == auto_out_r_bits_id ? 3'h5 : _GEN_138;
  assign _GEN_140 = 4'h9 == auto_out_r_bits_id ? 3'h0 : _GEN_139;
  assign _GEN_141 = 4'ha == auto_out_r_bits_id ? 3'h7 : _GEN_140;
  assign _GEN_142 = 4'hb == auto_out_r_bits_id ? 3'h3 : _GEN_141;
  assign _GEN_143 = 4'hc == auto_out_r_bits_id ? 3'h2 : _GEN_142;
  assign _GEN_144 = 4'hd == auto_out_r_bits_id ? 3'h3 : _GEN_143;
  assign _GEN_145 = 4'he == auto_out_r_bits_id ? 3'h2 : _GEN_144;
  assign _GEN_146 = 4'hf == auto_out_r_bits_id ? 3'h5 : _GEN_145;
  assign _T_1292_7 = Queue_45_io_enq_ready;
  assign _T_1292_6 = Queue_44_io_enq_ready;
  assign _T_1292_5 = Queue_43_io_enq_ready;
  assign _T_1292_4 = Queue_42_io_enq_ready;
  assign _T_1292_3 = Queue_41_io_enq_ready;
  assign _T_1292_2 = Queue_40_io_enq_ready;
  assign _T_1292_1 = Queue_39_io_enq_ready;
  assign _T_1292_0 = Queue_38_io_enq_ready;
  assign _GEN_148 = 3'h1 == _GEN_146 ? _T_1292_1 : _T_1292_0;
  assign _GEN_149 = 3'h2 == _GEN_146 ? _T_1292_2 : _GEN_148;
  assign _GEN_150 = 3'h3 == _GEN_146 ? _T_1292_3 : _GEN_149;
  assign _GEN_151 = 3'h4 == _GEN_146 ? _T_1292_4 : _GEN_150;
  assign _GEN_152 = 3'h5 == _GEN_146 ? _T_1292_5 : _GEN_151;
  assign _GEN_153 = 3'h6 == _GEN_146 ? _T_1292_6 : _GEN_152;
  assign _T_1288 = _T_1231 + 32'h2;
  assign _T_1289 = _T_1280[1:0];
  assign _GEN_171 = {{30'd0}, _T_1289};
  assign _T_1294 = 8'h1 << _GEN_146;
  assign _T_1296 = _T_1294[0];
  assign _T_1297 = _T_1294[1];
  assign _T_1298 = _T_1294[2];
  assign _T_1299 = _T_1294[3];
  assign _T_1300 = _T_1294[4];
  assign _T_1301 = _T_1294[5];
  assign _T_1302 = _T_1294[6];
  assign _T_1303 = _T_1294[7];
  assign _T_1314 = Queue_38_io_deq_bits_timestamp <= _T_1231;
  assign _T_1315 = _T_1314 | _T_1230;
  assign _T_1316 = Queue_38_io_deq_valid & _T_1315;
  assign _T_1312_ready = Queue_46_io_enq_ready;
  assign _T_1362 = _T_1361 == 1'h0;
  assign _T_1356 = Queue_45_io_deq_bits_timestamp <= _T_1231;
  assign _T_1357 = _T_1356 | _T_1230;
  assign _T_1358 = Queue_45_io_deq_valid & _T_1357;
  assign _T_1350 = Queue_44_io_deq_bits_timestamp <= _T_1231;
  assign _T_1351 = _T_1350 | _T_1230;
  assign _T_1352 = Queue_44_io_deq_valid & _T_1351;
  assign _T_1344 = Queue_43_io_deq_bits_timestamp <= _T_1231;
  assign _T_1345 = _T_1344 | _T_1230;
  assign _T_1346 = Queue_43_io_deq_valid & _T_1345;
  assign _T_1338 = Queue_42_io_deq_bits_timestamp <= _T_1231;
  assign _T_1339 = _T_1338 | _T_1230;
  assign _T_1340 = Queue_42_io_deq_valid & _T_1339;
  assign _T_1332 = Queue_41_io_deq_bits_timestamp <= _T_1231;
  assign _T_1333 = _T_1332 | _T_1230;
  assign _T_1334 = Queue_41_io_deq_valid & _T_1333;
  assign _T_1326 = Queue_40_io_deq_bits_timestamp <= _T_1231;
  assign _T_1327 = _T_1326 | _T_1230;
  assign _T_1328 = Queue_40_io_deq_valid & _T_1327;
  assign _T_1320 = Queue_39_io_deq_bits_timestamp <= _T_1231;
  assign _T_1321 = _T_1320 | _T_1230;
  assign _T_1322 = Queue_39_io_deq_valid & _T_1321;
  assign _T_1370 = {_T_1358,_T_1352,_T_1346,_T_1340,_T_1334,_T_1328,_T_1322,_T_1316};
  assign _T_1378 = ~ _T_1377;
  assign _T_1379 = _T_1370 & _T_1378;
  assign _T_1380 = {_T_1379,_T_1358,_T_1352,_T_1346,_T_1340,_T_1334,_T_1328,_T_1322,_T_1316};
  assign _T_1381 = _T_1380[15:1];
  assign _GEN_172 = {{1'd0}, _T_1381};
  assign _T_1382 = _T_1380 | _GEN_172;
  assign _T_1383 = _T_1382[15:2];
  assign _GEN_173 = {{2'd0}, _T_1383};
  assign _T_1384 = _T_1382 | _GEN_173;
  assign _T_1385 = _T_1384[15:4];
  assign _GEN_174 = {{4'd0}, _T_1385};
  assign _T_1386 = _T_1384 | _GEN_174;
  assign _T_1388 = _T_1386[15:1];
  assign _T_1389 = {_T_1377, 8'h0};
  assign _GEN_175 = {{1'd0}, _T_1388};
  assign _T_1390 = _GEN_175 | _T_1389;
  assign _T_1391 = _T_1390[15:8];
  assign _T_1392 = _T_1390[7:0];
  assign _T_1393 = _T_1391 & _T_1392;
  assign _T_1394 = ~ _T_1393;
  assign _T_1409 = _T_1394[0];
  assign _T_1510_0 = _T_1362 ? _T_1409 : _T_1508_0;
  assign _T_1511 = _T_1312_ready & _T_1510_0;
  assign _T_1410 = _T_1394[1];
  assign _T_1510_1 = _T_1362 ? _T_1410 : _T_1508_1;
  assign _T_1512 = _T_1312_ready & _T_1510_1;
  assign _T_1411 = _T_1394[2];
  assign _T_1510_2 = _T_1362 ? _T_1411 : _T_1508_2;
  assign _T_1513 = _T_1312_ready & _T_1510_2;
  assign _T_1412 = _T_1394[3];
  assign _T_1510_3 = _T_1362 ? _T_1412 : _T_1508_3;
  assign _T_1514 = _T_1312_ready & _T_1510_3;
  assign _T_1413 = _T_1394[4];
  assign _T_1510_4 = _T_1362 ? _T_1413 : _T_1508_4;
  assign _T_1515 = _T_1312_ready & _T_1510_4;
  assign _T_1414 = _T_1394[5];
  assign _T_1510_5 = _T_1362 ? _T_1414 : _T_1508_5;
  assign _T_1516 = _T_1312_ready & _T_1510_5;
  assign _T_1415 = _T_1394[6];
  assign _T_1510_6 = _T_1362 ? _T_1415 : _T_1508_6;
  assign _T_1517 = _T_1312_ready & _T_1510_6;
  assign _T_1416 = _T_1394[7];
  assign _T_1510_7 = _T_1362 ? _T_1416 : _T_1508_7;
  assign _T_1518 = _T_1312_ready & _T_1510_7;
  assign _T_1363 = _T_1362 & _T_1312_ready;
  assign _T_1372 = _T_1370 == _T_1370;
  assign _T_1374 = _T_1372 | reset;
  assign _T_1375 = _T_1374 == 1'h0;
  assign _T_1395 = _T_1370 != 8'h0;
  assign _T_1396 = _T_1363 & _T_1395;
  assign _T_1397 = _T_1394 & _T_1370;
  assign _T_1398 = {_T_1397, 1'h0};
  assign _T_1399 = _T_1398[7:0];
  assign _T_1400 = _T_1397 | _T_1399;
  assign _T_1401 = {_T_1400, 2'h0};
  assign _T_1402 = _T_1401[7:0];
  assign _T_1403 = _T_1400 | _T_1402;
  assign _T_1404 = {_T_1403, 4'h0};
  assign _T_1405 = _T_1404[7:0];
  assign _T_1406 = _T_1403 | _T_1405;
  assign _T_1418 = _T_1409 & _T_1316;
  assign _T_1419 = _T_1410 & _T_1322;
  assign _T_1420 = _T_1411 & _T_1328;
  assign _T_1421 = _T_1412 & _T_1334;
  assign _T_1422 = _T_1413 & _T_1340;
  assign _T_1423 = _T_1414 & _T_1346;
  assign _T_1424 = _T_1415 & _T_1352;
  assign _T_1425 = _T_1416 & _T_1358;
  assign _T_1428 = _T_1418 | _T_1419;
  assign _T_1429 = _T_1428 | _T_1420;
  assign _T_1430 = _T_1429 | _T_1421;
  assign _T_1431 = _T_1430 | _T_1422;
  assign _T_1432 = _T_1431 | _T_1423;
  assign _T_1433 = _T_1432 | _T_1424;
  assign _T_1434 = _T_1433 | _T_1425;
  assign _T_1436 = _T_1418 == 1'h0;
  assign _T_1439 = _T_1419 == 1'h0;
  assign _T_1440 = _T_1436 | _T_1439;
  assign _T_1441 = _T_1428 == 1'h0;
  assign _T_1442 = _T_1420 == 1'h0;
  assign _T_1443 = _T_1441 | _T_1442;
  assign _T_1444 = _T_1429 == 1'h0;
  assign _T_1445 = _T_1421 == 1'h0;
  assign _T_1446 = _T_1444 | _T_1445;
  assign _T_1447 = _T_1430 == 1'h0;
  assign _T_1448 = _T_1422 == 1'h0;
  assign _T_1449 = _T_1447 | _T_1448;
  assign _T_1450 = _T_1431 == 1'h0;
  assign _T_1451 = _T_1423 == 1'h0;
  assign _T_1452 = _T_1450 | _T_1451;
  assign _T_1453 = _T_1432 == 1'h0;
  assign _T_1454 = _T_1424 == 1'h0;
  assign _T_1455 = _T_1453 | _T_1454;
  assign _T_1456 = _T_1433 == 1'h0;
  assign _T_1457 = _T_1425 == 1'h0;
  assign _T_1458 = _T_1456 | _T_1457;
  assign _T_1460 = _T_1440 & _T_1443;
  assign _T_1461 = _T_1460 & _T_1446;
  assign _T_1462 = _T_1461 & _T_1449;
  assign _T_1463 = _T_1462 & _T_1452;
  assign _T_1464 = _T_1463 & _T_1455;
  assign _T_1465 = _T_1464 & _T_1458;
  assign _T_1467 = _T_1465 | reset;
  assign _T_1468 = _T_1467 == 1'h0;
  assign _T_1469 = _T_1316 | _T_1322;
  assign _T_1470 = _T_1469 | _T_1328;
  assign _T_1471 = _T_1470 | _T_1334;
  assign _T_1472 = _T_1471 | _T_1340;
  assign _T_1473 = _T_1472 | _T_1346;
  assign _T_1474 = _T_1473 | _T_1352;
  assign _T_1475 = _T_1474 | _T_1358;
  assign _T_1476 = _T_1475 == 1'h0;
  assign _T_1484 = _T_1476 | _T_1434;
  assign _T_1486 = _T_1484 | reset;
  assign _T_1487 = _T_1486 == 1'h0;
  assign _T_1526 = _T_1508_0 ? _T_1316 : 1'h0;
  assign _T_1527 = _T_1508_1 ? _T_1322 : 1'h0;
  assign _T_1534 = _T_1526 | _T_1527;
  assign _T_1528 = _T_1508_2 ? _T_1328 : 1'h0;
  assign _T_1535 = _T_1534 | _T_1528;
  assign _T_1529 = _T_1508_3 ? _T_1334 : 1'h0;
  assign _T_1536 = _T_1535 | _T_1529;
  assign _T_1530 = _T_1508_4 ? _T_1340 : 1'h0;
  assign _T_1537 = _T_1536 | _T_1530;
  assign _T_1531 = _T_1508_5 ? _T_1346 : 1'h0;
  assign _T_1538 = _T_1537 | _T_1531;
  assign _T_1532 = _T_1508_6 ? _T_1352 : 1'h0;
  assign _T_1539 = _T_1538 | _T_1532;
  assign _T_1533 = _T_1508_7 ? _T_1358 : 1'h0;
  assign _T_1540 = _T_1539 | _T_1533;
  assign _T_1542 = _T_1362 ? _T_1475 : _T_1540;
  assign _T_1503 = _T_1312_ready & _T_1542;
  assign _T_1505 = _T_1361 - _T_1503;
  assign _T_1509_0 = _T_1362 ? _T_1418 : _T_1508_0;
  assign _T_1509_1 = _T_1362 ? _T_1419 : _T_1508_1;
  assign _T_1509_2 = _T_1362 ? _T_1420 : _T_1508_2;
  assign _T_1509_3 = _T_1362 ? _T_1421 : _T_1508_3;
  assign _T_1509_4 = _T_1362 ? _T_1422 : _T_1508_4;
  assign _T_1509_5 = _T_1362 ? _T_1423 : _T_1508_5;
  assign _T_1509_6 = _T_1362 ? _T_1424 : _T_1508_6;
  assign _T_1509_7 = _T_1362 ? _T_1425 : _T_1508_7;
  assign _T_1313_bits_resp = Queue_38_io_deq_bits_data_resp;
  assign _T_1313_bits_last = Queue_38_io_deq_bits_data_last;
  assign _T_1313_bits_id = Queue_38_io_deq_bits_data_id;
  assign _T_1313_bits_data = Queue_38_io_deq_bits_data_data;
  assign _T_1545 = {_T_1313_bits_id,_T_1313_bits_data,_T_1313_bits_resp,_T_1313_bits_last};
  assign _T_1546 = _T_1509_0 ? _T_1545 : 39'h0;
  assign _T_1319_bits_resp = Queue_39_io_deq_bits_data_resp;
  assign _T_1319_bits_last = Queue_39_io_deq_bits_data_last;
  assign _T_1319_bits_id = Queue_39_io_deq_bits_data_id;
  assign _T_1319_bits_data = Queue_39_io_deq_bits_data_data;
  assign _T_1549 = {_T_1319_bits_id,_T_1319_bits_data,_T_1319_bits_resp,_T_1319_bits_last};
  assign _T_1550 = _T_1509_1 ? _T_1549 : 39'h0;
  assign _T_1325_bits_resp = Queue_40_io_deq_bits_data_resp;
  assign _T_1325_bits_last = Queue_40_io_deq_bits_data_last;
  assign _T_1325_bits_id = Queue_40_io_deq_bits_data_id;
  assign _T_1325_bits_data = Queue_40_io_deq_bits_data_data;
  assign _T_1553 = {_T_1325_bits_id,_T_1325_bits_data,_T_1325_bits_resp,_T_1325_bits_last};
  assign _T_1554 = _T_1509_2 ? _T_1553 : 39'h0;
  assign _T_1331_bits_resp = Queue_41_io_deq_bits_data_resp;
  assign _T_1331_bits_last = Queue_41_io_deq_bits_data_last;
  assign _T_1331_bits_id = Queue_41_io_deq_bits_data_id;
  assign _T_1331_bits_data = Queue_41_io_deq_bits_data_data;
  assign _T_1557 = {_T_1331_bits_id,_T_1331_bits_data,_T_1331_bits_resp,_T_1331_bits_last};
  assign _T_1558 = _T_1509_3 ? _T_1557 : 39'h0;
  assign _T_1337_bits_resp = Queue_42_io_deq_bits_data_resp;
  assign _T_1337_bits_last = Queue_42_io_deq_bits_data_last;
  assign _T_1337_bits_id = Queue_42_io_deq_bits_data_id;
  assign _T_1337_bits_data = Queue_42_io_deq_bits_data_data;
  assign _T_1561 = {_T_1337_bits_id,_T_1337_bits_data,_T_1337_bits_resp,_T_1337_bits_last};
  assign _T_1562 = _T_1509_4 ? _T_1561 : 39'h0;
  assign _T_1343_bits_resp = Queue_43_io_deq_bits_data_resp;
  assign _T_1343_bits_last = Queue_43_io_deq_bits_data_last;
  assign _T_1343_bits_id = Queue_43_io_deq_bits_data_id;
  assign _T_1343_bits_data = Queue_43_io_deq_bits_data_data;
  assign _T_1565 = {_T_1343_bits_id,_T_1343_bits_data,_T_1343_bits_resp,_T_1343_bits_last};
  assign _T_1566 = _T_1509_5 ? _T_1565 : 39'h0;
  assign _T_1349_bits_resp = Queue_44_io_deq_bits_data_resp;
  assign _T_1349_bits_last = Queue_44_io_deq_bits_data_last;
  assign _T_1349_bits_id = Queue_44_io_deq_bits_data_id;
  assign _T_1349_bits_data = Queue_44_io_deq_bits_data_data;
  assign _T_1569 = {_T_1349_bits_id,_T_1349_bits_data,_T_1349_bits_resp,_T_1349_bits_last};
  assign _T_1570 = _T_1509_6 ? _T_1569 : 39'h0;
  assign _T_1355_bits_resp = Queue_45_io_deq_bits_data_resp;
  assign _T_1355_bits_last = Queue_45_io_deq_bits_data_last;
  assign _T_1355_bits_id = Queue_45_io_deq_bits_data_id;
  assign _T_1355_bits_data = Queue_45_io_deq_bits_data_data;
  assign _T_1573 = {_T_1355_bits_id,_T_1355_bits_data,_T_1355_bits_resp,_T_1355_bits_last};
  assign _T_1574 = _T_1509_7 ? _T_1573 : 39'h0;
  assign _T_1575 = _T_1546 | _T_1550;
  assign _T_1576 = _T_1575 | _T_1554;
  assign _T_1577 = _T_1576 | _T_1558;
  assign _T_1578 = _T_1577 | _T_1562;
  assign _T_1579 = _T_1578 | _T_1566;
  assign _T_1580 = _T_1579 | _T_1570;
  assign _T_1581 = _T_1580 | _T_1574;
  assign auto_in_aw_ready = Queue_io_enq_ready & _T_65;
  assign auto_in_w_ready = _GEN_48 & _T_4_valid;
  assign auto_in_b_valid = Queue_37_io_deq_valid;
  assign auto_in_b_bits_id = Queue_37_io_deq_bits_id;
  assign auto_in_b_bits_resp = Queue_37_io_deq_bits_resp;
  assign auto_in_ar_ready = _GEN_104 & _T_536;
  assign auto_in_r_valid = Queue_46_io_deq_valid;
  assign auto_in_r_bits_id = Queue_46_io_deq_bits_id;
  assign auto_in_r_bits_data = Queue_46_io_deq_bits_data;
  assign auto_in_r_bits_resp = Queue_46_io_deq_bits_resp;
  assign auto_in_r_bits_last = Queue_46_io_deq_bits_last;
  assign auto_out_aw_valid = Queue_11_io_deq_valid;
  assign auto_out_aw_bits_id = Queue_11_io_deq_bits_id;
  assign auto_out_aw_bits_addr = Queue_11_io_deq_bits_addr;
  assign auto_out_aw_bits_len = Queue_11_io_deq_bits_len;
  assign auto_out_aw_bits_size = Queue_11_io_deq_bits_size;
  assign auto_out_aw_bits_burst = Queue_11_io_deq_bits_burst;
  assign auto_out_w_valid = _T_414_valid & _GEN_80;
  assign auto_out_w_bits_data = 3'h7 == _T_414_bits ? _T_451_7_data : _GEN_67;
  assign auto_out_w_bits_strb = 3'h7 == _T_414_bits ? _T_451_7_strb : _GEN_68;
  assign auto_out_w_bits_last = 3'h7 == _T_414_bits ? _T_451_7_last : _GEN_69;
  assign auto_out_b_ready = 3'h7 == _GEN_121 ? _T_950_7 : _GEN_128;
  assign auto_out_ar_valid = Queue_28_io_deq_valid;
  assign auto_out_ar_bits_id = Queue_28_io_deq_bits_id;
  assign auto_out_ar_bits_addr = Queue_28_io_deq_bits_addr;
  assign auto_out_ar_bits_len = Queue_28_io_deq_bits_len;
  assign auto_out_ar_bits_size = Queue_28_io_deq_bits_size;
  assign auto_out_ar_bits_burst = Queue_28_io_deq_bits_burst;
  assign auto_out_r_ready = 3'h7 == _GEN_146 ? _T_1292_7 : _GEN_153;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_aw_valid & _T_65;
  assign Queue_io_enq_bits = 4'hf == auto_in_aw_bits_id ? 3'h5 : _GEN_14;
  assign Queue_io_deq_ready = _T_419 & auto_in_w_valid;
  assign MaxPeriodFibonacciLFSR__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR__EVAL_9 = 1'h1;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_63 & _T_75;
  assign Queue_1_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_1_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_1_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_1_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_1_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_1_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_1_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_1_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_1_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_1_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_1_io_deq_ready = _T_290 & _T_94;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = _T_63 & _T_76;
  assign Queue_2_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_2_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_2_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_2_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_2_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_2_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_2_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_2_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_2_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_2_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_2_io_deq_ready = _T_291 & _T_100;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = _T_63 & _T_77;
  assign Queue_3_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_3_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_3_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_3_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_3_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_3_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_3_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_3_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_3_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_3_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_3_io_deq_ready = _T_292 & _T_106;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = _T_63 & _T_78;
  assign Queue_4_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_4_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_4_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_4_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_4_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_4_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_4_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_4_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_4_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_4_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_4_io_deq_ready = _T_293 & _T_112;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_5_io_enq_valid = _T_63 & _T_79;
  assign Queue_5_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_5_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_5_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_5_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_5_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_5_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_5_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_5_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_5_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_5_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_5_io_deq_ready = _T_294 & _T_118;
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_6_io_enq_valid = _T_63 & _T_80;
  assign Queue_6_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_6_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_6_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_6_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_6_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_6_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_6_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_6_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_6_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_6_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_6_io_deq_ready = _T_295 & _T_124;
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_7_io_enq_valid = _T_63 & _T_81;
  assign Queue_7_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_7_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_7_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_7_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_7_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_7_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_7_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_7_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_7_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_7_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_7_io_deq_ready = _T_296 & _T_130;
  assign Queue_8_clock = clock;
  assign Queue_8_reset = reset;
  assign Queue_8_io_enq_valid = _T_63 & _T_82;
  assign Queue_8_io_enq_bits_data_id = auto_in_aw_bits_id;
  assign Queue_8_io_enq_bits_data_addr = auto_in_aw_bits_addr;
  assign Queue_8_io_enq_bits_data_len = auto_in_aw_bits_len;
  assign Queue_8_io_enq_bits_data_size = auto_in_aw_bits_size;
  assign Queue_8_io_enq_bits_data_burst = auto_in_aw_bits_burst;
  assign Queue_8_io_enq_bits_data_lock = auto_in_aw_bits_lock;
  assign Queue_8_io_enq_bits_data_cache = auto_in_aw_bits_cache;
  assign Queue_8_io_enq_bits_data_prot = auto_in_aw_bits_prot;
  assign Queue_8_io_enq_bits_data_qos = auto_in_aw_bits_qos;
  assign Queue_8_io_enq_bits_timestamp = _T_67 + _GEN_156;
  assign Queue_8_io_deq_ready = _T_297 & _T_136;
  assign Queue_9_clock = clock;
  assign Queue_9_reset = reset;
  assign Queue_9_io_enq_valid = _T_141 ? _T_254 : _T_319;
  assign Queue_9_io_enq_bits_id = _T_400[59:56];
  assign Queue_9_io_enq_bits_addr = _T_400[55:25];
  assign Queue_9_io_enq_bits_len = _T_400[24:17];
  assign Queue_9_io_enq_bits_size = _T_400[16:14];
  assign Queue_9_io_enq_bits_burst = _T_400[13:12];
  assign Queue_9_io_deq_ready = Queue_10_io_enq_ready & _T_413_ready;
  assign Queue_10_clock = clock;
  assign Queue_10_reset = reset;
  assign Queue_10_io_enq_valid = _T_412_valid & _T_413_ready;
  assign Queue_10_io_enq_bits = 4'hf == _T_412_bits_id ? 3'h5 : _GEN_39;
  assign Queue_10_io_deq_ready = _T_452 & auto_out_w_ready;
  assign Queue_11_clock = clock;
  assign Queue_11_reset = reset;
  assign Queue_11_io_enq_valid = _T_412_valid & Queue_10_io_enq_ready;
  assign Queue_11_io_enq_bits_id = Queue_9_io_deq_bits_id;
  assign Queue_11_io_enq_bits_addr = Queue_9_io_deq_bits_addr;
  assign Queue_11_io_enq_bits_len = Queue_9_io_deq_bits_len;
  assign Queue_11_io_enq_bits_size = Queue_9_io_deq_bits_size;
  assign Queue_11_io_enq_bits_burst = Queue_9_io_deq_bits_burst;
  assign Queue_11_io_deq_ready = auto_out_aw_ready;
  assign Queue_12_clock = clock;
  assign Queue_12_reset = reset;
  assign Queue_12_io_enq_valid = _T_433 & _T_425;
  assign Queue_12_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_12_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_12_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_12_io_deq_ready = _T_466 & _T_458;
  assign Queue_13_clock = clock;
  assign Queue_13_reset = reset;
  assign Queue_13_io_enq_valid = _T_433 & _T_426;
  assign Queue_13_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_13_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_13_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_13_io_deq_ready = _T_466 & _T_459;
  assign Queue_14_clock = clock;
  assign Queue_14_reset = reset;
  assign Queue_14_io_enq_valid = _T_433 & _T_427;
  assign Queue_14_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_14_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_14_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_14_io_deq_ready = _T_466 & _T_460;
  assign Queue_15_clock = clock;
  assign Queue_15_reset = reset;
  assign Queue_15_io_enq_valid = _T_433 & _T_428;
  assign Queue_15_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_15_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_15_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_15_io_deq_ready = _T_466 & _T_461;
  assign Queue_16_clock = clock;
  assign Queue_16_reset = reset;
  assign Queue_16_io_enq_valid = _T_433 & _T_429;
  assign Queue_16_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_16_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_16_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_16_io_deq_ready = _T_466 & _T_462;
  assign Queue_17_clock = clock;
  assign Queue_17_reset = reset;
  assign Queue_17_io_enq_valid = _T_433 & _T_430;
  assign Queue_17_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_17_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_17_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_17_io_deq_ready = _T_466 & _T_463;
  assign Queue_18_clock = clock;
  assign Queue_18_reset = reset;
  assign Queue_18_io_enq_valid = _T_433 & _T_431;
  assign Queue_18_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_18_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_18_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_18_io_deq_ready = _T_466 & _T_464;
  assign Queue_19_clock = clock;
  assign Queue_19_reset = reset;
  assign Queue_19_io_enq_valid = _T_433 & _T_432;
  assign Queue_19_io_enq_bits_data = auto_in_w_bits_data;
  assign Queue_19_io_enq_bits_strb = auto_in_w_bits_strb;
  assign Queue_19_io_enq_bits_last = auto_in_w_bits_last;
  assign Queue_19_io_deq_ready = _T_466 & _T_465;
  assign MaxPeriodFibonacciLFSR_1__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR_1__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR_1__EVAL_9 = 1'h1;
  assign Queue_20_clock = clock;
  assign Queue_20_reset = reset;
  assign Queue_20_io_enq_valid = _T_537 & _T_549;
  assign Queue_20_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_20_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_20_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_20_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_20_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_20_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_20_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_20_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_20_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_20_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_20_io_deq_ready = _T_764 & _T_568;
  assign Queue_21_clock = clock;
  assign Queue_21_reset = reset;
  assign Queue_21_io_enq_valid = _T_537 & _T_550;
  assign Queue_21_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_21_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_21_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_21_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_21_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_21_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_21_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_21_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_21_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_21_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_21_io_deq_ready = _T_765 & _T_574;
  assign Queue_22_clock = clock;
  assign Queue_22_reset = reset;
  assign Queue_22_io_enq_valid = _T_537 & _T_551;
  assign Queue_22_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_22_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_22_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_22_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_22_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_22_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_22_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_22_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_22_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_22_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_22_io_deq_ready = _T_766 & _T_580;
  assign Queue_23_clock = clock;
  assign Queue_23_reset = reset;
  assign Queue_23_io_enq_valid = _T_537 & _T_552;
  assign Queue_23_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_23_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_23_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_23_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_23_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_23_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_23_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_23_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_23_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_23_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_23_io_deq_ready = _T_767 & _T_586;
  assign Queue_24_clock = clock;
  assign Queue_24_reset = reset;
  assign Queue_24_io_enq_valid = _T_537 & _T_553;
  assign Queue_24_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_24_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_24_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_24_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_24_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_24_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_24_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_24_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_24_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_24_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_24_io_deq_ready = _T_768 & _T_592;
  assign Queue_25_clock = clock;
  assign Queue_25_reset = reset;
  assign Queue_25_io_enq_valid = _T_537 & _T_554;
  assign Queue_25_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_25_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_25_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_25_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_25_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_25_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_25_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_25_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_25_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_25_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_25_io_deq_ready = _T_769 & _T_598;
  assign Queue_26_clock = clock;
  assign Queue_26_reset = reset;
  assign Queue_26_io_enq_valid = _T_537 & _T_555;
  assign Queue_26_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_26_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_26_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_26_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_26_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_26_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_26_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_26_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_26_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_26_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_26_io_deq_ready = _T_770 & _T_604;
  assign Queue_27_clock = clock;
  assign Queue_27_reset = reset;
  assign Queue_27_io_enq_valid = _T_537 & _T_556;
  assign Queue_27_io_enq_bits_data_id = auto_in_ar_bits_id;
  assign Queue_27_io_enq_bits_data_addr = auto_in_ar_bits_addr;
  assign Queue_27_io_enq_bits_data_len = auto_in_ar_bits_len;
  assign Queue_27_io_enq_bits_data_size = auto_in_ar_bits_size;
  assign Queue_27_io_enq_bits_data_burst = auto_in_ar_bits_burst;
  assign Queue_27_io_enq_bits_data_lock = auto_in_ar_bits_lock;
  assign Queue_27_io_enq_bits_data_cache = auto_in_ar_bits_cache;
  assign Queue_27_io_enq_bits_data_prot = auto_in_ar_bits_prot;
  assign Queue_27_io_enq_bits_data_qos = auto_in_ar_bits_qos;
  assign Queue_27_io_enq_bits_timestamp = _T_541 + _GEN_161;
  assign Queue_27_io_deq_ready = _T_771 & _T_610;
  assign Queue_28_clock = clock;
  assign Queue_28_reset = reset;
  assign Queue_28_io_enq_valid = _T_615 ? _T_728 : _T_793;
  assign Queue_28_io_enq_bits_id = _T_874[59:56];
  assign Queue_28_io_enq_bits_addr = _T_874[55:25];
  assign Queue_28_io_enq_bits_len = _T_874[24:17];
  assign Queue_28_io_enq_bits_size = _T_874[16:14];
  assign Queue_28_io_enq_bits_burst = _T_874[13:12];
  assign Queue_28_io_deq_ready = auto_out_ar_ready;
  assign MaxPeriodFibonacciLFSR_2__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR_2__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR_2__EVAL_9 = 1'h1;
  assign Queue_29_clock = clock;
  assign Queue_29_reset = reset;
  assign Queue_29_io_enq_valid = auto_out_b_valid & _T_954;
  assign Queue_29_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_29_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_29_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_29_io_deq_ready = _T_1169 & _T_973;
  assign Queue_30_clock = clock;
  assign Queue_30_reset = reset;
  assign Queue_30_io_enq_valid = auto_out_b_valid & _T_955;
  assign Queue_30_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_30_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_30_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_30_io_deq_ready = _T_1170 & _T_979;
  assign Queue_31_clock = clock;
  assign Queue_31_reset = reset;
  assign Queue_31_io_enq_valid = auto_out_b_valid & _T_956;
  assign Queue_31_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_31_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_31_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_31_io_deq_ready = _T_1171 & _T_985;
  assign Queue_32_clock = clock;
  assign Queue_32_reset = reset;
  assign Queue_32_io_enq_valid = auto_out_b_valid & _T_957;
  assign Queue_32_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_32_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_32_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_32_io_deq_ready = _T_1172 & _T_991;
  assign Queue_33_clock = clock;
  assign Queue_33_reset = reset;
  assign Queue_33_io_enq_valid = auto_out_b_valid & _T_958;
  assign Queue_33_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_33_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_33_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_33_io_deq_ready = _T_1173 & _T_997;
  assign Queue_34_clock = clock;
  assign Queue_34_reset = reset;
  assign Queue_34_io_enq_valid = auto_out_b_valid & _T_959;
  assign Queue_34_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_34_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_34_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_34_io_deq_ready = _T_1174 & _T_1003;
  assign Queue_35_clock = clock;
  assign Queue_35_reset = reset;
  assign Queue_35_io_enq_valid = auto_out_b_valid & _T_960;
  assign Queue_35_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_35_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_35_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_35_io_deq_ready = _T_1175 & _T_1009;
  assign Queue_36_clock = clock;
  assign Queue_36_reset = reset;
  assign Queue_36_io_enq_valid = auto_out_b_valid & _T_961;
  assign Queue_36_io_enq_bits_data_id = auto_out_b_bits_id;
  assign Queue_36_io_enq_bits_data_resp = auto_out_b_bits_resp;
  assign Queue_36_io_enq_bits_timestamp = _T_946 + _GEN_166;
  assign Queue_36_io_deq_ready = _T_1176 & _T_1015;
  assign Queue_37_clock = clock;
  assign Queue_37_reset = reset;
  assign Queue_37_io_enq_valid = _T_1020 ? _T_1133 : _T_1198;
  assign Queue_37_io_enq_bits_id = _T_1223[5:2];
  assign Queue_37_io_enq_bits_resp = _T_1223[1:0];
  assign Queue_37_io_deq_ready = auto_in_b_ready;
  assign MaxPeriodFibonacciLFSR_3__EVAL_15 = clock;
  assign MaxPeriodFibonacciLFSR_3__EVAL_13 = reset;
  assign MaxPeriodFibonacciLFSR_3__EVAL_9 = 1'h1;
  assign Queue_38_clock = clock;
  assign Queue_38_reset = reset;
  assign Queue_38_io_enq_valid = auto_out_r_valid & _T_1296;
  assign Queue_38_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_38_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_38_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_38_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_38_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_38_io_deq_ready = _T_1511 & _T_1315;
  assign Queue_39_clock = clock;
  assign Queue_39_reset = reset;
  assign Queue_39_io_enq_valid = auto_out_r_valid & _T_1297;
  assign Queue_39_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_39_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_39_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_39_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_39_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_39_io_deq_ready = _T_1512 & _T_1321;
  assign Queue_40_clock = clock;
  assign Queue_40_reset = reset;
  assign Queue_40_io_enq_valid = auto_out_r_valid & _T_1298;
  assign Queue_40_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_40_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_40_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_40_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_40_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_40_io_deq_ready = _T_1513 & _T_1327;
  assign Queue_41_clock = clock;
  assign Queue_41_reset = reset;
  assign Queue_41_io_enq_valid = auto_out_r_valid & _T_1299;
  assign Queue_41_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_41_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_41_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_41_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_41_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_41_io_deq_ready = _T_1514 & _T_1333;
  assign Queue_42_clock = clock;
  assign Queue_42_reset = reset;
  assign Queue_42_io_enq_valid = auto_out_r_valid & _T_1300;
  assign Queue_42_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_42_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_42_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_42_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_42_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_42_io_deq_ready = _T_1515 & _T_1339;
  assign Queue_43_clock = clock;
  assign Queue_43_reset = reset;
  assign Queue_43_io_enq_valid = auto_out_r_valid & _T_1301;
  assign Queue_43_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_43_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_43_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_43_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_43_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_43_io_deq_ready = _T_1516 & _T_1345;
  assign Queue_44_clock = clock;
  assign Queue_44_reset = reset;
  assign Queue_44_io_enq_valid = auto_out_r_valid & _T_1302;
  assign Queue_44_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_44_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_44_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_44_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_44_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_44_io_deq_ready = _T_1517 & _T_1351;
  assign Queue_45_clock = clock;
  assign Queue_45_reset = reset;
  assign Queue_45_io_enq_valid = auto_out_r_valid & _T_1303;
  assign Queue_45_io_enq_bits_data_id = auto_out_r_bits_id;
  assign Queue_45_io_enq_bits_data_data = auto_out_r_bits_data;
  assign Queue_45_io_enq_bits_data_resp = auto_out_r_bits_resp;
  assign Queue_45_io_enq_bits_data_last = auto_out_r_bits_last;
  assign Queue_45_io_enq_bits_timestamp = _T_1288 + _GEN_171;
  assign Queue_45_io_deq_ready = _T_1518 & _T_1357;
  assign Queue_46_clock = clock;
  assign Queue_46_reset = reset;
  assign Queue_46_io_enq_valid = _T_1362 ? _T_1475 : _T_1540;
  assign Queue_46_io_enq_bits_id = _T_1581[38:35];
  assign Queue_46_io_enq_bits_data = _T_1581[34:3];
  assign Queue_46_io_enq_bits_resp = _T_1581[2:1];
  assign Queue_46_io_enq_bits_last = _T_1581[0];
  assign Queue_46_io_deq_ready = auto_in_r_ready;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_140 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_156 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_287_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_287_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_287_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_287_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_287_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_287_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_287_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_287_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_484 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_614 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_630 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_761_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_761_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_761_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_761_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_761_4 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_761_5 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_761_6 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_761_7 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_889 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1019 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1035 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1166_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1166_1 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1166_2 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1166_3 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1166_4 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_1166_5 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_1166_6 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1166_7 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_1231 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_1361 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_1377 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_1508_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_1508_1 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_1508_2 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_1508_3 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1508_4 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_1508_5 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_1508_6 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1508_7 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_10 <= 32'h0;
    end else begin
      _T_10 <= _T_12;
    end
    if (reset) begin
      _T_140 <= 1'h0;
    end else begin
      if (_T_142) begin
        _T_140 <= 1'h0;
      end else begin
        _T_140 <= _T_284;
      end
    end
    if (reset) begin
      _T_156 <= 8'hff;
    end else begin
      if (_T_175) begin
        _T_156 <= _T_185;
      end
    end
    if (reset) begin
      _T_287_0 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_0 <= _T_197;
      end
    end
    if (reset) begin
      _T_287_1 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_1 <= _T_198;
      end
    end
    if (reset) begin
      _T_287_2 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_2 <= _T_199;
      end
    end
    if (reset) begin
      _T_287_3 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_3 <= _T_200;
      end
    end
    if (reset) begin
      _T_287_4 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_4 <= _T_201;
      end
    end
    if (reset) begin
      _T_287_5 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_5 <= _T_202;
      end
    end
    if (reset) begin
      _T_287_6 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_6 <= _T_203;
      end
    end
    if (reset) begin
      _T_287_7 <= 1'h0;
    end else begin
      if (_T_141) begin
        _T_287_7 <= _T_204;
      end
    end
    if (reset) begin
      _T_484 <= 32'h0;
    end else begin
      _T_484 <= _T_486;
    end
    if (reset) begin
      _T_614 <= 1'h0;
    end else begin
      if (_T_616) begin
        _T_614 <= 1'h0;
      end else begin
        _T_614 <= _T_758;
      end
    end
    if (reset) begin
      _T_630 <= 8'hff;
    end else begin
      if (_T_649) begin
        _T_630 <= _T_659;
      end
    end
    if (reset) begin
      _T_761_0 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_0 <= _T_671;
      end
    end
    if (reset) begin
      _T_761_1 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_1 <= _T_672;
      end
    end
    if (reset) begin
      _T_761_2 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_2 <= _T_673;
      end
    end
    if (reset) begin
      _T_761_3 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_3 <= _T_674;
      end
    end
    if (reset) begin
      _T_761_4 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_4 <= _T_675;
      end
    end
    if (reset) begin
      _T_761_5 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_5 <= _T_676;
      end
    end
    if (reset) begin
      _T_761_6 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_6 <= _T_677;
      end
    end
    if (reset) begin
      _T_761_7 <= 1'h0;
    end else begin
      if (_T_615) begin
        _T_761_7 <= _T_678;
      end
    end
    if (reset) begin
      _T_889 <= 32'h0;
    end else begin
      _T_889 <= _T_891;
    end
    if (reset) begin
      _T_1019 <= 1'h0;
    end else begin
      if (_T_1021) begin
        _T_1019 <= 1'h0;
      end else begin
        _T_1019 <= _T_1163;
      end
    end
    if (reset) begin
      _T_1035 <= 8'hff;
    end else begin
      if (_T_1054) begin
        _T_1035 <= _T_1064;
      end
    end
    if (reset) begin
      _T_1166_0 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_0 <= _T_1076;
      end
    end
    if (reset) begin
      _T_1166_1 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_1 <= _T_1077;
      end
    end
    if (reset) begin
      _T_1166_2 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_2 <= _T_1078;
      end
    end
    if (reset) begin
      _T_1166_3 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_3 <= _T_1079;
      end
    end
    if (reset) begin
      _T_1166_4 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_4 <= _T_1080;
      end
    end
    if (reset) begin
      _T_1166_5 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_5 <= _T_1081;
      end
    end
    if (reset) begin
      _T_1166_6 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_6 <= _T_1082;
      end
    end
    if (reset) begin
      _T_1166_7 <= 1'h0;
    end else begin
      if (_T_1020) begin
        _T_1166_7 <= _T_1083;
      end
    end
    if (reset) begin
      _T_1231 <= 32'h0;
    end else begin
      _T_1231 <= _T_1233;
    end
    if (reset) begin
      _T_1361 <= 1'h0;
    end else begin
      if (_T_1363) begin
        _T_1361 <= 1'h0;
      end else begin
        _T_1361 <= _T_1505;
      end
    end
    if (reset) begin
      _T_1377 <= 8'hff;
    end else begin
      if (_T_1396) begin
        _T_1377 <= _T_1406;
      end
    end
    if (reset) begin
      _T_1508_0 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_0 <= _T_1418;
      end
    end
    if (reset) begin
      _T_1508_1 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_1 <= _T_1419;
      end
    end
    if (reset) begin
      _T_1508_2 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_2 <= _T_1420;
      end
    end
    if (reset) begin
      _T_1508_3 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_3 <= _T_1421;
      end
    end
    if (reset) begin
      _T_1508_4 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_4 <= _T_1422;
      end
    end
    if (reset) begin
      _T_1508_5 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_5 <= _T_1423;
      end
    end
    if (reset) begin
      _T_1508_6 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_6 <= _T_1424;
      end
    end
    if (reset) begin
      _T_1508_7 <= 1'h0;
    end else begin
      if (_T_1362) begin
        _T_1508_7 <= _T_1425;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_154) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_247) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_266) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_721) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_721) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_740) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_740) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1033) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1145) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1375) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1375) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1468) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1468) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1487) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
