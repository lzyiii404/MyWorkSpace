//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_162(
  input  [7:0]  _EVAL,
  output [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  output        _EVAL_4,
  input  [29:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  output [2:0]  _EVAL_8,
  output [7:0]  _EVAL_9,
  output        _EVAL_10,
  input  [2:0]  _EVAL_11,
  output [29:0] _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [1:0]  _EVAL_17,
  output [2:0]  _EVAL_18,
  input  [3:0]  _EVAL_19,
  output        _EVAL_20,
  output [1:0]  _EVAL_21,
  input         _EVAL_22
);
  reg  _EVAL_23 [0:1];
  reg [31:0] _RAND_0;
  wire  _EVAL_23__EVAL_24_data;
  wire  _EVAL_23__EVAL_24_addr;
  wire  _EVAL_23__EVAL_25_data;
  wire  _EVAL_23__EVAL_25_addr;
  wire  _EVAL_23__EVAL_25_mask;
  wire  _EVAL_23__EVAL_25_en;
  reg [7:0] _EVAL_31 [0:1];
  reg [31:0] _RAND_1;
  wire [7:0] _EVAL_31__EVAL_32_data;
  wire  _EVAL_31__EVAL_32_addr;
  wire [7:0] _EVAL_31__EVAL_33_data;
  wire  _EVAL_31__EVAL_33_addr;
  wire  _EVAL_31__EVAL_33_mask;
  wire  _EVAL_31__EVAL_33_en;
  reg  _EVAL_34 [0:1];
  reg [31:0] _RAND_2;
  wire  _EVAL_34__EVAL_35_data;
  wire  _EVAL_34__EVAL_35_addr;
  wire  _EVAL_34__EVAL_36_data;
  wire  _EVAL_34__EVAL_36_addr;
  wire  _EVAL_34__EVAL_36_mask;
  wire  _EVAL_34__EVAL_36_en;
  reg [3:0] _EVAL_38 [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] _EVAL_38__EVAL_39_data;
  wire  _EVAL_38__EVAL_39_addr;
  wire [3:0] _EVAL_38__EVAL_40_data;
  wire  _EVAL_38__EVAL_40_addr;
  wire  _EVAL_38__EVAL_40_mask;
  wire  _EVAL_38__EVAL_40_en;
  reg [29:0] _EVAL_42 [0:1];
  reg [31:0] _RAND_4;
  wire [29:0] _EVAL_42__EVAL_43_data;
  wire  _EVAL_42__EVAL_43_addr;
  wire [29:0] _EVAL_42__EVAL_44_data;
  wire  _EVAL_42__EVAL_44_addr;
  wire  _EVAL_42__EVAL_44_mask;
  wire  _EVAL_42__EVAL_44_en;
  reg [3:0] _EVAL_47 [0:1];
  reg [31:0] _RAND_5;
  wire [3:0] _EVAL_47__EVAL_48_data;
  wire  _EVAL_47__EVAL_48_addr;
  wire [3:0] _EVAL_47__EVAL_49_data;
  wire  _EVAL_47__EVAL_49_addr;
  wire  _EVAL_47__EVAL_49_mask;
  wire  _EVAL_47__EVAL_49_en;
  reg [2:0] _EVAL_57 [0:1];
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire [2:0] _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  reg [2:0] _EVAL_61 [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] _EVAL_61__EVAL_62_data;
  wire  _EVAL_61__EVAL_62_addr;
  wire [2:0] _EVAL_61__EVAL_63_data;
  wire  _EVAL_61__EVAL_63_addr;
  wire  _EVAL_61__EVAL_63_mask;
  wire  _EVAL_61__EVAL_63_en;
  reg [1:0] _EVAL_64 [0:1];
  reg [31:0] _RAND_8;
  wire [1:0] _EVAL_64__EVAL_65_data;
  wire  _EVAL_64__EVAL_65_addr;
  wire [1:0] _EVAL_64__EVAL_66_data;
  wire  _EVAL_64__EVAL_66_addr;
  wire  _EVAL_64__EVAL_66_mask;
  wire  _EVAL_64__EVAL_66_en;
  reg  _EVAL_26;
  reg [31:0] _RAND_9;
  reg  _EVAL_52;
  reg [31:0] _RAND_10;
  reg  _EVAL_53;
  reg [31:0] _RAND_11;
  wire  _EVAL_46;
  wire  _EVAL_60;
  wire  _EVAL_54;
  wire  _EVAL_30;
  wire  _EVAL_37;
  wire  _EVAL_51;
  wire  _EVAL_55;
  wire  _EVAL_27;
  wire  _EVAL_50;
  assign _EVAL_23__EVAL_24_addr = _EVAL_52;
  assign _EVAL_23__EVAL_24_data = _EVAL_23[_EVAL_23__EVAL_24_addr];
  assign _EVAL_23__EVAL_25_data = _EVAL_7;
  assign _EVAL_23__EVAL_25_addr = _EVAL_26;
  assign _EVAL_23__EVAL_25_mask = 1'h1;
  assign _EVAL_23__EVAL_25_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_31__EVAL_32_addr = _EVAL_52;
  assign _EVAL_31__EVAL_32_data = _EVAL_31[_EVAL_31__EVAL_32_addr];
  assign _EVAL_31__EVAL_33_data = _EVAL;
  assign _EVAL_31__EVAL_33_addr = _EVAL_26;
  assign _EVAL_31__EVAL_33_mask = 1'h1;
  assign _EVAL_31__EVAL_33_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_34__EVAL_35_addr = _EVAL_52;
  assign _EVAL_34__EVAL_35_data = _EVAL_34[_EVAL_34__EVAL_35_addr];
  assign _EVAL_34__EVAL_36_data = _EVAL_14;
  assign _EVAL_34__EVAL_36_addr = _EVAL_26;
  assign _EVAL_34__EVAL_36_mask = 1'h1;
  assign _EVAL_34__EVAL_36_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_38__EVAL_39_addr = _EVAL_52;
  assign _EVAL_38__EVAL_39_data = _EVAL_38[_EVAL_38__EVAL_39_addr];
  assign _EVAL_38__EVAL_40_data = _EVAL_15;
  assign _EVAL_38__EVAL_40_addr = _EVAL_26;
  assign _EVAL_38__EVAL_40_mask = 1'h1;
  assign _EVAL_38__EVAL_40_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_42__EVAL_43_addr = _EVAL_52;
  assign _EVAL_42__EVAL_43_data = _EVAL_42[_EVAL_42__EVAL_43_addr];
  assign _EVAL_42__EVAL_44_data = _EVAL_5;
  assign _EVAL_42__EVAL_44_addr = _EVAL_26;
  assign _EVAL_42__EVAL_44_mask = 1'h1;
  assign _EVAL_42__EVAL_44_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_47__EVAL_48_addr = _EVAL_52;
  assign _EVAL_47__EVAL_48_data = _EVAL_47[_EVAL_47__EVAL_48_addr];
  assign _EVAL_47__EVAL_49_data = _EVAL_19;
  assign _EVAL_47__EVAL_49_addr = _EVAL_26;
  assign _EVAL_47__EVAL_49_mask = 1'h1;
  assign _EVAL_47__EVAL_49_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_57__EVAL_58_addr = _EVAL_52;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_3;
  assign _EVAL_57__EVAL_59_addr = _EVAL_26;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_61__EVAL_62_addr = _EVAL_52;
  assign _EVAL_61__EVAL_62_data = _EVAL_61[_EVAL_61__EVAL_62_addr];
  assign _EVAL_61__EVAL_63_data = _EVAL_11;
  assign _EVAL_61__EVAL_63_addr = _EVAL_26;
  assign _EVAL_61__EVAL_63_mask = 1'h1;
  assign _EVAL_61__EVAL_63_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_64__EVAL_65_addr = _EVAL_52;
  assign _EVAL_64__EVAL_65_data = _EVAL_64[_EVAL_64__EVAL_65_addr];
  assign _EVAL_64__EVAL_66_data = _EVAL_17;
  assign _EVAL_64__EVAL_66_addr = _EVAL_26;
  assign _EVAL_64__EVAL_66_mask = 1'h1;
  assign _EVAL_64__EVAL_66_en = _EVAL_10 & _EVAL_6;
  assign _EVAL_46 = _EVAL_10 & _EVAL_6;
  assign _EVAL_60 = _EVAL_26 + 1'h1;
  assign _EVAL_54 = _EVAL_1 & _EVAL_20;
  assign _EVAL_30 = _EVAL_52 + 1'h1;
  assign _EVAL_37 = _EVAL_46 != _EVAL_54;
  assign _EVAL_51 = _EVAL_26 == _EVAL_52;
  assign _EVAL_55 = _EVAL_53 == 1'h0;
  assign _EVAL_27 = _EVAL_51 & _EVAL_55;
  assign _EVAL_50 = _EVAL_51 & _EVAL_53;
  assign _EVAL_21 = _EVAL_64__EVAL_65_data;
  assign _EVAL_12 = _EVAL_42__EVAL_43_data;
  assign _EVAL_8 = _EVAL_57__EVAL_58_data;
  assign _EVAL_4 = _EVAL_23__EVAL_24_data;
  assign _EVAL_0 = _EVAL_38__EVAL_39_data;
  assign _EVAL_13 = _EVAL_34__EVAL_35_data;
  assign _EVAL_10 = _EVAL_50 == 1'h0;
  assign _EVAL_20 = _EVAL_27 == 1'h0;
  assign _EVAL_18 = _EVAL_61__EVAL_62_data;
  assign _EVAL_16 = _EVAL_47__EVAL_48_data;
  assign _EVAL_9 = _EVAL_31__EVAL_32_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_23[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_31[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_34[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_38[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_42[initvar] = _RAND_4[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_47[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_6[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_61[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_64[initvar] = _RAND_8[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_26 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_52 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_53 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if(_EVAL_23__EVAL_25_en & _EVAL_23__EVAL_25_mask) begin
      _EVAL_23[_EVAL_23__EVAL_25_addr] <= _EVAL_23__EVAL_25_data;
    end
    if(_EVAL_31__EVAL_33_en & _EVAL_31__EVAL_33_mask) begin
      _EVAL_31[_EVAL_31__EVAL_33_addr] <= _EVAL_31__EVAL_33_data;
    end
    if(_EVAL_34__EVAL_36_en & _EVAL_34__EVAL_36_mask) begin
      _EVAL_34[_EVAL_34__EVAL_36_addr] <= _EVAL_34__EVAL_36_data;
    end
    if(_EVAL_38__EVAL_40_en & _EVAL_38__EVAL_40_mask) begin
      _EVAL_38[_EVAL_38__EVAL_40_addr] <= _EVAL_38__EVAL_40_data;
    end
    if(_EVAL_42__EVAL_44_en & _EVAL_42__EVAL_44_mask) begin
      _EVAL_42[_EVAL_42__EVAL_44_addr] <= _EVAL_42__EVAL_44_data;
    end
    if(_EVAL_47__EVAL_49_en & _EVAL_47__EVAL_49_mask) begin
      _EVAL_47[_EVAL_47__EVAL_49_addr] <= _EVAL_47__EVAL_49_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if(_EVAL_61__EVAL_63_en & _EVAL_61__EVAL_63_mask) begin
      _EVAL_61[_EVAL_61__EVAL_63_addr] <= _EVAL_61__EVAL_63_data;
    end
    if(_EVAL_64__EVAL_66_en & _EVAL_64__EVAL_66_mask) begin
      _EVAL_64[_EVAL_64__EVAL_66_addr] <= _EVAL_64__EVAL_66_data;
    end
    if (_EVAL_22) begin
      _EVAL_26 <= 1'h0;
    end else begin
      if (_EVAL_46) begin
        _EVAL_26 <= _EVAL_60;
      end
    end
    if (_EVAL_22) begin
      _EVAL_52 <= 1'h0;
    end else begin
      if (_EVAL_54) begin
        _EVAL_52 <= _EVAL_30;
      end
    end
    if (_EVAL_22) begin
      _EVAL_53 <= 1'h0;
    end else begin
      if (_EVAL_37) begin
        _EVAL_53 <= _EVAL_46;
      end
    end
  end
endmodule
