//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_178_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [29:0] _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [6:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [6:0]  _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [1:0] _EVAL_50;
  reg [31:0] _RAND_0;
  reg [5:0] _EVAL_55;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_60;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_72;
  reg [31:0] _RAND_3;
  reg [5:0] _EVAL_94;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_110;
  reg [31:0] _RAND_5;
  reg [3:0] _EVAL_121;
  reg [31:0] _RAND_6;
  reg  _EVAL_127;
  reg [31:0] _RAND_7;
  reg [5:0] _EVAL_131;
  reg [31:0] _RAND_8;
  reg  _EVAL_188;
  reg [31:0] _RAND_9;
  reg [29:0] _EVAL_214;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_250;
  reg [31:0] _RAND_11;
  reg [6:0] _EVAL_286;
  reg [31:0] _RAND_12;
  reg [72:0] _EVAL_308;
  reg [95:0] _RAND_13;
  reg [5:0] _EVAL_329;
  reg [31:0] _RAND_14;
  reg [6:0] _EVAL_344;
  reg [31:0] _RAND_15;
  reg [31:0] _EVAL_369;
  reg [31:0] _RAND_16;
  wire  _EVAL_227;
  wire  _EVAL_235;
  wire  _EVAL_260;
  wire [1:0] _EVAL_204;
  wire [1:0] _EVAL_350;
  wire  _EVAL_201;
  wire  _EVAL_33;
  wire  _EVAL_141;
  wire  _EVAL_347;
  wire  _EVAL_62;
  wire  _EVAL_129;
  wire  _EVAL_160;
  wire  _EVAL_186;
  wire  _EVAL_300;
  wire [30:0] _EVAL_42;
  wire [30:0] _EVAL_314;
  wire [30:0] _EVAL_198;
  wire [72:0] _EVAL_156;
  wire  _EVAL_179;
  wire [29:0] _EVAL_137;
  wire [30:0] _EVAL_164;
  wire [30:0] _EVAL_138;
  wire [30:0] _EVAL_229;
  wire  _EVAL_120;
  wire [29:0] _EVAL_338;
  wire [30:0] _EVAL_193;
  wire [30:0] _EVAL_54;
  wire [30:0] _EVAL_46;
  wire  _EVAL_133;
  wire  _EVAL_84;
  wire [29:0] _EVAL_199;
  wire [30:0] _EVAL_118;
  wire [30:0] _EVAL_108;
  wire [30:0] _EVAL_64;
  wire  _EVAL_358;
  wire  _EVAL_35;
  wire  _EVAL_68;
  wire  _EVAL_48;
  wire [29:0] _EVAL_298;
  wire [30:0] _EVAL_21;
  wire [30:0] _EVAL_348;
  wire [30:0] _EVAL_371;
  wire  _EVAL_187;
  wire  _EVAL_213;
  wire [22:0] _EVAL_145;
  wire [7:0] _EVAL_124;
  wire [7:0] _EVAL_155;
  wire [29:0] _EVAL_75;
  wire [29:0] _EVAL_109;
  wire  _EVAL_244;
  wire  _EVAL_232;
  wire  _EVAL_243;
  wire  _EVAL_172;
  wire  _EVAL_40;
  wire  _EVAL_26;
  wire  _EVAL_271;
  wire  _EVAL_102;
  wire  _EVAL_328;
  wire  _EVAL_276;
  wire  _EVAL_125;
  wire  _EVAL_246;
  wire  _EVAL_242;
  wire  _EVAL_299;
  wire  _EVAL_159;
  wire  _EVAL_364;
  wire  _EVAL_116;
  wire  _EVAL_85;
  wire  _EVAL_65;
  wire  _EVAL_67;
  wire  _EVAL_281;
  wire  _EVAL_146;
  wire  _EVAL_210;
  wire  _EVAL_253;
  wire  _EVAL_177;
  wire  _EVAL_190;
  wire  _EVAL_66;
  wire  _EVAL_20;
  wire  _EVAL_161;
  wire  _EVAL_206;
  wire  _EVAL_189;
  wire  _EVAL_366;
  wire  _EVAL_273;
  wire  _EVAL_95;
  wire [3:0] _EVAL_104;
  wire  _EVAL_359;
  wire  _EVAL_325;
  wire  _EVAL_140;
  wire  _EVAL_221;
  wire  _EVAL_88;
  wire [29:0] _EVAL_368;
  wire [30:0] _EVAL_165;
  wire [30:0] _EVAL_277;
  wire [30:0] _EVAL_290;
  wire  _EVAL_24;
  wire  _EVAL_245;
  wire  _EVAL_256;
  wire  _EVAL_289;
  wire [127:0] _EVAL_167;
  wire [127:0] _EVAL_360;
  wire  _EVAL_291;
  wire  _EVAL_261;
  wire  _EVAL_153;
  wire  _EVAL_247;
  wire  _EVAL_27;
  wire  _EVAL_123;
  wire  _EVAL_119;
  wire  _EVAL_252;
  wire  _EVAL_296;
  wire  _EVAL_309;
  wire  _EVAL_112;
  wire  _EVAL_239;
  wire [29:0] _EVAL_173;
  wire [30:0] _EVAL_219;
  wire [30:0] _EVAL_354;
  wire [30:0] _EVAL_211;
  wire  _EVAL_351;
  wire  _EVAL_362;
  wire  _EVAL_316;
  wire  _EVAL_320;
  wire [72:0] _EVAL_195;
  wire [72:0] _EVAL_32;
  wire [72:0] _EVAL_113;
  wire  _EVAL_324;
  wire [3:0] _EVAL_321;
  wire  _EVAL_236;
  wire  _EVAL_43;
  wire  _EVAL_134;
  wire  _EVAL_80;
  wire [22:0] _EVAL_30;
  wire  _EVAL_275;
  wire  _EVAL_220;
  wire  _EVAL_310;
  wire  _EVAL_332;
  wire [3:0] _EVAL_31;
  wire  _EVAL_349;
  wire [2:0] _EVAL_53;
  wire  _EVAL_56;
  wire  _EVAL_79;
  wire  _EVAL_36;
  wire  _EVAL_343;
  wire  _EVAL_86;
  wire  _EVAL_122;
  wire  _EVAL_197;
  wire  _EVAL_228;
  wire  _EVAL_258;
  wire  _EVAL_264;
  wire  _EVAL_287;
  wire  _EVAL_139;
  wire  _EVAL_106;
  wire  _EVAL_342;
  wire  _EVAL_370;
  wire  _EVAL_234;
  wire  _EVAL_337;
  wire  _EVAL_183;
  wire  _EVAL_185;
  wire  _EVAL_158;
  wire  _EVAL_238;
  wire [3:0] _EVAL_44;
  wire  _EVAL_175;
  wire [2:0] _EVAL_295;
  wire  _EVAL_69;
  wire  _EVAL_365;
  wire  _EVAL_361;
  wire  _EVAL_203;
  wire  _EVAL_22;
  wire  _EVAL_38;
  wire  _EVAL_307;
  wire  _EVAL_111;
  wire  _EVAL_315;
  wire  _EVAL_126;
  wire [3:0] _EVAL_345;
  wire [5:0] _EVAL_168;
  wire  _EVAL_249;
  wire  _EVAL_34;
  wire  _EVAL_319;
  wire  _EVAL_92;
  wire  _EVAL_143;
  wire  _EVAL_226;
  wire  _EVAL_100;
  wire [127:0] _EVAL_170;
  wire [127:0] _EVAL_341;
  wire [72:0] _EVAL_99;
  wire  _EVAL_233;
  wire  _EVAL_41;
  wire  _EVAL_294;
  wire  _EVAL_334;
  wire  _EVAL_200;
  wire  _EVAL_115;
  wire  _EVAL_335;
  wire  _EVAL_28;
  wire  _EVAL_231;
  wire  _EVAL_194;
  wire [7:0] _EVAL_81;
  wire [7:0] _EVAL_346;
  wire [5:0] _EVAL_171;
  wire [5:0] _EVAL_78;
  wire  _EVAL_262;
  wire  _EVAL_71;
  wire  _EVAL_23;
  wire  _EVAL_87;
  wire  _EVAL_230;
  wire  _EVAL_279;
  wire  _EVAL_304;
  wire  _EVAL_306;
  wire  _EVAL_322;
  wire  _EVAL_148;
  wire  _EVAL_292;
  wire  _EVAL_254;
  wire  _EVAL_58;
  wire  _EVAL_103;
  wire  _EVAL_278;
  wire  _EVAL_19;
  wire  _EVAL_248;
  wire  _EVAL_301;
  wire  _EVAL_136;
  wire  _EVAL_149;
  wire  _EVAL_333;
  wire  _EVAL_89;
  wire [3:0] _EVAL_303;
  wire  _EVAL_178;
  wire  _EVAL_152;
  wire  _EVAL_51;
  wire  _EVAL_218;
  wire  _EVAL_96;
  wire  _EVAL_326;
  wire  _EVAL_293;
  wire  _EVAL_207;
  wire  _EVAL_356;
  wire  _EVAL_147;
  wire  _EVAL_285;
  wire  _EVAL_205;
  wire  _EVAL_169;
  wire [5:0] _EVAL_70;
  wire  _EVAL_61;
  wire [72:0] _EVAL_59;
  wire  _EVAL_265;
  wire  _EVAL_114;
  wire  _EVAL_162;
  wire  _EVAL_202;
  wire  _EVAL_107;
  wire  _EVAL_284;
  wire  _EVAL_340;
  wire  _EVAL_318;
  wire  _EVAL_154;
  wire  _EVAL_355;
  wire  _EVAL_45;
  wire  _EVAL_176;
  wire  _EVAL_331;
  wire  _EVAL_151;
  wire  _EVAL_317;
  wire [5:0] _EVAL_191;
  wire  _EVAL_29;
  wire  _EVAL_93;
  wire  _EVAL_257;
  wire  _EVAL_174;
  wire  _EVAL_47;
  wire  _EVAL_327;
  wire  _EVAL_222;
  wire  _EVAL_77;
  wire  _EVAL_181;
  wire  _EVAL_101;
  wire  _EVAL_269;
  wire  _EVAL_150;
  wire  _EVAL_357;
  wire  _EVAL_237;
  wire  _EVAL_132;
  wire  _EVAL_240;
  wire  _EVAL_268;
  wire  _EVAL_263;
  wire  _EVAL_25;
  wire  _EVAL_223;
  wire  _EVAL_330;
  wire  _EVAL_217;
  wire  _EVAL_182;
  wire  _EVAL_272;
  wire  _EVAL_255;
  wire [72:0] _EVAL_117;
  wire  _EVAL_288;
  wire  _EVAL_130;
  wire  _EVAL_363;
  wire  _EVAL_212;
  wire  _EVAL_336;
  wire  _EVAL_76;
  wire  _EVAL_37;
  wire  _EVAL_39;
  wire  _EVAL_311;
  wire  _EVAL_266;
  wire  _EVAL_57;
  wire  _EVAL_73;
  wire  _EVAL_302;
  wire  _EVAL_208;
  wire  _EVAL_352;
  wire  _EVAL_209;
  wire  _EVAL_142;
  wire [5:0] _EVAL_180;
  wire  _EVAL_323;
  wire  _EVAL_282;
  wire  _EVAL_241;
  wire  _EVAL_283;
  wire  _EVAL_251;
  wire  _EVAL_82;
  wire [72:0] _EVAL_305;
  wire  _EVAL_192;
  wire  _EVAL_297;
  wire  _EVAL_128;
  wire  _EVAL_353;
  wire  _EVAL_367;
  wire  _EVAL_98;
  wire  _EVAL_215;
  wire [31:0] _EVAL_224;
  wire  _EVAL_91;
  wire  _EVAL_280;
  wire  _EVAL_196;
  wire  _EVAL_52;
  wire  _EVAL_157;
  wire  _EVAL_166;
  wire  _EVAL_259;
  wire  _EVAL_312;
  wire  _EVAL_63;
  wire  _EVAL_83;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_227 = _EVAL_329 == 6'h0;
  assign _EVAL_235 = _EVAL_16 >= 4'h2;
  assign _EVAL_260 = _EVAL_16[0];
  assign _EVAL_204 = 2'h1 << _EVAL_260;
  assign _EVAL_350 = _EVAL_204 | 2'h1;
  assign _EVAL_201 = _EVAL_350[1];
  assign _EVAL_33 = _EVAL_9[1];
  assign _EVAL_141 = _EVAL_201 & _EVAL_33;
  assign _EVAL_347 = _EVAL_235 | _EVAL_141;
  assign _EVAL_62 = _EVAL_1 == _EVAL_127;
  assign _EVAL_129 = _EVAL_1 == 1'h0;
  assign _EVAL_160 = _EVAL_129 | _EVAL_10;
  assign _EVAL_186 = _EVAL_6 <= 3'h6;
  assign _EVAL_300 = _EVAL_186 | _EVAL_10;
  assign _EVAL_42 = {1'b0,$signed(_EVAL_9)};
  assign _EVAL_314 = $signed(_EVAL_42) & $signed(-31'sh5000);
  assign _EVAL_198 = $signed(_EVAL_314);
  assign _EVAL_156 = _EVAL_308 >> _EVAL_13;
  assign _EVAL_179 = _EVAL_3 == 3'h0;
  assign _EVAL_137 = _EVAL_9 ^ 30'h3000;
  assign _EVAL_164 = {1'b0,$signed(_EVAL_137)};
  assign _EVAL_138 = $signed(_EVAL_164) & $signed(-31'sh1000);
  assign _EVAL_229 = $signed(_EVAL_138);
  assign _EVAL_120 = $signed(_EVAL_229) == $signed(31'sh0);
  assign _EVAL_338 = _EVAL_9 ^ 30'hc000000;
  assign _EVAL_193 = {1'b0,$signed(_EVAL_338)};
  assign _EVAL_54 = $signed(_EVAL_193) & $signed(-31'sh4000000);
  assign _EVAL_46 = $signed(_EVAL_54);
  assign _EVAL_133 = $signed(_EVAL_46) == $signed(31'sh0);
  assign _EVAL_84 = _EVAL_120 | _EVAL_133;
  assign _EVAL_199 = _EVAL_9 ^ 30'h2000000;
  assign _EVAL_118 = {1'b0,$signed(_EVAL_199)};
  assign _EVAL_108 = $signed(_EVAL_118) & $signed(-31'sh10000);
  assign _EVAL_64 = $signed(_EVAL_108);
  assign _EVAL_358 = $signed(_EVAL_64) == $signed(31'sh0);
  assign _EVAL_35 = _EVAL_84 | _EVAL_358;
  assign _EVAL_68 = $signed(_EVAL_198) == $signed(31'sh0);
  assign _EVAL_48 = _EVAL_35 | _EVAL_68;
  assign _EVAL_298 = _EVAL_9 ^ 30'h1800000;
  assign _EVAL_21 = {1'b0,$signed(_EVAL_298)};
  assign _EVAL_348 = $signed(_EVAL_21) & $signed(-31'sh8000);
  assign _EVAL_371 = $signed(_EVAL_348);
  assign _EVAL_187 = $signed(_EVAL_371) == $signed(31'sh0);
  assign _EVAL_213 = _EVAL_48 | _EVAL_187;
  assign _EVAL_145 = 23'hff << _EVAL_16;
  assign _EVAL_124 = _EVAL_145[7:0];
  assign _EVAL_155 = ~ _EVAL_124;
  assign _EVAL_75 = {{22'd0}, _EVAL_155};
  assign _EVAL_109 = _EVAL_9 & _EVAL_75;
  assign _EVAL_244 = _EVAL_6 == 3'h5;
  assign _EVAL_232 = _EVAL_7 & _EVAL_244;
  assign _EVAL_243 = _EVAL_0 == _EVAL_50;
  assign _EVAL_172 = _EVAL_308 != 73'h0;
  assign _EVAL_40 = _EVAL_172 == 1'h0;
  assign _EVAL_26 = plusarg_reader_out == 32'h0;
  assign _EVAL_271 = _EVAL_40 | _EVAL_26;
  assign _EVAL_102 = _EVAL_369 < plusarg_reader_out;
  assign _EVAL_328 = _EVAL_271 | _EVAL_102;
  assign _EVAL_276 = _EVAL_328 | _EVAL_10;
  assign _EVAL_125 = _EVAL_62 | _EVAL_10;
  assign _EVAL_246 = _EVAL_13 == 7'h40;
  assign _EVAL_242 = 4'h6 == _EVAL_16;
  assign _EVAL_299 = _EVAL_246 ? _EVAL_242 : 1'h0;
  assign _EVAL_159 = _EVAL_299 | _EVAL_10;
  assign _EVAL_364 = _EVAL_159 == 1'h0;
  assign _EVAL_116 = _EVAL_350[0];
  assign _EVAL_85 = _EVAL_9[0];
  assign _EVAL_65 = _EVAL_33 & _EVAL_85;
  assign _EVAL_67 = _EVAL_116 & _EVAL_65;
  assign _EVAL_281 = _EVAL_347 | _EVAL_67;
  assign _EVAL_146 = _EVAL_85 == 1'h0;
  assign _EVAL_210 = _EVAL_33 & _EVAL_146;
  assign _EVAL_253 = _EVAL_116 & _EVAL_210;
  assign _EVAL_177 = _EVAL_347 | _EVAL_253;
  assign _EVAL_190 = _EVAL_33 == 1'h0;
  assign _EVAL_66 = _EVAL_201 & _EVAL_190;
  assign _EVAL_20 = _EVAL_235 | _EVAL_66;
  assign _EVAL_161 = _EVAL_190 & _EVAL_85;
  assign _EVAL_206 = _EVAL_116 & _EVAL_161;
  assign _EVAL_189 = _EVAL_20 | _EVAL_206;
  assign _EVAL_366 = _EVAL_190 & _EVAL_146;
  assign _EVAL_273 = _EVAL_116 & _EVAL_366;
  assign _EVAL_95 = _EVAL_20 | _EVAL_273;
  assign _EVAL_104 = {_EVAL_281,_EVAL_177,_EVAL_189,_EVAL_95};
  assign _EVAL_359 = _EVAL_3 == _EVAL_60;
  assign _EVAL_325 = _EVAL_0 != 2'h2;
  assign _EVAL_140 = _EVAL_325 | _EVAL_10;
  assign _EVAL_221 = _EVAL_140 == 1'h0;
  assign _EVAL_88 = _EVAL_3 <= 3'h2;
  assign _EVAL_368 = _EVAL_9 ^ 30'h20000000;
  assign _EVAL_165 = {1'b0,$signed(_EVAL_368)};
  assign _EVAL_277 = $signed(_EVAL_165) & $signed(-31'sh2000);
  assign _EVAL_290 = $signed(_EVAL_277);
  assign _EVAL_24 = $signed(_EVAL_290) == $signed(31'sh0);
  assign _EVAL_245 = _EVAL & _EVAL_15;
  assign _EVAL_256 = _EVAL_55 == 6'h0;
  assign _EVAL_289 = _EVAL_245 & _EVAL_256;
  assign _EVAL_167 = 128'h1 << _EVAL_13;
  assign _EVAL_360 = _EVAL_289 ? _EVAL_167 : 128'h0;
  assign _EVAL_291 = _EVAL_5[2];
  assign _EVAL_261 = _EVAL_291 == 1'h0;
  assign _EVAL_153 = _EVAL_156[0];
  assign _EVAL_247 = _EVAL_153 == 1'h0;
  assign _EVAL_27 = _EVAL_247 | _EVAL_10;
  assign _EVAL_123 = _EVAL_27 == 1'h0;
  assign _EVAL_119 = _EVAL_8 == _EVAL_104;
  assign _EVAL_252 = _EVAL_119 | _EVAL_10;
  assign _EVAL_296 = _EVAL_252 == 1'h0;
  assign _EVAL_309 = _EVAL_133 | _EVAL_358;
  assign _EVAL_112 = _EVAL_309 | _EVAL_68;
  assign _EVAL_239 = _EVAL_112 | _EVAL_187;
  assign _EVAL_173 = _EVAL_9 ^ 30'h1900000;
  assign _EVAL_219 = {1'b0,$signed(_EVAL_173)};
  assign _EVAL_354 = $signed(_EVAL_219) & $signed(-31'sh2000);
  assign _EVAL_211 = $signed(_EVAL_354);
  assign _EVAL_351 = $signed(_EVAL_211) == $signed(31'sh0);
  assign _EVAL_362 = _EVAL_239 | _EVAL_351;
  assign _EVAL_316 = _EVAL_13 == _EVAL_286;
  assign _EVAL_320 = _EVAL_316 | _EVAL_10;
  assign _EVAL_195 = _EVAL_360[72:0];
  assign _EVAL_32 = _EVAL_195 | _EVAL_308;
  assign _EVAL_113 = _EVAL_32 >> _EVAL_17;
  assign _EVAL_324 = _EVAL_113[0];
  assign _EVAL_321 = ~ _EVAL_8;
  assign _EVAL_236 = _EVAL_321 == 4'h0;
  assign _EVAL_43 = _EVAL_236 | _EVAL_10;
  assign _EVAL_134 = _EVAL_3 <= 3'h4;
  assign _EVAL_80 = _EVAL_134 | _EVAL_10;
  assign _EVAL_30 = 23'hff << _EVAL_14;
  assign _EVAL_275 = _EVAL_5 == 3'h4;
  assign _EVAL_220 = _EVAL_17 == 7'h48;
  assign _EVAL_310 = _EVAL_17 == 7'h40;
  assign _EVAL_332 = _EVAL_220 | _EVAL_310;
  assign _EVAL_31 = _EVAL_17[6:3];
  assign _EVAL_349 = _EVAL_31 == 4'h8;
  assign _EVAL_53 = _EVAL_17[2:0];
  assign _EVAL_56 = 3'h1 <= _EVAL_53;
  assign _EVAL_79 = _EVAL_349 & _EVAL_56;
  assign _EVAL_36 = _EVAL_332 | _EVAL_79;
  assign _EVAL_343 = _EVAL_17 == 7'h20;
  assign _EVAL_86 = _EVAL_36 | _EVAL_343;
  assign _EVAL_122 = _EVAL_31 == 4'h0;
  assign _EVAL_197 = _EVAL_86 | _EVAL_122;
  assign _EVAL_228 = _EVAL_31 == 4'h1;
  assign _EVAL_258 = _EVAL_197 | _EVAL_228;
  assign _EVAL_264 = _EVAL_31 == 4'h2;
  assign _EVAL_287 = _EVAL_258 | _EVAL_264;
  assign _EVAL_139 = _EVAL_31 == 4'h3;
  assign _EVAL_106 = _EVAL_287 | _EVAL_139;
  assign _EVAL_342 = _EVAL_43 == 1'h0;
  assign _EVAL_370 = _EVAL_213 | _EVAL_351;
  assign _EVAL_234 = _EVAL_16 == _EVAL_72;
  assign _EVAL_337 = _EVAL_109 == 30'h0;
  assign _EVAL_183 = _EVAL_16 <= 4'h8;
  assign _EVAL_185 = _EVAL_183 & _EVAL_120;
  assign _EVAL_158 = _EVAL_13 == 7'h48;
  assign _EVAL_238 = _EVAL_158 | _EVAL_246;
  assign _EVAL_44 = _EVAL_13[6:3];
  assign _EVAL_175 = _EVAL_44 == 4'h8;
  assign _EVAL_295 = _EVAL_13[2:0];
  assign _EVAL_69 = 3'h1 <= _EVAL_295;
  assign _EVAL_365 = _EVAL_175 & _EVAL_69;
  assign _EVAL_361 = _EVAL_238 | _EVAL_365;
  assign _EVAL_203 = _EVAL_13 == 7'h20;
  assign _EVAL_22 = _EVAL_361 | _EVAL_203;
  assign _EVAL_38 = _EVAL_44 == 4'h0;
  assign _EVAL_307 = _EVAL_22 | _EVAL_38;
  assign _EVAL_111 = _EVAL_44 == 4'h1;
  assign _EVAL_315 = _EVAL_307 | _EVAL_111;
  assign _EVAL_126 = _EVAL_10 == 1'h0;
  assign _EVAL_345 = ~ _EVAL_104;
  assign _EVAL_168 = _EVAL_329 - 6'h1;
  assign _EVAL_249 = _EVAL_9 == _EVAL_214;
  assign _EVAL_34 = _EVAL_12 & _EVAL_7;
  assign _EVAL_319 = _EVAL_131 == 6'h0;
  assign _EVAL_92 = _EVAL_34 & _EVAL_319;
  assign _EVAL_143 = _EVAL_6 == 3'h6;
  assign _EVAL_226 = _EVAL_143 == 1'h0;
  assign _EVAL_100 = _EVAL_92 & _EVAL_226;
  assign _EVAL_170 = 128'h1 << _EVAL_17;
  assign _EVAL_341 = _EVAL_100 ? _EVAL_170 : 128'h0;
  assign _EVAL_99 = _EVAL_341[72:0];
  assign _EVAL_233 = _EVAL_195 != _EVAL_99;
  assign _EVAL_41 = _EVAL_195 != 73'h0;
  assign _EVAL_294 = _EVAL_41 == 1'h0;
  assign _EVAL_334 = _EVAL_233 | _EVAL_294;
  assign _EVAL_200 = _EVAL_334 | _EVAL_10;
  assign _EVAL_115 = _EVAL_200 == 1'h0;
  assign _EVAL_335 = _EVAL_18 == 1'h0;
  assign _EVAL_28 = _EVAL_335 | _EVAL_10;
  assign _EVAL_231 = _EVAL_28 == 1'h0;
  assign _EVAL_194 = _EVAL_6[0];
  assign _EVAL_81 = _EVAL_30[7:0];
  assign _EVAL_346 = ~ _EVAL_81;
  assign _EVAL_171 = _EVAL_346[7:2];
  assign _EVAL_78 = _EVAL_131 - 6'h1;
  assign _EVAL_262 = _EVAL_235 | _EVAL_10;
  assign _EVAL_71 = _EVAL_5 == 3'h5;
  assign _EVAL_23 = _EVAL_14 == _EVAL_121;
  assign _EVAL_87 = _EVAL_5 == 3'h3;
  assign _EVAL_230 = _EVAL_3 != 3'h0;
  assign _EVAL_279 = _EVAL_230 | _EVAL_10;
  assign _EVAL_304 = _EVAL_279 == 1'h0;
  assign _EVAL_306 = _EVAL_6 == _EVAL_110;
  assign _EVAL_322 = _EVAL_306 | _EVAL_10;
  assign _EVAL_148 = _EVAL_129 | _EVAL_4;
  assign _EVAL_292 = _EVAL_14 >= 4'h2;
  assign _EVAL_254 = _EVAL_292 | _EVAL_10;
  assign _EVAL_58 = _EVAL_5 == 3'h6;
  assign _EVAL_103 = _EVAL_243 | _EVAL_10;
  assign _EVAL_278 = _EVAL_5 == 3'h1;
  assign _EVAL_19 = _EVAL_5 == 3'h7;
  assign _EVAL_248 = _EVAL_15 & _EVAL_19;
  assign _EVAL_301 = _EVAL_15 & _EVAL_278;
  assign _EVAL_136 = _EVAL_6 == 3'h1;
  assign _EVAL_149 = _EVAL_80 == 1'h0;
  assign _EVAL_333 = _EVAL_5 == 3'h0;
  assign _EVAL_89 = _EVAL_15 & _EVAL_333;
  assign _EVAL_303 = _EVAL_8 & _EVAL_345;
  assign _EVAL_178 = _EVAL_16 <= 4'h6;
  assign _EVAL_152 = _EVAL_362 | _EVAL_24;
  assign _EVAL_51 = _EVAL_178 & _EVAL_152;
  assign _EVAL_218 = _EVAL_185 | _EVAL_51;
  assign _EVAL_96 = _EVAL_218 | _EVAL_10;
  assign _EVAL_326 = _EVAL_44 == 4'h2;
  assign _EVAL_293 = _EVAL_315 | _EVAL_326;
  assign _EVAL_207 = _EVAL_44 == 4'h3;
  assign _EVAL_356 = _EVAL_293 | _EVAL_207;
  assign _EVAL_147 = _EVAL_356 | _EVAL_10;
  assign _EVAL_285 = _EVAL_245 & _EVAL_227;
  assign _EVAL_205 = _EVAL_94 == 6'h0;
  assign _EVAL_169 = _EVAL_88 | _EVAL_10;
  assign _EVAL_70 = _EVAL_155[7:2];
  assign _EVAL_61 = _EVAL_15 & _EVAL_58;
  assign _EVAL_59 = _EVAL_308 | _EVAL_195;
  assign _EVAL_265 = _EVAL_227 == 1'h0;
  assign _EVAL_114 = _EVAL_262 == 1'h0;
  assign _EVAL_162 = _EVAL_249 | _EVAL_10;
  assign _EVAL_202 = _EVAL_4 == 1'h0;
  assign _EVAL_107 = _EVAL_202 | _EVAL_10;
  assign _EVAL_284 = _EVAL_6 == 3'h4;
  assign _EVAL_340 = _EVAL_7 & _EVAL_284;
  assign _EVAL_318 = _EVAL_6 == 3'h0;
  assign _EVAL_154 = _EVAL_359 | _EVAL_10;
  assign _EVAL_355 = _EVAL_154 == 1'h0;
  assign _EVAL_45 = _EVAL_103 == 1'h0;
  assign _EVAL_176 = _EVAL_234 | _EVAL_10;
  assign _EVAL_331 = _EVAL_205 == 1'h0;
  assign _EVAL_151 = _EVAL_7 & _EVAL_331;
  assign _EVAL_317 = _EVAL_324 | _EVAL_10;
  assign _EVAL_191 = _EVAL_55 - 6'h1;
  assign _EVAL_29 = _EVAL_6 == 3'h2;
  assign _EVAL_93 = _EVAL_125 == 1'h0;
  assign _EVAL_257 = _EVAL_0 == 2'h0;
  assign _EVAL_174 = _EVAL_257 | _EVAL_10;
  assign _EVAL_47 = _EVAL_174 == 1'h0;
  assign _EVAL_327 = _EVAL_322 == 1'h0;
  assign _EVAL_222 = _EVAL_106 | _EVAL_10;
  assign _EVAL_77 = _EVAL_337 | _EVAL_10;
  assign _EVAL_181 = _EVAL_303 == 4'h0;
  assign _EVAL_101 = _EVAL_181 | _EVAL_10;
  assign _EVAL_269 = _EVAL_176 == 1'h0;
  assign _EVAL_150 = _EVAL_169 == 1'h0;
  assign _EVAL_357 = _EVAL_0 <= 2'h2;
  assign _EVAL_237 = _EVAL_357 | _EVAL_10;
  assign _EVAL_132 = _EVAL_5 == _EVAL_250;
  assign _EVAL_240 = _EVAL_132 | _EVAL_10;
  assign _EVAL_268 = _EVAL_317 == 1'h0;
  assign _EVAL_263 = _EVAL_16 <= 4'h2;
  assign _EVAL_25 = _EVAL_370 | _EVAL_24;
  assign _EVAL_223 = _EVAL_263 & _EVAL_25;
  assign _EVAL_330 = _EVAL_223 | _EVAL_10;
  assign _EVAL_217 = _EVAL_17 == _EVAL_344;
  assign _EVAL_182 = _EVAL_217 | _EVAL_10;
  assign _EVAL_272 = _EVAL_182 == 1'h0;
  assign _EVAL_255 = _EVAL_245 | _EVAL_34;
  assign _EVAL_117 = ~ _EVAL_99;
  assign _EVAL_288 = _EVAL_3 <= 3'h3;
  assign _EVAL_130 = _EVAL_288 | _EVAL_10;
  assign _EVAL_363 = _EVAL_130 == 1'h0;
  assign _EVAL_212 = _EVAL_34 & _EVAL_205;
  assign _EVAL_336 = _EVAL_179 | _EVAL_10;
  assign _EVAL_76 = _EVAL_15 & _EVAL_265;
  assign _EVAL_37 = _EVAL_330 == 1'h0;
  assign _EVAL_39 = _EVAL_107 == 1'h0;
  assign _EVAL_311 = _EVAL_23 | _EVAL_10;
  assign _EVAL_266 = _EVAL_311 == 1'h0;
  assign _EVAL_57 = _EVAL_336 == 1'h0;
  assign _EVAL_73 = _EVAL_96 == 1'h0;
  assign _EVAL_302 = _EVAL_254 == 1'h0;
  assign _EVAL_208 = _EVAL_11 == _EVAL_188;
  assign _EVAL_352 = _EVAL_300 == 1'h0;
  assign _EVAL_209 = _EVAL_222 == 1'h0;
  assign _EVAL_142 = _EVAL_240 == 1'h0;
  assign _EVAL_180 = _EVAL_94 - 6'h1;
  assign _EVAL_323 = _EVAL_148 | _EVAL_10;
  assign _EVAL_282 = _EVAL_7 & _EVAL_29;
  assign _EVAL_241 = _EVAL_15 & _EVAL_275;
  assign _EVAL_283 = _EVAL_185 | _EVAL_10;
  assign _EVAL_251 = _EVAL_283 == 1'h0;
  assign _EVAL_82 = _EVAL_7 & _EVAL_143;
  assign _EVAL_305 = _EVAL_59 & _EVAL_117;
  assign _EVAL_192 = _EVAL_237 == 1'h0;
  assign _EVAL_297 = _EVAL_208 | _EVAL_10;
  assign _EVAL_128 = _EVAL_297 == 1'h0;
  assign _EVAL_353 = _EVAL_7 & _EVAL_318;
  assign _EVAL_367 = _EVAL_15 & _EVAL_71;
  assign _EVAL_98 = _EVAL_101 == 1'h0;
  assign _EVAL_215 = _EVAL_320 == 1'h0;
  assign _EVAL_224 = _EVAL_369 + 32'h1;
  assign _EVAL_91 = _EVAL_77 == 1'h0;
  assign _EVAL_280 = _EVAL_162 == 1'h0;
  assign _EVAL_196 = _EVAL_160 == 1'h0;
  assign _EVAL_52 = _EVAL_5 == 3'h2;
  assign _EVAL_157 = _EVAL_15 & _EVAL_52;
  assign _EVAL_166 = _EVAL_7 & _EVAL_136;
  assign _EVAL_259 = _EVAL_15 & _EVAL_87;
  assign _EVAL_312 = _EVAL_276 == 1'h0;
  assign _EVAL_63 = _EVAL_147 == 1'h0;
  assign _EVAL_83 = _EVAL_323 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_50 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_55 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_60 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_72 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_94 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_110 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_121 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_127 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_131 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_188 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_214 = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_250 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_286 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {3{`RANDOM}};
  _EVAL_308 = _RAND_13[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_329 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_344 = _RAND_15[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_369 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_212) begin
      _EVAL_50 <= _EVAL_0;
    end
    if (_EVAL_10) begin
      _EVAL_55 <= 6'h0;
    end else begin
      if (_EVAL_245) begin
        if (_EVAL_256) begin
          if (_EVAL_261) begin
            _EVAL_55 <= _EVAL_70;
          end else begin
            _EVAL_55 <= 6'h0;
          end
        end else begin
          _EVAL_55 <= _EVAL_191;
        end
      end
    end
    if (_EVAL_285) begin
      _EVAL_60 <= _EVAL_3;
    end
    if (_EVAL_285) begin
      _EVAL_72 <= _EVAL_16;
    end
    if (_EVAL_10) begin
      _EVAL_94 <= 6'h0;
    end else begin
      if (_EVAL_34) begin
        if (_EVAL_205) begin
          if (_EVAL_194) begin
            _EVAL_94 <= _EVAL_171;
          end else begin
            _EVAL_94 <= 6'h0;
          end
        end else begin
          _EVAL_94 <= _EVAL_180;
        end
      end
    end
    if (_EVAL_212) begin
      _EVAL_110 <= _EVAL_6;
    end
    if (_EVAL_212) begin
      _EVAL_121 <= _EVAL_14;
    end
    if (_EVAL_212) begin
      _EVAL_127 <= _EVAL_1;
    end
    if (_EVAL_10) begin
      _EVAL_131 <= 6'h0;
    end else begin
      if (_EVAL_34) begin
        if (_EVAL_319) begin
          if (_EVAL_194) begin
            _EVAL_131 <= _EVAL_171;
          end else begin
            _EVAL_131 <= 6'h0;
          end
        end else begin
          _EVAL_131 <= _EVAL_78;
        end
      end
    end
    if (_EVAL_212) begin
      _EVAL_188 <= _EVAL_11;
    end
    if (_EVAL_285) begin
      _EVAL_214 <= _EVAL_9;
    end
    if (_EVAL_285) begin
      _EVAL_250 <= _EVAL_5;
    end
    if (_EVAL_285) begin
      _EVAL_286 <= _EVAL_13;
    end
    if (_EVAL_10) begin
      _EVAL_308 <= 73'h0;
    end else begin
      _EVAL_308 <= _EVAL_305;
    end
    if (_EVAL_10) begin
      _EVAL_329 <= 6'h0;
    end else begin
      if (_EVAL_245) begin
        if (_EVAL_227) begin
          if (_EVAL_261) begin
            _EVAL_329 <= _EVAL_70;
          end else begin
            _EVAL_329 <= 6'h0;
          end
        end else begin
          _EVAL_329 <= _EVAL_168;
        end
      end
    end
    if (_EVAL_212) begin
      _EVAL_344 <= _EVAL_17;
    end
    if (_EVAL_10) begin
      _EVAL_369 <= 32'h0;
    end else begin
      if (_EVAL_255) begin
        _EVAL_369 <= 32'h0;
      end else begin
        _EVAL_369 <= _EVAL_224;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4645064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e64c3d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34d41986)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c61394d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ba81fa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b5c8fe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7caac78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3b92f33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2058f3bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a132dd3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(592353b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ca0a2ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92f95045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6047a1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10c9bd8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(671c84e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8718fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d9f5fcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0b8ae53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c4263e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c6c13f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab7f8219)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e339569f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce453341)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f52f086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4caa620)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82949b3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5eba59f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1971885e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b76c8f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0bd2fa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2892e64c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ca59507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e73a0a7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59823d0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b92eaa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81a1e1dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e786411)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4062e79d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c11e18d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d46fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21354a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10f02908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ed50d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61f93f48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(647a3394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(855f92df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e0a8b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53b01d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a3608a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(987d8041)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23fe0f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d203979e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb67f91c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c39e3c5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cf478f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e4a163e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f2f2c05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4e16682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0bb5159)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(416d051f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf9649d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1f35aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5df7a53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a57df908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8492c9fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df842e5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33de6758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a673afc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(794f9eb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6078bcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5941f18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3896140e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fd92a9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b10a1ff8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f7d807)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fd496a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b042ba99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf28b11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40e19c23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2eb9a0a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c17a3ff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd942d88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecaf81c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8df262eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc5ddf3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f13b1e9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5819069f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a215ca0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba11ab2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
