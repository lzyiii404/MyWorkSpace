//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_185(
  output [11:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [11:0] _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [2:0]  _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input  [27:0] _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  output [1:0]  _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_68,
  input  [3:0]  _EVAL_69,
  input         _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  input         _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  input         _EVAL_77,
  input         _EVAL_78,
  input  [1:0]  _EVAL_79,
  input         _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input  [31:0] _EVAL_84,
  input         _EVAL_85,
  input  [2:0]  _EVAL_86,
  input         _EVAL_87,
  input         _EVAL_88,
  input         _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_92,
  input         _EVAL_93,
  input         _EVAL_94,
  input         _EVAL_95,
  input         _EVAL_96,
  input         _EVAL_97,
  input         _EVAL_98,
  input         _EVAL_99,
  input         _EVAL_100,
  input         _EVAL_101,
  input         _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  input         _EVAL_108,
  input         _EVAL_109,
  input         _EVAL_110,
  input         _EVAL_111,
  input         _EVAL_112,
  input         _EVAL_113,
  input         _EVAL_114,
  input         _EVAL_115,
  input         _EVAL_116,
  input         _EVAL_117,
  input         _EVAL_118,
  input         _EVAL_119,
  input         _EVAL_120,
  input         _EVAL_121,
  input         _EVAL_122,
  input         _EVAL_123,
  input         _EVAL_124,
  input         _EVAL_125,
  input         _EVAL_126,
  input         _EVAL_127,
  input         _EVAL_128,
  input         _EVAL_129,
  output [31:0] _EVAL_130,
  input         _EVAL_131,
  input         _EVAL_132,
  input         _EVAL_133,
  input         _EVAL_134,
  input         _EVAL_135,
  input         _EVAL_136,
  input         _EVAL_137,
  output        _EVAL_138,
  input         _EVAL_139,
  input         _EVAL_140,
  input         _EVAL_141,
  input         _EVAL_142,
  input  [2:0]  _EVAL_143,
  input         _EVAL_144
);
  wire  LevelGateway_54__EVAL;
  wire  LevelGateway_54__EVAL_0;
  wire  LevelGateway_54__EVAL_1;
  wire  LevelGateway_54__EVAL_2;
  wire  LevelGateway_54__EVAL_3;
  wire  LevelGateway_54__EVAL_4;
  wire  LevelGateway_65__EVAL;
  wire  LevelGateway_65__EVAL_0;
  wire  LevelGateway_65__EVAL_1;
  wire  LevelGateway_65__EVAL_2;
  wire  LevelGateway_65__EVAL_3;
  wire  LevelGateway_65__EVAL_4;
  wire  LevelGateway__EVAL;
  wire  LevelGateway__EVAL_0;
  wire  LevelGateway__EVAL_1;
  wire  LevelGateway__EVAL_2;
  wire  LevelGateway__EVAL_3;
  wire  LevelGateway__EVAL_4;
  wire  LevelGateway_16__EVAL;
  wire  LevelGateway_16__EVAL_0;
  wire  LevelGateway_16__EVAL_1;
  wire  LevelGateway_16__EVAL_2;
  wire  LevelGateway_16__EVAL_3;
  wire  LevelGateway_16__EVAL_4;
  wire  LevelGateway_34__EVAL;
  wire  LevelGateway_34__EVAL_0;
  wire  LevelGateway_34__EVAL_1;
  wire  LevelGateway_34__EVAL_2;
  wire  LevelGateway_34__EVAL_3;
  wire  LevelGateway_34__EVAL_4;
  wire  LevelGateway_92__EVAL;
  wire  LevelGateway_92__EVAL_0;
  wire  LevelGateway_92__EVAL_1;
  wire  LevelGateway_92__EVAL_2;
  wire  LevelGateway_92__EVAL_3;
  wire  LevelGateway_92__EVAL_4;
  wire  LevelGateway_39__EVAL;
  wire  LevelGateway_39__EVAL_0;
  wire  LevelGateway_39__EVAL_1;
  wire  LevelGateway_39__EVAL_2;
  wire  LevelGateway_39__EVAL_3;
  wire  LevelGateway_39__EVAL_4;
  wire  LevelGateway_120__EVAL;
  wire  LevelGateway_120__EVAL_0;
  wire  LevelGateway_120__EVAL_1;
  wire  LevelGateway_120__EVAL_2;
  wire  LevelGateway_120__EVAL_3;
  wire  LevelGateway_120__EVAL_4;
  wire  LevelGateway_76__EVAL;
  wire  LevelGateway_76__EVAL_0;
  wire  LevelGateway_76__EVAL_1;
  wire  LevelGateway_76__EVAL_2;
  wire  LevelGateway_76__EVAL_3;
  wire  LevelGateway_76__EVAL_4;
  wire  LevelGateway_82__EVAL;
  wire  LevelGateway_82__EVAL_0;
  wire  LevelGateway_82__EVAL_1;
  wire  LevelGateway_82__EVAL_2;
  wire  LevelGateway_82__EVAL_3;
  wire  LevelGateway_82__EVAL_4;
  wire  LevelGateway_118__EVAL;
  wire  LevelGateway_118__EVAL_0;
  wire  LevelGateway_118__EVAL_1;
  wire  LevelGateway_118__EVAL_2;
  wire  LevelGateway_118__EVAL_3;
  wire  LevelGateway_118__EVAL_4;
  wire  LevelGateway_104__EVAL;
  wire  LevelGateway_104__EVAL_0;
  wire  LevelGateway_104__EVAL_1;
  wire  LevelGateway_104__EVAL_2;
  wire  LevelGateway_104__EVAL_3;
  wire  LevelGateway_104__EVAL_4;
  wire  LevelGateway_112__EVAL;
  wire  LevelGateway_112__EVAL_0;
  wire  LevelGateway_112__EVAL_1;
  wire  LevelGateway_112__EVAL_2;
  wire  LevelGateway_112__EVAL_3;
  wire  LevelGateway_112__EVAL_4;
  wire  LevelGateway_50__EVAL;
  wire  LevelGateway_50__EVAL_0;
  wire  LevelGateway_50__EVAL_1;
  wire  LevelGateway_50__EVAL_2;
  wire  LevelGateway_50__EVAL_3;
  wire  LevelGateway_50__EVAL_4;
  wire  LevelGateway_96__EVAL;
  wire  LevelGateway_96__EVAL_0;
  wire  LevelGateway_96__EVAL_1;
  wire  LevelGateway_96__EVAL_2;
  wire  LevelGateway_96__EVAL_3;
  wire  LevelGateway_96__EVAL_4;
  wire  LevelGateway_108__EVAL;
  wire  LevelGateway_108__EVAL_0;
  wire  LevelGateway_108__EVAL_1;
  wire  LevelGateway_108__EVAL_2;
  wire  LevelGateway_108__EVAL_3;
  wire  LevelGateway_108__EVAL_4;
  wire  LevelGateway_101__EVAL;
  wire  LevelGateway_101__EVAL_0;
  wire  LevelGateway_101__EVAL_1;
  wire  LevelGateway_101__EVAL_2;
  wire  LevelGateway_101__EVAL_3;
  wire  LevelGateway_101__EVAL_4;
  wire  LevelGateway_79__EVAL;
  wire  LevelGateway_79__EVAL_0;
  wire  LevelGateway_79__EVAL_1;
  wire  LevelGateway_79__EVAL_2;
  wire  LevelGateway_79__EVAL_3;
  wire  LevelGateway_79__EVAL_4;
  wire  LevelGateway_42__EVAL;
  wire  LevelGateway_42__EVAL_0;
  wire  LevelGateway_42__EVAL_1;
  wire  LevelGateway_42__EVAL_2;
  wire  LevelGateway_42__EVAL_3;
  wire  LevelGateway_42__EVAL_4;
  wire  LevelGateway_55__EVAL;
  wire  LevelGateway_55__EVAL_0;
  wire  LevelGateway_55__EVAL_1;
  wire  LevelGateway_55__EVAL_2;
  wire  LevelGateway_55__EVAL_3;
  wire  LevelGateway_55__EVAL_4;
  wire  LevelGateway_109__EVAL;
  wire  LevelGateway_109__EVAL_0;
  wire  LevelGateway_109__EVAL_1;
  wire  LevelGateway_109__EVAL_2;
  wire  LevelGateway_109__EVAL_3;
  wire  LevelGateway_109__EVAL_4;
  wire  LevelGateway_105__EVAL;
  wire  LevelGateway_105__EVAL_0;
  wire  LevelGateway_105__EVAL_1;
  wire  LevelGateway_105__EVAL_2;
  wire  LevelGateway_105__EVAL_3;
  wire  LevelGateway_105__EVAL_4;
  wire  LevelGateway_63__EVAL;
  wire  LevelGateway_63__EVAL_0;
  wire  LevelGateway_63__EVAL_1;
  wire  LevelGateway_63__EVAL_2;
  wire  LevelGateway_63__EVAL_3;
  wire  LevelGateway_63__EVAL_4;
  wire  LevelGateway_14__EVAL;
  wire  LevelGateway_14__EVAL_0;
  wire  LevelGateway_14__EVAL_1;
  wire  LevelGateway_14__EVAL_2;
  wire  LevelGateway_14__EVAL_3;
  wire  LevelGateway_14__EVAL_4;
  wire  LevelGateway_44__EVAL;
  wire  LevelGateway_44__EVAL_0;
  wire  LevelGateway_44__EVAL_1;
  wire  LevelGateway_44__EVAL_2;
  wire  LevelGateway_44__EVAL_3;
  wire  LevelGateway_44__EVAL_4;
  wire  LevelGateway_123__EVAL;
  wire  LevelGateway_123__EVAL_0;
  wire  LevelGateway_123__EVAL_1;
  wire  LevelGateway_123__EVAL_2;
  wire  LevelGateway_123__EVAL_3;
  wire  LevelGateway_123__EVAL_4;
  wire  LevelGateway_70__EVAL;
  wire  LevelGateway_70__EVAL_0;
  wire  LevelGateway_70__EVAL_1;
  wire  LevelGateway_70__EVAL_2;
  wire  LevelGateway_70__EVAL_3;
  wire  LevelGateway_70__EVAL_4;
  wire  LevelGateway_122__EVAL;
  wire  LevelGateway_122__EVAL_0;
  wire  LevelGateway_122__EVAL_1;
  wire  LevelGateway_122__EVAL_2;
  wire  LevelGateway_122__EVAL_3;
  wire  LevelGateway_122__EVAL_4;
  wire  LevelGateway_4__EVAL;
  wire  LevelGateway_4__EVAL_0;
  wire  LevelGateway_4__EVAL_1;
  wire  LevelGateway_4__EVAL_2;
  wire  LevelGateway_4__EVAL_3;
  wire  LevelGateway_4__EVAL_4;
  wire  LevelGateway_5__EVAL;
  wire  LevelGateway_5__EVAL_0;
  wire  LevelGateway_5__EVAL_1;
  wire  LevelGateway_5__EVAL_2;
  wire  LevelGateway_5__EVAL_3;
  wire  LevelGateway_5__EVAL_4;
  wire  LevelGateway_37__EVAL;
  wire  LevelGateway_37__EVAL_0;
  wire  LevelGateway_37__EVAL_1;
  wire  LevelGateway_37__EVAL_2;
  wire  LevelGateway_37__EVAL_3;
  wire  LevelGateway_37__EVAL_4;
  wire  LevelGateway_25__EVAL;
  wire  LevelGateway_25__EVAL_0;
  wire  LevelGateway_25__EVAL_1;
  wire  LevelGateway_25__EVAL_2;
  wire  LevelGateway_25__EVAL_3;
  wire  LevelGateway_25__EVAL_4;
  wire  LevelGateway_114__EVAL;
  wire  LevelGateway_114__EVAL_0;
  wire  LevelGateway_114__EVAL_1;
  wire  LevelGateway_114__EVAL_2;
  wire  LevelGateway_114__EVAL_3;
  wire  LevelGateway_114__EVAL_4;
  wire  LevelGateway_56__EVAL;
  wire  LevelGateway_56__EVAL_0;
  wire  LevelGateway_56__EVAL_1;
  wire  LevelGateway_56__EVAL_2;
  wire  LevelGateway_56__EVAL_3;
  wire  LevelGateway_56__EVAL_4;
  wire  LevelGateway_71__EVAL;
  wire  LevelGateway_71__EVAL_0;
  wire  LevelGateway_71__EVAL_1;
  wire  LevelGateway_71__EVAL_2;
  wire  LevelGateway_71__EVAL_3;
  wire  LevelGateway_71__EVAL_4;
  wire  LevelGateway_64__EVAL;
  wire  LevelGateway_64__EVAL_0;
  wire  LevelGateway_64__EVAL_1;
  wire  LevelGateway_64__EVAL_2;
  wire  LevelGateway_64__EVAL_3;
  wire  LevelGateway_64__EVAL_4;
  wire [31:0] Queue__EVAL;
  wire [13:0] Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire [13:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire [23:0] Queue__EVAL_6;
  wire [31:0] Queue__EVAL_7;
  wire [23:0] Queue__EVAL_8;
  wire  Queue__EVAL_9;
  wire [3:0] Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire  Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire [3:0] Queue__EVAL_14;
  wire  LevelGateway_73__EVAL;
  wire  LevelGateway_73__EVAL_0;
  wire  LevelGateway_73__EVAL_1;
  wire  LevelGateway_73__EVAL_2;
  wire  LevelGateway_73__EVAL_3;
  wire  LevelGateway_73__EVAL_4;
  wire  LevelGateway_99__EVAL;
  wire  LevelGateway_99__EVAL_0;
  wire  LevelGateway_99__EVAL_1;
  wire  LevelGateway_99__EVAL_2;
  wire  LevelGateway_99__EVAL_3;
  wire  LevelGateway_99__EVAL_4;
  wire  LevelGateway_115__EVAL;
  wire  LevelGateway_115__EVAL_0;
  wire  LevelGateway_115__EVAL_1;
  wire  LevelGateway_115__EVAL_2;
  wire  LevelGateway_115__EVAL_3;
  wire  LevelGateway_115__EVAL_4;
  wire  LevelGateway_94__EVAL;
  wire  LevelGateway_94__EVAL_0;
  wire  LevelGateway_94__EVAL_1;
  wire  LevelGateway_94__EVAL_2;
  wire  LevelGateway_94__EVAL_3;
  wire  LevelGateway_94__EVAL_4;
  wire  LevelGateway_49__EVAL;
  wire  LevelGateway_49__EVAL_0;
  wire  LevelGateway_49__EVAL_1;
  wire  LevelGateway_49__EVAL_2;
  wire  LevelGateway_49__EVAL_3;
  wire  LevelGateway_49__EVAL_4;
  wire  LevelGateway_48__EVAL;
  wire  LevelGateway_48__EVAL_0;
  wire  LevelGateway_48__EVAL_1;
  wire  LevelGateway_48__EVAL_2;
  wire  LevelGateway_48__EVAL_3;
  wire  LevelGateway_48__EVAL_4;
  wire  LevelGateway_62__EVAL;
  wire  LevelGateway_62__EVAL_0;
  wire  LevelGateway_62__EVAL_1;
  wire  LevelGateway_62__EVAL_2;
  wire  LevelGateway_62__EVAL_3;
  wire  LevelGateway_62__EVAL_4;
  wire  LevelGateway_103__EVAL;
  wire  LevelGateway_103__EVAL_0;
  wire  LevelGateway_103__EVAL_1;
  wire  LevelGateway_103__EVAL_2;
  wire  LevelGateway_103__EVAL_3;
  wire  LevelGateway_103__EVAL_4;
  wire  LevelGateway_15__EVAL;
  wire  LevelGateway_15__EVAL_0;
  wire  LevelGateway_15__EVAL_1;
  wire  LevelGateway_15__EVAL_2;
  wire  LevelGateway_15__EVAL_3;
  wire  LevelGateway_15__EVAL_4;
  wire  LevelGateway_102__EVAL;
  wire  LevelGateway_102__EVAL_0;
  wire  LevelGateway_102__EVAL_1;
  wire  LevelGateway_102__EVAL_2;
  wire  LevelGateway_102__EVAL_3;
  wire  LevelGateway_102__EVAL_4;
  wire  LevelGateway_83__EVAL;
  wire  LevelGateway_83__EVAL_0;
  wire  LevelGateway_83__EVAL_1;
  wire  LevelGateway_83__EVAL_2;
  wire  LevelGateway_83__EVAL_3;
  wire  LevelGateway_83__EVAL_4;
  wire  LevelGateway_95__EVAL;
  wire  LevelGateway_95__EVAL_0;
  wire  LevelGateway_95__EVAL_1;
  wire  LevelGateway_95__EVAL_2;
  wire  LevelGateway_95__EVAL_3;
  wire  LevelGateway_95__EVAL_4;
  wire  LevelGateway_38__EVAL;
  wire  LevelGateway_38__EVAL_0;
  wire  LevelGateway_38__EVAL_1;
  wire  LevelGateway_38__EVAL_2;
  wire  LevelGateway_38__EVAL_3;
  wire  LevelGateway_38__EVAL_4;
  wire  LevelGateway_29__EVAL;
  wire  LevelGateway_29__EVAL_0;
  wire  LevelGateway_29__EVAL_1;
  wire  LevelGateway_29__EVAL_2;
  wire  LevelGateway_29__EVAL_3;
  wire  LevelGateway_29__EVAL_4;
  wire  LevelGateway_35__EVAL;
  wire  LevelGateway_35__EVAL_0;
  wire  LevelGateway_35__EVAL_1;
  wire  LevelGateway_35__EVAL_2;
  wire  LevelGateway_35__EVAL_3;
  wire  LevelGateway_35__EVAL_4;
  wire  LevelGateway_9__EVAL;
  wire  LevelGateway_9__EVAL_0;
  wire  LevelGateway_9__EVAL_1;
  wire  LevelGateway_9__EVAL_2;
  wire  LevelGateway_9__EVAL_3;
  wire  LevelGateway_9__EVAL_4;
  wire  LevelGateway_86__EVAL;
  wire  LevelGateway_86__EVAL_0;
  wire  LevelGateway_86__EVAL_1;
  wire  LevelGateway_86__EVAL_2;
  wire  LevelGateway_86__EVAL_3;
  wire  LevelGateway_86__EVAL_4;
  wire  LevelGateway_100__EVAL;
  wire  LevelGateway_100__EVAL_0;
  wire  LevelGateway_100__EVAL_1;
  wire  LevelGateway_100__EVAL_2;
  wire  LevelGateway_100__EVAL_3;
  wire  LevelGateway_100__EVAL_4;
  wire  LevelGateway_69__EVAL;
  wire  LevelGateway_69__EVAL_0;
  wire  LevelGateway_69__EVAL_1;
  wire  LevelGateway_69__EVAL_2;
  wire  LevelGateway_69__EVAL_3;
  wire  LevelGateway_69__EVAL_4;
  wire  LevelGateway_81__EVAL;
  wire  LevelGateway_81__EVAL_0;
  wire  LevelGateway_81__EVAL_1;
  wire  LevelGateway_81__EVAL_2;
  wire  LevelGateway_81__EVAL_3;
  wire  LevelGateway_81__EVAL_4;
  wire  LevelGateway_75__EVAL;
  wire  LevelGateway_75__EVAL_0;
  wire  LevelGateway_75__EVAL_1;
  wire  LevelGateway_75__EVAL_2;
  wire  LevelGateway_75__EVAL_3;
  wire  LevelGateway_75__EVAL_4;
  wire  LevelGateway_66__EVAL;
  wire  LevelGateway_66__EVAL_0;
  wire  LevelGateway_66__EVAL_1;
  wire  LevelGateway_66__EVAL_2;
  wire  LevelGateway_66__EVAL_3;
  wire  LevelGateway_66__EVAL_4;
  wire  LevelGateway_10__EVAL;
  wire  LevelGateway_10__EVAL_0;
  wire  LevelGateway_10__EVAL_1;
  wire  LevelGateway_10__EVAL_2;
  wire  LevelGateway_10__EVAL_3;
  wire  LevelGateway_10__EVAL_4;
  wire  LevelGateway_91__EVAL;
  wire  LevelGateway_91__EVAL_0;
  wire  LevelGateway_91__EVAL_1;
  wire  LevelGateway_91__EVAL_2;
  wire  LevelGateway_91__EVAL_3;
  wire  LevelGateway_91__EVAL_4;
  wire  LevelGateway_67__EVAL;
  wire  LevelGateway_67__EVAL_0;
  wire  LevelGateway_67__EVAL_1;
  wire  LevelGateway_67__EVAL_2;
  wire  LevelGateway_67__EVAL_3;
  wire  LevelGateway_67__EVAL_4;
  wire  LevelGateway_27__EVAL;
  wire  LevelGateway_27__EVAL_0;
  wire  LevelGateway_27__EVAL_1;
  wire  LevelGateway_27__EVAL_2;
  wire  LevelGateway_27__EVAL_3;
  wire  LevelGateway_27__EVAL_4;
  wire  LevelGateway_89__EVAL;
  wire  LevelGateway_89__EVAL_0;
  wire  LevelGateway_89__EVAL_1;
  wire  LevelGateway_89__EVAL_2;
  wire  LevelGateway_89__EVAL_3;
  wire  LevelGateway_89__EVAL_4;
  wire  LevelGateway_12__EVAL;
  wire  LevelGateway_12__EVAL_0;
  wire  LevelGateway_12__EVAL_1;
  wire  LevelGateway_12__EVAL_2;
  wire  LevelGateway_12__EVAL_3;
  wire  LevelGateway_12__EVAL_4;
  wire  LevelGateway_28__EVAL;
  wire  LevelGateway_28__EVAL_0;
  wire  LevelGateway_28__EVAL_1;
  wire  LevelGateway_28__EVAL_2;
  wire  LevelGateway_28__EVAL_3;
  wire  LevelGateway_28__EVAL_4;
  wire  LevelGateway_58__EVAL;
  wire  LevelGateway_58__EVAL_0;
  wire  LevelGateway_58__EVAL_1;
  wire  LevelGateway_58__EVAL_2;
  wire  LevelGateway_58__EVAL_3;
  wire  LevelGateway_58__EVAL_4;
  wire  LevelGateway_6__EVAL;
  wire  LevelGateway_6__EVAL_0;
  wire  LevelGateway_6__EVAL_1;
  wire  LevelGateway_6__EVAL_2;
  wire  LevelGateway_6__EVAL_3;
  wire  LevelGateway_6__EVAL_4;
  wire  LevelGateway_98__EVAL;
  wire  LevelGateway_98__EVAL_0;
  wire  LevelGateway_98__EVAL_1;
  wire  LevelGateway_98__EVAL_2;
  wire  LevelGateway_98__EVAL_3;
  wire  LevelGateway_98__EVAL_4;
  wire  LevelGateway_107__EVAL;
  wire  LevelGateway_107__EVAL_0;
  wire  LevelGateway_107__EVAL_1;
  wire  LevelGateway_107__EVAL_2;
  wire  LevelGateway_107__EVAL_3;
  wire  LevelGateway_107__EVAL_4;
  wire  LevelGateway_93__EVAL;
  wire  LevelGateway_93__EVAL_0;
  wire  LevelGateway_93__EVAL_1;
  wire  LevelGateway_93__EVAL_2;
  wire  LevelGateway_93__EVAL_3;
  wire  LevelGateway_93__EVAL_4;
  wire  LevelGateway_126__EVAL;
  wire  LevelGateway_126__EVAL_0;
  wire  LevelGateway_126__EVAL_1;
  wire  LevelGateway_126__EVAL_2;
  wire  LevelGateway_126__EVAL_3;
  wire  LevelGateway_126__EVAL_4;
  wire  LevelGateway_97__EVAL;
  wire  LevelGateway_97__EVAL_0;
  wire  LevelGateway_97__EVAL_1;
  wire  LevelGateway_97__EVAL_2;
  wire  LevelGateway_97__EVAL_3;
  wire  LevelGateway_97__EVAL_4;
  wire  LevelGateway_57__EVAL;
  wire  LevelGateway_57__EVAL_0;
  wire  LevelGateway_57__EVAL_1;
  wire  LevelGateway_57__EVAL_2;
  wire  LevelGateway_57__EVAL_3;
  wire  LevelGateway_57__EVAL_4;
  wire  LevelGateway_72__EVAL;
  wire  LevelGateway_72__EVAL_0;
  wire  LevelGateway_72__EVAL_1;
  wire  LevelGateway_72__EVAL_2;
  wire  LevelGateway_72__EVAL_3;
  wire  LevelGateway_72__EVAL_4;
  wire [2:0] PLICFanIn__EVAL;
  wire [2:0] PLICFanIn__EVAL_0;
  wire [2:0] PLICFanIn__EVAL_1;
  wire [2:0] PLICFanIn__EVAL_2;
  wire [2:0] PLICFanIn__EVAL_3;
  wire [2:0] PLICFanIn__EVAL_4;
  wire [2:0] PLICFanIn__EVAL_5;
  wire [2:0] PLICFanIn__EVAL_6;
  wire [2:0] PLICFanIn__EVAL_7;
  wire [2:0] PLICFanIn__EVAL_8;
  wire [2:0] PLICFanIn__EVAL_9;
  wire [2:0] PLICFanIn__EVAL_10;
  wire [2:0] PLICFanIn__EVAL_11;
  wire [2:0] PLICFanIn__EVAL_12;
  wire [2:0] PLICFanIn__EVAL_13;
  wire [2:0] PLICFanIn__EVAL_14;
  wire [2:0] PLICFanIn__EVAL_15;
  wire [2:0] PLICFanIn__EVAL_16;
  wire [2:0] PLICFanIn__EVAL_17;
  wire [2:0] PLICFanIn__EVAL_18;
  wire [2:0] PLICFanIn__EVAL_19;
  wire [2:0] PLICFanIn__EVAL_20;
  wire [2:0] PLICFanIn__EVAL_21;
  wire [2:0] PLICFanIn__EVAL_22;
  wire [2:0] PLICFanIn__EVAL_23;
  wire [2:0] PLICFanIn__EVAL_24;
  wire [2:0] PLICFanIn__EVAL_25;
  wire [2:0] PLICFanIn__EVAL_26;
  wire [2:0] PLICFanIn__EVAL_27;
  wire [2:0] PLICFanIn__EVAL_28;
  wire [2:0] PLICFanIn__EVAL_29;
  wire [2:0] PLICFanIn__EVAL_30;
  wire [2:0] PLICFanIn__EVAL_31;
  wire [2:0] PLICFanIn__EVAL_32;
  wire [2:0] PLICFanIn__EVAL_33;
  wire [2:0] PLICFanIn__EVAL_34;
  wire [2:0] PLICFanIn__EVAL_35;
  wire [6:0] PLICFanIn__EVAL_36;
  wire [2:0] PLICFanIn__EVAL_37;
  wire [2:0] PLICFanIn__EVAL_38;
  wire [2:0] PLICFanIn__EVAL_39;
  wire [2:0] PLICFanIn__EVAL_40;
  wire [2:0] PLICFanIn__EVAL_41;
  wire [2:0] PLICFanIn__EVAL_42;
  wire [2:0] PLICFanIn__EVAL_43;
  wire [2:0] PLICFanIn__EVAL_44;
  wire [2:0] PLICFanIn__EVAL_45;
  wire [2:0] PLICFanIn__EVAL_46;
  wire [2:0] PLICFanIn__EVAL_47;
  wire [2:0] PLICFanIn__EVAL_48;
  wire [2:0] PLICFanIn__EVAL_49;
  wire [2:0] PLICFanIn__EVAL_50;
  wire [2:0] PLICFanIn__EVAL_51;
  wire [2:0] PLICFanIn__EVAL_52;
  wire [2:0] PLICFanIn__EVAL_53;
  wire [2:0] PLICFanIn__EVAL_54;
  wire [2:0] PLICFanIn__EVAL_55;
  wire [2:0] PLICFanIn__EVAL_56;
  wire [2:0] PLICFanIn__EVAL_57;
  wire [2:0] PLICFanIn__EVAL_58;
  wire [2:0] PLICFanIn__EVAL_59;
  wire [2:0] PLICFanIn__EVAL_60;
  wire [2:0] PLICFanIn__EVAL_61;
  wire [2:0] PLICFanIn__EVAL_62;
  wire [2:0] PLICFanIn__EVAL_63;
  wire [2:0] PLICFanIn__EVAL_64;
  wire [2:0] PLICFanIn__EVAL_65;
  wire [2:0] PLICFanIn__EVAL_66;
  wire [2:0] PLICFanIn__EVAL_67;
  wire [2:0] PLICFanIn__EVAL_68;
  wire [2:0] PLICFanIn__EVAL_69;
  wire [2:0] PLICFanIn__EVAL_70;
  wire [2:0] PLICFanIn__EVAL_71;
  wire [2:0] PLICFanIn__EVAL_72;
  wire [2:0] PLICFanIn__EVAL_73;
  wire [2:0] PLICFanIn__EVAL_74;
  wire [2:0] PLICFanIn__EVAL_75;
  wire [2:0] PLICFanIn__EVAL_76;
  wire [2:0] PLICFanIn__EVAL_77;
  wire [2:0] PLICFanIn__EVAL_78;
  wire [2:0] PLICFanIn__EVAL_79;
  wire [2:0] PLICFanIn__EVAL_80;
  wire [2:0] PLICFanIn__EVAL_81;
  wire [2:0] PLICFanIn__EVAL_82;
  wire [2:0] PLICFanIn__EVAL_83;
  wire [2:0] PLICFanIn__EVAL_84;
  wire [2:0] PLICFanIn__EVAL_85;
  wire [2:0] PLICFanIn__EVAL_86;
  wire [2:0] PLICFanIn__EVAL_87;
  wire [2:0] PLICFanIn__EVAL_88;
  wire [2:0] PLICFanIn__EVAL_89;
  wire [2:0] PLICFanIn__EVAL_90;
  wire [2:0] PLICFanIn__EVAL_91;
  wire [2:0] PLICFanIn__EVAL_92;
  wire [2:0] PLICFanIn__EVAL_93;
  wire [2:0] PLICFanIn__EVAL_94;
  wire [2:0] PLICFanIn__EVAL_95;
  wire [2:0] PLICFanIn__EVAL_96;
  wire [2:0] PLICFanIn__EVAL_97;
  wire [2:0] PLICFanIn__EVAL_98;
  wire [2:0] PLICFanIn__EVAL_99;
  wire [2:0] PLICFanIn__EVAL_100;
  wire [2:0] PLICFanIn__EVAL_101;
  wire [2:0] PLICFanIn__EVAL_102;
  wire [2:0] PLICFanIn__EVAL_103;
  wire [2:0] PLICFanIn__EVAL_104;
  wire [2:0] PLICFanIn__EVAL_105;
  wire [2:0] PLICFanIn__EVAL_106;
  wire [2:0] PLICFanIn__EVAL_107;
  wire [2:0] PLICFanIn__EVAL_108;
  wire [2:0] PLICFanIn__EVAL_109;
  wire [2:0] PLICFanIn__EVAL_110;
  wire [2:0] PLICFanIn__EVAL_111;
  wire [2:0] PLICFanIn__EVAL_112;
  wire [126:0] PLICFanIn__EVAL_113;
  wire [2:0] PLICFanIn__EVAL_114;
  wire [2:0] PLICFanIn__EVAL_115;
  wire [2:0] PLICFanIn__EVAL_116;
  wire [2:0] PLICFanIn__EVAL_117;
  wire [2:0] PLICFanIn__EVAL_118;
  wire [2:0] PLICFanIn__EVAL_119;
  wire [2:0] PLICFanIn__EVAL_120;
  wire [2:0] PLICFanIn__EVAL_121;
  wire [2:0] PLICFanIn__EVAL_122;
  wire [2:0] PLICFanIn__EVAL_123;
  wire [2:0] PLICFanIn__EVAL_124;
  wire [2:0] PLICFanIn__EVAL_125;
  wire [2:0] PLICFanIn__EVAL_126;
  wire [2:0] PLICFanIn__EVAL_127;
  wire [2:0] PLICFanIn__EVAL_128;
  wire  LevelGateway_43__EVAL;
  wire  LevelGateway_43__EVAL_0;
  wire  LevelGateway_43__EVAL_1;
  wire  LevelGateway_43__EVAL_2;
  wire  LevelGateway_43__EVAL_3;
  wire  LevelGateway_43__EVAL_4;
  wire  LevelGateway_30__EVAL;
  wire  LevelGateway_30__EVAL_0;
  wire  LevelGateway_30__EVAL_1;
  wire  LevelGateway_30__EVAL_2;
  wire  LevelGateway_30__EVAL_3;
  wire  LevelGateway_30__EVAL_4;
  wire  LevelGateway_7__EVAL;
  wire  LevelGateway_7__EVAL_0;
  wire  LevelGateway_7__EVAL_1;
  wire  LevelGateway_7__EVAL_2;
  wire  LevelGateway_7__EVAL_3;
  wire  LevelGateway_7__EVAL_4;
  wire  LevelGateway_68__EVAL;
  wire  LevelGateway_68__EVAL_0;
  wire  LevelGateway_68__EVAL_1;
  wire  LevelGateway_68__EVAL_2;
  wire  LevelGateway_68__EVAL_3;
  wire  LevelGateway_68__EVAL_4;
  wire  LevelGateway_84__EVAL;
  wire  LevelGateway_84__EVAL_0;
  wire  LevelGateway_84__EVAL_1;
  wire  LevelGateway_84__EVAL_2;
  wire  LevelGateway_84__EVAL_3;
  wire  LevelGateway_84__EVAL_4;
  wire  LevelGateway_116__EVAL;
  wire  LevelGateway_116__EVAL_0;
  wire  LevelGateway_116__EVAL_1;
  wire  LevelGateway_116__EVAL_2;
  wire  LevelGateway_116__EVAL_3;
  wire  LevelGateway_116__EVAL_4;
  wire  LevelGateway_53__EVAL;
  wire  LevelGateway_53__EVAL_0;
  wire  LevelGateway_53__EVAL_1;
  wire  LevelGateway_53__EVAL_2;
  wire  LevelGateway_53__EVAL_3;
  wire  LevelGateway_53__EVAL_4;
  wire  LevelGateway_88__EVAL;
  wire  LevelGateway_88__EVAL_0;
  wire  LevelGateway_88__EVAL_1;
  wire  LevelGateway_88__EVAL_2;
  wire  LevelGateway_88__EVAL_3;
  wire  LevelGateway_88__EVAL_4;
  wire  LevelGateway_13__EVAL;
  wire  LevelGateway_13__EVAL_0;
  wire  LevelGateway_13__EVAL_1;
  wire  LevelGateway_13__EVAL_2;
  wire  LevelGateway_13__EVAL_3;
  wire  LevelGateway_13__EVAL_4;
  wire  LevelGateway_117__EVAL;
  wire  LevelGateway_117__EVAL_0;
  wire  LevelGateway_117__EVAL_1;
  wire  LevelGateway_117__EVAL_2;
  wire  LevelGateway_117__EVAL_3;
  wire  LevelGateway_117__EVAL_4;
  wire  LevelGateway_3__EVAL;
  wire  LevelGateway_3__EVAL_0;
  wire  LevelGateway_3__EVAL_1;
  wire  LevelGateway_3__EVAL_2;
  wire  LevelGateway_3__EVAL_3;
  wire  LevelGateway_3__EVAL_4;
  wire  LevelGateway_47__EVAL;
  wire  LevelGateway_47__EVAL_0;
  wire  LevelGateway_47__EVAL_1;
  wire  LevelGateway_47__EVAL_2;
  wire  LevelGateway_47__EVAL_3;
  wire  LevelGateway_47__EVAL_4;
  wire  LevelGateway_85__EVAL;
  wire  LevelGateway_85__EVAL_0;
  wire  LevelGateway_85__EVAL_1;
  wire  LevelGateway_85__EVAL_2;
  wire  LevelGateway_85__EVAL_3;
  wire  LevelGateway_85__EVAL_4;
  wire  LevelGateway_46__EVAL;
  wire  LevelGateway_46__EVAL_0;
  wire  LevelGateway_46__EVAL_1;
  wire  LevelGateway_46__EVAL_2;
  wire  LevelGateway_46__EVAL_3;
  wire  LevelGateway_46__EVAL_4;
  wire  LevelGateway_60__EVAL;
  wire  LevelGateway_60__EVAL_0;
  wire  LevelGateway_60__EVAL_1;
  wire  LevelGateway_60__EVAL_2;
  wire  LevelGateway_60__EVAL_3;
  wire  LevelGateway_60__EVAL_4;
  wire  LevelGateway_20__EVAL;
  wire  LevelGateway_20__EVAL_0;
  wire  LevelGateway_20__EVAL_1;
  wire  LevelGateway_20__EVAL_2;
  wire  LevelGateway_20__EVAL_3;
  wire  LevelGateway_20__EVAL_4;
  wire  LevelGateway_17__EVAL;
  wire  LevelGateway_17__EVAL_0;
  wire  LevelGateway_17__EVAL_1;
  wire  LevelGateway_17__EVAL_2;
  wire  LevelGateway_17__EVAL_3;
  wire  LevelGateway_17__EVAL_4;
  wire  LevelGateway_59__EVAL;
  wire  LevelGateway_59__EVAL_0;
  wire  LevelGateway_59__EVAL_1;
  wire  LevelGateway_59__EVAL_2;
  wire  LevelGateway_59__EVAL_3;
  wire  LevelGateway_59__EVAL_4;
  wire  LevelGateway_124__EVAL;
  wire  LevelGateway_124__EVAL_0;
  wire  LevelGateway_124__EVAL_1;
  wire  LevelGateway_124__EVAL_2;
  wire  LevelGateway_124__EVAL_3;
  wire  LevelGateway_124__EVAL_4;
  wire  LevelGateway_61__EVAL;
  wire  LevelGateway_61__EVAL_0;
  wire  LevelGateway_61__EVAL_1;
  wire  LevelGateway_61__EVAL_2;
  wire  LevelGateway_61__EVAL_3;
  wire  LevelGateway_61__EVAL_4;
  wire  LevelGateway_2__EVAL;
  wire  LevelGateway_2__EVAL_0;
  wire  LevelGateway_2__EVAL_1;
  wire  LevelGateway_2__EVAL_2;
  wire  LevelGateway_2__EVAL_3;
  wire  LevelGateway_2__EVAL_4;
  wire  LevelGateway_40__EVAL;
  wire  LevelGateway_40__EVAL_0;
  wire  LevelGateway_40__EVAL_1;
  wire  LevelGateway_40__EVAL_2;
  wire  LevelGateway_40__EVAL_3;
  wire  LevelGateway_40__EVAL_4;
  wire  LevelGateway_33__EVAL;
  wire  LevelGateway_33__EVAL_0;
  wire  LevelGateway_33__EVAL_1;
  wire  LevelGateway_33__EVAL_2;
  wire  LevelGateway_33__EVAL_3;
  wire  LevelGateway_33__EVAL_4;
  wire  LevelGateway_21__EVAL;
  wire  LevelGateway_21__EVAL_0;
  wire  LevelGateway_21__EVAL_1;
  wire  LevelGateway_21__EVAL_2;
  wire  LevelGateway_21__EVAL_3;
  wire  LevelGateway_21__EVAL_4;
  wire  LevelGateway_26__EVAL;
  wire  LevelGateway_26__EVAL_0;
  wire  LevelGateway_26__EVAL_1;
  wire  LevelGateway_26__EVAL_2;
  wire  LevelGateway_26__EVAL_3;
  wire  LevelGateway_26__EVAL_4;
  wire  LevelGateway_110__EVAL;
  wire  LevelGateway_110__EVAL_0;
  wire  LevelGateway_110__EVAL_1;
  wire  LevelGateway_110__EVAL_2;
  wire  LevelGateway_110__EVAL_3;
  wire  LevelGateway_110__EVAL_4;
  wire  LevelGateway_90__EVAL;
  wire  LevelGateway_90__EVAL_0;
  wire  LevelGateway_90__EVAL_1;
  wire  LevelGateway_90__EVAL_2;
  wire  LevelGateway_90__EVAL_3;
  wire  LevelGateway_90__EVAL_4;
  wire  LevelGateway_119__EVAL;
  wire  LevelGateway_119__EVAL_0;
  wire  LevelGateway_119__EVAL_1;
  wire  LevelGateway_119__EVAL_2;
  wire  LevelGateway_119__EVAL_3;
  wire  LevelGateway_119__EVAL_4;
  wire  LevelGateway_23__EVAL;
  wire  LevelGateway_23__EVAL_0;
  wire  LevelGateway_23__EVAL_1;
  wire  LevelGateway_23__EVAL_2;
  wire  LevelGateway_23__EVAL_3;
  wire  LevelGateway_23__EVAL_4;
  wire  LevelGateway_80__EVAL;
  wire  LevelGateway_80__EVAL_0;
  wire  LevelGateway_80__EVAL_1;
  wire  LevelGateway_80__EVAL_2;
  wire  LevelGateway_80__EVAL_3;
  wire  LevelGateway_80__EVAL_4;
  wire  LevelGateway_41__EVAL;
  wire  LevelGateway_41__EVAL_0;
  wire  LevelGateway_41__EVAL_1;
  wire  LevelGateway_41__EVAL_2;
  wire  LevelGateway_41__EVAL_3;
  wire  LevelGateway_41__EVAL_4;
  wire  LevelGateway_78__EVAL;
  wire  LevelGateway_78__EVAL_0;
  wire  LevelGateway_78__EVAL_1;
  wire  LevelGateway_78__EVAL_2;
  wire  LevelGateway_78__EVAL_3;
  wire  LevelGateway_78__EVAL_4;
  wire  LevelGateway_121__EVAL;
  wire  LevelGateway_121__EVAL_0;
  wire  LevelGateway_121__EVAL_1;
  wire  LevelGateway_121__EVAL_2;
  wire  LevelGateway_121__EVAL_3;
  wire  LevelGateway_121__EVAL_4;
  wire  LevelGateway_31__EVAL;
  wire  LevelGateway_31__EVAL_0;
  wire  LevelGateway_31__EVAL_1;
  wire  LevelGateway_31__EVAL_2;
  wire  LevelGateway_31__EVAL_3;
  wire  LevelGateway_31__EVAL_4;
  wire  LevelGateway_19__EVAL;
  wire  LevelGateway_19__EVAL_0;
  wire  LevelGateway_19__EVAL_1;
  wire  LevelGateway_19__EVAL_2;
  wire  LevelGateway_19__EVAL_3;
  wire  LevelGateway_19__EVAL_4;
  wire  LevelGateway_113__EVAL;
  wire  LevelGateway_113__EVAL_0;
  wire  LevelGateway_113__EVAL_1;
  wire  LevelGateway_113__EVAL_2;
  wire  LevelGateway_113__EVAL_3;
  wire  LevelGateway_113__EVAL_4;
  wire  LevelGateway_111__EVAL;
  wire  LevelGateway_111__EVAL_0;
  wire  LevelGateway_111__EVAL_1;
  wire  LevelGateway_111__EVAL_2;
  wire  LevelGateway_111__EVAL_3;
  wire  LevelGateway_111__EVAL_4;
  wire  LevelGateway_77__EVAL;
  wire  LevelGateway_77__EVAL_0;
  wire  LevelGateway_77__EVAL_1;
  wire  LevelGateway_77__EVAL_2;
  wire  LevelGateway_77__EVAL_3;
  wire  LevelGateway_77__EVAL_4;
  wire  LevelGateway_11__EVAL;
  wire  LevelGateway_11__EVAL_0;
  wire  LevelGateway_11__EVAL_1;
  wire  LevelGateway_11__EVAL_2;
  wire  LevelGateway_11__EVAL_3;
  wire  LevelGateway_11__EVAL_4;
  wire  LevelGateway_36__EVAL;
  wire  LevelGateway_36__EVAL_0;
  wire  LevelGateway_36__EVAL_1;
  wire  LevelGateway_36__EVAL_2;
  wire  LevelGateway_36__EVAL_3;
  wire  LevelGateway_36__EVAL_4;
  wire  LevelGateway_24__EVAL;
  wire  LevelGateway_24__EVAL_0;
  wire  LevelGateway_24__EVAL_1;
  wire  LevelGateway_24__EVAL_2;
  wire  LevelGateway_24__EVAL_3;
  wire  LevelGateway_24__EVAL_4;
  wire  LevelGateway_125__EVAL;
  wire  LevelGateway_125__EVAL_0;
  wire  LevelGateway_125__EVAL_1;
  wire  LevelGateway_125__EVAL_2;
  wire  LevelGateway_125__EVAL_3;
  wire  LevelGateway_125__EVAL_4;
  wire  LevelGateway_45__EVAL;
  wire  LevelGateway_45__EVAL_0;
  wire  LevelGateway_45__EVAL_1;
  wire  LevelGateway_45__EVAL_2;
  wire  LevelGateway_45__EVAL_3;
  wire  LevelGateway_45__EVAL_4;
  wire  LevelGateway_106__EVAL;
  wire  LevelGateway_106__EVAL_0;
  wire  LevelGateway_106__EVAL_1;
  wire  LevelGateway_106__EVAL_2;
  wire  LevelGateway_106__EVAL_3;
  wire  LevelGateway_106__EVAL_4;
  wire  LevelGateway_8__EVAL;
  wire  LevelGateway_8__EVAL_0;
  wire  LevelGateway_8__EVAL_1;
  wire  LevelGateway_8__EVAL_2;
  wire  LevelGateway_8__EVAL_3;
  wire  LevelGateway_8__EVAL_4;
  wire  LevelGateway_1__EVAL;
  wire  LevelGateway_1__EVAL_0;
  wire  LevelGateway_1__EVAL_1;
  wire  LevelGateway_1__EVAL_2;
  wire  LevelGateway_1__EVAL_3;
  wire  LevelGateway_1__EVAL_4;
  wire  LevelGateway_52__EVAL;
  wire  LevelGateway_52__EVAL_0;
  wire  LevelGateway_52__EVAL_1;
  wire  LevelGateway_52__EVAL_2;
  wire  LevelGateway_52__EVAL_3;
  wire  LevelGateway_52__EVAL_4;
  wire  LevelGateway_87__EVAL;
  wire  LevelGateway_87__EVAL_0;
  wire  LevelGateway_87__EVAL_1;
  wire  LevelGateway_87__EVAL_2;
  wire  LevelGateway_87__EVAL_3;
  wire  LevelGateway_87__EVAL_4;
  wire  LevelGateway_74__EVAL;
  wire  LevelGateway_74__EVAL_0;
  wire  LevelGateway_74__EVAL_1;
  wire  LevelGateway_74__EVAL_2;
  wire  LevelGateway_74__EVAL_3;
  wire  LevelGateway_74__EVAL_4;
  wire  LevelGateway_18__EVAL;
  wire  LevelGateway_18__EVAL_0;
  wire  LevelGateway_18__EVAL_1;
  wire  LevelGateway_18__EVAL_2;
  wire  LevelGateway_18__EVAL_3;
  wire  LevelGateway_18__EVAL_4;
  wire  LevelGateway_22__EVAL;
  wire  LevelGateway_22__EVAL_0;
  wire  LevelGateway_22__EVAL_1;
  wire  LevelGateway_22__EVAL_2;
  wire  LevelGateway_22__EVAL_3;
  wire  LevelGateway_22__EVAL_4;
  wire  LevelGateway_51__EVAL;
  wire  LevelGateway_51__EVAL_0;
  wire  LevelGateway_51__EVAL_1;
  wire  LevelGateway_51__EVAL_2;
  wire  LevelGateway_51__EVAL_3;
  wire  LevelGateway_51__EVAL_4;
  wire  LevelGateway_32__EVAL;
  wire  LevelGateway_32__EVAL_0;
  wire  LevelGateway_32__EVAL_1;
  wire  LevelGateway_32__EVAL_2;
  wire  LevelGateway_32__EVAL_3;
  wire  LevelGateway_32__EVAL_4;
  reg [2:0] _EVAL_147;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_155;
  reg [31:0] _RAND_1;
  reg  _EVAL_163;
  reg [31:0] _RAND_2;
  reg  _EVAL_176;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_188;
  reg [31:0] _RAND_4;
  reg  _EVAL_194;
  reg [31:0] _RAND_5;
  reg  _EVAL_200;
  reg [31:0] _RAND_6;
  reg  _EVAL_212;
  reg [31:0] _RAND_7;
  reg  _EVAL_217;
  reg [31:0] _RAND_8;
  reg  _EVAL_222;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_247;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_251;
  reg [31:0] _RAND_11;
  reg  _EVAL_269;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_285;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_286;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_293;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_304;
  reg [31:0] _RAND_16;
  reg  _EVAL_306;
  reg [31:0] _RAND_17;
  reg [2:0] _EVAL_331;
  reg [31:0] _RAND_18;
  reg [2:0] _EVAL_354;
  reg [31:0] _RAND_19;
  reg [7:0] _EVAL_366;
  reg [31:0] _RAND_20;
  reg  _EVAL_371;
  reg [31:0] _RAND_21;
  reg  _EVAL_387;
  reg [31:0] _RAND_22;
  reg [2:0] _EVAL_410;
  reg [31:0] _RAND_23;
  reg  _EVAL_421;
  reg [31:0] _RAND_24;
  reg  _EVAL_427;
  reg [31:0] _RAND_25;
  reg [2:0] _EVAL_444;
  reg [31:0] _RAND_26;
  reg  _EVAL_448;
  reg [31:0] _RAND_27;
  reg  _EVAL_449;
  reg [31:0] _RAND_28;
  reg  _EVAL_462;
  reg [31:0] _RAND_29;
  reg  _EVAL_480;
  reg [31:0] _RAND_30;
  reg [2:0] _EVAL_481;
  reg [31:0] _RAND_31;
  reg [2:0] _EVAL_485;
  reg [31:0] _RAND_32;
  reg  _EVAL_492;
  reg [31:0] _RAND_33;
  reg  _EVAL_497;
  reg [31:0] _RAND_34;
  reg [2:0] _EVAL_512;
  reg [31:0] _RAND_35;
  reg  _EVAL_519;
  reg [31:0] _RAND_36;
  reg [2:0] _EVAL_548;
  reg [31:0] _RAND_37;
  reg  _EVAL_552;
  reg [31:0] _RAND_38;
  reg  _EVAL_569;
  reg [31:0] _RAND_39;
  reg  _EVAL_581;
  reg [31:0] _RAND_40;
  reg  _EVAL_614;
  reg [31:0] _RAND_41;
  reg [2:0] _EVAL_648;
  reg [31:0] _RAND_42;
  reg [2:0] _EVAL_663;
  reg [31:0] _RAND_43;
  reg  _EVAL_673;
  reg [31:0] _RAND_44;
  reg [2:0] _EVAL_675;
  reg [31:0] _RAND_45;
  reg  _EVAL_690;
  reg [31:0] _RAND_46;
  reg  _EVAL_715;
  reg [31:0] _RAND_47;
  reg  _EVAL_730;
  reg [31:0] _RAND_48;
  reg [2:0] _EVAL_739;
  reg [31:0] _RAND_49;
  reg  _EVAL_741;
  reg [31:0] _RAND_50;
  reg [2:0] _EVAL_750;
  reg [31:0] _RAND_51;
  reg [2:0] _EVAL_757;
  reg [31:0] _RAND_52;
  reg [2:0] _EVAL_762;
  reg [31:0] _RAND_53;
  reg [2:0] _EVAL_765;
  reg [31:0] _RAND_54;
  reg [2:0] _EVAL_768;
  reg [31:0] _RAND_55;
  reg  _EVAL_770;
  reg [31:0] _RAND_56;
  reg [2:0] _EVAL_835;
  reg [31:0] _RAND_57;
  reg  _EVAL_880;
  reg [31:0] _RAND_58;
  reg [2:0] _EVAL_902;
  reg [31:0] _RAND_59;
  reg  _EVAL_912;
  reg [31:0] _RAND_60;
  reg  _EVAL_947;
  reg [31:0] _RAND_61;
  reg  _EVAL_989;
  reg [31:0] _RAND_62;
  reg [2:0] _EVAL_1035;
  reg [31:0] _RAND_63;
  reg  _EVAL_1073;
  reg [31:0] _RAND_64;
  reg [2:0] _EVAL_1088;
  reg [31:0] _RAND_65;
  reg  _EVAL_1121;
  reg [31:0] _RAND_66;
  reg [2:0] _EVAL_1122;
  reg [31:0] _RAND_67;
  reg [2:0] _EVAL_1127;
  reg [31:0] _RAND_68;
  reg [2:0] _EVAL_1142;
  reg [31:0] _RAND_69;
  reg [2:0] _EVAL_1151;
  reg [31:0] _RAND_70;
  reg [2:0] _EVAL_1156;
  reg [31:0] _RAND_71;
  reg [7:0] _EVAL_1162;
  reg [31:0] _RAND_72;
  reg [2:0] _EVAL_1168;
  reg [31:0] _RAND_73;
  reg [2:0] _EVAL_1176;
  reg [31:0] _RAND_74;
  reg  _EVAL_1206;
  reg [31:0] _RAND_75;
  reg [2:0] _EVAL_1212;
  reg [31:0] _RAND_76;
  reg [2:0] _EVAL_1239;
  reg [31:0] _RAND_77;
  reg [2:0] _EVAL_1253;
  reg [31:0] _RAND_78;
  reg  _EVAL_1261;
  reg [31:0] _RAND_79;
  reg [2:0] _EVAL_1266;
  reg [31:0] _RAND_80;
  reg  _EVAL_1267;
  reg [31:0] _RAND_81;
  reg  _EVAL_1270;
  reg [31:0] _RAND_82;
  reg [2:0] _EVAL_1280;
  reg [31:0] _RAND_83;
  reg  _EVAL_1313;
  reg [31:0] _RAND_84;
  reg  _EVAL_1315;
  reg [31:0] _RAND_85;
  reg [2:0] _EVAL_1351;
  reg [31:0] _RAND_86;
  reg [2:0] _EVAL_1365;
  reg [31:0] _RAND_87;
  reg [2:0] _EVAL_1390;
  reg [31:0] _RAND_88;
  reg [2:0] _EVAL_1433;
  reg [31:0] _RAND_89;
  reg [2:0] _EVAL_1438;
  reg [31:0] _RAND_90;
  reg [2:0] _EVAL_1444;
  reg [31:0] _RAND_91;
  reg  _EVAL_1456;
  reg [31:0] _RAND_92;
  reg  _EVAL_1471;
  reg [31:0] _RAND_93;
  reg  _EVAL_1496;
  reg [31:0] _RAND_94;
  reg  _EVAL_1521;
  reg [31:0] _RAND_95;
  reg [2:0] _EVAL_1526;
  reg [31:0] _RAND_96;
  reg  _EVAL_1536;
  reg [31:0] _RAND_97;
  reg  _EVAL_1556;
  reg [31:0] _RAND_98;
  reg [2:0] _EVAL_1562;
  reg [31:0] _RAND_99;
  reg  _EVAL_1580;
  reg [31:0] _RAND_100;
  reg  _EVAL_1587;
  reg [31:0] _RAND_101;
  reg  _EVAL_1597;
  reg [31:0] _RAND_102;
  reg  _EVAL_1599;
  reg [31:0] _RAND_103;
  reg [7:0] _EVAL_1639;
  reg [31:0] _RAND_104;
  reg [2:0] _EVAL_1660;
  reg [31:0] _RAND_105;
  reg [2:0] _EVAL_1680;
  reg [31:0] _RAND_106;
  reg [7:0] _EVAL_1697;
  reg [31:0] _RAND_107;
  reg [6:0] _EVAL_1698;
  reg [31:0] _RAND_108;
  reg  _EVAL_1708;
  reg [31:0] _RAND_109;
  reg  _EVAL_1709;
  reg [31:0] _RAND_110;
  reg [2:0] _EVAL_1738;
  reg [31:0] _RAND_111;
  reg  _EVAL_1753;
  reg [31:0] _RAND_112;
  reg [7:0] _EVAL_1776;
  reg [31:0] _RAND_113;
  reg [2:0] _EVAL_1783;
  reg [31:0] _RAND_114;
  reg [2:0] _EVAL_1786;
  reg [31:0] _RAND_115;
  reg  _EVAL_1788;
  reg [31:0] _RAND_116;
  reg [2:0] _EVAL_1801;
  reg [31:0] _RAND_117;
  reg [2:0] _EVAL_1819;
  reg [31:0] _RAND_118;
  reg [2:0] _EVAL_1870;
  reg [31:0] _RAND_119;
  reg  _EVAL_1917;
  reg [31:0] _RAND_120;
  reg  _EVAL_1929;
  reg [31:0] _RAND_121;
  reg  _EVAL_1930;
  reg [31:0] _RAND_122;
  reg  _EVAL_1938;
  reg [31:0] _RAND_123;
  reg [2:0] _EVAL_1962;
  reg [31:0] _RAND_124;
  reg  _EVAL_1979;
  reg [31:0] _RAND_125;
  reg [2:0] _EVAL_1980;
  reg [31:0] _RAND_126;
  reg [7:0] _EVAL_2018;
  reg [31:0] _RAND_127;
  reg [2:0] _EVAL_2035;
  reg [31:0] _RAND_128;
  reg  _EVAL_2050;
  reg [31:0] _RAND_129;
  reg [2:0] _EVAL_2055;
  reg [31:0] _RAND_130;
  reg [7:0] _EVAL_2073;
  reg [31:0] _RAND_131;
  reg [2:0] _EVAL_2110;
  reg [31:0] _RAND_132;
  reg [2:0] _EVAL_2111;
  reg [31:0] _RAND_133;
  reg [2:0] _EVAL_2121;
  reg [31:0] _RAND_134;
  reg  _EVAL_2128;
  reg [31:0] _RAND_135;
  reg  _EVAL_2133;
  reg [31:0] _RAND_136;
  reg  _EVAL_2155;
  reg [31:0] _RAND_137;
  reg  _EVAL_2159;
  reg [31:0] _RAND_138;
  reg [7:0] _EVAL_2188;
  reg [31:0] _RAND_139;
  reg  _EVAL_2202;
  reg [31:0] _RAND_140;
  reg  _EVAL_2209;
  reg [31:0] _RAND_141;
  reg  _EVAL_2214;
  reg [31:0] _RAND_142;
  reg [2:0] _EVAL_2231;
  reg [31:0] _RAND_143;
  reg  _EVAL_2254;
  reg [31:0] _RAND_144;
  reg [2:0] _EVAL_2256;
  reg [31:0] _RAND_145;
  reg [2:0] _EVAL_2290;
  reg [31:0] _RAND_146;
  reg [2:0] _EVAL_2306;
  reg [31:0] _RAND_147;
  reg [2:0] _EVAL_2311;
  reg [31:0] _RAND_148;
  reg [2:0] _EVAL_2334;
  reg [31:0] _RAND_149;
  reg [2:0] _EVAL_2336;
  reg [31:0] _RAND_150;
  reg  _EVAL_2341;
  reg [31:0] _RAND_151;
  reg [2:0] _EVAL_2356;
  reg [31:0] _RAND_152;
  reg [2:0] _EVAL_2481;
  reg [31:0] _RAND_153;
  reg [2:0] _EVAL_2484;
  reg [31:0] _RAND_154;
  reg  _EVAL_2485;
  reg [31:0] _RAND_155;
  reg [2:0] _EVAL_2491;
  reg [31:0] _RAND_156;
  reg [2:0] _EVAL_2500;
  reg [31:0] _RAND_157;
  reg  _EVAL_2507;
  reg [31:0] _RAND_158;
  reg [2:0] _EVAL_2536;
  reg [31:0] _RAND_159;
  reg  _EVAL_2582;
  reg [31:0] _RAND_160;
  reg [2:0] _EVAL_2584;
  reg [31:0] _RAND_161;
  reg [2:0] _EVAL_2646;
  reg [31:0] _RAND_162;
  reg  _EVAL_2648;
  reg [31:0] _RAND_163;
  reg [2:0] _EVAL_2653;
  reg [31:0] _RAND_164;
  reg  _EVAL_2666;
  reg [31:0] _RAND_165;
  reg [2:0] _EVAL_2677;
  reg [31:0] _RAND_166;
  reg  _EVAL_2684;
  reg [31:0] _RAND_167;
  reg  _EVAL_2688;
  reg [31:0] _RAND_168;
  reg  _EVAL_2701;
  reg [31:0] _RAND_169;
  reg [2:0] _EVAL_2720;
  reg [31:0] _RAND_170;
  reg [7:0] _EVAL_2754;
  reg [31:0] _RAND_171;
  reg [2:0] _EVAL_2760;
  reg [31:0] _RAND_172;
  reg  _EVAL_2803;
  reg [31:0] _RAND_173;
  reg  _EVAL_2807;
  reg [31:0] _RAND_174;
  reg  _EVAL_2809;
  reg [31:0] _RAND_175;
  reg [2:0] _EVAL_2810;
  reg [31:0] _RAND_176;
  reg  _EVAL_2826;
  reg [31:0] _RAND_177;
  reg  _EVAL_2838;
  reg [31:0] _RAND_178;
  reg  _EVAL_2850;
  reg [31:0] _RAND_179;
  reg [2:0] _EVAL_2851;
  reg [31:0] _RAND_180;
  reg  _EVAL_2870;
  reg [31:0] _RAND_181;
  reg [2:0] _EVAL_2881;
  reg [31:0] _RAND_182;
  reg [2:0] _EVAL_2937;
  reg [31:0] _RAND_183;
  reg  _EVAL_2938;
  reg [31:0] _RAND_184;
  reg  _EVAL_2942;
  reg [31:0] _RAND_185;
  reg  _EVAL_2953;
  reg [31:0] _RAND_186;
  reg [2:0] _EVAL_2958;
  reg [31:0] _RAND_187;
  reg [2:0] _EVAL_2965;
  reg [31:0] _RAND_188;
  reg  _EVAL_2972;
  reg [31:0] _RAND_189;
  reg [2:0] _EVAL_3008;
  reg [31:0] _RAND_190;
  reg [2:0] _EVAL_3014;
  reg [31:0] _RAND_191;
  reg  _EVAL_3023;
  reg [31:0] _RAND_192;
  reg  _EVAL_3025;
  reg [31:0] _RAND_193;
  reg  _EVAL_3039;
  reg [31:0] _RAND_194;
  reg [2:0] _EVAL_3056;
  reg [31:0] _RAND_195;
  reg [2:0] _EVAL_3102;
  reg [31:0] _RAND_196;
  reg [2:0] _EVAL_3113;
  reg [31:0] _RAND_197;
  reg [2:0] _EVAL_3118;
  reg [31:0] _RAND_198;
  reg  _EVAL_3137;
  reg [31:0] _RAND_199;
  reg  _EVAL_3167;
  reg [31:0] _RAND_200;
  reg  _EVAL_3192;
  reg [31:0] _RAND_201;
  reg [2:0] _EVAL_3195;
  reg [31:0] _RAND_202;
  reg  _EVAL_3199;
  reg [31:0] _RAND_203;
  reg [2:0] _EVAL_3204;
  reg [31:0] _RAND_204;
  reg [2:0] _EVAL_3216;
  reg [31:0] _RAND_205;
  reg  _EVAL_3222;
  reg [31:0] _RAND_206;
  reg [6:0] _EVAL_3235;
  reg [31:0] _RAND_207;
  reg [2:0] _EVAL_3242;
  reg [31:0] _RAND_208;
  reg  _EVAL_3245;
  reg [31:0] _RAND_209;
  reg [2:0] _EVAL_3267;
  reg [31:0] _RAND_210;
  reg [2:0] _EVAL_3274;
  reg [31:0] _RAND_211;
  reg  _EVAL_3279;
  reg [31:0] _RAND_212;
  reg  _EVAL_3283;
  reg [31:0] _RAND_213;
  reg  _EVAL_3296;
  reg [31:0] _RAND_214;
  reg  _EVAL_3299;
  reg [31:0] _RAND_215;
  reg [2:0] _EVAL_3312;
  reg [31:0] _RAND_216;
  reg [2:0] _EVAL_3315;
  reg [31:0] _RAND_217;
  reg  _EVAL_3317;
  reg [31:0] _RAND_218;
  reg [2:0] _EVAL_3331;
  reg [31:0] _RAND_219;
  reg [2:0] _EVAL_3336;
  reg [31:0] _RAND_220;
  reg  _EVAL_3359;
  reg [31:0] _RAND_221;
  reg  _EVAL_3361;
  reg [31:0] _RAND_222;
  reg [2:0] _EVAL_3383;
  reg [31:0] _RAND_223;
  reg  _EVAL_3407;
  reg [31:0] _RAND_224;
  reg  _EVAL_3419;
  reg [31:0] _RAND_225;
  reg [7:0] _EVAL_3421;
  reg [31:0] _RAND_226;
  reg [7:0] _EVAL_3488;
  reg [31:0] _RAND_227;
  reg  _EVAL_3505;
  reg [31:0] _RAND_228;
  reg  _EVAL_3527;
  reg [31:0] _RAND_229;
  reg  _EVAL_3551;
  reg [31:0] _RAND_230;
  reg [2:0] _EVAL_3552;
  reg [31:0] _RAND_231;
  reg [2:0] _EVAL_3554;
  reg [31:0] _RAND_232;
  reg [2:0] _EVAL_3563;
  reg [31:0] _RAND_233;
  reg [2:0] _EVAL_3571;
  reg [31:0] _RAND_234;
  reg [2:0] _EVAL_3573;
  reg [31:0] _RAND_235;
  reg [2:0] _EVAL_3591;
  reg [31:0] _RAND_236;
  reg [2:0] _EVAL_3608;
  reg [31:0] _RAND_237;
  reg [7:0] _EVAL_3623;
  reg [31:0] _RAND_238;
  reg  _EVAL_3636;
  reg [31:0] _RAND_239;
  reg [2:0] _EVAL_3644;
  reg [31:0] _RAND_240;
  reg [2:0] _EVAL_3645;
  reg [31:0] _RAND_241;
  reg  _EVAL_3713;
  reg [31:0] _RAND_242;
  reg  _EVAL_3715;
  reg [31:0] _RAND_243;
  reg  _EVAL_3720;
  reg [31:0] _RAND_244;
  reg [2:0] _EVAL_3721;
  reg [31:0] _RAND_245;
  reg  _EVAL_3728;
  reg [31:0] _RAND_246;
  reg [2:0] _EVAL_3731;
  reg [31:0] _RAND_247;
  reg [2:0] _EVAL_3733;
  reg [31:0] _RAND_248;
  reg [2:0] _EVAL_3740;
  reg [31:0] _RAND_249;
  reg [7:0] _EVAL_3743;
  reg [31:0] _RAND_250;
  reg  _EVAL_3750;
  reg [31:0] _RAND_251;
  reg  _EVAL_3757;
  reg [31:0] _RAND_252;
  reg  _EVAL_3759;
  reg [31:0] _RAND_253;
  reg [2:0] _EVAL_3768;
  reg [31:0] _RAND_254;
  reg  _EVAL_3783;
  reg [31:0] _RAND_255;
  reg  _EVAL_3788;
  reg [31:0] _RAND_256;
  reg [2:0] _EVAL_3801;
  reg [31:0] _RAND_257;
  reg [2:0] _EVAL_3804;
  reg [31:0] _RAND_258;
  reg [2:0] _EVAL_3843;
  reg [31:0] _RAND_259;
  reg  _EVAL_3850;
  reg [31:0] _RAND_260;
  reg [7:0] _EVAL_3870;
  reg [31:0] _RAND_261;
  reg  _EVAL_3899;
  reg [31:0] _RAND_262;
  reg [2:0] _EVAL_3909;
  reg [31:0] _RAND_263;
  reg [7:0] _EVAL_3913;
  reg [31:0] _RAND_264;
  reg [2:0] _EVAL_3943;
  reg [31:0] _RAND_265;
  reg  _EVAL_3964;
  reg [31:0] _RAND_266;
  reg  _EVAL_3996;
  reg [31:0] _RAND_267;
  reg [2:0] _EVAL_4013;
  reg [31:0] _RAND_268;
  reg  _EVAL_4034;
  reg [31:0] _RAND_269;
  reg [2:0] _EVAL_4050;
  reg [31:0] _RAND_270;
  reg  _EVAL_4063;
  reg [31:0] _RAND_271;
  reg [2:0] _EVAL_4066;
  reg [31:0] _RAND_272;
  wire [25:0] _EVAL_910;
  wire  _EVAL_2134;
  wire  _EVAL_1716;
  wire  _EVAL_3673;
  wire  _EVAL_1141;
  wire  _EVAL_2526;
  wire  _EVAL_2033;
  wire  _EVAL_2718;
  wire  _EVAL_2486;
  wire  _EVAL_640;
  wire  _EVAL_3992;
  wire  _EVAL_397;
  wire  _EVAL_2460;
  wire  _EVAL_3606;
  wire [9:0] _EVAL_1450;
  wire [1023:0] _EVAL_2999;
  wire  _EVAL_2866;
  wire  _EVAL_3344;
  wire [23:0] _EVAL_3888;
  wire  _EVAL_2267;
  wire  _EVAL_1644;
  wire  _EVAL_915;
  wire [7:0] _EVAL_287;
  wire  _EVAL_2436;
  wire [7:0] _EVAL_3655;
  wire  _EVAL_4053;
  wire [7:0] _EVAL_2619;
  wire  _EVAL_1637;
  wire [7:0] _EVAL_352;
  wire [31:0] _EVAL_2124;
  wire [2:0] _EVAL_3165;
  wire  _EVAL_591;
  wire  _EVAL_532;
  wire  _EVAL_886;
  wire  _EVAL_3851;
  wire  _EVAL_3050;
  wire  _EVAL_1440;
  wire  _EVAL_3081;
  wire  _EVAL_4052;
  wire  _EVAL_2575;
  wire  _EVAL_964;
  wire  _EVAL_2656;
  wire  _EVAL_3526;
  wire  _EVAL_3146;
  wire  _EVAL_1023;
  wire  _EVAL_3602;
  wire  _EVAL_2966;
  wire  _EVAL_742;
  wire  _EVAL_1018;
  wire  _EVAL_3758;
  wire  _EVAL_368;
  wire  _EVAL_1362;
  wire  _EVAL_870;
  wire  _EVAL_2716;
  wire  _EVAL_3097;
  wire  _EVAL_841;
  wire  _EVAL_3044;
  wire  _EVAL_3226;
  wire  _EVAL_584;
  wire  _EVAL_3400;
  wire  _EVAL_1014;
  wire  _EVAL_1838;
  wire  _EVAL_1891;
  wire  _EVAL_907;
  wire  _EVAL_1425;
  wire  _EVAL_1185;
  wire  _EVAL_1489;
  wire  _EVAL_2265;
  wire  _EVAL_3179;
  wire  _EVAL_2269;
  wire  _EVAL_922;
  wire  _EVAL_1991;
  wire  _EVAL_2441;
  wire  _EVAL_3002;
  wire  _EVAL_350;
  wire  _EVAL_3718;
  wire  _EVAL_443;
  wire  _EVAL_2448;
  wire  _EVAL_2777;
  wire  _EVAL_2361;
  wire  _EVAL_373;
  wire  _EVAL_3550;
  wire  _EVAL_2496;
  wire  _EVAL_2308;
  wire  _EVAL_1421;
  wire  _EVAL_3500;
  wire  _EVAL_1163;
  wire  _EVAL_700;
  wire  _EVAL_1301;
  wire  _EVAL_4011;
  wire  _EVAL_942;
  wire  _EVAL_3177;
  wire  _EVAL_1859;
  wire  _EVAL_1672;
  wire  _EVAL_2434;
  wire  _EVAL_2841;
  wire  _EVAL_3802;
  wire  _EVAL_3883;
  wire  _EVAL_1080;
  wire  _EVAL_2192;
  wire  _EVAL_2510;
  wire  _EVAL_2970;
  wire  _EVAL_165;
  wire  _EVAL_2863;
  wire  _EVAL_3127;
  wire  _EVAL_3494;
  wire  _EVAL_3590;
  wire  _EVAL_1282;
  wire  _EVAL_3839;
  wire  _EVAL_2801;
  wire  _EVAL_2771;
  wire  _EVAL_711;
  wire  _EVAL_1939;
  wire  _EVAL_159;
  wire  _EVAL_1321;
  wire  _EVAL_1987;
  wire  _EVAL_1387;
  wire  _EVAL_3800;
  wire  _EVAL_1198;
  wire  _EVAL_1713;
  wire  _EVAL_1366;
  wire  _EVAL_2153;
  wire  _EVAL_2347;
  wire  _EVAL_3428;
  wire  _EVAL_562;
  wire  _EVAL_529;
  wire  _EVAL_3072;
  wire  _EVAL_1583;
  wire  _EVAL_854;
  wire  _EVAL_3382;
  wire  _EVAL_249;
  wire  _EVAL_775;
  wire  _EVAL_1108;
  wire  _EVAL_1059;
  wire  _EVAL_1779;
  wire  _EVAL_3523;
  wire  _EVAL_2314;
  wire  _EVAL_988;
  wire  _EVAL_1167;
  wire  _EVAL_2633;
  wire  _EVAL_277;
  wire  _EVAL_652;
  wire  _EVAL_2989;
  wire  _EVAL_878;
  wire  _EVAL_888;
  wire  _EVAL_4025;
  wire  _EVAL_2868;
  wire  _EVAL_3605;
  wire  _EVAL_1594;
  wire  _EVAL_459;
  wire  _EVAL_1170;
  wire  _EVAL_1189;
  wire  _EVAL_1565;
  wire  _EVAL_3941;
  wire  _EVAL_3866;
  wire  _EVAL_1810;
  wire  _EVAL_3232;
  wire  _EVAL_1318;
  wire  _EVAL_4015;
  wire  _EVAL_1849;
  wire  _EVAL_3174;
  wire  _EVAL_945;
  wire  _EVAL_559;
  wire  _EVAL_148;
  wire  _EVAL_1736;
  wire  _EVAL_1173;
  wire  _EVAL_684;
  wire  _EVAL_2318;
  wire  _EVAL_2220;
  wire  _EVAL_491;
  wire  _EVAL_3412;
  wire  _EVAL_1292;
  wire  _EVAL_1483;
  wire  _EVAL_3556;
  wire  _EVAL_1574;
  wire  _EVAL_3828;
  wire  _EVAL_517;
  wire  _EVAL_583;
  wire  _EVAL_3125;
  wire  _EVAL_3995;
  wire  _EVAL_2670;
  wire  _EVAL_3247;
  wire  _EVAL_2299;
  wire  _EVAL_3811;
  wire  _EVAL_1231;
  wire  _EVAL_3722;
  wire  _EVAL_3109;
  wire  _EVAL_2435;
  wire  _EVAL_4021;
  wire  _EVAL_2781;
  wire  _EVAL_2088;
  wire  _EVAL_2440;
  wire  _EVAL_1418;
  wire  _EVAL_2832;
  wire  _EVAL_3042;
  wire  _EVAL_537;
  wire  _EVAL_898;
  wire  _EVAL_1727;
  wire  _EVAL_1734;
  wire  _EVAL_3172;
  wire  _EVAL_460;
  wire  _EVAL_1407;
  wire  _EVAL_3147;
  wire  _EVAL_2451;
  wire  _EVAL_3841;
  wire  _EVAL_2847;
  wire  _EVAL_1777;
  wire  _EVAL_2790;
  wire  _EVAL_2234;
  wire  _EVAL_1676;
  wire  _EVAL_626;
  wire  _EVAL_3059;
  wire  _EVAL_2184;
  wire  _EVAL_429;
  wire  _EVAL_390;
  wire  _EVAL_2158;
  wire  _EVAL_826;
  wire  _EVAL_2107;
  wire  _EVAL_1847;
  wire [6:0] _EVAL_2616;
  wire [127:0] _EVAL_1635;
  wire  _EVAL_1805;
  wire  _EVAL_1077;
  wire  _EVAL_1531;
  wire  _EVAL_1886;
  wire  _EVAL_378;
  wire  _EVAL_4026;
  wire  _EVAL_3215;
  wire  _EVAL_2232;
  wire  _EVAL_632;
  wire  _EVAL_3688;
  wire  _EVAL_2917;
  wire [9:0] _EVAL_3878;
  wire [18:0] _EVAL_3760;
  wire [27:0] _EVAL_618;
  wire [31:0] _EVAL_2860;
  wire [9:0] _EVAL_716;
  wire [18:0] _EVAL_2797;
  wire [27:0] _EVAL_2226;
  wire [31:0] _EVAL_1293;
  wire [9:0] _EVAL_1590;
  wire [18:0] _EVAL_3587;
  wire [27:0] _EVAL_267;
  wire [31:0] _EVAL_521;
  wire [9:0] _EVAL_760;
  wire [18:0] _EVAL_1227;
  wire [27:0] _EVAL_1511;
  wire [31:0] _EVAL_1721;
  wire [31:0] _EVAL_2362;
  wire [31:0] _EVAL_3259;
  wire [31:0] _EVAL_3026;
  wire [31:0] _EVAL_4029;
  wire [3:0] _EVAL_1970;
  wire [31:0] _EVAL_1286;
  wire [31:0] _EVAL_1710;
  wire [31:0] _EVAL_197;
  wire [31:0] _EVAL_837;
  wire [31:0] _EVAL_2355;
  wire [31:0] _EVAL_2915;
  wire [31:0] _EVAL_3944;
  wire [31:0] _EVAL_334;
  wire [31:0] _EVAL_3837;
  wire [31:0] _EVAL_2623;
  wire [31:0] _EVAL_1750;
  wire [31:0] _EVAL_2612;
  wire [31:0] _EVAL_1305;
  wire [31:0] _EVAL_923;
  wire [31:0] _EVAL_2975;
  wire [31:0] _EVAL_1114;
  wire [31:0] _EVAL_2025;
  wire [31:0] _EVAL_423;
  wire [31:0] _EVAL_1943;
  wire [31:0] _EVAL_2968;
  wire [31:0] _EVAL_2113;
  wire [31:0] _EVAL_1430;
  wire [31:0] _EVAL_3957;
  wire [31:0] _EVAL_2094;
  wire [31:0] _EVAL_1380;
  wire [31:0] _EVAL_1608;
  wire [31:0] _EVAL_2749;
  wire [31:0] _EVAL_2190;
  wire [31:0] _EVAL_1804;
  wire [31:0] _EVAL_3219;
  wire [31:0] _EVAL_325;
  wire [31:0] _EVAL_2281;
  wire [31:0] _EVAL_811;
  wire [31:0] _EVAL_3627;
  wire [31:0] _EVAL_1273;
  wire [31:0] _EVAL_3301;
  wire [31:0] _EVAL_2502;
  wire [31:0] _EVAL_3017;
  wire [31:0] _EVAL_1625;
  wire [31:0] _EVAL_1722;
  wire [31:0] _EVAL_3466;
  wire [31:0] _EVAL_276;
  wire [31:0] _EVAL_2561;
  wire [31:0] _EVAL_2882;
  wire [31:0] _EVAL_389;
  wire [31:0] _EVAL_3540;
  wire [31:0] _EVAL_2090;
  wire [31:0] _EVAL_2065;
  wire [31:0] _EVAL_2982;
  wire [31:0] _EVAL_1402;
  wire [31:0] _EVAL_1339;
  wire [31:0] _EVAL_2531;
  wire [31:0] _EVAL_1752;
  wire [31:0] _EVAL_3815;
  wire [31:0] _EVAL_2853;
  wire [31:0] _EVAL_2100;
  wire [31:0] _EVAL_2081;
  wire [31:0] _EVAL_1774;
  wire [31:0] _EVAL_1795;
  wire [31:0] _EVAL_3798;
  wire [31:0] _EVAL_940;
  wire [31:0] _EVAL_1137;
  wire [31:0] _EVAL_709;
  wire [31:0] _EVAL_2802;
  wire [31:0] _EVAL_2141;
  wire [31:0] _EVAL_409;
  wire [31:0] _EVAL_794;
  wire [31:0] _EVAL_891;
  wire [31:0] _EVAL_3950;
  wire [31:0] _EVAL_3928;
  wire [31:0] _EVAL_1186;
  wire [31:0] _EVAL_2119;
  wire [31:0] _EVAL_218;
  wire [31:0] _EVAL_1934;
  wire [31:0] _EVAL_1466;
  wire [31:0] _EVAL_3867;
  wire [31:0] _EVAL_2389;
  wire [31:0] _EVAL_836;
  wire [31:0] _EVAL_2092;
  wire [31:0] _EVAL_1448;
  wire [31:0] _EVAL_2026;
  wire [31:0] _EVAL_2912;
  wire [31:0] _EVAL_3030;
  wire [31:0] _EVAL_2766;
  wire [31:0] _EVAL_1578;
  wire  _EVAL_585;
  wire  _EVAL_3586;
  wire  _EVAL_1487;
  wire  _EVAL_1626;
  wire  _EVAL_2628;
  wire  _EVAL_294;
  wire  _EVAL_2578;
  wire  _EVAL_2956;
  wire  _EVAL_2610;
  wire  _EVAL_3418;
  wire  _EVAL_1667;
  wire  _EVAL_1973;
  wire  _EVAL_3593;
  wire  _EVAL_1820;
  wire  _EVAL_725;
  wire  _EVAL_364;
  wire  _EVAL_3152;
  wire  _EVAL_3617;
  wire  _EVAL_2140;
  wire  _EVAL_2252;
  wire  _EVAL_3504;
  wire  _EVAL_318;
  wire  _EVAL_3181;
  wire  _EVAL_3936;
  wire  _EVAL_2130;
  wire  _EVAL_822;
  wire  _EVAL_1515;
  wire  _EVAL_617;
  wire  _EVAL_2514;
  wire  _EVAL_2543;
  wire  _EVAL_943;
  wire  _EVAL_1852;
  wire  _EVAL_2057;
  wire  _EVAL_3820;
  wire  _EVAL_3860;
  wire  _EVAL_1765;
  wire  _EVAL_2122;
  wire  _EVAL_339;
  wire  _EVAL_1416;
  wire  _EVAL_3323;
  wire  _EVAL_881;
  wire  _EVAL_4039;
  wire  _EVAL_2535;
  wire  _EVAL_262;
  wire  _EVAL_1055;
  wire  _EVAL_2625;
  wire  _EVAL_3159;
  wire  _EVAL_3233;
  wire  _EVAL_1572;
  wire  _EVAL_3358;
  wire  _EVAL_237;
  wire  _EVAL_472;
  wire  _EVAL_2003;
  wire  _EVAL_2007;
  wire  _EVAL_3300;
  wire  _EVAL_178;
  wire  _EVAL_2066;
  wire  _EVAL_1399;
  wire  _EVAL_1601;
  wire  _EVAL_2432;
  wire  _EVAL_3729;
  wire  _EVAL_1132;
  wire  _EVAL_2659;
  wire  _EVAL_555;
  wire  _EVAL_808;
  wire  _EVAL_1965;
  wire  _EVAL_2410;
  wire  _EVAL_2763;
  wire  _EVAL_2102;
  wire  _EVAL_3776;
  wire  _EVAL_3401;
  wire  _EVAL_2796;
  wire  _EVAL_840;
  wire  _EVAL_1097;
  wire  _EVAL_1945;
  wire  _EVAL_2932;
  wire  _EVAL_2060;
  wire  _EVAL_1946;
  wire  _EVAL_1952;
  wire  _EVAL_2000;
  wire  _EVAL_3994;
  wire  _EVAL_1669;
  wire  _EVAL_1931;
  wire  _EVAL_511;
  wire [31:0] _EVAL_1875;
  wire [31:0] _EVAL_3564;
  wire [31:0] _EVAL_3258;
  wire [31:0] _EVAL_516;
  wire [31:0] _EVAL_2147;
  wire [31:0] _EVAL_928;
  wire [31:0] _EVAL_254;
  wire [31:0] _EVAL_1130;
  wire [31:0] _EVAL_2063;
  wire [31:0] _EVAL_3911;
  wire [31:0] _EVAL_2867;
  wire [31:0] _EVAL_3898;
  wire [31:0] _EVAL_4038;
  wire [31:0] _EVAL_3158;
  wire [31:0] _EVAL_1052;
  wire [31:0] _EVAL_1329;
  wire [31:0] _EVAL_3364;
  wire [31:0] _EVAL_1959;
  wire [31:0] _EVAL_2228;
  wire [31:0] _EVAL_1051;
  wire [31:0] _EVAL_3646;
  wire [31:0] _EVAL_1061;
  wire [31:0] _EVAL_3060;
  wire [31:0] _EVAL_1866;
  wire [31:0] _EVAL_3831;
  wire [31:0] _EVAL_703;
  wire [31:0] _EVAL_225;
  wire [31:0] _EVAL_1985;
  wire [31:0] _EVAL_2877;
  wire [31:0] _EVAL_1468;
  wire [31:0] _EVAL_1741;
  wire [31:0] _EVAL_2459;
  wire [31:0] _EVAL_1393;
  wire [31:0] _EVAL_1323;
  wire [31:0] _EVAL_149;
  wire [31:0] _EVAL_1343;
  wire [31:0] _EVAL_2513;
  wire [31:0] _EVAL_2148;
  wire [31:0] _EVAL_329;
  wire [31:0] _EVAL_3385;
  wire [31:0] _EVAL_2640;
  wire [31:0] _EVAL_3772;
  wire [31:0] _EVAL_2095;
  wire [31:0] _EVAL_461;
  wire [31:0] _EVAL_542;
  wire [31:0] _EVAL_3614;
  wire [31:0] _EVAL_1654;
  wire [31:0] _EVAL_1376;
  wire [31:0] _EVAL_2728;
  wire  _EVAL_1907;
  wire  _EVAL_1328;
  wire [6:0] _EVAL_1332;
  wire  _EVAL_3082;
  wire  _EVAL_1811;
  wire  _EVAL_1352;
  wire  _EVAL_3907;
  wire  _EVAL_2056;
  wire  _EVAL_1458;
  wire  _EVAL_1717;
  wire  _EVAL_348;
  wire  _EVAL_2104;
  wire  _EVAL_3231;
  wire  _EVAL_3370;
  wire  _EVAL_722;
  wire  _EVAL_3881;
  wire  _EVAL_2310;
  wire  _EVAL_2848;
  wire  _EVAL_3671;
  wire  _EVAL_3595;
  wire  _EVAL_3534;
  wire  _EVAL_1236;
  wire  _EVAL_2861;
  wire  _EVAL_2524;
  wire  _EVAL_2001;
  wire  _EVAL_829;
  wire  _EVAL_1634;
  wire  _EVAL_2079;
  wire  _EVAL_416;
  wire  _EVAL_4001;
  wire [7:0] _EVAL_2288;
  wire  _EVAL_189;
  wire  _EVAL_1294;
  wire  _EVAL_3499;
  wire  _EVAL_195;
  wire  _EVAL_2940;
  wire  _EVAL_3094;
  wire  _EVAL_3584;
  wire  _EVAL_873;
  wire  _EVAL_3756;
  wire  _EVAL_3061;
  wire  _EVAL_1229;
  wire  _EVAL_2571;
  wire  _EVAL_2415;
  wire  _EVAL_1915;
  wire  _EVAL_1958;
  wire  _EVAL_1201;
  wire [7:0] _EVAL_638;
  wire  _EVAL_1856;
  wire  _EVAL_2208;
  wire  _EVAL_938;
  wire  _EVAL_1699;
  wire  _EVAL_464;
  wire  _EVAL_2869;
  wire  _EVAL_824;
  wire  _EVAL_3755;
  wire  _EVAL_2745;
  wire  _EVAL_2573;
  wire  _EVAL_1475;
  wire  _EVAL_1785;
  wire  _EVAL_1452;
  wire  _EVAL_1992;
  wire  _EVAL_846;
  wire  _EVAL_2835;
  wire  _EVAL_2856;
  wire  _EVAL_362;
  wire  _EVAL_533;
  wire  _EVAL_2660;
  wire  _EVAL_3424;
  wire  _EVAL_2118;
  wire  _EVAL_3348;
  wire  _EVAL_1790;
  wire  _EVAL_2464;
  wire  _EVAL_3379;
  wire  _EVAL_3134;
  wire  _EVAL_3665;
  wire  _EVAL_3439;
  wire  _EVAL_736;
  wire  _EVAL_2713;
  wire  _EVAL_1877;
  wire  _EVAL_2054;
  wire  _EVAL_3895;
  wire  _EVAL_3415;
  wire  _EVAL_660;
  wire  _EVAL_2052;
  wire  _EVAL_3404;
  wire  _EVAL_2006;
  wire  _EVAL_1355;
  wire [7:0] _EVAL_3372;
  wire  _EVAL_187;
  wire  _EVAL_2528;
  wire  _EVAL_4020;
  wire  _EVAL_2171;
  wire  _EVAL_3594;
  wire [7:0] _EVAL_695;
  wire  _EVAL_2335;
  wire  _EVAL_2865;
  wire  _EVAL_979;
  wire  _EVAL_3932;
  wire  _EVAL_3961;
  wire  _EVAL_1780;
  wire  _EVAL_2555;
  wire  _EVAL_3240;
  wire  _EVAL_2156;
  wire [7:0] _EVAL_3055;
  wire  _EVAL_3454;
  wire  _EVAL_2664;
  wire  _EVAL_3930;
  wire  _EVAL_2615;
  wire  _EVAL_3546;
  wire  _EVAL_2782;
  wire  _EVAL_704;
  wire  _EVAL_3292;
  wire  _EVAL_3256;
  wire  _EVAL_4054;
  wire  _EVAL_1944;
  wire  _EVAL_3325;
  wire  _EVAL_3816;
  wire  _EVAL_2204;
  wire  _EVAL_1839;
  wire  _EVAL_1533;
  wire  _EVAL_3520;
  wire  _EVAL_3918;
  wire  _EVAL_3908;
  wire  _EVAL_1462;
  wire  _EVAL_3390;
  wire  _EVAL_3705;
  wire  _EVAL_1887;
  wire  _EVAL_1107;
  wire  _EVAL_985;
  wire  _EVAL_2183;
  wire  _EVAL_3018;
  wire  _EVAL_1232;
  wire  _EVAL_2572;
  wire  _EVAL_2969;
  wire  _EVAL_3434;
  wire  _EVAL_622;
  wire  _EVAL_2333;
  wire  _EVAL_1021;
  wire  _EVAL_3817;
  wire  _EVAL_1486;
  wire  _EVAL_2907;
  wire  _EVAL_1196;
  wire  _EVAL_1265;
  wire  _EVAL_428;
  wire  _EVAL_828;
  wire  _EVAL_3156;
  wire  _EVAL_320;
  wire [7:0] _EVAL_1552;
  wire [7:0] _EVAL_2287;
  wire [15:0] _EVAL_1746;
  wire [31:0] _EVAL_3239;
  wire  _EVAL_226;
  wire  _EVAL_2746;
  wire  _EVAL_3078;
  wire  _EVAL_1009;
  wire  _EVAL_146;
  wire  _EVAL_2048;
  wire  _EVAL_1181;
  wire [7:0] _EVAL_2047;
  wire  _EVAL_845;
  wire  _EVAL_3884;
  wire  _EVAL_3318;
  wire  _EVAL_438;
  wire  _EVAL_1503;
  wire  _EVAL_263;
  wire  _EVAL_3641;
  wire  _EVAL_3508;
  wire  _EVAL_653;
  wire  _EVAL_207;
  wire  _EVAL_3423;
  wire  _EVAL_921;
  wire  _EVAL_1289;
  wire [13:0] _EVAL_291;
  wire  _EVAL_236;
  wire  _EVAL_1516;
  wire  _EVAL_3220;
  wire  _EVAL_1326;
  wire  _EVAL_271;
  wire  _EVAL_607;
  wire  _EVAL_1337;
  wire  _EVAL_1309;
  wire  _EVAL_1706;
  wire  _EVAL_1881;
  wire  _EVAL_3098;
  wire  _EVAL_1548;
  wire  _EVAL_2248;
  wire  _EVAL_2559;
  wire  _EVAL_2354;
  wire  _EVAL_2515;
  wire  _EVAL_3642;
  wire  _EVAL_3282;
  wire  _EVAL_1704;
  wire  _EVAL_2463;
  wire  _EVAL_245;
  wire  _EVAL_1549;
  wire  _EVAL_1914;
  wire  _EVAL_3679;
  wire  _EVAL_3959;
  wire  _EVAL_1853;
  wire  _EVAL_2346;
  wire  _EVAL_3074;
  wire  _EVAL_3234;
  wire  _EVAL_1731;
  wire  _EVAL_1164;
  wire  _EVAL_917;
  wire  _EVAL_1855;
  wire  _EVAL_455;
  wire  _EVAL_507;
  wire  _EVAL_1368;
  wire  _EVAL_466;
  wire  _EVAL_353;
  wire  _EVAL_2852;
  wire  _EVAL_2947;
  wire  _EVAL_3459;
  wire  _EVAL_248;
  wire  _EVAL_3628;
  wire  _EVAL_1876;
  wire  _EVAL_2553;
  wire  _EVAL_2845;
  wire  _EVAL_1613;
  wire  _EVAL_1259;
  wire  _EVAL_809;
  wire  _EVAL_2825;
  wire  _EVAL_4056;
  wire  _EVAL_303;
  wire  _EVAL_3443;
  wire  _EVAL_514;
  wire  _EVAL_3509;
  wire  _EVAL_2008;
  wire  _EVAL_3680;
  wire  _EVAL_851;
  wire  _EVAL_3690;
  wire  _EVAL_930;
  wire  _EVAL_3489;
  wire  _EVAL_3726;
  wire  _EVAL_1880;
  wire  _EVAL_2146;
  wire  _EVAL_2624;
  wire  _EVAL_401;
  wire  _EVAL_2279;
  wire  _EVAL_2574;
  wire  _EVAL_753;
  wire  _EVAL_2779;
  wire  _EVAL_1222;
  wire  _EVAL_2730;
  wire  _EVAL_1241;
  wire  _EVAL_3069;
  wire  _EVAL_3221;
  wire  _EVAL_1085;
  wire  _EVAL_795;
  wire  _EVAL_3919;
  wire  _EVAL_1525;
  wire  _EVAL_899;
  wire  _EVAL_926;
  wire  _EVAL_3043;
  wire  _EVAL_415;
  wire  _EVAL_323;
  wire  _EVAL_1956;
  wire  _EVAL_3803;
  wire  _EVAL_1843;
  wire  _EVAL_1890;
  wire  _EVAL_2391;
  wire  _EVAL_509;
  wire  _EVAL_2858;
  wire  _EVAL_3431;
  wire  _EVAL_1986;
  wire  _EVAL_4068;
  wire  _EVAL_2477;
  wire  _EVAL_1500;
  wire  _EVAL_2443;
  wire  _EVAL_3335;
  wire  _EVAL_2548;
  wire  _EVAL_3252;
  wire  _EVAL_3053;
  wire  _EVAL_265;
  wire  _EVAL_1397;
  wire  _EVAL_1537;
  wire  _EVAL_2902;
  wire  _EVAL_488;
  wire  _EVAL_3852;
  wire  _EVAL_3675;
  wire  _EVAL_1648;
  wire  _EVAL_2742;
  wire  _EVAL_540;
  wire  _EVAL_1264;
  wire  _EVAL_1283;
  wire  _EVAL_574;
  wire  _EVAL_2750;
  wire  _EVAL_1298;
  wire  _EVAL_2366;
  wire  _EVAL_2631;
  wire  _EVAL_1230;
  wire  _EVAL_2303;
  wire  _EVAL_1002;
  wire  _EVAL_565;
  wire  _EVAL_2595;
  wire  _EVAL_3122;
  wire  _EVAL_1215;
  wire  _EVAL_3088;
  wire  _EVAL_792;
  wire  _EVAL_2696;
  wire [62:0] _EVAL_3497;
  wire [127:0] _EVAL_1469;
  wire [31:0] _EVAL_1584;
  wire [6:0] _EVAL_666;
  wire [127:0] _EVAL_553;
  wire  _EVAL_3970;
  wire  _EVAL_1990;
  wire  _EVAL_3166;
  wire  _EVAL_2136;
  wire  _EVAL_2277;
  wire  _EVAL_515;
  wire  _EVAL_527;
  wire  _EVAL_2532;
  wire  _EVAL_3117;
  wire  _EVAL_3689;
  wire  _EVAL_1408;
  wire  _EVAL_436;
  wire  _EVAL_274;
  wire  _EVAL_1136;
  wire  _EVAL_377;
  wire  _EVAL_748;
  wire  _EVAL_1707;
  wire  _EVAL_939;
  wire  _EVAL_2125;
  wire  _EVAL_2959;
  wire  _EVAL_2157;
  wire  _EVAL_3037;
  wire  _EVAL_3744;
  wire  _EVAL_1793;
  wire  _EVAL_590;
  wire  _EVAL_1873;
  wire  _EVAL_1512;
  wire  _EVAL_4017;
  wire  _EVAL_973;
  wire  _EVAL_257;
  wire  _EVAL_800;
  wire  _EVAL_2251;
  wire  _EVAL_2446;
  wire  _EVAL_1177;
  wire  _EVAL_4044;
  wire  _EVAL_3096;
  wire  _EVAL_3864;
  wire  _EVAL_821;
  wire  _EVAL_727;
  wire  _EVAL_2317;
  wire  _EVAL_2106;
  wire  _EVAL_1888;
  wire  _EVAL_592;
  wire  _EVAL_1148;
  wire  _EVAL_1913;
  wire  _EVAL_229;
  wire  _EVAL_525;
  wire  _EVAL_3409;
  wire  _EVAL_3510;
  wire  _EVAL_2291;
  wire  _EVAL_375;
  wire  _EVAL_1432;
  wire  _EVAL_1257;
  wire  _EVAL_3476;
  wire  _EVAL_3136;
  wire  _EVAL_586;
  wire  _EVAL_3269;
  wire  _EVAL_3529;
  wire  _EVAL_4032;
  wire  _EVAL_4041;
  wire  _EVAL_4040;
  wire  _EVAL_2731;
  wire  _EVAL_2662;
  wire  _EVAL_4043;
  wire  _EVAL_3273;
  wire [6:0] _EVAL_3432;
  wire  _EVAL_1064;
  wire  _EVAL_3265;
  wire  _EVAL_3549;
  wire  _EVAL_2565;
  wire  _EVAL_1502;
  wire  _EVAL_3981;
  wire  _EVAL_3203;
  wire  _EVAL_220;
  wire  _EVAL_1414;
  wire  _EVAL_3873;
  wire  _EVAL_1922;
  wire  _EVAL_3882;
  wire  _EVAL_4062;
  wire  _EVAL_3847;
  wire  _EVAL_1764;
  wire  _EVAL_2480;
  wire  _EVAL_2697;
  wire  _EVAL_3707;
  wire  _EVAL_2233;
  wire  _EVAL_3588;
  wire  _EVAL_710;
  wire  _EVAL_2770;
  wire  _EVAL_847;
  wire  _EVAL_1202;
  wire  _EVAL_3429;
  wire  _EVAL_2567;
  wire  _EVAL_1069;
  wire  _EVAL_2189;
  wire  _EVAL_2388;
  wire  _EVAL_2705;
  wire  _EVAL_2823;
  wire  _EVAL_2503;
  wire  _EVAL_1124;
  wire  _EVAL_3011;
  wire  _EVAL_2320;
  wire  _EVAL_1100;
  wire  _EVAL_927;
  wire  _EVAL_3436;
  wire  _EVAL_2981;
  wire  _EVAL_2467;
  wire  _EVAL_3880;
  wire [7:0] _EVAL_2115;
  wire [15:0] _EVAL_2629;
  wire [31:0] _EVAL_1473;
  wire [7:0] _EVAL_946;
  wire [7:0] _EVAL_2872;
  wire [15:0] _EVAL_3380;
  wire [31:0] _EVAL_1674;
  wire [7:0] _EVAL_594;
  wire [6:0] _EVAL_2883;
  wire [14:0] _EVAL_3972;
  wire [30:0] _EVAL_3999;
  wire [126:0] _EVAL_3572;
  wire  _EVAL_1730;
  wire  _EVAL_3334;
  wire  _EVAL_1439;
  wire  _EVAL_732;
  wire  _EVAL_308;
  wire  _EVAL_2237;
  wire  _EVAL_1068;
  wire  _EVAL_1948;
  wire  _EVAL_987;
  wire  _EVAL_3620;
  wire  _EVAL_1763;
  wire  _EVAL_1235;
  wire  _EVAL_759;
  wire  _EVAL_1297;
  wire  _EVAL_1650;
  wire  _EVAL_219;
  wire  _EVAL_1768;
  wire  _EVAL_260;
  wire  _EVAL_2743;
  wire  _EVAL_1582;
  wire  _EVAL_2627;
  wire  _EVAL_3682;
  wire  _EVAL_1204;
  wire  _EVAL_1837;
  wire  _EVAL_335;
  wire  _EVAL_2449;
  wire  _EVAL_1392;
  wire  _EVAL_1541;
  wire  _EVAL_2139;
  wire  _EVAL_2644;
  wire  _EVAL_1237;
  wire  _EVAL_561;
  wire  _EVAL_679;
  wire  _EVAL_3844;
  wire  _EVAL_2545;
  wire  _EVAL_2447;
  wire  _EVAL_1957;
  wire  _EVAL_3287;
  wire  _EVAL_326;
  wire  _EVAL_4070;
  wire  _EVAL_954;
  wire  _EVAL_1213;
  wire  _EVAL_1216;
  wire  _EVAL_3615;
  wire  _EVAL_612;
  wire  _EVAL_3101;
  wire  _EVAL_896;
  wire  _EVAL_412;
  wire  _EVAL_3169;
  wire  _EVAL_1325;
  wire  _EVAL_3350;
  wire  _EVAL_2126;
  wire  _EVAL_3185;
  wire  _EVAL_203;
  wire  _EVAL_2325;
  wire  _EVAL_315;
  wire  _EVAL_355;
  wire  _EVAL_3879;
  wire  _EVAL_2242;
  wire  _EVAL_3041;
  wire  _EVAL_2669;
  wire  _EVAL_1564;
  wire  _EVAL_2455;
  wire  _EVAL_1936;
  wire  _EVAL_2129;
  wire  _EVAL_1833;
  wire  _EVAL_2468;
  wire  _EVAL_1072;
  wire  _EVAL_2097;
  wire  _EVAL_2023;
  wire  _EVAL_1677;
  wire  _EVAL_3991;
  wire  _EVAL_1919;
  wire  _EVAL_1243;
  wire  _EVAL_2144;
  wire  _EVAL_3945;
  wire  _EVAL_2454;
  wire  _EVAL_3784;
  wire  _EVAL_342;
  wire  _EVAL_3661;
  wire  _EVAL_606;
  wire  _EVAL_2690;
  wire  _EVAL_2520;
  wire  _EVAL_1013;
  wire  _EVAL_3293;
  wire  _EVAL_3659;
  wire  _EVAL_3100;
  wire  _EVAL_3709;
  wire  _EVAL_981;
  wire  _EVAL_1182;
  wire  _EVAL_2642;
  wire  _EVAL_3853;
  wire  _EVAL_3024;
  wire  _EVAL_994;
  wire  _EVAL_2103;
  wire  _EVAL_2682;
  wire  _EVAL_2229;
  wire  _EVAL_4009;
  wire  _EVAL_3142;
  wire  _EVAL_3266;
  wire  _EVAL_1096;
  wire  _EVAL_1557;
  wire  _EVAL_1492;
  wire  _EVAL_691;
  wire  _EVAL_2167;
  wire  _EVAL_3923;
  wire  _EVAL_1211;
  wire  _EVAL_2426;
  wire  _EVAL_2828;
  wire  _EVAL_1200;
  wire  _EVAL_3460;
  wire  _EVAL_2302;
  wire  _EVAL_3903;
  wire  _EVAL_1892;
  wire  _EVAL_1841;
  wire  _EVAL_380;
  wire  _EVAL_3832;
  wire  _EVAL_3490;
  wire  _EVAL_2788;
  wire  _EVAL_252;
  wire  _EVAL_720;
  wire  _EVAL_420;
  wire  _EVAL_734;
  wire  _EVAL_3868;
  wire  _EVAL_3662;
  wire  _EVAL_773;
  wire  _EVAL_1226;
  wire  _EVAL_2554;
  wire  _EVAL_231;
  wire  _EVAL_3667;
  wire  _EVAL_1400;
  wire  _EVAL_1602;
  wire  _EVAL_3823;
  wire  _EVAL_1338;
  wire [31:0] _EVAL_3244;
  wire [31:0] _EVAL_2301;
  wire [31:0] _EVAL_1171;
  wire [31:0] _EVAL_1802;
  wire  _EVAL_2011;
  wire  _EVAL_2944;
  wire  _EVAL_3579;
  wire  _EVAL_2886;
  wire  _EVAL_1427;
  wire  _EVAL_2143;
  wire  _EVAL_1671;
  wire  _EVAL_3687;
  wire  _EVAL_1240;
  wire  _EVAL_3012;
  wire  _EVAL_1611;
  wire  _EVAL_3618;
  wire  _EVAL_3625;
  wire  _EVAL_2539;
  wire  _EVAL_2939;
  wire  _EVAL_3337;
  wire  _EVAL_2187;
  wire  _EVAL_2210;
  wire  _EVAL_925;
  wire  _EVAL_3213;
  wire  _EVAL_3887;
  wire  _EVAL_345;
  wire  _EVAL_667;
  wire  _EVAL_2607;
  wire  _EVAL_2304;
  wire  _EVAL_1067;
  wire  _EVAL_3765;
  wire  _EVAL_3184;
  wire  _EVAL_2910;
  wire  _EVAL_167;
  wire  _EVAL_1370;
  wire  _EVAL_879;
  wire  _EVAL_2557;
  wire  _EVAL_1682;
  wire  _EVAL_2899;
  wire  _EVAL_2494;
  wire  _EVAL_3539;
  wire  _EVAL_1955;
  wire  _EVAL_963;
  wire  _EVAL_3371;
  wire  _EVAL_3091;
  wire  _EVAL_1617;
  wire  _EVAL_3940;
  wire  _EVAL_316;
  wire  _EVAL_1357;
  wire  _EVAL_310;
  wire  _EVAL_2421;
  wire  _EVAL_2378;
  wire  _EVAL_372;
  wire  _EVAL_3006;
  wire  _EVAL_865;
  wire  _EVAL_1751;
  wire  _EVAL_812;
  wire  _EVAL_3822;
  wire  _EVAL_2533;
  wire  _EVAL_2952;
  wire  _EVAL_2416;
  wire  _EVAL_2579;
  wire  _EVAL_3825;
  wire  _EVAL_1424;
  wire  _EVAL_2818;
  wire  _EVAL_1614;
  wire  _EVAL_1858;
  wire  _EVAL_2971;
  wire  _EVAL_2137;
  wire  _EVAL_313;
  wire  _EVAL_3107;
  wire  _EVAL_1225;
  wire  _EVAL_295;
  wire  _EVAL_3384;
  wire  _EVAL_830;
  wire  _EVAL_3157;
  wire  _EVAL_1027;
  wire  _EVAL_1131;
  wire  _EVAL_832;
  wire  _EVAL_1558;
  wire  _EVAL_557;
  wire  _EVAL_2686;
  wire  _EVAL_2854;
  wire  _EVAL_1816;
  wire  _EVAL_3547;
  wire  _EVAL_3589;
  wire  _EVAL_1210;
  wire  _EVAL_3064;
  wire  _EVAL_1835;
  wire  _EVAL_360;
  wire  _EVAL_1723;
  wire  _EVAL_4064;
  wire  _EVAL_221;
  wire  _EVAL_3946;
  wire  _EVAL_712;
  wire  _EVAL_971;
  wire  _EVAL_1161;
  wire  _EVAL_723;
  wire  _EVAL_956;
  wire  _EVAL_731;
  wire  _EVAL_539;
  wire  _EVAL_505;
  wire  _EVAL_1633;
  wire  _EVAL_875;
  wire  _EVAL_1019;
  wire  _EVAL_3374;
  wire  _EVAL_1527;
  wire  _EVAL_1120;
  wire  _EVAL_2608;
  wire  _EVAL_1555;
  wire  _EVAL_1784;
  wire  _EVAL_381;
  wire  _EVAL_1454;
  wire  _EVAL_1113;
  wire  _EVAL_3952;
  wire  _EVAL_1848;
  wire  _EVAL_190;
  wire  _EVAL_2893;
  wire  _EVAL_2225;
  wire  _EVAL_1509;
  wire  _EVAL_820;
  wire  _EVAL_242;
  wire  _EVAL_571;
  wire  _EVAL_2169;
  wire  _EVAL_199;
  wire  _EVAL_2131;
  wire  _EVAL_2365;
  wire  _EVAL_2482;
  wire  _EVAL_2651;
  wire  _EVAL_3338;
  wire  _EVAL_1655;
  wire  _EVAL_2889;
  wire  _EVAL_1350;
  wire  _EVAL_1740;
  wire  _EVAL_815;
  wire  _EVAL_788;
  wire  _EVAL_1070;
  wire  _EVAL_1771;
  wire  _EVAL_346;
  wire  _EVAL_1076;
  wire  _EVAL_476;
  wire  _EVAL_2698;
  wire  _EVAL_1386;
  wire  _EVAL_363;
  wire  _EVAL_2382;
  wire  _EVAL_268;
  wire  _EVAL_2827;
  wire  _EVAL_3047;
  wire  _EVAL_2005;
  wire  _EVAL_866;
  wire  _EVAL_793;
  wire  _EVAL_3553;
  wire [127:0] _EVAL_3469;
  wire [127:0] _EVAL_3491;
  wire  _EVAL_3263;
  wire  _EVAL_2430;
  wire  _EVAL_631;
  wire  _EVAL_2963;
  wire  _EVAL_1081;
  wire  _EVAL_1756;
  wire  _EVAL_3896;
  wire  _EVAL_3769;
  wire  _EVAL_3150;
  wire  _EVAL_3065;
  wire  _EVAL_2017;
  wire  _EVAL_2058;
  wire  _EVAL_1062;
  wire  _EVAL_1690;
  wire  _EVAL_780;
  wire  _EVAL_395;
  wire  _EVAL_1175;
  wire  _EVAL_3099;
  wire  _EVAL_2601;
  wire  _EVAL_1999;
  wire  _EVAL_2911;
  wire  _EVAL_3632;
  wire  _EVAL_3388;
  wire [126:0] _EVAL_2527;
  wire  _EVAL_3799;
  wire  _EVAL_3921;
  wire  _EVAL_3198;
  wire  _EVAL_2438;
  wire  _EVAL_1506;
  wire  _EVAL_1550;
  wire  _EVAL_2589;
  wire  _EVAL_1242;
  wire  _EVAL_807;
  wire  _EVAL_1773;
  wire  _EVAL_2059;
  wire  _EVAL_3112;
  wire  _EVAL_2330;
  wire  _EVAL_796;
  wire  _EVAL_1066;
  wire  _EVAL_2715;
  wire  _EVAL_1205;
  wire  _EVAL_3353;
  wire  _EVAL_3314;
  wire  _EVAL_1477;
  wire  _EVAL_1485;
  wire  _EVAL_3566;
  wire  _EVAL_1769;
  wire  _EVAL_1899;
  wire  _EVAL_1571;
  wire  _EVAL_4028;
  wire  _EVAL_2739;
  wire  _EVAL_1815;
  wire  _EVAL_1737;
  wire  _EVAL_3433;
  wire  _EVAL_2511;
  wire  _EVAL_1291;
  wire  _EVAL_682;
  wire  _EVAL_3515;
  wire  _EVAL_3629;
  wire  _EVAL_2309;
  wire  _EVAL_2903;
  wire  _EVAL_3890;
  wire  _EVAL_3329;
  wire  _EVAL_2142;
  wire  _EVAL_1094;
  wire  _EVAL_2358;
  wire  _EVAL_1287;
  wire  _EVAL_1135;
  wire  _EVAL_867;
  wire  _EVAL_2150;
  wire  _EVAL_3683;
  wire  _EVAL_1927;
  wire  _EVAL_3486;
  wire  _EVAL_2206;
  wire  _EVAL_1109;
  wire  _EVAL_3028;
  wire  _EVAL_3681;
  wire  _EVAL_1725;
  wire  _EVAL_2084;
  wire  _EVAL_3135;
  wire  _EVAL_1015;
  wire  _EVAL_3045;
  wire  _EVAL_2791;
  wire  _EVAL_3993;
  wire  _EVAL_2120;
  wire  _EVAL_1540;
  wire  _EVAL_1585;
  wire  _EVAL_3663;
  wire  _EVAL_1966;
  wire  _EVAL_3519;
  wire  _EVAL_1596;
  wire  _EVAL_1434;
  wire  _EVAL_2257;
  wire  _EVAL_447;
  wire  _EVAL_1758;
  wire  _EVAL_3410;
  wire  _EVAL_1063;
  wire  _EVAL_1144;
  wire  _EVAL_2885;
  wire  _EVAL_2117;
  wire  _EVAL_1333;
  wire  _EVAL_2786;
  wire  _EVAL_2163;
  wire  _EVAL_1827;
  wire  _EVAL_473;
  wire  _EVAL_2767;
  wire  _EVAL_2704;
  wire  _EVAL_968;
  wire  _EVAL_479;
  wire  _EVAL_2764;
  wire  _EVAL_864;
  wire  _EVAL_3013;
  wire  _EVAL_1640;
  wire  _EVAL_3710;
  wire  _EVAL_1190;
  wire  _EVAL_2639;
  wire  _EVAL_3186;
  wire  _EVAL_171;
  wire  _EVAL_3677;
  wire  _EVAL_2588;
  wire  _EVAL_718;
  wire  _EVAL_1472;
  wire  _EVAL_2913;
  wire  _EVAL_797;
  wire  _EVAL_3749;
  wire  _EVAL_2593;
  wire  _EVAL_2425;
  wire  _EVAL_3351;
  wire  _EVAL_450;
  wire  _EVAL_1799;
  wire  _EVAL_2316;
  wire  _EVAL_3139;
  wire  _EVAL_3426;
  wire  _EVAL_2064;
  wire  _EVAL_2404;
  wire  _EVAL_2597;
  wire  _EVAL_986;
  wire  _EVAL_3719;
  wire  _EVAL_4010;
  wire  _EVAL_3997;
  wire  _EVAL_2408;
  wire  _EVAL_1178;
  wire  _EVAL_1465;
  wire  _EVAL_1845;
  wire  _EVAL_299;
  wire  _EVAL_2109;
  wire  _EVAL_2037;
  wire  _EVAL_391;
  wire  _EVAL_1449;
  wire  _EVAL_3774;
  wire  _EVAL_341;
  wire  _EVAL_2581;
  wire  _EVAL_1311;
  wire  _EVAL_3796;
  wire  _EVAL_1093;
  wire  _EVAL_2654;
  wire  _EVAL_3456;
  wire  _EVAL_3842;
  wire  _EVAL_1728;
  wire  _EVAL_2411;
  wire  _EVAL_2015;
  wire  _EVAL_2563;
  wire  _EVAL_1559;
  wire  _EVAL_1246;
  wire  _EVAL_1244;
  wire  _EVAL_1042;
  wire  _EVAL_3751;
  wire  _EVAL_3650;
  wire  _EVAL_2070;
  wire  _EVAL_2806;
  wire [7:0] _EVAL_3020;
  wire  _EVAL_3724;
  wire  _EVAL_2590;
  wire  _EVAL_3284;
  wire  _EVAL_1378;
  wire  _EVAL_3214;
  wire  _EVAL_570;
  wire  _EVAL_3998;
  wire  _EVAL_2218;
  wire  _EVAL_706;
  wire [31:0] _EVAL_4027;
  wire [7:0] _EVAL_688;
  wire  _EVAL_2099;
  wire  _EVAL_541;
  wire  _EVAL_1139;
  wire  _EVAL_1157;
  wire  _EVAL_2909;
  wire  _EVAL_1218;
  wire  _EVAL_4061;
  wire  _EVAL_3191;
  wire  _EVAL_3281;
  wire  _EVAL_1251;
  wire  _EVAL_2278;
  wire  _EVAL_214;
  wire  _EVAL_3892;
  wire  _EVAL_3005;
  wire  _EVAL_2898;
  wire  _EVAL_1461;
  wire  _EVAL_3543;
  wire  _EVAL_3275;
  wire  _EVAL_1998;
  wire  _EVAL_2751;
  wire  _EVAL_2785;
  wire  _EVAL_3649;
  wire  _EVAL_1632;
  wire  _EVAL_3669;
  wire  _EVAL_1874;
  wire  _EVAL_1082;
  wire  _EVAL_3766;
  wire  _EVAL_3070;
  wire  _EVAL_1479;
  wire  _EVAL_2737;
  wire  _EVAL_457;
  wire  _EVAL_1134;
  wire  _EVAL_3738;
  wire  _EVAL_3356;
  wire  _EVAL_2603;
  wire  _EVAL_3495;
  wire  _EVAL_1403;
  wire  _EVAL_1591;
  wire  _EVAL_1510;
  wire  _EVAL_3583;
  wire  _EVAL_298;
  wire  _EVAL_2160;
  wire  _EVAL_2261;
  wire  _EVAL_1453;
  wire  _EVAL_1197;
  wire  _EVAL_1863;
  wire  _EVAL_2198;
  wire  _EVAL_2844;
  wire  _EVAL_1187;
  wire  _EVAL_608;
  wire  _EVAL_816;
  wire  _EVAL_3103;
  wire  _EVAL_359;
  wire  _EVAL_182;
  wire  _EVAL_1918;
  wire  _EVAL_651;
  wire  _EVAL_3939;
  wire  _EVAL_1663;
  wire  _EVAL_3764;
  wire  _EVAL_2776;
  wire  _EVAL_1446;
  wire  _EVAL_1025;
  wire  _EVAL_2729;
  wire  _EVAL_1159;
  wire  _EVAL_3581;
  wire [7:0] _EVAL_1861;
  wire  _EVAL_975;
  wire  _EVAL_2439;
  wire  _EVAL_2663;
  wire  _EVAL_576;
  wire  _EVAL_1271;
  wire  _EVAL_1842;
  wire  _EVAL_2744;
  wire [2:0] _EVAL_3965;
  SiFive__EVAL_182 LevelGateway_54 (
    ._EVAL(LevelGateway_54__EVAL),
    ._EVAL_0(LevelGateway_54__EVAL_0),
    ._EVAL_1(LevelGateway_54__EVAL_1),
    ._EVAL_2(LevelGateway_54__EVAL_2),
    ._EVAL_3(LevelGateway_54__EVAL_3),
    ._EVAL_4(LevelGateway_54__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_65 (
    ._EVAL(LevelGateway_65__EVAL),
    ._EVAL_0(LevelGateway_65__EVAL_0),
    ._EVAL_1(LevelGateway_65__EVAL_1),
    ._EVAL_2(LevelGateway_65__EVAL_2),
    ._EVAL_3(LevelGateway_65__EVAL_3),
    ._EVAL_4(LevelGateway_65__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway (
    ._EVAL(LevelGateway__EVAL),
    ._EVAL_0(LevelGateway__EVAL_0),
    ._EVAL_1(LevelGateway__EVAL_1),
    ._EVAL_2(LevelGateway__EVAL_2),
    ._EVAL_3(LevelGateway__EVAL_3),
    ._EVAL_4(LevelGateway__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_16 (
    ._EVAL(LevelGateway_16__EVAL),
    ._EVAL_0(LevelGateway_16__EVAL_0),
    ._EVAL_1(LevelGateway_16__EVAL_1),
    ._EVAL_2(LevelGateway_16__EVAL_2),
    ._EVAL_3(LevelGateway_16__EVAL_3),
    ._EVAL_4(LevelGateway_16__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_34 (
    ._EVAL(LevelGateway_34__EVAL),
    ._EVAL_0(LevelGateway_34__EVAL_0),
    ._EVAL_1(LevelGateway_34__EVAL_1),
    ._EVAL_2(LevelGateway_34__EVAL_2),
    ._EVAL_3(LevelGateway_34__EVAL_3),
    ._EVAL_4(LevelGateway_34__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_92 (
    ._EVAL(LevelGateway_92__EVAL),
    ._EVAL_0(LevelGateway_92__EVAL_0),
    ._EVAL_1(LevelGateway_92__EVAL_1),
    ._EVAL_2(LevelGateway_92__EVAL_2),
    ._EVAL_3(LevelGateway_92__EVAL_3),
    ._EVAL_4(LevelGateway_92__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_39 (
    ._EVAL(LevelGateway_39__EVAL),
    ._EVAL_0(LevelGateway_39__EVAL_0),
    ._EVAL_1(LevelGateway_39__EVAL_1),
    ._EVAL_2(LevelGateway_39__EVAL_2),
    ._EVAL_3(LevelGateway_39__EVAL_3),
    ._EVAL_4(LevelGateway_39__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_120 (
    ._EVAL(LevelGateway_120__EVAL),
    ._EVAL_0(LevelGateway_120__EVAL_0),
    ._EVAL_1(LevelGateway_120__EVAL_1),
    ._EVAL_2(LevelGateway_120__EVAL_2),
    ._EVAL_3(LevelGateway_120__EVAL_3),
    ._EVAL_4(LevelGateway_120__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_76 (
    ._EVAL(LevelGateway_76__EVAL),
    ._EVAL_0(LevelGateway_76__EVAL_0),
    ._EVAL_1(LevelGateway_76__EVAL_1),
    ._EVAL_2(LevelGateway_76__EVAL_2),
    ._EVAL_3(LevelGateway_76__EVAL_3),
    ._EVAL_4(LevelGateway_76__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_82 (
    ._EVAL(LevelGateway_82__EVAL),
    ._EVAL_0(LevelGateway_82__EVAL_0),
    ._EVAL_1(LevelGateway_82__EVAL_1),
    ._EVAL_2(LevelGateway_82__EVAL_2),
    ._EVAL_3(LevelGateway_82__EVAL_3),
    ._EVAL_4(LevelGateway_82__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_118 (
    ._EVAL(LevelGateway_118__EVAL),
    ._EVAL_0(LevelGateway_118__EVAL_0),
    ._EVAL_1(LevelGateway_118__EVAL_1),
    ._EVAL_2(LevelGateway_118__EVAL_2),
    ._EVAL_3(LevelGateway_118__EVAL_3),
    ._EVAL_4(LevelGateway_118__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_104 (
    ._EVAL(LevelGateway_104__EVAL),
    ._EVAL_0(LevelGateway_104__EVAL_0),
    ._EVAL_1(LevelGateway_104__EVAL_1),
    ._EVAL_2(LevelGateway_104__EVAL_2),
    ._EVAL_3(LevelGateway_104__EVAL_3),
    ._EVAL_4(LevelGateway_104__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_112 (
    ._EVAL(LevelGateway_112__EVAL),
    ._EVAL_0(LevelGateway_112__EVAL_0),
    ._EVAL_1(LevelGateway_112__EVAL_1),
    ._EVAL_2(LevelGateway_112__EVAL_2),
    ._EVAL_3(LevelGateway_112__EVAL_3),
    ._EVAL_4(LevelGateway_112__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_50 (
    ._EVAL(LevelGateway_50__EVAL),
    ._EVAL_0(LevelGateway_50__EVAL_0),
    ._EVAL_1(LevelGateway_50__EVAL_1),
    ._EVAL_2(LevelGateway_50__EVAL_2),
    ._EVAL_3(LevelGateway_50__EVAL_3),
    ._EVAL_4(LevelGateway_50__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_96 (
    ._EVAL(LevelGateway_96__EVAL),
    ._EVAL_0(LevelGateway_96__EVAL_0),
    ._EVAL_1(LevelGateway_96__EVAL_1),
    ._EVAL_2(LevelGateway_96__EVAL_2),
    ._EVAL_3(LevelGateway_96__EVAL_3),
    ._EVAL_4(LevelGateway_96__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_108 (
    ._EVAL(LevelGateway_108__EVAL),
    ._EVAL_0(LevelGateway_108__EVAL_0),
    ._EVAL_1(LevelGateway_108__EVAL_1),
    ._EVAL_2(LevelGateway_108__EVAL_2),
    ._EVAL_3(LevelGateway_108__EVAL_3),
    ._EVAL_4(LevelGateway_108__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_101 (
    ._EVAL(LevelGateway_101__EVAL),
    ._EVAL_0(LevelGateway_101__EVAL_0),
    ._EVAL_1(LevelGateway_101__EVAL_1),
    ._EVAL_2(LevelGateway_101__EVAL_2),
    ._EVAL_3(LevelGateway_101__EVAL_3),
    ._EVAL_4(LevelGateway_101__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_79 (
    ._EVAL(LevelGateway_79__EVAL),
    ._EVAL_0(LevelGateway_79__EVAL_0),
    ._EVAL_1(LevelGateway_79__EVAL_1),
    ._EVAL_2(LevelGateway_79__EVAL_2),
    ._EVAL_3(LevelGateway_79__EVAL_3),
    ._EVAL_4(LevelGateway_79__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_42 (
    ._EVAL(LevelGateway_42__EVAL),
    ._EVAL_0(LevelGateway_42__EVAL_0),
    ._EVAL_1(LevelGateway_42__EVAL_1),
    ._EVAL_2(LevelGateway_42__EVAL_2),
    ._EVAL_3(LevelGateway_42__EVAL_3),
    ._EVAL_4(LevelGateway_42__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_55 (
    ._EVAL(LevelGateway_55__EVAL),
    ._EVAL_0(LevelGateway_55__EVAL_0),
    ._EVAL_1(LevelGateway_55__EVAL_1),
    ._EVAL_2(LevelGateway_55__EVAL_2),
    ._EVAL_3(LevelGateway_55__EVAL_3),
    ._EVAL_4(LevelGateway_55__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_109 (
    ._EVAL(LevelGateway_109__EVAL),
    ._EVAL_0(LevelGateway_109__EVAL_0),
    ._EVAL_1(LevelGateway_109__EVAL_1),
    ._EVAL_2(LevelGateway_109__EVAL_2),
    ._EVAL_3(LevelGateway_109__EVAL_3),
    ._EVAL_4(LevelGateway_109__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_105 (
    ._EVAL(LevelGateway_105__EVAL),
    ._EVAL_0(LevelGateway_105__EVAL_0),
    ._EVAL_1(LevelGateway_105__EVAL_1),
    ._EVAL_2(LevelGateway_105__EVAL_2),
    ._EVAL_3(LevelGateway_105__EVAL_3),
    ._EVAL_4(LevelGateway_105__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_63 (
    ._EVAL(LevelGateway_63__EVAL),
    ._EVAL_0(LevelGateway_63__EVAL_0),
    ._EVAL_1(LevelGateway_63__EVAL_1),
    ._EVAL_2(LevelGateway_63__EVAL_2),
    ._EVAL_3(LevelGateway_63__EVAL_3),
    ._EVAL_4(LevelGateway_63__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_14 (
    ._EVAL(LevelGateway_14__EVAL),
    ._EVAL_0(LevelGateway_14__EVAL_0),
    ._EVAL_1(LevelGateway_14__EVAL_1),
    ._EVAL_2(LevelGateway_14__EVAL_2),
    ._EVAL_3(LevelGateway_14__EVAL_3),
    ._EVAL_4(LevelGateway_14__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_44 (
    ._EVAL(LevelGateway_44__EVAL),
    ._EVAL_0(LevelGateway_44__EVAL_0),
    ._EVAL_1(LevelGateway_44__EVAL_1),
    ._EVAL_2(LevelGateway_44__EVAL_2),
    ._EVAL_3(LevelGateway_44__EVAL_3),
    ._EVAL_4(LevelGateway_44__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_123 (
    ._EVAL(LevelGateway_123__EVAL),
    ._EVAL_0(LevelGateway_123__EVAL_0),
    ._EVAL_1(LevelGateway_123__EVAL_1),
    ._EVAL_2(LevelGateway_123__EVAL_2),
    ._EVAL_3(LevelGateway_123__EVAL_3),
    ._EVAL_4(LevelGateway_123__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_70 (
    ._EVAL(LevelGateway_70__EVAL),
    ._EVAL_0(LevelGateway_70__EVAL_0),
    ._EVAL_1(LevelGateway_70__EVAL_1),
    ._EVAL_2(LevelGateway_70__EVAL_2),
    ._EVAL_3(LevelGateway_70__EVAL_3),
    ._EVAL_4(LevelGateway_70__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_122 (
    ._EVAL(LevelGateway_122__EVAL),
    ._EVAL_0(LevelGateway_122__EVAL_0),
    ._EVAL_1(LevelGateway_122__EVAL_1),
    ._EVAL_2(LevelGateway_122__EVAL_2),
    ._EVAL_3(LevelGateway_122__EVAL_3),
    ._EVAL_4(LevelGateway_122__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_4 (
    ._EVAL(LevelGateway_4__EVAL),
    ._EVAL_0(LevelGateway_4__EVAL_0),
    ._EVAL_1(LevelGateway_4__EVAL_1),
    ._EVAL_2(LevelGateway_4__EVAL_2),
    ._EVAL_3(LevelGateway_4__EVAL_3),
    ._EVAL_4(LevelGateway_4__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_5 (
    ._EVAL(LevelGateway_5__EVAL),
    ._EVAL_0(LevelGateway_5__EVAL_0),
    ._EVAL_1(LevelGateway_5__EVAL_1),
    ._EVAL_2(LevelGateway_5__EVAL_2),
    ._EVAL_3(LevelGateway_5__EVAL_3),
    ._EVAL_4(LevelGateway_5__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_37 (
    ._EVAL(LevelGateway_37__EVAL),
    ._EVAL_0(LevelGateway_37__EVAL_0),
    ._EVAL_1(LevelGateway_37__EVAL_1),
    ._EVAL_2(LevelGateway_37__EVAL_2),
    ._EVAL_3(LevelGateway_37__EVAL_3),
    ._EVAL_4(LevelGateway_37__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_25 (
    ._EVAL(LevelGateway_25__EVAL),
    ._EVAL_0(LevelGateway_25__EVAL_0),
    ._EVAL_1(LevelGateway_25__EVAL_1),
    ._EVAL_2(LevelGateway_25__EVAL_2),
    ._EVAL_3(LevelGateway_25__EVAL_3),
    ._EVAL_4(LevelGateway_25__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_114 (
    ._EVAL(LevelGateway_114__EVAL),
    ._EVAL_0(LevelGateway_114__EVAL_0),
    ._EVAL_1(LevelGateway_114__EVAL_1),
    ._EVAL_2(LevelGateway_114__EVAL_2),
    ._EVAL_3(LevelGateway_114__EVAL_3),
    ._EVAL_4(LevelGateway_114__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_56 (
    ._EVAL(LevelGateway_56__EVAL),
    ._EVAL_0(LevelGateway_56__EVAL_0),
    ._EVAL_1(LevelGateway_56__EVAL_1),
    ._EVAL_2(LevelGateway_56__EVAL_2),
    ._EVAL_3(LevelGateway_56__EVAL_3),
    ._EVAL_4(LevelGateway_56__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_71 (
    ._EVAL(LevelGateway_71__EVAL),
    ._EVAL_0(LevelGateway_71__EVAL_0),
    ._EVAL_1(LevelGateway_71__EVAL_1),
    ._EVAL_2(LevelGateway_71__EVAL_2),
    ._EVAL_3(LevelGateway_71__EVAL_3),
    ._EVAL_4(LevelGateway_71__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_64 (
    ._EVAL(LevelGateway_64__EVAL),
    ._EVAL_0(LevelGateway_64__EVAL_0),
    ._EVAL_1(LevelGateway_64__EVAL_1),
    ._EVAL_2(LevelGateway_64__EVAL_2),
    ._EVAL_3(LevelGateway_64__EVAL_3),
    ._EVAL_4(LevelGateway_64__EVAL_4)
  );
  SiFive__EVAL_184 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14)
  );
  SiFive__EVAL_182 LevelGateway_73 (
    ._EVAL(LevelGateway_73__EVAL),
    ._EVAL_0(LevelGateway_73__EVAL_0),
    ._EVAL_1(LevelGateway_73__EVAL_1),
    ._EVAL_2(LevelGateway_73__EVAL_2),
    ._EVAL_3(LevelGateway_73__EVAL_3),
    ._EVAL_4(LevelGateway_73__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_99 (
    ._EVAL(LevelGateway_99__EVAL),
    ._EVAL_0(LevelGateway_99__EVAL_0),
    ._EVAL_1(LevelGateway_99__EVAL_1),
    ._EVAL_2(LevelGateway_99__EVAL_2),
    ._EVAL_3(LevelGateway_99__EVAL_3),
    ._EVAL_4(LevelGateway_99__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_115 (
    ._EVAL(LevelGateway_115__EVAL),
    ._EVAL_0(LevelGateway_115__EVAL_0),
    ._EVAL_1(LevelGateway_115__EVAL_1),
    ._EVAL_2(LevelGateway_115__EVAL_2),
    ._EVAL_3(LevelGateway_115__EVAL_3),
    ._EVAL_4(LevelGateway_115__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_94 (
    ._EVAL(LevelGateway_94__EVAL),
    ._EVAL_0(LevelGateway_94__EVAL_0),
    ._EVAL_1(LevelGateway_94__EVAL_1),
    ._EVAL_2(LevelGateway_94__EVAL_2),
    ._EVAL_3(LevelGateway_94__EVAL_3),
    ._EVAL_4(LevelGateway_94__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_49 (
    ._EVAL(LevelGateway_49__EVAL),
    ._EVAL_0(LevelGateway_49__EVAL_0),
    ._EVAL_1(LevelGateway_49__EVAL_1),
    ._EVAL_2(LevelGateway_49__EVAL_2),
    ._EVAL_3(LevelGateway_49__EVAL_3),
    ._EVAL_4(LevelGateway_49__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_48 (
    ._EVAL(LevelGateway_48__EVAL),
    ._EVAL_0(LevelGateway_48__EVAL_0),
    ._EVAL_1(LevelGateway_48__EVAL_1),
    ._EVAL_2(LevelGateway_48__EVAL_2),
    ._EVAL_3(LevelGateway_48__EVAL_3),
    ._EVAL_4(LevelGateway_48__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_62 (
    ._EVAL(LevelGateway_62__EVAL),
    ._EVAL_0(LevelGateway_62__EVAL_0),
    ._EVAL_1(LevelGateway_62__EVAL_1),
    ._EVAL_2(LevelGateway_62__EVAL_2),
    ._EVAL_3(LevelGateway_62__EVAL_3),
    ._EVAL_4(LevelGateway_62__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_103 (
    ._EVAL(LevelGateway_103__EVAL),
    ._EVAL_0(LevelGateway_103__EVAL_0),
    ._EVAL_1(LevelGateway_103__EVAL_1),
    ._EVAL_2(LevelGateway_103__EVAL_2),
    ._EVAL_3(LevelGateway_103__EVAL_3),
    ._EVAL_4(LevelGateway_103__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_15 (
    ._EVAL(LevelGateway_15__EVAL),
    ._EVAL_0(LevelGateway_15__EVAL_0),
    ._EVAL_1(LevelGateway_15__EVAL_1),
    ._EVAL_2(LevelGateway_15__EVAL_2),
    ._EVAL_3(LevelGateway_15__EVAL_3),
    ._EVAL_4(LevelGateway_15__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_102 (
    ._EVAL(LevelGateway_102__EVAL),
    ._EVAL_0(LevelGateway_102__EVAL_0),
    ._EVAL_1(LevelGateway_102__EVAL_1),
    ._EVAL_2(LevelGateway_102__EVAL_2),
    ._EVAL_3(LevelGateway_102__EVAL_3),
    ._EVAL_4(LevelGateway_102__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_83 (
    ._EVAL(LevelGateway_83__EVAL),
    ._EVAL_0(LevelGateway_83__EVAL_0),
    ._EVAL_1(LevelGateway_83__EVAL_1),
    ._EVAL_2(LevelGateway_83__EVAL_2),
    ._EVAL_3(LevelGateway_83__EVAL_3),
    ._EVAL_4(LevelGateway_83__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_95 (
    ._EVAL(LevelGateway_95__EVAL),
    ._EVAL_0(LevelGateway_95__EVAL_0),
    ._EVAL_1(LevelGateway_95__EVAL_1),
    ._EVAL_2(LevelGateway_95__EVAL_2),
    ._EVAL_3(LevelGateway_95__EVAL_3),
    ._EVAL_4(LevelGateway_95__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_38 (
    ._EVAL(LevelGateway_38__EVAL),
    ._EVAL_0(LevelGateway_38__EVAL_0),
    ._EVAL_1(LevelGateway_38__EVAL_1),
    ._EVAL_2(LevelGateway_38__EVAL_2),
    ._EVAL_3(LevelGateway_38__EVAL_3),
    ._EVAL_4(LevelGateway_38__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_29 (
    ._EVAL(LevelGateway_29__EVAL),
    ._EVAL_0(LevelGateway_29__EVAL_0),
    ._EVAL_1(LevelGateway_29__EVAL_1),
    ._EVAL_2(LevelGateway_29__EVAL_2),
    ._EVAL_3(LevelGateway_29__EVAL_3),
    ._EVAL_4(LevelGateway_29__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_35 (
    ._EVAL(LevelGateway_35__EVAL),
    ._EVAL_0(LevelGateway_35__EVAL_0),
    ._EVAL_1(LevelGateway_35__EVAL_1),
    ._EVAL_2(LevelGateway_35__EVAL_2),
    ._EVAL_3(LevelGateway_35__EVAL_3),
    ._EVAL_4(LevelGateway_35__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_9 (
    ._EVAL(LevelGateway_9__EVAL),
    ._EVAL_0(LevelGateway_9__EVAL_0),
    ._EVAL_1(LevelGateway_9__EVAL_1),
    ._EVAL_2(LevelGateway_9__EVAL_2),
    ._EVAL_3(LevelGateway_9__EVAL_3),
    ._EVAL_4(LevelGateway_9__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_86 (
    ._EVAL(LevelGateway_86__EVAL),
    ._EVAL_0(LevelGateway_86__EVAL_0),
    ._EVAL_1(LevelGateway_86__EVAL_1),
    ._EVAL_2(LevelGateway_86__EVAL_2),
    ._EVAL_3(LevelGateway_86__EVAL_3),
    ._EVAL_4(LevelGateway_86__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_100 (
    ._EVAL(LevelGateway_100__EVAL),
    ._EVAL_0(LevelGateway_100__EVAL_0),
    ._EVAL_1(LevelGateway_100__EVAL_1),
    ._EVAL_2(LevelGateway_100__EVAL_2),
    ._EVAL_3(LevelGateway_100__EVAL_3),
    ._EVAL_4(LevelGateway_100__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_69 (
    ._EVAL(LevelGateway_69__EVAL),
    ._EVAL_0(LevelGateway_69__EVAL_0),
    ._EVAL_1(LevelGateway_69__EVAL_1),
    ._EVAL_2(LevelGateway_69__EVAL_2),
    ._EVAL_3(LevelGateway_69__EVAL_3),
    ._EVAL_4(LevelGateway_69__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_81 (
    ._EVAL(LevelGateway_81__EVAL),
    ._EVAL_0(LevelGateway_81__EVAL_0),
    ._EVAL_1(LevelGateway_81__EVAL_1),
    ._EVAL_2(LevelGateway_81__EVAL_2),
    ._EVAL_3(LevelGateway_81__EVAL_3),
    ._EVAL_4(LevelGateway_81__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_75 (
    ._EVAL(LevelGateway_75__EVAL),
    ._EVAL_0(LevelGateway_75__EVAL_0),
    ._EVAL_1(LevelGateway_75__EVAL_1),
    ._EVAL_2(LevelGateway_75__EVAL_2),
    ._EVAL_3(LevelGateway_75__EVAL_3),
    ._EVAL_4(LevelGateway_75__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_66 (
    ._EVAL(LevelGateway_66__EVAL),
    ._EVAL_0(LevelGateway_66__EVAL_0),
    ._EVAL_1(LevelGateway_66__EVAL_1),
    ._EVAL_2(LevelGateway_66__EVAL_2),
    ._EVAL_3(LevelGateway_66__EVAL_3),
    ._EVAL_4(LevelGateway_66__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_10 (
    ._EVAL(LevelGateway_10__EVAL),
    ._EVAL_0(LevelGateway_10__EVAL_0),
    ._EVAL_1(LevelGateway_10__EVAL_1),
    ._EVAL_2(LevelGateway_10__EVAL_2),
    ._EVAL_3(LevelGateway_10__EVAL_3),
    ._EVAL_4(LevelGateway_10__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_91 (
    ._EVAL(LevelGateway_91__EVAL),
    ._EVAL_0(LevelGateway_91__EVAL_0),
    ._EVAL_1(LevelGateway_91__EVAL_1),
    ._EVAL_2(LevelGateway_91__EVAL_2),
    ._EVAL_3(LevelGateway_91__EVAL_3),
    ._EVAL_4(LevelGateway_91__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_67 (
    ._EVAL(LevelGateway_67__EVAL),
    ._EVAL_0(LevelGateway_67__EVAL_0),
    ._EVAL_1(LevelGateway_67__EVAL_1),
    ._EVAL_2(LevelGateway_67__EVAL_2),
    ._EVAL_3(LevelGateway_67__EVAL_3),
    ._EVAL_4(LevelGateway_67__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_27 (
    ._EVAL(LevelGateway_27__EVAL),
    ._EVAL_0(LevelGateway_27__EVAL_0),
    ._EVAL_1(LevelGateway_27__EVAL_1),
    ._EVAL_2(LevelGateway_27__EVAL_2),
    ._EVAL_3(LevelGateway_27__EVAL_3),
    ._EVAL_4(LevelGateway_27__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_89 (
    ._EVAL(LevelGateway_89__EVAL),
    ._EVAL_0(LevelGateway_89__EVAL_0),
    ._EVAL_1(LevelGateway_89__EVAL_1),
    ._EVAL_2(LevelGateway_89__EVAL_2),
    ._EVAL_3(LevelGateway_89__EVAL_3),
    ._EVAL_4(LevelGateway_89__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_12 (
    ._EVAL(LevelGateway_12__EVAL),
    ._EVAL_0(LevelGateway_12__EVAL_0),
    ._EVAL_1(LevelGateway_12__EVAL_1),
    ._EVAL_2(LevelGateway_12__EVAL_2),
    ._EVAL_3(LevelGateway_12__EVAL_3),
    ._EVAL_4(LevelGateway_12__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_28 (
    ._EVAL(LevelGateway_28__EVAL),
    ._EVAL_0(LevelGateway_28__EVAL_0),
    ._EVAL_1(LevelGateway_28__EVAL_1),
    ._EVAL_2(LevelGateway_28__EVAL_2),
    ._EVAL_3(LevelGateway_28__EVAL_3),
    ._EVAL_4(LevelGateway_28__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_58 (
    ._EVAL(LevelGateway_58__EVAL),
    ._EVAL_0(LevelGateway_58__EVAL_0),
    ._EVAL_1(LevelGateway_58__EVAL_1),
    ._EVAL_2(LevelGateway_58__EVAL_2),
    ._EVAL_3(LevelGateway_58__EVAL_3),
    ._EVAL_4(LevelGateway_58__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_6 (
    ._EVAL(LevelGateway_6__EVAL),
    ._EVAL_0(LevelGateway_6__EVAL_0),
    ._EVAL_1(LevelGateway_6__EVAL_1),
    ._EVAL_2(LevelGateway_6__EVAL_2),
    ._EVAL_3(LevelGateway_6__EVAL_3),
    ._EVAL_4(LevelGateway_6__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_98 (
    ._EVAL(LevelGateway_98__EVAL),
    ._EVAL_0(LevelGateway_98__EVAL_0),
    ._EVAL_1(LevelGateway_98__EVAL_1),
    ._EVAL_2(LevelGateway_98__EVAL_2),
    ._EVAL_3(LevelGateway_98__EVAL_3),
    ._EVAL_4(LevelGateway_98__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_107 (
    ._EVAL(LevelGateway_107__EVAL),
    ._EVAL_0(LevelGateway_107__EVAL_0),
    ._EVAL_1(LevelGateway_107__EVAL_1),
    ._EVAL_2(LevelGateway_107__EVAL_2),
    ._EVAL_3(LevelGateway_107__EVAL_3),
    ._EVAL_4(LevelGateway_107__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_93 (
    ._EVAL(LevelGateway_93__EVAL),
    ._EVAL_0(LevelGateway_93__EVAL_0),
    ._EVAL_1(LevelGateway_93__EVAL_1),
    ._EVAL_2(LevelGateway_93__EVAL_2),
    ._EVAL_3(LevelGateway_93__EVAL_3),
    ._EVAL_4(LevelGateway_93__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_126 (
    ._EVAL(LevelGateway_126__EVAL),
    ._EVAL_0(LevelGateway_126__EVAL_0),
    ._EVAL_1(LevelGateway_126__EVAL_1),
    ._EVAL_2(LevelGateway_126__EVAL_2),
    ._EVAL_3(LevelGateway_126__EVAL_3),
    ._EVAL_4(LevelGateway_126__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_97 (
    ._EVAL(LevelGateway_97__EVAL),
    ._EVAL_0(LevelGateway_97__EVAL_0),
    ._EVAL_1(LevelGateway_97__EVAL_1),
    ._EVAL_2(LevelGateway_97__EVAL_2),
    ._EVAL_3(LevelGateway_97__EVAL_3),
    ._EVAL_4(LevelGateway_97__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_57 (
    ._EVAL(LevelGateway_57__EVAL),
    ._EVAL_0(LevelGateway_57__EVAL_0),
    ._EVAL_1(LevelGateway_57__EVAL_1),
    ._EVAL_2(LevelGateway_57__EVAL_2),
    ._EVAL_3(LevelGateway_57__EVAL_3),
    ._EVAL_4(LevelGateway_57__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_72 (
    ._EVAL(LevelGateway_72__EVAL),
    ._EVAL_0(LevelGateway_72__EVAL_0),
    ._EVAL_1(LevelGateway_72__EVAL_1),
    ._EVAL_2(LevelGateway_72__EVAL_2),
    ._EVAL_3(LevelGateway_72__EVAL_3),
    ._EVAL_4(LevelGateway_72__EVAL_4)
  );
  SiFive__EVAL_183 PLICFanIn (
    ._EVAL(PLICFanIn__EVAL),
    ._EVAL_0(PLICFanIn__EVAL_0),
    ._EVAL_1(PLICFanIn__EVAL_1),
    ._EVAL_2(PLICFanIn__EVAL_2),
    ._EVAL_3(PLICFanIn__EVAL_3),
    ._EVAL_4(PLICFanIn__EVAL_4),
    ._EVAL_5(PLICFanIn__EVAL_5),
    ._EVAL_6(PLICFanIn__EVAL_6),
    ._EVAL_7(PLICFanIn__EVAL_7),
    ._EVAL_8(PLICFanIn__EVAL_8),
    ._EVAL_9(PLICFanIn__EVAL_9),
    ._EVAL_10(PLICFanIn__EVAL_10),
    ._EVAL_11(PLICFanIn__EVAL_11),
    ._EVAL_12(PLICFanIn__EVAL_12),
    ._EVAL_13(PLICFanIn__EVAL_13),
    ._EVAL_14(PLICFanIn__EVAL_14),
    ._EVAL_15(PLICFanIn__EVAL_15),
    ._EVAL_16(PLICFanIn__EVAL_16),
    ._EVAL_17(PLICFanIn__EVAL_17),
    ._EVAL_18(PLICFanIn__EVAL_18),
    ._EVAL_19(PLICFanIn__EVAL_19),
    ._EVAL_20(PLICFanIn__EVAL_20),
    ._EVAL_21(PLICFanIn__EVAL_21),
    ._EVAL_22(PLICFanIn__EVAL_22),
    ._EVAL_23(PLICFanIn__EVAL_23),
    ._EVAL_24(PLICFanIn__EVAL_24),
    ._EVAL_25(PLICFanIn__EVAL_25),
    ._EVAL_26(PLICFanIn__EVAL_26),
    ._EVAL_27(PLICFanIn__EVAL_27),
    ._EVAL_28(PLICFanIn__EVAL_28),
    ._EVAL_29(PLICFanIn__EVAL_29),
    ._EVAL_30(PLICFanIn__EVAL_30),
    ._EVAL_31(PLICFanIn__EVAL_31),
    ._EVAL_32(PLICFanIn__EVAL_32),
    ._EVAL_33(PLICFanIn__EVAL_33),
    ._EVAL_34(PLICFanIn__EVAL_34),
    ._EVAL_35(PLICFanIn__EVAL_35),
    ._EVAL_36(PLICFanIn__EVAL_36),
    ._EVAL_37(PLICFanIn__EVAL_37),
    ._EVAL_38(PLICFanIn__EVAL_38),
    ._EVAL_39(PLICFanIn__EVAL_39),
    ._EVAL_40(PLICFanIn__EVAL_40),
    ._EVAL_41(PLICFanIn__EVAL_41),
    ._EVAL_42(PLICFanIn__EVAL_42),
    ._EVAL_43(PLICFanIn__EVAL_43),
    ._EVAL_44(PLICFanIn__EVAL_44),
    ._EVAL_45(PLICFanIn__EVAL_45),
    ._EVAL_46(PLICFanIn__EVAL_46),
    ._EVAL_47(PLICFanIn__EVAL_47),
    ._EVAL_48(PLICFanIn__EVAL_48),
    ._EVAL_49(PLICFanIn__EVAL_49),
    ._EVAL_50(PLICFanIn__EVAL_50),
    ._EVAL_51(PLICFanIn__EVAL_51),
    ._EVAL_52(PLICFanIn__EVAL_52),
    ._EVAL_53(PLICFanIn__EVAL_53),
    ._EVAL_54(PLICFanIn__EVAL_54),
    ._EVAL_55(PLICFanIn__EVAL_55),
    ._EVAL_56(PLICFanIn__EVAL_56),
    ._EVAL_57(PLICFanIn__EVAL_57),
    ._EVAL_58(PLICFanIn__EVAL_58),
    ._EVAL_59(PLICFanIn__EVAL_59),
    ._EVAL_60(PLICFanIn__EVAL_60),
    ._EVAL_61(PLICFanIn__EVAL_61),
    ._EVAL_62(PLICFanIn__EVAL_62),
    ._EVAL_63(PLICFanIn__EVAL_63),
    ._EVAL_64(PLICFanIn__EVAL_64),
    ._EVAL_65(PLICFanIn__EVAL_65),
    ._EVAL_66(PLICFanIn__EVAL_66),
    ._EVAL_67(PLICFanIn__EVAL_67),
    ._EVAL_68(PLICFanIn__EVAL_68),
    ._EVAL_69(PLICFanIn__EVAL_69),
    ._EVAL_70(PLICFanIn__EVAL_70),
    ._EVAL_71(PLICFanIn__EVAL_71),
    ._EVAL_72(PLICFanIn__EVAL_72),
    ._EVAL_73(PLICFanIn__EVAL_73),
    ._EVAL_74(PLICFanIn__EVAL_74),
    ._EVAL_75(PLICFanIn__EVAL_75),
    ._EVAL_76(PLICFanIn__EVAL_76),
    ._EVAL_77(PLICFanIn__EVAL_77),
    ._EVAL_78(PLICFanIn__EVAL_78),
    ._EVAL_79(PLICFanIn__EVAL_79),
    ._EVAL_80(PLICFanIn__EVAL_80),
    ._EVAL_81(PLICFanIn__EVAL_81),
    ._EVAL_82(PLICFanIn__EVAL_82),
    ._EVAL_83(PLICFanIn__EVAL_83),
    ._EVAL_84(PLICFanIn__EVAL_84),
    ._EVAL_85(PLICFanIn__EVAL_85),
    ._EVAL_86(PLICFanIn__EVAL_86),
    ._EVAL_87(PLICFanIn__EVAL_87),
    ._EVAL_88(PLICFanIn__EVAL_88),
    ._EVAL_89(PLICFanIn__EVAL_89),
    ._EVAL_90(PLICFanIn__EVAL_90),
    ._EVAL_91(PLICFanIn__EVAL_91),
    ._EVAL_92(PLICFanIn__EVAL_92),
    ._EVAL_93(PLICFanIn__EVAL_93),
    ._EVAL_94(PLICFanIn__EVAL_94),
    ._EVAL_95(PLICFanIn__EVAL_95),
    ._EVAL_96(PLICFanIn__EVAL_96),
    ._EVAL_97(PLICFanIn__EVAL_97),
    ._EVAL_98(PLICFanIn__EVAL_98),
    ._EVAL_99(PLICFanIn__EVAL_99),
    ._EVAL_100(PLICFanIn__EVAL_100),
    ._EVAL_101(PLICFanIn__EVAL_101),
    ._EVAL_102(PLICFanIn__EVAL_102),
    ._EVAL_103(PLICFanIn__EVAL_103),
    ._EVAL_104(PLICFanIn__EVAL_104),
    ._EVAL_105(PLICFanIn__EVAL_105),
    ._EVAL_106(PLICFanIn__EVAL_106),
    ._EVAL_107(PLICFanIn__EVAL_107),
    ._EVAL_108(PLICFanIn__EVAL_108),
    ._EVAL_109(PLICFanIn__EVAL_109),
    ._EVAL_110(PLICFanIn__EVAL_110),
    ._EVAL_111(PLICFanIn__EVAL_111),
    ._EVAL_112(PLICFanIn__EVAL_112),
    ._EVAL_113(PLICFanIn__EVAL_113),
    ._EVAL_114(PLICFanIn__EVAL_114),
    ._EVAL_115(PLICFanIn__EVAL_115),
    ._EVAL_116(PLICFanIn__EVAL_116),
    ._EVAL_117(PLICFanIn__EVAL_117),
    ._EVAL_118(PLICFanIn__EVAL_118),
    ._EVAL_119(PLICFanIn__EVAL_119),
    ._EVAL_120(PLICFanIn__EVAL_120),
    ._EVAL_121(PLICFanIn__EVAL_121),
    ._EVAL_122(PLICFanIn__EVAL_122),
    ._EVAL_123(PLICFanIn__EVAL_123),
    ._EVAL_124(PLICFanIn__EVAL_124),
    ._EVAL_125(PLICFanIn__EVAL_125),
    ._EVAL_126(PLICFanIn__EVAL_126),
    ._EVAL_127(PLICFanIn__EVAL_127),
    ._EVAL_128(PLICFanIn__EVAL_128)
  );
  SiFive__EVAL_182 LevelGateway_43 (
    ._EVAL(LevelGateway_43__EVAL),
    ._EVAL_0(LevelGateway_43__EVAL_0),
    ._EVAL_1(LevelGateway_43__EVAL_1),
    ._EVAL_2(LevelGateway_43__EVAL_2),
    ._EVAL_3(LevelGateway_43__EVAL_3),
    ._EVAL_4(LevelGateway_43__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_30 (
    ._EVAL(LevelGateway_30__EVAL),
    ._EVAL_0(LevelGateway_30__EVAL_0),
    ._EVAL_1(LevelGateway_30__EVAL_1),
    ._EVAL_2(LevelGateway_30__EVAL_2),
    ._EVAL_3(LevelGateway_30__EVAL_3),
    ._EVAL_4(LevelGateway_30__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_7 (
    ._EVAL(LevelGateway_7__EVAL),
    ._EVAL_0(LevelGateway_7__EVAL_0),
    ._EVAL_1(LevelGateway_7__EVAL_1),
    ._EVAL_2(LevelGateway_7__EVAL_2),
    ._EVAL_3(LevelGateway_7__EVAL_3),
    ._EVAL_4(LevelGateway_7__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_68 (
    ._EVAL(LevelGateway_68__EVAL),
    ._EVAL_0(LevelGateway_68__EVAL_0),
    ._EVAL_1(LevelGateway_68__EVAL_1),
    ._EVAL_2(LevelGateway_68__EVAL_2),
    ._EVAL_3(LevelGateway_68__EVAL_3),
    ._EVAL_4(LevelGateway_68__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_84 (
    ._EVAL(LevelGateway_84__EVAL),
    ._EVAL_0(LevelGateway_84__EVAL_0),
    ._EVAL_1(LevelGateway_84__EVAL_1),
    ._EVAL_2(LevelGateway_84__EVAL_2),
    ._EVAL_3(LevelGateway_84__EVAL_3),
    ._EVAL_4(LevelGateway_84__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_116 (
    ._EVAL(LevelGateway_116__EVAL),
    ._EVAL_0(LevelGateway_116__EVAL_0),
    ._EVAL_1(LevelGateway_116__EVAL_1),
    ._EVAL_2(LevelGateway_116__EVAL_2),
    ._EVAL_3(LevelGateway_116__EVAL_3),
    ._EVAL_4(LevelGateway_116__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_53 (
    ._EVAL(LevelGateway_53__EVAL),
    ._EVAL_0(LevelGateway_53__EVAL_0),
    ._EVAL_1(LevelGateway_53__EVAL_1),
    ._EVAL_2(LevelGateway_53__EVAL_2),
    ._EVAL_3(LevelGateway_53__EVAL_3),
    ._EVAL_4(LevelGateway_53__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_88 (
    ._EVAL(LevelGateway_88__EVAL),
    ._EVAL_0(LevelGateway_88__EVAL_0),
    ._EVAL_1(LevelGateway_88__EVAL_1),
    ._EVAL_2(LevelGateway_88__EVAL_2),
    ._EVAL_3(LevelGateway_88__EVAL_3),
    ._EVAL_4(LevelGateway_88__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_13 (
    ._EVAL(LevelGateway_13__EVAL),
    ._EVAL_0(LevelGateway_13__EVAL_0),
    ._EVAL_1(LevelGateway_13__EVAL_1),
    ._EVAL_2(LevelGateway_13__EVAL_2),
    ._EVAL_3(LevelGateway_13__EVAL_3),
    ._EVAL_4(LevelGateway_13__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_117 (
    ._EVAL(LevelGateway_117__EVAL),
    ._EVAL_0(LevelGateway_117__EVAL_0),
    ._EVAL_1(LevelGateway_117__EVAL_1),
    ._EVAL_2(LevelGateway_117__EVAL_2),
    ._EVAL_3(LevelGateway_117__EVAL_3),
    ._EVAL_4(LevelGateway_117__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_3 (
    ._EVAL(LevelGateway_3__EVAL),
    ._EVAL_0(LevelGateway_3__EVAL_0),
    ._EVAL_1(LevelGateway_3__EVAL_1),
    ._EVAL_2(LevelGateway_3__EVAL_2),
    ._EVAL_3(LevelGateway_3__EVAL_3),
    ._EVAL_4(LevelGateway_3__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_47 (
    ._EVAL(LevelGateway_47__EVAL),
    ._EVAL_0(LevelGateway_47__EVAL_0),
    ._EVAL_1(LevelGateway_47__EVAL_1),
    ._EVAL_2(LevelGateway_47__EVAL_2),
    ._EVAL_3(LevelGateway_47__EVAL_3),
    ._EVAL_4(LevelGateway_47__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_85 (
    ._EVAL(LevelGateway_85__EVAL),
    ._EVAL_0(LevelGateway_85__EVAL_0),
    ._EVAL_1(LevelGateway_85__EVAL_1),
    ._EVAL_2(LevelGateway_85__EVAL_2),
    ._EVAL_3(LevelGateway_85__EVAL_3),
    ._EVAL_4(LevelGateway_85__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_46 (
    ._EVAL(LevelGateway_46__EVAL),
    ._EVAL_0(LevelGateway_46__EVAL_0),
    ._EVAL_1(LevelGateway_46__EVAL_1),
    ._EVAL_2(LevelGateway_46__EVAL_2),
    ._EVAL_3(LevelGateway_46__EVAL_3),
    ._EVAL_4(LevelGateway_46__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_60 (
    ._EVAL(LevelGateway_60__EVAL),
    ._EVAL_0(LevelGateway_60__EVAL_0),
    ._EVAL_1(LevelGateway_60__EVAL_1),
    ._EVAL_2(LevelGateway_60__EVAL_2),
    ._EVAL_3(LevelGateway_60__EVAL_3),
    ._EVAL_4(LevelGateway_60__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_20 (
    ._EVAL(LevelGateway_20__EVAL),
    ._EVAL_0(LevelGateway_20__EVAL_0),
    ._EVAL_1(LevelGateway_20__EVAL_1),
    ._EVAL_2(LevelGateway_20__EVAL_2),
    ._EVAL_3(LevelGateway_20__EVAL_3),
    ._EVAL_4(LevelGateway_20__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_17 (
    ._EVAL(LevelGateway_17__EVAL),
    ._EVAL_0(LevelGateway_17__EVAL_0),
    ._EVAL_1(LevelGateway_17__EVAL_1),
    ._EVAL_2(LevelGateway_17__EVAL_2),
    ._EVAL_3(LevelGateway_17__EVAL_3),
    ._EVAL_4(LevelGateway_17__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_59 (
    ._EVAL(LevelGateway_59__EVAL),
    ._EVAL_0(LevelGateway_59__EVAL_0),
    ._EVAL_1(LevelGateway_59__EVAL_1),
    ._EVAL_2(LevelGateway_59__EVAL_2),
    ._EVAL_3(LevelGateway_59__EVAL_3),
    ._EVAL_4(LevelGateway_59__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_124 (
    ._EVAL(LevelGateway_124__EVAL),
    ._EVAL_0(LevelGateway_124__EVAL_0),
    ._EVAL_1(LevelGateway_124__EVAL_1),
    ._EVAL_2(LevelGateway_124__EVAL_2),
    ._EVAL_3(LevelGateway_124__EVAL_3),
    ._EVAL_4(LevelGateway_124__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_61 (
    ._EVAL(LevelGateway_61__EVAL),
    ._EVAL_0(LevelGateway_61__EVAL_0),
    ._EVAL_1(LevelGateway_61__EVAL_1),
    ._EVAL_2(LevelGateway_61__EVAL_2),
    ._EVAL_3(LevelGateway_61__EVAL_3),
    ._EVAL_4(LevelGateway_61__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_2 (
    ._EVAL(LevelGateway_2__EVAL),
    ._EVAL_0(LevelGateway_2__EVAL_0),
    ._EVAL_1(LevelGateway_2__EVAL_1),
    ._EVAL_2(LevelGateway_2__EVAL_2),
    ._EVAL_3(LevelGateway_2__EVAL_3),
    ._EVAL_4(LevelGateway_2__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_40 (
    ._EVAL(LevelGateway_40__EVAL),
    ._EVAL_0(LevelGateway_40__EVAL_0),
    ._EVAL_1(LevelGateway_40__EVAL_1),
    ._EVAL_2(LevelGateway_40__EVAL_2),
    ._EVAL_3(LevelGateway_40__EVAL_3),
    ._EVAL_4(LevelGateway_40__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_33 (
    ._EVAL(LevelGateway_33__EVAL),
    ._EVAL_0(LevelGateway_33__EVAL_0),
    ._EVAL_1(LevelGateway_33__EVAL_1),
    ._EVAL_2(LevelGateway_33__EVAL_2),
    ._EVAL_3(LevelGateway_33__EVAL_3),
    ._EVAL_4(LevelGateway_33__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_21 (
    ._EVAL(LevelGateway_21__EVAL),
    ._EVAL_0(LevelGateway_21__EVAL_0),
    ._EVAL_1(LevelGateway_21__EVAL_1),
    ._EVAL_2(LevelGateway_21__EVAL_2),
    ._EVAL_3(LevelGateway_21__EVAL_3),
    ._EVAL_4(LevelGateway_21__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_26 (
    ._EVAL(LevelGateway_26__EVAL),
    ._EVAL_0(LevelGateway_26__EVAL_0),
    ._EVAL_1(LevelGateway_26__EVAL_1),
    ._EVAL_2(LevelGateway_26__EVAL_2),
    ._EVAL_3(LevelGateway_26__EVAL_3),
    ._EVAL_4(LevelGateway_26__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_110 (
    ._EVAL(LevelGateway_110__EVAL),
    ._EVAL_0(LevelGateway_110__EVAL_0),
    ._EVAL_1(LevelGateway_110__EVAL_1),
    ._EVAL_2(LevelGateway_110__EVAL_2),
    ._EVAL_3(LevelGateway_110__EVAL_3),
    ._EVAL_4(LevelGateway_110__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_90 (
    ._EVAL(LevelGateway_90__EVAL),
    ._EVAL_0(LevelGateway_90__EVAL_0),
    ._EVAL_1(LevelGateway_90__EVAL_1),
    ._EVAL_2(LevelGateway_90__EVAL_2),
    ._EVAL_3(LevelGateway_90__EVAL_3),
    ._EVAL_4(LevelGateway_90__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_119 (
    ._EVAL(LevelGateway_119__EVAL),
    ._EVAL_0(LevelGateway_119__EVAL_0),
    ._EVAL_1(LevelGateway_119__EVAL_1),
    ._EVAL_2(LevelGateway_119__EVAL_2),
    ._EVAL_3(LevelGateway_119__EVAL_3),
    ._EVAL_4(LevelGateway_119__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_23 (
    ._EVAL(LevelGateway_23__EVAL),
    ._EVAL_0(LevelGateway_23__EVAL_0),
    ._EVAL_1(LevelGateway_23__EVAL_1),
    ._EVAL_2(LevelGateway_23__EVAL_2),
    ._EVAL_3(LevelGateway_23__EVAL_3),
    ._EVAL_4(LevelGateway_23__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_80 (
    ._EVAL(LevelGateway_80__EVAL),
    ._EVAL_0(LevelGateway_80__EVAL_0),
    ._EVAL_1(LevelGateway_80__EVAL_1),
    ._EVAL_2(LevelGateway_80__EVAL_2),
    ._EVAL_3(LevelGateway_80__EVAL_3),
    ._EVAL_4(LevelGateway_80__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_41 (
    ._EVAL(LevelGateway_41__EVAL),
    ._EVAL_0(LevelGateway_41__EVAL_0),
    ._EVAL_1(LevelGateway_41__EVAL_1),
    ._EVAL_2(LevelGateway_41__EVAL_2),
    ._EVAL_3(LevelGateway_41__EVAL_3),
    ._EVAL_4(LevelGateway_41__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_78 (
    ._EVAL(LevelGateway_78__EVAL),
    ._EVAL_0(LevelGateway_78__EVAL_0),
    ._EVAL_1(LevelGateway_78__EVAL_1),
    ._EVAL_2(LevelGateway_78__EVAL_2),
    ._EVAL_3(LevelGateway_78__EVAL_3),
    ._EVAL_4(LevelGateway_78__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_121 (
    ._EVAL(LevelGateway_121__EVAL),
    ._EVAL_0(LevelGateway_121__EVAL_0),
    ._EVAL_1(LevelGateway_121__EVAL_1),
    ._EVAL_2(LevelGateway_121__EVAL_2),
    ._EVAL_3(LevelGateway_121__EVAL_3),
    ._EVAL_4(LevelGateway_121__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_31 (
    ._EVAL(LevelGateway_31__EVAL),
    ._EVAL_0(LevelGateway_31__EVAL_0),
    ._EVAL_1(LevelGateway_31__EVAL_1),
    ._EVAL_2(LevelGateway_31__EVAL_2),
    ._EVAL_3(LevelGateway_31__EVAL_3),
    ._EVAL_4(LevelGateway_31__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_19 (
    ._EVAL(LevelGateway_19__EVAL),
    ._EVAL_0(LevelGateway_19__EVAL_0),
    ._EVAL_1(LevelGateway_19__EVAL_1),
    ._EVAL_2(LevelGateway_19__EVAL_2),
    ._EVAL_3(LevelGateway_19__EVAL_3),
    ._EVAL_4(LevelGateway_19__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_113 (
    ._EVAL(LevelGateway_113__EVAL),
    ._EVAL_0(LevelGateway_113__EVAL_0),
    ._EVAL_1(LevelGateway_113__EVAL_1),
    ._EVAL_2(LevelGateway_113__EVAL_2),
    ._EVAL_3(LevelGateway_113__EVAL_3),
    ._EVAL_4(LevelGateway_113__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_111 (
    ._EVAL(LevelGateway_111__EVAL),
    ._EVAL_0(LevelGateway_111__EVAL_0),
    ._EVAL_1(LevelGateway_111__EVAL_1),
    ._EVAL_2(LevelGateway_111__EVAL_2),
    ._EVAL_3(LevelGateway_111__EVAL_3),
    ._EVAL_4(LevelGateway_111__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_77 (
    ._EVAL(LevelGateway_77__EVAL),
    ._EVAL_0(LevelGateway_77__EVAL_0),
    ._EVAL_1(LevelGateway_77__EVAL_1),
    ._EVAL_2(LevelGateway_77__EVAL_2),
    ._EVAL_3(LevelGateway_77__EVAL_3),
    ._EVAL_4(LevelGateway_77__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_11 (
    ._EVAL(LevelGateway_11__EVAL),
    ._EVAL_0(LevelGateway_11__EVAL_0),
    ._EVAL_1(LevelGateway_11__EVAL_1),
    ._EVAL_2(LevelGateway_11__EVAL_2),
    ._EVAL_3(LevelGateway_11__EVAL_3),
    ._EVAL_4(LevelGateway_11__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_36 (
    ._EVAL(LevelGateway_36__EVAL),
    ._EVAL_0(LevelGateway_36__EVAL_0),
    ._EVAL_1(LevelGateway_36__EVAL_1),
    ._EVAL_2(LevelGateway_36__EVAL_2),
    ._EVAL_3(LevelGateway_36__EVAL_3),
    ._EVAL_4(LevelGateway_36__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_24 (
    ._EVAL(LevelGateway_24__EVAL),
    ._EVAL_0(LevelGateway_24__EVAL_0),
    ._EVAL_1(LevelGateway_24__EVAL_1),
    ._EVAL_2(LevelGateway_24__EVAL_2),
    ._EVAL_3(LevelGateway_24__EVAL_3),
    ._EVAL_4(LevelGateway_24__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_125 (
    ._EVAL(LevelGateway_125__EVAL),
    ._EVAL_0(LevelGateway_125__EVAL_0),
    ._EVAL_1(LevelGateway_125__EVAL_1),
    ._EVAL_2(LevelGateway_125__EVAL_2),
    ._EVAL_3(LevelGateway_125__EVAL_3),
    ._EVAL_4(LevelGateway_125__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_45 (
    ._EVAL(LevelGateway_45__EVAL),
    ._EVAL_0(LevelGateway_45__EVAL_0),
    ._EVAL_1(LevelGateway_45__EVAL_1),
    ._EVAL_2(LevelGateway_45__EVAL_2),
    ._EVAL_3(LevelGateway_45__EVAL_3),
    ._EVAL_4(LevelGateway_45__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_106 (
    ._EVAL(LevelGateway_106__EVAL),
    ._EVAL_0(LevelGateway_106__EVAL_0),
    ._EVAL_1(LevelGateway_106__EVAL_1),
    ._EVAL_2(LevelGateway_106__EVAL_2),
    ._EVAL_3(LevelGateway_106__EVAL_3),
    ._EVAL_4(LevelGateway_106__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_8 (
    ._EVAL(LevelGateway_8__EVAL),
    ._EVAL_0(LevelGateway_8__EVAL_0),
    ._EVAL_1(LevelGateway_8__EVAL_1),
    ._EVAL_2(LevelGateway_8__EVAL_2),
    ._EVAL_3(LevelGateway_8__EVAL_3),
    ._EVAL_4(LevelGateway_8__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_1 (
    ._EVAL(LevelGateway_1__EVAL),
    ._EVAL_0(LevelGateway_1__EVAL_0),
    ._EVAL_1(LevelGateway_1__EVAL_1),
    ._EVAL_2(LevelGateway_1__EVAL_2),
    ._EVAL_3(LevelGateway_1__EVAL_3),
    ._EVAL_4(LevelGateway_1__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_52 (
    ._EVAL(LevelGateway_52__EVAL),
    ._EVAL_0(LevelGateway_52__EVAL_0),
    ._EVAL_1(LevelGateway_52__EVAL_1),
    ._EVAL_2(LevelGateway_52__EVAL_2),
    ._EVAL_3(LevelGateway_52__EVAL_3),
    ._EVAL_4(LevelGateway_52__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_87 (
    ._EVAL(LevelGateway_87__EVAL),
    ._EVAL_0(LevelGateway_87__EVAL_0),
    ._EVAL_1(LevelGateway_87__EVAL_1),
    ._EVAL_2(LevelGateway_87__EVAL_2),
    ._EVAL_3(LevelGateway_87__EVAL_3),
    ._EVAL_4(LevelGateway_87__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_74 (
    ._EVAL(LevelGateway_74__EVAL),
    ._EVAL_0(LevelGateway_74__EVAL_0),
    ._EVAL_1(LevelGateway_74__EVAL_1),
    ._EVAL_2(LevelGateway_74__EVAL_2),
    ._EVAL_3(LevelGateway_74__EVAL_3),
    ._EVAL_4(LevelGateway_74__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_18 (
    ._EVAL(LevelGateway_18__EVAL),
    ._EVAL_0(LevelGateway_18__EVAL_0),
    ._EVAL_1(LevelGateway_18__EVAL_1),
    ._EVAL_2(LevelGateway_18__EVAL_2),
    ._EVAL_3(LevelGateway_18__EVAL_3),
    ._EVAL_4(LevelGateway_18__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_22 (
    ._EVAL(LevelGateway_22__EVAL),
    ._EVAL_0(LevelGateway_22__EVAL_0),
    ._EVAL_1(LevelGateway_22__EVAL_1),
    ._EVAL_2(LevelGateway_22__EVAL_2),
    ._EVAL_3(LevelGateway_22__EVAL_3),
    ._EVAL_4(LevelGateway_22__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_51 (
    ._EVAL(LevelGateway_51__EVAL),
    ._EVAL_0(LevelGateway_51__EVAL_0),
    ._EVAL_1(LevelGateway_51__EVAL_1),
    ._EVAL_2(LevelGateway_51__EVAL_2),
    ._EVAL_3(LevelGateway_51__EVAL_3),
    ._EVAL_4(LevelGateway_51__EVAL_4)
  );
  SiFive__EVAL_182 LevelGateway_32 (
    ._EVAL(LevelGateway_32__EVAL),
    ._EVAL_0(LevelGateway_32__EVAL_0),
    ._EVAL_1(LevelGateway_32__EVAL_1),
    ._EVAL_2(LevelGateway_32__EVAL_2),
    ._EVAL_3(LevelGateway_32__EVAL_3),
    ._EVAL_4(LevelGateway_32__EVAL_4)
  );
  assign _EVAL_910 = _EVAL_51[27:2];
  assign _EVAL_2134 = Queue__EVAL_12 & _EVAL_59;
  assign _EVAL_1716 = Queue__EVAL_13 == 1'h0;
  assign _EVAL_3673 = _EVAL_2134 & _EVAL_1716;
  assign _EVAL_1141 = Queue__EVAL_6[19];
  assign _EVAL_2526 = Queue__EVAL_6[11];
  assign _EVAL_2033 = Queue__EVAL_6[10];
  assign _EVAL_2718 = Queue__EVAL_6[6];
  assign _EVAL_2486 = Queue__EVAL_6[5];
  assign _EVAL_640 = Queue__EVAL_6[4];
  assign _EVAL_3992 = Queue__EVAL_6[3];
  assign _EVAL_397 = Queue__EVAL_6[2];
  assign _EVAL_2460 = Queue__EVAL_6[1];
  assign _EVAL_3606 = Queue__EVAL_6[0];
  assign _EVAL_1450 = {_EVAL_1141,_EVAL_2526,_EVAL_2033,_EVAL_2718,_EVAL_2486,_EVAL_640,_EVAL_3992,_EVAL_397,_EVAL_2460,_EVAL_3606};
  assign _EVAL_2999 = 1024'h1 << _EVAL_1450;
  assign _EVAL_2866 = _EVAL_2999[21];
  assign _EVAL_3344 = _EVAL_3673 & _EVAL_2866;
  assign _EVAL_3888 = Queue__EVAL_6 & 24'hf7f380;
  assign _EVAL_2267 = _EVAL_3888 == 24'h0;
  assign _EVAL_1644 = _EVAL_3344 & _EVAL_2267;
  assign _EVAL_915 = Queue__EVAL_10[3];
  assign _EVAL_287 = _EVAL_915 ? 8'hff : 8'h0;
  assign _EVAL_2436 = Queue__EVAL_10[2];
  assign _EVAL_3655 = _EVAL_2436 ? 8'hff : 8'h0;
  assign _EVAL_4053 = Queue__EVAL_10[1];
  assign _EVAL_2619 = _EVAL_4053 ? 8'hff : 8'h0;
  assign _EVAL_1637 = Queue__EVAL_10[0];
  assign _EVAL_352 = _EVAL_1637 ? 8'hff : 8'h0;
  assign _EVAL_2124 = {_EVAL_287,_EVAL_3655,_EVAL_2619,_EVAL_352};
  assign _EVAL_3165 = _EVAL_2124[2:0];
  assign _EVAL_591 = _EVAL_3165 == 3'h7;
  assign _EVAL_532 = _EVAL_1644 & _EVAL_591;
  assign _EVAL_886 = _EVAL_2999[97];
  assign _EVAL_3851 = _EVAL_3673 & _EVAL_886;
  assign _EVAL_3050 = _EVAL_3851 & _EVAL_2267;
  assign _EVAL_1440 = 10'h34 == _EVAL_1450;
  assign _EVAL_3081 = 10'h35 == _EVAL_1450;
  assign _EVAL_4052 = 10'h36 == _EVAL_1450;
  assign _EVAL_2575 = 10'h37 == _EVAL_1450;
  assign _EVAL_964 = 10'h38 == _EVAL_1450;
  assign _EVAL_2656 = 10'h39 == _EVAL_1450;
  assign _EVAL_3526 = 10'h3a == _EVAL_1450;
  assign _EVAL_3146 = 10'h3b == _EVAL_1450;
  assign _EVAL_1023 = 10'h3c == _EVAL_1450;
  assign _EVAL_3602 = 10'h3d == _EVAL_1450;
  assign _EVAL_2966 = 10'h3e == _EVAL_1450;
  assign _EVAL_742 = 10'h3f == _EVAL_1450;
  assign _EVAL_1018 = 10'h40 == _EVAL_1450;
  assign _EVAL_3758 = 10'h41 == _EVAL_1450;
  assign _EVAL_368 = 10'h42 == _EVAL_1450;
  assign _EVAL_1362 = 10'h43 == _EVAL_1450;
  assign _EVAL_870 = 10'h44 == _EVAL_1450;
  assign _EVAL_2716 = 10'h45 == _EVAL_1450;
  assign _EVAL_3097 = 10'h46 == _EVAL_1450;
  assign _EVAL_841 = 10'h47 == _EVAL_1450;
  assign _EVAL_3044 = 10'h48 == _EVAL_1450;
  assign _EVAL_3226 = 10'h49 == _EVAL_1450;
  assign _EVAL_584 = 10'h4a == _EVAL_1450;
  assign _EVAL_3400 = 10'h4b == _EVAL_1450;
  assign _EVAL_1014 = 10'h4c == _EVAL_1450;
  assign _EVAL_1838 = 10'h4d == _EVAL_1450;
  assign _EVAL_1891 = 10'h4e == _EVAL_1450;
  assign _EVAL_907 = 10'h4f == _EVAL_1450;
  assign _EVAL_1425 = 10'h50 == _EVAL_1450;
  assign _EVAL_1185 = 10'h51 == _EVAL_1450;
  assign _EVAL_1489 = 10'h52 == _EVAL_1450;
  assign _EVAL_2265 = 10'h53 == _EVAL_1450;
  assign _EVAL_3179 = 10'h54 == _EVAL_1450;
  assign _EVAL_2269 = 10'h55 == _EVAL_1450;
  assign _EVAL_922 = 10'h56 == _EVAL_1450;
  assign _EVAL_1991 = 10'h57 == _EVAL_1450;
  assign _EVAL_2441 = 10'h58 == _EVAL_1450;
  assign _EVAL_3002 = 10'h59 == _EVAL_1450;
  assign _EVAL_350 = 10'h5a == _EVAL_1450;
  assign _EVAL_3718 = 10'h5b == _EVAL_1450;
  assign _EVAL_443 = 10'h5c == _EVAL_1450;
  assign _EVAL_2448 = 10'h5d == _EVAL_1450;
  assign _EVAL_2777 = 10'h5e == _EVAL_1450;
  assign _EVAL_2361 = 10'h5f == _EVAL_1450;
  assign _EVAL_373 = 10'h60 == _EVAL_1450;
  assign _EVAL_3550 = 10'h61 == _EVAL_1450;
  assign _EVAL_2496 = 10'h62 == _EVAL_1450;
  assign _EVAL_2308 = 10'h63 == _EVAL_1450;
  assign _EVAL_1421 = 10'h64 == _EVAL_1450;
  assign _EVAL_3500 = 10'h65 == _EVAL_1450;
  assign _EVAL_1163 = 10'h66 == _EVAL_1450;
  assign _EVAL_700 = 10'h67 == _EVAL_1450;
  assign _EVAL_1301 = 10'h68 == _EVAL_1450;
  assign _EVAL_4011 = 10'h69 == _EVAL_1450;
  assign _EVAL_942 = 10'h6a == _EVAL_1450;
  assign _EVAL_3177 = 10'h6b == _EVAL_1450;
  assign _EVAL_1859 = 10'h6c == _EVAL_1450;
  assign _EVAL_1672 = 10'h6d == _EVAL_1450;
  assign _EVAL_2434 = 10'h6e == _EVAL_1450;
  assign _EVAL_2841 = 10'h6f == _EVAL_1450;
  assign _EVAL_3802 = 10'h70 == _EVAL_1450;
  assign _EVAL_3883 = 10'h71 == _EVAL_1450;
  assign _EVAL_1080 = 10'h72 == _EVAL_1450;
  assign _EVAL_2192 = 10'h73 == _EVAL_1450;
  assign _EVAL_2510 = 10'h74 == _EVAL_1450;
  assign _EVAL_2970 = 10'h75 == _EVAL_1450;
  assign _EVAL_165 = 10'h76 == _EVAL_1450;
  assign _EVAL_2863 = 10'h77 == _EVAL_1450;
  assign _EVAL_3127 = 10'h78 == _EVAL_1450;
  assign _EVAL_3494 = 10'h79 == _EVAL_1450;
  assign _EVAL_3590 = 10'h7a == _EVAL_1450;
  assign _EVAL_1282 = 10'h7b == _EVAL_1450;
  assign _EVAL_3839 = 10'h7c == _EVAL_1450;
  assign _EVAL_2801 = 10'h7d == _EVAL_1450;
  assign _EVAL_2771 = 10'h7e == _EVAL_1450;
  assign _EVAL_711 = 10'h7f == _EVAL_1450;
  assign _EVAL_1939 = 10'h80 == _EVAL_1450;
  assign _EVAL_159 = 10'h81 == _EVAL_1450;
  assign _EVAL_1321 = 10'h82 == _EVAL_1450;
  assign _EVAL_1987 = 10'h83 == _EVAL_1450;
  assign _EVAL_1387 = 10'h100 == _EVAL_1450;
  assign _EVAL_3800 = 10'h101 == _EVAL_1450;
  assign _EVAL_1198 = 10'h102 == _EVAL_1450;
  assign _EVAL_1713 = 10'h103 == _EVAL_1450;
  assign _EVAL_1366 = 10'h200 == _EVAL_1450;
  assign _EVAL_2153 = 10'h201 == _EVAL_1450;
  assign _EVAL_2347 = _EVAL_2153 ? _EVAL_2267 : 1'h1;
  assign _EVAL_3428 = _EVAL_1366 ? _EVAL_2267 : _EVAL_2347;
  assign _EVAL_562 = _EVAL_1713 ? _EVAL_2267 : _EVAL_3428;
  assign _EVAL_529 = _EVAL_1198 ? _EVAL_2267 : _EVAL_562;
  assign _EVAL_3072 = _EVAL_3800 ? _EVAL_2267 : _EVAL_529;
  assign _EVAL_1583 = _EVAL_1387 ? _EVAL_2267 : _EVAL_3072;
  assign _EVAL_854 = _EVAL_1987 ? _EVAL_2267 : _EVAL_1583;
  assign _EVAL_3382 = _EVAL_1321 ? _EVAL_2267 : _EVAL_854;
  assign _EVAL_249 = _EVAL_159 ? _EVAL_2267 : _EVAL_3382;
  assign _EVAL_775 = _EVAL_1939 ? _EVAL_2267 : _EVAL_249;
  assign _EVAL_1108 = _EVAL_711 ? _EVAL_2267 : _EVAL_775;
  assign _EVAL_1059 = _EVAL_2771 ? _EVAL_2267 : _EVAL_1108;
  assign _EVAL_1779 = _EVAL_2801 ? _EVAL_2267 : _EVAL_1059;
  assign _EVAL_3523 = _EVAL_3839 ? _EVAL_2267 : _EVAL_1779;
  assign _EVAL_2314 = _EVAL_1282 ? _EVAL_2267 : _EVAL_3523;
  assign _EVAL_988 = _EVAL_3590 ? _EVAL_2267 : _EVAL_2314;
  assign _EVAL_1167 = _EVAL_3494 ? _EVAL_2267 : _EVAL_988;
  assign _EVAL_2633 = _EVAL_3127 ? _EVAL_2267 : _EVAL_1167;
  assign _EVAL_277 = _EVAL_2863 ? _EVAL_2267 : _EVAL_2633;
  assign _EVAL_652 = _EVAL_165 ? _EVAL_2267 : _EVAL_277;
  assign _EVAL_2989 = _EVAL_2970 ? _EVAL_2267 : _EVAL_652;
  assign _EVAL_878 = _EVAL_2510 ? _EVAL_2267 : _EVAL_2989;
  assign _EVAL_888 = _EVAL_2192 ? _EVAL_2267 : _EVAL_878;
  assign _EVAL_4025 = _EVAL_1080 ? _EVAL_2267 : _EVAL_888;
  assign _EVAL_2868 = _EVAL_3883 ? _EVAL_2267 : _EVAL_4025;
  assign _EVAL_3605 = _EVAL_3802 ? _EVAL_2267 : _EVAL_2868;
  assign _EVAL_1594 = _EVAL_2841 ? _EVAL_2267 : _EVAL_3605;
  assign _EVAL_459 = _EVAL_2434 ? _EVAL_2267 : _EVAL_1594;
  assign _EVAL_1170 = _EVAL_1672 ? _EVAL_2267 : _EVAL_459;
  assign _EVAL_1189 = _EVAL_1859 ? _EVAL_2267 : _EVAL_1170;
  assign _EVAL_1565 = _EVAL_3177 ? _EVAL_2267 : _EVAL_1189;
  assign _EVAL_3941 = _EVAL_942 ? _EVAL_2267 : _EVAL_1565;
  assign _EVAL_3866 = _EVAL_4011 ? _EVAL_2267 : _EVAL_3941;
  assign _EVAL_1810 = _EVAL_1301 ? _EVAL_2267 : _EVAL_3866;
  assign _EVAL_3232 = _EVAL_700 ? _EVAL_2267 : _EVAL_1810;
  assign _EVAL_1318 = _EVAL_1163 ? _EVAL_2267 : _EVAL_3232;
  assign _EVAL_4015 = _EVAL_3500 ? _EVAL_2267 : _EVAL_1318;
  assign _EVAL_1849 = _EVAL_1421 ? _EVAL_2267 : _EVAL_4015;
  assign _EVAL_3174 = _EVAL_2308 ? _EVAL_2267 : _EVAL_1849;
  assign _EVAL_945 = _EVAL_2496 ? _EVAL_2267 : _EVAL_3174;
  assign _EVAL_559 = _EVAL_3550 ? _EVAL_2267 : _EVAL_945;
  assign _EVAL_148 = _EVAL_373 ? _EVAL_2267 : _EVAL_559;
  assign _EVAL_1736 = _EVAL_2361 ? _EVAL_2267 : _EVAL_148;
  assign _EVAL_1173 = _EVAL_2777 ? _EVAL_2267 : _EVAL_1736;
  assign _EVAL_684 = _EVAL_2448 ? _EVAL_2267 : _EVAL_1173;
  assign _EVAL_2318 = _EVAL_443 ? _EVAL_2267 : _EVAL_684;
  assign _EVAL_2220 = _EVAL_3718 ? _EVAL_2267 : _EVAL_2318;
  assign _EVAL_491 = _EVAL_350 ? _EVAL_2267 : _EVAL_2220;
  assign _EVAL_3412 = _EVAL_3002 ? _EVAL_2267 : _EVAL_491;
  assign _EVAL_1292 = _EVAL_2441 ? _EVAL_2267 : _EVAL_3412;
  assign _EVAL_1483 = _EVAL_1991 ? _EVAL_2267 : _EVAL_1292;
  assign _EVAL_3556 = _EVAL_922 ? _EVAL_2267 : _EVAL_1483;
  assign _EVAL_1574 = _EVAL_2269 ? _EVAL_2267 : _EVAL_3556;
  assign _EVAL_3828 = _EVAL_3179 ? _EVAL_2267 : _EVAL_1574;
  assign _EVAL_517 = _EVAL_2265 ? _EVAL_2267 : _EVAL_3828;
  assign _EVAL_583 = _EVAL_1489 ? _EVAL_2267 : _EVAL_517;
  assign _EVAL_3125 = _EVAL_1185 ? _EVAL_2267 : _EVAL_583;
  assign _EVAL_3995 = _EVAL_1425 ? _EVAL_2267 : _EVAL_3125;
  assign _EVAL_2670 = _EVAL_907 ? _EVAL_2267 : _EVAL_3995;
  assign _EVAL_3247 = _EVAL_1891 ? _EVAL_2267 : _EVAL_2670;
  assign _EVAL_2299 = _EVAL_1838 ? _EVAL_2267 : _EVAL_3247;
  assign _EVAL_3811 = _EVAL_1014 ? _EVAL_2267 : _EVAL_2299;
  assign _EVAL_1231 = _EVAL_3400 ? _EVAL_2267 : _EVAL_3811;
  assign _EVAL_3722 = _EVAL_584 ? _EVAL_2267 : _EVAL_1231;
  assign _EVAL_3109 = _EVAL_3226 ? _EVAL_2267 : _EVAL_3722;
  assign _EVAL_2435 = _EVAL_3044 ? _EVAL_2267 : _EVAL_3109;
  assign _EVAL_4021 = _EVAL_841 ? _EVAL_2267 : _EVAL_2435;
  assign _EVAL_2781 = _EVAL_3097 ? _EVAL_2267 : _EVAL_4021;
  assign _EVAL_2088 = _EVAL_2716 ? _EVAL_2267 : _EVAL_2781;
  assign _EVAL_2440 = _EVAL_870 ? _EVAL_2267 : _EVAL_2088;
  assign _EVAL_1418 = _EVAL_1362 ? _EVAL_2267 : _EVAL_2440;
  assign _EVAL_2832 = _EVAL_368 ? _EVAL_2267 : _EVAL_1418;
  assign _EVAL_3042 = _EVAL_3758 ? _EVAL_2267 : _EVAL_2832;
  assign _EVAL_537 = _EVAL_1018 ? _EVAL_2267 : _EVAL_3042;
  assign _EVAL_898 = _EVAL_742 ? _EVAL_2267 : _EVAL_537;
  assign _EVAL_1727 = _EVAL_2966 ? _EVAL_2267 : _EVAL_898;
  assign _EVAL_1734 = _EVAL_3602 ? _EVAL_2267 : _EVAL_1727;
  assign _EVAL_3172 = _EVAL_1023 ? _EVAL_2267 : _EVAL_1734;
  assign _EVAL_460 = _EVAL_3146 ? _EVAL_2267 : _EVAL_3172;
  assign _EVAL_1407 = _EVAL_3526 ? _EVAL_2267 : _EVAL_460;
  assign _EVAL_3147 = _EVAL_2656 ? _EVAL_2267 : _EVAL_1407;
  assign _EVAL_2451 = _EVAL_964 ? _EVAL_2267 : _EVAL_3147;
  assign _EVAL_3841 = _EVAL_2575 ? _EVAL_2267 : _EVAL_2451;
  assign _EVAL_2847 = _EVAL_4052 ? _EVAL_2267 : _EVAL_3841;
  assign _EVAL_1777 = _EVAL_3081 ? _EVAL_2267 : _EVAL_2847;
  assign _EVAL_2790 = _EVAL_1440 ? _EVAL_2267 : _EVAL_1777;
  assign _EVAL_2234 = _EVAL_2999[83];
  assign _EVAL_1676 = _EVAL_3673 & _EVAL_2234;
  assign _EVAL_626 = _EVAL_1676 & _EVAL_2267;
  assign _EVAL_3059 = _EVAL_2134 & Queue__EVAL_13;
  assign _EVAL_2184 = _EVAL_2999[6];
  assign _EVAL_429 = _EVAL_2999[39];
  assign _EVAL_390 = _EVAL_2999[513];
  assign _EVAL_2158 = _EVAL_3059 & _EVAL_390;
  assign _EVAL_826 = _EVAL_2158 & _EVAL_2267;
  assign _EVAL_2107 = _EVAL_2124 != 32'h0;
  assign _EVAL_1847 = _EVAL_826 & _EVAL_2107;
  assign _EVAL_2616 = _EVAL_1847 ? _EVAL_3235 : 7'h0;
  assign _EVAL_1635 = 128'h1 << _EVAL_2616;
  assign _EVAL_1805 = _EVAL_1635[46];
  assign _EVAL_1077 = _EVAL_1805 | LevelGateway_45__EVAL_3;
  assign _EVAL_1531 = _EVAL_2999[512];
  assign _EVAL_1886 = _EVAL_2999[103];
  assign _EVAL_378 = _EVAL_1635[18];
  assign _EVAL_4026 = _EVAL_378 == 1'h0;
  assign _EVAL_3215 = _EVAL_2999[126];
  assign _EVAL_2232 = _EVAL_3673 & _EVAL_3215;
  assign _EVAL_632 = _EVAL_2232 & _EVAL_2267;
  assign _EVAL_3688 = _EVAL_1635[88];
  assign _EVAL_2917 = _EVAL_3688 == 1'h0;
  assign _EVAL_3878 = {_EVAL_200,_EVAL_2807,_EVAL_1788,_EVAL_3759,_EVAL_163,_EVAL_2826,_EVAL_371,_EVAL_2209,_EVAL_2133,1'h0};
  assign _EVAL_3760 = {_EVAL_269,_EVAL_2128,_EVAL_581,_EVAL_1556,_EVAL_1121,_EVAL_3636,_EVAL_3750,_EVAL_1979,_EVAL_673,_EVAL_3878};
  assign _EVAL_618 = {_EVAL_448,_EVAL_387,_EVAL_306,_EVAL_614,_EVAL_2214,_EVAL_217,_EVAL_1708,_EVAL_3192,_EVAL_2666,_EVAL_3760};
  assign _EVAL_2860 = {_EVAL_3222,_EVAL_1597,_EVAL_3317,_EVAL_3505,_EVAL_618};
  assign _EVAL_716 = {_EVAL_3407,_EVAL_1929,_EVAL_989,_EVAL_2684,_EVAL_427,_EVAL_1456,_EVAL_492,_EVAL_1315,_EVAL_462,_EVAL_2507};
  assign _EVAL_2797 = {_EVAL_3720,_EVAL_222,_EVAL_2485,_EVAL_1709,_EVAL_3715,_EVAL_3025,_EVAL_690,_EVAL_3899,_EVAL_2155,_EVAL_716};
  assign _EVAL_2226 = {_EVAL_3137,_EVAL_1206,_EVAL_3527,_EVAL_2254,_EVAL_2688,_EVAL_2582,_EVAL_2803,_EVAL_2050,_EVAL_1313,_EVAL_2797};
  assign _EVAL_1293 = {_EVAL_1073,_EVAL_2870,_EVAL_2341,_EVAL_2648,_EVAL_2226};
  assign _EVAL_1590 = {_EVAL_497,_EVAL_3039,_EVAL_552,_EVAL_3023,_EVAL_2701,_EVAL_421,_EVAL_3359,_EVAL_4034,_EVAL_947,_EVAL_1587};
  assign _EVAL_3587 = {_EVAL_3299,_EVAL_1536,_EVAL_1580,_EVAL_2850,_EVAL_880,_EVAL_212,_EVAL_1930,_EVAL_3361,_EVAL_2159,_EVAL_1590};
  assign _EVAL_267 = {_EVAL_3757,_EVAL_3996,_EVAL_1270,_EVAL_2972,_EVAL_2809,_EVAL_3245,_EVAL_3551,_EVAL_3728,_EVAL_1261,_EVAL_3587};
  assign _EVAL_521 = {_EVAL_2953,_EVAL_3788,_EVAL_3783,_EVAL_3279,_EVAL_267};
  assign _EVAL_760 = {_EVAL_3199,_EVAL_3964,_EVAL_194,_EVAL_3283,_EVAL_912,_EVAL_3296,_EVAL_770,_EVAL_2838,_EVAL_730,_EVAL_1521};
  assign _EVAL_1227 = {_EVAL_1917,_EVAL_480,_EVAL_1496,_EVAL_715,_EVAL_1267,_EVAL_176,_EVAL_2942,_EVAL_3419,_EVAL_569,_EVAL_760};
  assign _EVAL_1511 = {_EVAL_1599,_EVAL_2938,_EVAL_741,_EVAL_2202,_EVAL_4063,_EVAL_519,_EVAL_1938,_EVAL_3167,_EVAL_1753,_EVAL_1227};
  assign _EVAL_1721 = {_EVAL_3713,_EVAL_3850,_EVAL_449,_EVAL_1471,_EVAL_1511};
  assign _EVAL_2362 = {_EVAL_3743,_EVAL_3421,_EVAL_1639,_EVAL_1698,1'h0};
  assign _EVAL_3259 = {_EVAL_366,_EVAL_3870,_EVAL_3913,_EVAL_3488};
  assign _EVAL_3026 = {_EVAL_1776,_EVAL_2754,_EVAL_2073,_EVAL_1162};
  assign _EVAL_4029 = {_EVAL_3623,_EVAL_1697,_EVAL_2188,_EVAL_2018};
  assign _EVAL_1970 = {1'h0,_EVAL_663};
  assign _EVAL_1286 = {{28'd0}, _EVAL_1970};
  assign _EVAL_1710 = {{25'd0}, _EVAL_3235};
  assign _EVAL_197 = _EVAL_2153 ? _EVAL_1710 : 32'h0;
  assign _EVAL_837 = _EVAL_1366 ? _EVAL_1286 : _EVAL_197;
  assign _EVAL_2355 = _EVAL_1713 ? _EVAL_4029 : _EVAL_837;
  assign _EVAL_2915 = _EVAL_1198 ? _EVAL_3026 : _EVAL_2355;
  assign _EVAL_3944 = _EVAL_3800 ? _EVAL_3259 : _EVAL_2915;
  assign _EVAL_334 = _EVAL_1387 ? _EVAL_2362 : _EVAL_3944;
  assign _EVAL_3837 = _EVAL_1987 ? _EVAL_1721 : _EVAL_334;
  assign _EVAL_2623 = _EVAL_1321 ? _EVAL_521 : _EVAL_3837;
  assign _EVAL_1750 = _EVAL_159 ? _EVAL_1293 : _EVAL_2623;
  assign _EVAL_2612 = _EVAL_1939 ? _EVAL_2860 : _EVAL_1750;
  assign _EVAL_1305 = _EVAL_711 ? {{29'd0}, _EVAL_3909} : _EVAL_2612;
  assign _EVAL_923 = _EVAL_2771 ? {{29'd0}, _EVAL_2334} : _EVAL_1305;
  assign _EVAL_2975 = _EVAL_2801 ? {{29'd0}, _EVAL_3591} : _EVAL_923;
  assign _EVAL_1114 = _EVAL_3839 ? {{29'd0}, _EVAL_1962} : _EVAL_2975;
  assign _EVAL_2025 = _EVAL_1282 ? {{29'd0}, _EVAL_1980} : _EVAL_1114;
  assign _EVAL_423 = _EVAL_3590 ? {{29'd0}, _EVAL_3204} : _EVAL_2025;
  assign _EVAL_1943 = _EVAL_3494 ? {{29'd0}, _EVAL_1351} : _EVAL_423;
  assign _EVAL_2968 = _EVAL_3127 ? {{29'd0}, _EVAL_648} : _EVAL_1943;
  assign _EVAL_2113 = _EVAL_2863 ? {{29'd0}, _EVAL_2290} : _EVAL_2968;
  assign _EVAL_1430 = _EVAL_165 ? {{29'd0}, _EVAL_3195} : _EVAL_2113;
  assign _EVAL_3957 = _EVAL_2970 ? {{29'd0}, _EVAL_188} : _EVAL_1430;
  assign _EVAL_2094 = _EVAL_2510 ? {{29'd0}, _EVAL_3118} : _EVAL_3957;
  assign _EVAL_1380 = _EVAL_2192 ? {{29'd0}, _EVAL_2306} : _EVAL_2094;
  assign _EVAL_1608 = _EVAL_1080 ? {{29'd0}, _EVAL_147} : _EVAL_1380;
  assign _EVAL_2749 = _EVAL_3883 ? {{29'd0}, _EVAL_1088} : _EVAL_1608;
  assign _EVAL_2190 = _EVAL_3802 ? {{29'd0}, _EVAL_2881} : _EVAL_2749;
  assign _EVAL_1804 = _EVAL_2841 ? {{29'd0}, _EVAL_1266} : _EVAL_2190;
  assign _EVAL_3219 = _EVAL_2434 ? {{29'd0}, _EVAL_3804} : _EVAL_1804;
  assign _EVAL_325 = _EVAL_1672 ? {{29'd0}, _EVAL_3943} : _EVAL_3219;
  assign _EVAL_2281 = _EVAL_1859 ? {{29'd0}, _EVAL_675} : _EVAL_325;
  assign _EVAL_811 = _EVAL_3177 ? {{29'd0}, _EVAL_2336} : _EVAL_2281;
  assign _EVAL_3627 = _EVAL_942 ? {{29'd0}, _EVAL_1239} : _EVAL_811;
  assign _EVAL_1273 = _EVAL_4011 ? {{29'd0}, _EVAL_2481} : _EVAL_3627;
  assign _EVAL_3301 = _EVAL_1301 ? {{29'd0}, _EVAL_2677} : _EVAL_1273;
  assign _EVAL_2502 = _EVAL_700 ? {{29'd0}, _EVAL_3645} : _EVAL_3301;
  assign _EVAL_3017 = _EVAL_1163 ? {{29'd0}, _EVAL_3267} : _EVAL_2502;
  assign _EVAL_1625 = _EVAL_3500 ? {{29'd0}, _EVAL_902} : _EVAL_3017;
  assign _EVAL_1722 = _EVAL_1421 ? {{29'd0}, _EVAL_2111} : _EVAL_1625;
  assign _EVAL_3466 = _EVAL_2308 ? {{29'd0}, _EVAL_3733} : _EVAL_1722;
  assign _EVAL_276 = _EVAL_2496 ? {{29'd0}, _EVAL_1168} : _EVAL_3466;
  assign _EVAL_2561 = _EVAL_3550 ? {{29'd0}, _EVAL_3242} : _EVAL_276;
  assign _EVAL_2882 = _EVAL_373 ? {{29'd0}, _EVAL_3731} : _EVAL_2561;
  assign _EVAL_389 = _EVAL_2361 ? {{29'd0}, _EVAL_768} : _EVAL_2882;
  assign _EVAL_3540 = _EVAL_2777 ? {{29'd0}, _EVAL_2055} : _EVAL_389;
  assign _EVAL_2090 = _EVAL_2448 ? {{29'd0}, _EVAL_410} : _EVAL_3540;
  assign _EVAL_2065 = _EVAL_443 ? {{29'd0}, _EVAL_1738} : _EVAL_2090;
  assign _EVAL_2982 = _EVAL_3718 ? {{29'd0}, _EVAL_2646} : _EVAL_2065;
  assign _EVAL_1402 = _EVAL_350 ? {{29'd0}, _EVAL_1151} : _EVAL_2982;
  assign _EVAL_1339 = _EVAL_3002 ? {{29'd0}, _EVAL_1660} : _EVAL_1402;
  assign _EVAL_2531 = _EVAL_2441 ? {{29'd0}, _EVAL_331} : _EVAL_1339;
  assign _EVAL_1752 = _EVAL_1991 ? {{29'd0}, _EVAL_1819} : _EVAL_2531;
  assign _EVAL_3815 = _EVAL_922 ? {{29'd0}, _EVAL_1127} : _EVAL_1752;
  assign _EVAL_2853 = _EVAL_2269 ? {{29'd0}, _EVAL_485} : _EVAL_3815;
  assign _EVAL_2100 = _EVAL_3179 ? {{29'd0}, _EVAL_765} : _EVAL_2853;
  assign _EVAL_2081 = _EVAL_2265 ? {{29'd0}, _EVAL_3315} : _EVAL_2100;
  assign _EVAL_1774 = _EVAL_1489 ? {{29'd0}, _EVAL_3768} : _EVAL_2081;
  assign _EVAL_1795 = _EVAL_1185 ? {{29'd0}, _EVAL_3801} : _EVAL_1774;
  assign _EVAL_3798 = _EVAL_1425 ? {{29'd0}, _EVAL_2256} : _EVAL_1795;
  assign _EVAL_940 = _EVAL_907 ? {{29'd0}, _EVAL_2356} : _EVAL_3798;
  assign _EVAL_1137 = _EVAL_1891 ? {{29'd0}, _EVAL_1212} : _EVAL_940;
  assign _EVAL_709 = _EVAL_1838 ? {{29'd0}, _EVAL_3331} : _EVAL_1137;
  assign _EVAL_2802 = _EVAL_1014 ? {{29'd0}, _EVAL_3552} : _EVAL_709;
  assign _EVAL_2141 = _EVAL_3400 ? {{29'd0}, _EVAL_3336} : _EVAL_2802;
  assign _EVAL_409 = _EVAL_584 ? {{29'd0}, _EVAL_2720} : _EVAL_2141;
  assign _EVAL_794 = _EVAL_3226 ? {{29'd0}, _EVAL_1390} : _EVAL_409;
  assign _EVAL_891 = _EVAL_3044 ? {{29'd0}, _EVAL_3312} : _EVAL_794;
  assign _EVAL_3950 = _EVAL_841 ? {{29'd0}, _EVAL_548} : _EVAL_891;
  assign _EVAL_3928 = _EVAL_3097 ? {{29'd0}, _EVAL_1680} : _EVAL_3950;
  assign _EVAL_1186 = _EVAL_2716 ? {{29'd0}, _EVAL_3563} : _EVAL_3928;
  assign _EVAL_2119 = _EVAL_870 ? {{29'd0}, _EVAL_757} : _EVAL_1186;
  assign _EVAL_218 = _EVAL_1362 ? {{29'd0}, _EVAL_1526} : _EVAL_2119;
  assign _EVAL_1934 = _EVAL_368 ? {{29'd0}, _EVAL_835} : _EVAL_218;
  assign _EVAL_1466 = _EVAL_3758 ? {{29'd0}, _EVAL_2035} : _EVAL_1934;
  assign _EVAL_3867 = _EVAL_1018 ? {{29'd0}, _EVAL_1253} : _EVAL_1466;
  assign _EVAL_2389 = _EVAL_742 ? {{29'd0}, _EVAL_3056} : _EVAL_3867;
  assign _EVAL_836 = _EVAL_2966 ? {{29'd0}, _EVAL_2231} : _EVAL_2389;
  assign _EVAL_2092 = _EVAL_3602 ? {{29'd0}, _EVAL_1365} : _EVAL_836;
  assign _EVAL_1448 = _EVAL_1023 ? {{29'd0}, _EVAL_1176} : _EVAL_2092;
  assign _EVAL_2026 = _EVAL_3146 ? {{29'd0}, _EVAL_1280} : _EVAL_1448;
  assign _EVAL_2912 = _EVAL_3526 ? {{29'd0}, _EVAL_2584} : _EVAL_2026;
  assign _EVAL_3030 = _EVAL_2656 ? {{29'd0}, _EVAL_3644} : _EVAL_2912;
  assign _EVAL_2766 = _EVAL_964 ? {{29'd0}, _EVAL_2500} : _EVAL_3030;
  assign _EVAL_1578 = _EVAL_2575 ? {{29'd0}, _EVAL_2958} : _EVAL_2766;
  assign _EVAL_585 = _EVAL_1635[29];
  assign _EVAL_3586 = _EVAL_585 | LevelGateway_28__EVAL_3;
  assign _EVAL_1487 = _EVAL_3673 & _EVAL_390;
  assign _EVAL_1626 = _EVAL_1635[85];
  assign _EVAL_2628 = _EVAL_1626 == 1'h0;
  assign _EVAL_294 = _EVAL_1635[49];
  assign _EVAL_2578 = _EVAL_294 | LevelGateway_48__EVAL_3;
  assign _EVAL_2956 = _EVAL_294 == 1'h0;
  assign _EVAL_2610 = _EVAL_2999[47];
  assign _EVAL_3418 = _EVAL_1635[104];
  assign _EVAL_1667 = _EVAL_1487 & _EVAL_2267;
  assign _EVAL_1973 = _EVAL_2124 == 32'hffffffff;
  assign _EVAL_3593 = _EVAL_1667 & _EVAL_1973;
  assign _EVAL_1820 = _EVAL_2999[90];
  assign _EVAL_725 = _EVAL_3673 & _EVAL_1820;
  assign _EVAL_364 = _EVAL_725 & _EVAL_2267;
  assign _EVAL_3152 = _EVAL_364 & _EVAL_591;
  assign _EVAL_3617 = _EVAL_1635[51];
  assign _EVAL_2140 = _EVAL_3617 == 1'h0;
  assign _EVAL_2252 = _EVAL_2999[68];
  assign _EVAL_3504 = _EVAL_3673 & _EVAL_2252;
  assign _EVAL_318 = _EVAL_2999[96];
  assign _EVAL_3181 = _EVAL_3673 & _EVAL_318;
  assign _EVAL_3936 = _EVAL_3181 & _EVAL_2267;
  assign _EVAL_2130 = _EVAL_3936 & _EVAL_591;
  assign _EVAL_822 = _EVAL_2999[117];
  assign _EVAL_1515 = _EVAL_2999[100];
  assign _EVAL_617 = _EVAL_3673 & _EVAL_1515;
  assign _EVAL_2514 = _EVAL_617 & _EVAL_2267;
  assign _EVAL_2543 = _EVAL_2999[18];
  assign _EVAL_943 = _EVAL_3673 & _EVAL_2543;
  assign _EVAL_1852 = _EVAL_943 & _EVAL_2267;
  assign _EVAL_2057 = _EVAL_1852 & _EVAL_591;
  assign _EVAL_3820 = _EVAL_2999[26];
  assign _EVAL_3860 = _EVAL_3673 & _EVAL_3820;
  assign _EVAL_1765 = _EVAL_3860 & _EVAL_2267;
  assign _EVAL_2122 = _EVAL_2999[61];
  assign _EVAL_339 = _EVAL_1635[118];
  assign _EVAL_1416 = 10'h6 == _EVAL_1450;
  assign _EVAL_3323 = 10'h7 == _EVAL_1450;
  assign _EVAL_881 = 10'h8 == _EVAL_1450;
  assign _EVAL_4039 = 10'h9 == _EVAL_1450;
  assign _EVAL_2535 = 10'ha == _EVAL_1450;
  assign _EVAL_262 = 10'hb == _EVAL_1450;
  assign _EVAL_1055 = 10'hc == _EVAL_1450;
  assign _EVAL_2625 = 10'hd == _EVAL_1450;
  assign _EVAL_3159 = 10'he == _EVAL_1450;
  assign _EVAL_3233 = 10'hf == _EVAL_1450;
  assign _EVAL_1572 = 10'h10 == _EVAL_1450;
  assign _EVAL_3358 = 10'h11 == _EVAL_1450;
  assign _EVAL_237 = 10'h12 == _EVAL_1450;
  assign _EVAL_472 = 10'h13 == _EVAL_1450;
  assign _EVAL_2003 = 10'h14 == _EVAL_1450;
  assign _EVAL_2007 = 10'h15 == _EVAL_1450;
  assign _EVAL_3300 = 10'h16 == _EVAL_1450;
  assign _EVAL_178 = 10'h17 == _EVAL_1450;
  assign _EVAL_2066 = 10'h18 == _EVAL_1450;
  assign _EVAL_1399 = 10'h19 == _EVAL_1450;
  assign _EVAL_1601 = 10'h1a == _EVAL_1450;
  assign _EVAL_2432 = 10'h1b == _EVAL_1450;
  assign _EVAL_3729 = 10'h1c == _EVAL_1450;
  assign _EVAL_1132 = 10'h1d == _EVAL_1450;
  assign _EVAL_2659 = 10'h1e == _EVAL_1450;
  assign _EVAL_555 = 10'h1f == _EVAL_1450;
  assign _EVAL_808 = 10'h20 == _EVAL_1450;
  assign _EVAL_1965 = 10'h21 == _EVAL_1450;
  assign _EVAL_2410 = 10'h22 == _EVAL_1450;
  assign _EVAL_2763 = 10'h23 == _EVAL_1450;
  assign _EVAL_2102 = 10'h24 == _EVAL_1450;
  assign _EVAL_3776 = 10'h25 == _EVAL_1450;
  assign _EVAL_3401 = 10'h26 == _EVAL_1450;
  assign _EVAL_2796 = 10'h27 == _EVAL_1450;
  assign _EVAL_840 = 10'h28 == _EVAL_1450;
  assign _EVAL_1097 = 10'h29 == _EVAL_1450;
  assign _EVAL_1945 = 10'h2a == _EVAL_1450;
  assign _EVAL_2932 = 10'h2b == _EVAL_1450;
  assign _EVAL_2060 = 10'h2c == _EVAL_1450;
  assign _EVAL_1946 = 10'h2d == _EVAL_1450;
  assign _EVAL_1952 = 10'h2e == _EVAL_1450;
  assign _EVAL_2000 = 10'h2f == _EVAL_1450;
  assign _EVAL_3994 = 10'h30 == _EVAL_1450;
  assign _EVAL_1669 = 10'h31 == _EVAL_1450;
  assign _EVAL_1931 = 10'h32 == _EVAL_1450;
  assign _EVAL_511 = 10'h33 == _EVAL_1450;
  assign _EVAL_1875 = _EVAL_4052 ? {{29'd0}, _EVAL_1438} : _EVAL_1578;
  assign _EVAL_3564 = _EVAL_3081 ? {{29'd0}, _EVAL_1783} : _EVAL_1875;
  assign _EVAL_3258 = _EVAL_1440 ? {{29'd0}, _EVAL_3216} : _EVAL_3564;
  assign _EVAL_516 = _EVAL_511 ? {{29'd0}, _EVAL_444} : _EVAL_3258;
  assign _EVAL_2147 = _EVAL_1931 ? {{29'd0}, _EVAL_2484} : _EVAL_516;
  assign _EVAL_928 = _EVAL_1669 ? {{29'd0}, _EVAL_3113} : _EVAL_2147;
  assign _EVAL_254 = _EVAL_3994 ? {{29'd0}, _EVAL_3014} : _EVAL_928;
  assign _EVAL_1130 = _EVAL_2000 ? {{29'd0}, _EVAL_2965} : _EVAL_254;
  assign _EVAL_2063 = _EVAL_1952 ? {{29'd0}, _EVAL_1433} : _EVAL_1130;
  assign _EVAL_3911 = _EVAL_1946 ? {{29'd0}, _EVAL_4013} : _EVAL_2063;
  assign _EVAL_2867 = _EVAL_2060 ? {{29'd0}, _EVAL_354} : _EVAL_3911;
  assign _EVAL_3898 = _EVAL_2932 ? {{29'd0}, _EVAL_293} : _EVAL_2867;
  assign _EVAL_4038 = _EVAL_1945 ? {{29'd0}, _EVAL_3721} : _EVAL_3898;
  assign _EVAL_3158 = _EVAL_1097 ? {{29'd0}, _EVAL_2121} : _EVAL_4038;
  assign _EVAL_1052 = _EVAL_840 ? {{29'd0}, _EVAL_512} : _EVAL_3158;
  assign _EVAL_1329 = _EVAL_2796 ? {{29'd0}, _EVAL_750} : _EVAL_1052;
  assign _EVAL_3364 = _EVAL_3401 ? {{29'd0}, _EVAL_3274} : _EVAL_1329;
  assign _EVAL_1959 = _EVAL_3776 ? {{29'd0}, _EVAL_762} : _EVAL_3364;
  assign _EVAL_2228 = _EVAL_2102 ? {{29'd0}, _EVAL_2810} : _EVAL_1959;
  assign _EVAL_1051 = _EVAL_2763 ? {{29'd0}, _EVAL_3554} : _EVAL_2228;
  assign _EVAL_3646 = _EVAL_2410 ? {{29'd0}, _EVAL_1035} : _EVAL_1051;
  assign _EVAL_1061 = _EVAL_1965 ? {{29'd0}, _EVAL_2851} : _EVAL_3646;
  assign _EVAL_3060 = _EVAL_808 ? {{29'd0}, _EVAL_1562} : _EVAL_1061;
  assign _EVAL_1866 = _EVAL_555 ? {{29'd0}, _EVAL_3608} : _EVAL_3060;
  assign _EVAL_3831 = _EVAL_2659 ? {{29'd0}, _EVAL_3843} : _EVAL_1866;
  assign _EVAL_703 = _EVAL_1132 ? {{29'd0}, _EVAL_3573} : _EVAL_3831;
  assign _EVAL_225 = _EVAL_3729 ? {{29'd0}, _EVAL_155} : _EVAL_703;
  assign _EVAL_1985 = _EVAL_2432 ? {{29'd0}, _EVAL_3008} : _EVAL_225;
  assign _EVAL_2877 = _EVAL_1601 ? {{29'd0}, _EVAL_2536} : _EVAL_1985;
  assign _EVAL_1468 = _EVAL_1399 ? {{29'd0}, _EVAL_247} : _EVAL_2877;
  assign _EVAL_1741 = _EVAL_2066 ? {{29'd0}, _EVAL_286} : _EVAL_1468;
  assign _EVAL_2459 = _EVAL_178 ? {{29'd0}, _EVAL_3740} : _EVAL_1741;
  assign _EVAL_1393 = _EVAL_3300 ? {{29'd0}, _EVAL_2311} : _EVAL_2459;
  assign _EVAL_1323 = _EVAL_2007 ? {{29'd0}, _EVAL_1122} : _EVAL_1393;
  assign _EVAL_149 = _EVAL_2003 ? {{29'd0}, _EVAL_3571} : _EVAL_1323;
  assign _EVAL_1343 = _EVAL_472 ? {{29'd0}, _EVAL_1142} : _EVAL_149;
  assign _EVAL_2513 = _EVAL_237 ? {{29'd0}, _EVAL_1786} : _EVAL_1343;
  assign _EVAL_2148 = _EVAL_3358 ? {{29'd0}, _EVAL_739} : _EVAL_2513;
  assign _EVAL_329 = _EVAL_1572 ? {{29'd0}, _EVAL_2937} : _EVAL_2148;
  assign _EVAL_3385 = _EVAL_3233 ? {{29'd0}, _EVAL_1870} : _EVAL_329;
  assign _EVAL_2640 = _EVAL_3159 ? {{29'd0}, _EVAL_2760} : _EVAL_3385;
  assign _EVAL_3772 = _EVAL_2625 ? {{29'd0}, _EVAL_1801} : _EVAL_2640;
  assign _EVAL_2095 = _EVAL_1055 ? {{29'd0}, _EVAL_2653} : _EVAL_3772;
  assign _EVAL_461 = _EVAL_262 ? {{29'd0}, _EVAL_3383} : _EVAL_2095;
  assign _EVAL_542 = _EVAL_2535 ? {{29'd0}, _EVAL_4050} : _EVAL_461;
  assign _EVAL_3614 = _EVAL_4039 ? {{29'd0}, _EVAL_2110} : _EVAL_542;
  assign _EVAL_1654 = _EVAL_881 ? {{29'd0}, _EVAL_2491} : _EVAL_3614;
  assign _EVAL_1376 = _EVAL_3323 ? {{29'd0}, _EVAL_481} : _EVAL_1654;
  assign _EVAL_2728 = _EVAL_1416 ? {{29'd0}, _EVAL_4066} : _EVAL_1376;
  assign _EVAL_1907 = _EVAL_2999[127];
  assign _EVAL_1328 = _EVAL_2999[256];
  assign _EVAL_1332 = _EVAL_2124[7:1];
  assign _EVAL_3082 = _EVAL_511 ? _EVAL_2267 : _EVAL_2790;
  assign _EVAL_1811 = _EVAL_1931 ? _EVAL_2267 : _EVAL_3082;
  assign _EVAL_1352 = _EVAL_1669 ? _EVAL_2267 : _EVAL_1811;
  assign _EVAL_3907 = _EVAL_3994 ? _EVAL_2267 : _EVAL_1352;
  assign _EVAL_2056 = _EVAL_2000 ? _EVAL_2267 : _EVAL_3907;
  assign _EVAL_1458 = _EVAL_1952 ? _EVAL_2267 : _EVAL_2056;
  assign _EVAL_1717 = _EVAL_1946 ? _EVAL_2267 : _EVAL_1458;
  assign _EVAL_348 = _EVAL_2060 ? _EVAL_2267 : _EVAL_1717;
  assign _EVAL_2104 = _EVAL_2932 ? _EVAL_2267 : _EVAL_348;
  assign _EVAL_3231 = _EVAL_1945 ? _EVAL_2267 : _EVAL_2104;
  assign _EVAL_3370 = _EVAL_1097 ? _EVAL_2267 : _EVAL_3231;
  assign _EVAL_722 = _EVAL_840 ? _EVAL_2267 : _EVAL_3370;
  assign _EVAL_3881 = _EVAL_2796 ? _EVAL_2267 : _EVAL_722;
  assign _EVAL_2310 = _EVAL_3401 ? _EVAL_2267 : _EVAL_3881;
  assign _EVAL_2848 = _EVAL_3776 ? _EVAL_2267 : _EVAL_2310;
  assign _EVAL_3671 = _EVAL_1635[52];
  assign _EVAL_3595 = _EVAL_3671 | LevelGateway_51__EVAL_3;
  assign _EVAL_3534 = _EVAL_3671 == 1'h0;
  assign _EVAL_1236 = _EVAL_2999[24];
  assign _EVAL_2861 = _EVAL_3673 & _EVAL_1236;
  assign _EVAL_2524 = _EVAL_2861 & _EVAL_2267;
  assign _EVAL_2001 = _EVAL_2524 & _EVAL_591;
  assign _EVAL_829 = _EVAL_2999[1];
  assign _EVAL_1634 = _EVAL_2999[48];
  assign _EVAL_2079 = _EVAL_3673 & _EVAL_1634;
  assign _EVAL_416 = _EVAL_2079 & _EVAL_2267;
  assign _EVAL_4001 = _EVAL_416 & _EVAL_591;
  assign _EVAL_2288 = {_EVAL_4063,_EVAL_519,_EVAL_1938,_EVAL_3167,_EVAL_1753,_EVAL_1917,_EVAL_480,_EVAL_1496};
  assign _EVAL_189 = _EVAL_1635[17];
  assign _EVAL_1294 = _EVAL_189 | LevelGateway_16__EVAL_3;
  assign _EVAL_3499 = _EVAL_1635[59];
  assign _EVAL_195 = _EVAL_3499 | LevelGateway_58__EVAL_3;
  assign _EVAL_2940 = _EVAL_2999[85];
  assign _EVAL_3094 = _EVAL_2999[33];
  assign _EVAL_3584 = _EVAL_3673 & _EVAL_3094;
  assign _EVAL_873 = _EVAL_2999[101];
  assign _EVAL_3756 = _EVAL_1635[70];
  assign _EVAL_3061 = _EVAL_1635[81];
  assign _EVAL_1229 = _EVAL_3061 | LevelGateway_80__EVAL_3;
  assign _EVAL_2571 = _EVAL_2999[84];
  assign _EVAL_2415 = _EVAL_3673 & _EVAL_2571;
  assign _EVAL_1915 = _EVAL_1635[7];
  assign _EVAL_1958 = _EVAL_1915 == 1'h0;
  assign _EVAL_1201 = _EVAL_2999[259];
  assign _EVAL_638 = _EVAL_2124[23:16];
  assign _EVAL_1856 = _EVAL_1635[68];
  assign _EVAL_2208 = _EVAL_1856 | LevelGateway_67__EVAL_3;
  assign _EVAL_938 = _EVAL_2999[17];
  assign _EVAL_1699 = _EVAL_3673 & _EVAL_938;
  assign _EVAL_464 = _EVAL_1699 & _EVAL_2267;
  assign _EVAL_2869 = _EVAL_464 & _EVAL_591;
  assign _EVAL_824 = _EVAL_2999[37];
  assign _EVAL_3755 = _EVAL_339 == 1'h0;
  assign _EVAL_2745 = _EVAL_1635[44];
  assign _EVAL_2573 = _EVAL_2745 == 1'h0;
  assign _EVAL_1475 = _EVAL_2999[80];
  assign _EVAL_1785 = _EVAL_1635[10];
  assign _EVAL_1452 = _EVAL_1785 == 1'h0;
  assign _EVAL_1992 = _EVAL_1635[75];
  assign _EVAL_846 = _EVAL_1992 == 1'h0;
  assign _EVAL_2835 = _EVAL_2999[79];
  assign _EVAL_2856 = _EVAL_2999[51];
  assign _EVAL_362 = _EVAL_3673 & _EVAL_2856;
  assign _EVAL_533 = _EVAL_362 & _EVAL_2267;
  assign _EVAL_2660 = _EVAL_533 & _EVAL_591;
  assign _EVAL_3424 = _EVAL_339 | LevelGateway_117__EVAL_3;
  assign _EVAL_2118 = _EVAL_2102 ? _EVAL_2267 : _EVAL_2848;
  assign _EVAL_3348 = _EVAL_2763 ? _EVAL_2267 : _EVAL_2118;
  assign _EVAL_1790 = _EVAL_2410 ? _EVAL_2267 : _EVAL_3348;
  assign _EVAL_2464 = _EVAL_1965 ? _EVAL_2267 : _EVAL_1790;
  assign _EVAL_3379 = _EVAL_808 ? _EVAL_2267 : _EVAL_2464;
  assign _EVAL_3134 = _EVAL_555 ? _EVAL_2267 : _EVAL_3379;
  assign _EVAL_3665 = _EVAL_2659 ? _EVAL_2267 : _EVAL_3134;
  assign _EVAL_3439 = _EVAL_1132 ? _EVAL_2267 : _EVAL_3665;
  assign _EVAL_736 = _EVAL_3729 ? _EVAL_2267 : _EVAL_3439;
  assign _EVAL_2713 = _EVAL_2999[64];
  assign _EVAL_1877 = _EVAL_3673 & _EVAL_2713;
  assign _EVAL_2054 = _EVAL_2999[111];
  assign _EVAL_3895 = _EVAL_3673 & _EVAL_2054;
  assign _EVAL_3415 = _EVAL_1877 & _EVAL_2267;
  assign _EVAL_660 = _EVAL_3415 & _EVAL_591;
  assign _EVAL_2052 = _EVAL_2999[107];
  assign _EVAL_3404 = _EVAL_3673 & _EVAL_2052;
  assign _EVAL_2006 = _EVAL_3404 & _EVAL_2267;
  assign _EVAL_1355 = _EVAL_2006 & _EVAL_591;
  assign _EVAL_3372 = _EVAL_2124[31:24];
  assign _EVAL_187 = _EVAL_3372 == 8'hff;
  assign _EVAL_2528 = _EVAL_2999[19];
  assign _EVAL_4020 = _EVAL_1635[99];
  assign _EVAL_2171 = _EVAL_3673 & _EVAL_1328;
  assign _EVAL_3594 = _EVAL_2171 & _EVAL_2267;
  assign _EVAL_695 = _EVAL_2124[15:8];
  assign _EVAL_2335 = _EVAL_695 == 8'hff;
  assign _EVAL_2865 = _EVAL_3594 & _EVAL_2335;
  assign _EVAL_979 = _EVAL_2999[29];
  assign _EVAL_3932 = _EVAL_2999[91];
  assign _EVAL_3961 = _EVAL_3673 & _EVAL_3932;
  assign _EVAL_1780 = _EVAL_1635[87];
  assign _EVAL_2555 = _EVAL_1780 == 1'h0;
  assign _EVAL_3240 = _EVAL_1635[105];
  assign _EVAL_2156 = _EVAL_3240 == 1'h0;
  assign _EVAL_3055 = _EVAL_2124[7:0];
  assign _EVAL_3454 = _EVAL_2999[63];
  assign _EVAL_2664 = _EVAL_3673 & _EVAL_3454;
  assign _EVAL_3930 = _EVAL_2664 & _EVAL_2267;
  assign _EVAL_2615 = _EVAL_1635[31];
  assign _EVAL_3546 = _EVAL_2615 | LevelGateway_30__EVAL_3;
  assign _EVAL_2782 = _EVAL_1635[94];
  assign _EVAL_704 = _EVAL_1635[11];
  assign _EVAL_3292 = _EVAL_704 | LevelGateway_10__EVAL_3;
  assign _EVAL_3256 = _EVAL_704 == 1'h0;
  assign _EVAL_4054 = _EVAL_2999[25];
  assign _EVAL_1944 = _EVAL_2999[30];
  assign _EVAL_3325 = _EVAL_2999[81];
  assign _EVAL_3816 = _EVAL_2999[124];
  assign _EVAL_2204 = _EVAL_3673 & _EVAL_3816;
  assign _EVAL_1839 = _EVAL_2204 & _EVAL_2267;
  assign _EVAL_1533 = _EVAL_2999[95];
  assign _EVAL_3520 = _EVAL_2999[34];
  assign _EVAL_3918 = _EVAL_3673 & _EVAL_3325;
  assign _EVAL_3908 = _EVAL_2999[76];
  assign _EVAL_1462 = _EVAL_1635[110];
  assign _EVAL_3390 = _EVAL_1462 | LevelGateway_109__EVAL_3;
  assign _EVAL_3705 = _EVAL_1635[63];
  assign _EVAL_1887 = _EVAL_3705 | LevelGateway_62__EVAL_3;
  assign _EVAL_1107 = _EVAL_2999[60];
  assign _EVAL_985 = _EVAL_2999[89];
  assign _EVAL_2183 = _EVAL_1635[90];
  assign _EVAL_3018 = _EVAL_2999[2];
  assign _EVAL_1232 = _EVAL_1765 & _EVAL_591;
  assign _EVAL_2572 = _EVAL_1635[74];
  assign _EVAL_2969 = _EVAL_2572 == 1'h0;
  assign _EVAL_3434 = _EVAL_1635[5];
  assign _EVAL_622 = _EVAL_3434 | LevelGateway_4__EVAL_3;
  assign _EVAL_2333 = _EVAL_1635[84];
  assign _EVAL_1021 = _EVAL_2333 | LevelGateway_83__EVAL_3;
  assign _EVAL_3817 = _EVAL_1635[24];
  assign _EVAL_1486 = _EVAL_3817 | LevelGateway_23__EVAL_3;
  assign _EVAL_2907 = _EVAL_3817 == 1'h0;
  assign _EVAL_1196 = _EVAL_1635[121];
  assign _EVAL_1265 = _EVAL_1196 | LevelGateway_120__EVAL_3;
  assign _EVAL_428 = _EVAL_1196 == 1'h0;
  assign _EVAL_828 = _EVAL_2999[102];
  assign _EVAL_3156 = _EVAL_3673 & _EVAL_828;
  assign _EVAL_320 = _EVAL_1780 | LevelGateway_86__EVAL_3;
  assign _EVAL_1552 = {_EVAL_2809,_EVAL_3245,_EVAL_3551,_EVAL_3728,_EVAL_1261,_EVAL_3299,_EVAL_1536,_EVAL_1580};
  assign _EVAL_2287 = {_EVAL_552,_EVAL_3023,_EVAL_2701,_EVAL_421,_EVAL_3359,_EVAL_4034,_EVAL_947,_EVAL_1587};
  assign _EVAL_1746 = {_EVAL_2850,_EVAL_880,_EVAL_212,_EVAL_1930,_EVAL_3361,_EVAL_2159,_EVAL_497,_EVAL_3039,_EVAL_2287};
  assign _EVAL_3239 = {_EVAL_2953,_EVAL_3788,_EVAL_3783,_EVAL_3279,_EVAL_3757,_EVAL_3996,_EVAL_1270,_EVAL_2972,_EVAL_1552,_EVAL_1746};
  assign _EVAL_226 = _EVAL_2999[122];
  assign _EVAL_2746 = _EVAL_1635[47];
  assign _EVAL_3078 = _EVAL_2746 == 1'h0;
  assign _EVAL_1009 = _EVAL_3673 & _EVAL_3520;
  assign _EVAL_146 = _EVAL_1009 & _EVAL_2267;
  assign _EVAL_2048 = _EVAL_146 & _EVAL_591;
  assign _EVAL_1181 = _EVAL_1635[76];
  assign _EVAL_2047 = Queue__EVAL[31:24];
  assign _EVAL_845 = _EVAL_2999[14];
  assign _EVAL_3884 = _EVAL_2999[116];
  assign _EVAL_3318 = _EVAL_2999[4];
  assign _EVAL_438 = _EVAL_3673 & _EVAL_3318;
  assign _EVAL_1503 = _EVAL_438 & _EVAL_2267;
  assign _EVAL_263 = _EVAL_1635[20];
  assign _EVAL_3641 = _EVAL_263 == 1'h0;
  assign _EVAL_3508 = _EVAL_2999[43];
  assign _EVAL_653 = _EVAL_3673 & _EVAL_3508;
  assign _EVAL_207 = _EVAL_653 & _EVAL_2267;
  assign _EVAL_3423 = _EVAL_2999[87];
  assign _EVAL_921 = _EVAL_3673 & _EVAL_3423;
  assign _EVAL_1289 = _EVAL_921 & _EVAL_2267;
  assign _EVAL_291 = Queue__EVAL_3;
  assign _EVAL_236 = _EVAL_2999[41];
  assign _EVAL_1516 = _EVAL_3673 & _EVAL_236;
  assign _EVAL_3220 = _EVAL_1516 & _EVAL_2267;
  assign _EVAL_1326 = _EVAL_2999[49];
  assign _EVAL_271 = _EVAL_3673 & _EVAL_2184;
  assign _EVAL_607 = _EVAL_271 & _EVAL_2267;
  assign _EVAL_1337 = _EVAL_607 & _EVAL_591;
  assign _EVAL_1309 = _EVAL_626 & _EVAL_591;
  assign _EVAL_1706 = _EVAL_2999[59];
  assign _EVAL_1881 = _EVAL_3673 & _EVAL_1706;
  assign _EVAL_3098 = _EVAL_1881 & _EVAL_2267;
  assign _EVAL_1548 = _EVAL_3098 & _EVAL_591;
  assign _EVAL_2248 = _EVAL_3673 & _EVAL_1201;
  assign _EVAL_2559 = _EVAL_2248 & _EVAL_2267;
  assign _EVAL_2354 = _EVAL_638 == 8'hff;
  assign _EVAL_2515 = _EVAL_2559 & _EVAL_2354;
  assign _EVAL_3642 = _EVAL_2999[74];
  assign _EVAL_3282 = _EVAL_3673 & _EVAL_3642;
  assign _EVAL_1704 = _EVAL_1635[36];
  assign _EVAL_2463 = _EVAL_1704 | LevelGateway_35__EVAL_3;
  assign _EVAL_245 = _EVAL_1635[25];
  assign _EVAL_1549 = _EVAL_1635[14];
  assign _EVAL_1914 = _EVAL_1549 | LevelGateway_13__EVAL_3;
  assign _EVAL_3679 = _EVAL_2999[58];
  assign _EVAL_3959 = _EVAL_3673 & _EVAL_3679;
  assign _EVAL_1853 = _EVAL_1635[117];
  assign _EVAL_2346 = _EVAL_1853 | LevelGateway_116__EVAL_3;
  assign _EVAL_3074 = _EVAL_3918 & _EVAL_2267;
  assign _EVAL_3234 = _EVAL_3074 & _EVAL_591;
  assign _EVAL_1731 = _EVAL_3673 & _EVAL_829;
  assign _EVAL_1164 = _EVAL_1731 & _EVAL_2267;
  assign _EVAL_917 = _EVAL_2745 | LevelGateway_43__EVAL_3;
  assign _EVAL_1855 = _EVAL_2615 == 1'h0;
  assign _EVAL_455 = _EVAL_2999[52];
  assign _EVAL_507 = _EVAL_3673 & _EVAL_455;
  assign _EVAL_1368 = _EVAL_507 & _EVAL_2267;
  assign _EVAL_466 = _EVAL_1368 & _EVAL_591;
  assign _EVAL_353 = _EVAL_2999[23];
  assign _EVAL_2852 = _EVAL_378 | LevelGateway_17__EVAL_3;
  assign _EVAL_2947 = _EVAL_2999[105];
  assign _EVAL_3459 = _EVAL_1635[38];
  assign _EVAL_248 = _EVAL_3459 | LevelGateway_37__EVAL_3;
  assign _EVAL_3628 = _EVAL_2999[38];
  assign _EVAL_1876 = _EVAL_3673 & _EVAL_1326;
  assign _EVAL_2553 = _EVAL_1876 & _EVAL_2267;
  assign _EVAL_2845 = _EVAL_2553 & _EVAL_591;
  assign _EVAL_1613 = _EVAL_2999[44];
  assign _EVAL_1259 = _EVAL_1626 | LevelGateway_84__EVAL_3;
  assign _EVAL_809 = _EVAL_3055 == 8'hff;
  assign _EVAL_2825 = _EVAL_2559 & _EVAL_809;
  assign _EVAL_4056 = _EVAL_3418 == 1'h0;
  assign _EVAL_303 = _EVAL_1181 | LevelGateway_75__EVAL_3;
  assign _EVAL_3443 = _EVAL_1181 == 1'h0;
  assign _EVAL_514 = _EVAL_1635[96];
  assign _EVAL_3509 = _EVAL_1635[6];
  assign _EVAL_2008 = _EVAL_1635[58];
  assign _EVAL_3680 = _EVAL_2008 == 1'h0;
  assign _EVAL_851 = _EVAL_2999[20];
  assign _EVAL_3690 = _EVAL_3673 & _EVAL_851;
  assign _EVAL_930 = _EVAL_3690 & _EVAL_2267;
  assign _EVAL_3489 = _EVAL_2999[108];
  assign _EVAL_3726 = _EVAL_930 & _EVAL_591;
  assign _EVAL_1880 = _EVAL_2999[10];
  assign _EVAL_2146 = _EVAL_1635[48];
  assign _EVAL_2624 = _EVAL_2146 | LevelGateway_47__EVAL_3;
  assign _EVAL_401 = _EVAL_2146 == 1'h0;
  assign _EVAL_2279 = _EVAL_1635[69];
  assign _EVAL_2574 = _EVAL_2279 == 1'h0;
  assign _EVAL_753 = _EVAL_2432 ? _EVAL_2267 : _EVAL_736;
  assign _EVAL_2779 = _EVAL_1601 ? _EVAL_2267 : _EVAL_753;
  assign _EVAL_1222 = _EVAL_1399 ? _EVAL_2267 : _EVAL_2779;
  assign _EVAL_2730 = _EVAL_2066 ? _EVAL_2267 : _EVAL_1222;
  assign _EVAL_1241 = _EVAL_178 ? _EVAL_2267 : _EVAL_2730;
  assign _EVAL_3069 = _EVAL_2999[22];
  assign _EVAL_3221 = _EVAL_3673 & _EVAL_979;
  assign _EVAL_1085 = _EVAL_3221 & _EVAL_2267;
  assign _EVAL_795 = _EVAL_1635[120];
  assign _EVAL_3919 = _EVAL_2999[67];
  assign _EVAL_1525 = _EVAL_3673 & _EVAL_3919;
  assign _EVAL_899 = _EVAL_1525 & _EVAL_2267;
  assign _EVAL_926 = _EVAL_2999[94];
  assign _EVAL_3043 = _EVAL_2999[118];
  assign _EVAL_415 = _EVAL_2999[258];
  assign _EVAL_323 = _EVAL_3673 & _EVAL_1944;
  assign _EVAL_1956 = _EVAL_323 & _EVAL_2267;
  assign _EVAL_3803 = _EVAL_1635[127];
  assign _EVAL_1843 = _EVAL_3803 == 1'h0;
  assign _EVAL_1890 = _EVAL_1635[41];
  assign _EVAL_2391 = _EVAL_1635[37];
  assign _EVAL_509 = _EVAL_2391 | LevelGateway_36__EVAL_3;
  assign _EVAL_2858 = _EVAL_1635[126];
  assign _EVAL_3431 = _EVAL_2858 | LevelGateway_125__EVAL_3;
  assign _EVAL_1986 = _EVAL_2858 == 1'h0;
  assign _EVAL_4068 = _EVAL_2572 | LevelGateway_73__EVAL_3;
  assign _EVAL_2477 = _EVAL_1635[114];
  assign _EVAL_1500 = _EVAL_2477 | LevelGateway_113__EVAL_3;
  assign _EVAL_2443 = _EVAL_2477 == 1'h0;
  assign _EVAL_3335 = _EVAL_1635[93];
  assign _EVAL_2548 = _EVAL_3335 | LevelGateway_92__EVAL_3;
  assign _EVAL_3252 = _EVAL_3335 == 1'h0;
  assign _EVAL_3053 = _EVAL_1635[27];
  assign _EVAL_265 = _EVAL_2999[5];
  assign _EVAL_1397 = _EVAL_3061 == 1'h0;
  assign _EVAL_1537 = _EVAL_1635[86];
  assign _EVAL_2902 = _EVAL_1537 | LevelGateway_85__EVAL_3;
  assign _EVAL_488 = _EVAL_1537 == 1'h0;
  assign _EVAL_3852 = _EVAL_3803 | LevelGateway_126__EVAL_3;
  assign _EVAL_3675 = _EVAL_795 | LevelGateway_119__EVAL_3;
  assign _EVAL_1648 = _EVAL_2999[112];
  assign _EVAL_2742 = _EVAL_2999[31];
  assign _EVAL_540 = _EVAL_1635[113];
  assign _EVAL_1264 = _EVAL_540 | LevelGateway_112__EVAL_3;
  assign _EVAL_1283 = _EVAL_1635[60];
  assign _EVAL_574 = _EVAL_1283 | LevelGateway_59__EVAL_3;
  assign _EVAL_2750 = _EVAL_1283 == 1'h0;
  assign _EVAL_1298 = _EVAL_3673 & _EVAL_2528;
  assign _EVAL_2366 = _EVAL_1298 & _EVAL_2267;
  assign _EVAL_2631 = _EVAL_3673 & _EVAL_2742;
  assign _EVAL_1230 = _EVAL_2999[11];
  assign _EVAL_2303 = _EVAL_2999[53];
  assign _EVAL_1002 = _EVAL_1635[101];
  assign _EVAL_565 = _EVAL_1002 == 1'h0;
  assign _EVAL_2595 = _EVAL_3673 & _EVAL_1107;
  assign _EVAL_3122 = _EVAL_2595 & _EVAL_2267;
  assign _EVAL_1215 = _EVAL_3122 & _EVAL_591;
  assign _EVAL_3088 = _EVAL_2999[8];
  assign _EVAL_792 = _EVAL_1332 == 7'h7f;
  assign _EVAL_2696 = _EVAL_3594 & _EVAL_792;
  assign _EVAL_3497 = {_EVAL_366,_EVAL_3870,_EVAL_3913,_EVAL_3488,_EVAL_3743,_EVAL_3421,_EVAL_1639,_EVAL_1698};
  assign _EVAL_1469 = {_EVAL_3623,_EVAL_1697,_EVAL_2188,_EVAL_2018,_EVAL_1776,_EVAL_2754,_EVAL_2073,_EVAL_1162,_EVAL_3497,1'h0};
  assign _EVAL_1584 = Queue__EVAL;
  assign _EVAL_666 = _EVAL_1584[6:0];
  assign _EVAL_553 = _EVAL_1469 >> _EVAL_666;
  assign _EVAL_3970 = _EVAL_553[0];
  assign _EVAL_1990 = _EVAL_3593 & _EVAL_3970;
  assign _EVAL_3166 = _EVAL_3673 & _EVAL_2947;
  assign _EVAL_2136 = _EVAL_1635[65];
  assign _EVAL_2277 = _EVAL_2136 | LevelGateway_64__EVAL_3;
  assign _EVAL_515 = _EVAL_2999[56];
  assign _EVAL_527 = _EVAL_3673 & _EVAL_515;
  assign _EVAL_2532 = _EVAL_527 & _EVAL_2267;
  assign _EVAL_3117 = _EVAL_2999[65];
  assign _EVAL_3689 = _EVAL_3673 & _EVAL_3117;
  assign _EVAL_1408 = _EVAL_3689 & _EVAL_2267;
  assign _EVAL_436 = _EVAL_1635[56];
  assign _EVAL_274 = _EVAL_436 | LevelGateway_55__EVAL_3;
  assign _EVAL_1136 = _EVAL_436 == 1'h0;
  assign _EVAL_377 = _EVAL_3673 & _EVAL_2610;
  assign _EVAL_748 = _EVAL_377 & _EVAL_2267;
  assign _EVAL_1707 = _EVAL_748 & _EVAL_591;
  assign _EVAL_939 = _EVAL_2999[104];
  assign _EVAL_2125 = _EVAL_3673 & _EVAL_939;
  assign _EVAL_2959 = _EVAL_2999[12];
  assign _EVAL_2157 = _EVAL_3673 & _EVAL_2959;
  assign _EVAL_3037 = _EVAL_2157 & _EVAL_2267;
  assign _EVAL_3744 = _EVAL_3037 & _EVAL_591;
  assign _EVAL_1793 = 10'h3 == _EVAL_1450;
  assign _EVAL_590 = 10'h4 == _EVAL_1450;
  assign _EVAL_1873 = 10'h5 == _EVAL_1450;
  assign _EVAL_1512 = _EVAL_3300 ? _EVAL_2267 : _EVAL_1241;
  assign _EVAL_4017 = _EVAL_2007 ? _EVAL_2267 : _EVAL_1512;
  assign _EVAL_973 = _EVAL_2003 ? _EVAL_2267 : _EVAL_4017;
  assign _EVAL_257 = _EVAL_472 ? _EVAL_2267 : _EVAL_973;
  assign _EVAL_800 = _EVAL_237 ? _EVAL_2267 : _EVAL_257;
  assign _EVAL_2251 = _EVAL_3358 ? _EVAL_2267 : _EVAL_800;
  assign _EVAL_2446 = _EVAL_1572 ? _EVAL_2267 : _EVAL_2251;
  assign _EVAL_1177 = _EVAL_3233 ? _EVAL_2267 : _EVAL_2446;
  assign _EVAL_4044 = _EVAL_3159 ? _EVAL_2267 : _EVAL_1177;
  assign _EVAL_3096 = _EVAL_2625 ? _EVAL_2267 : _EVAL_4044;
  assign _EVAL_3864 = _EVAL_1055 ? _EVAL_2267 : _EVAL_3096;
  assign _EVAL_821 = _EVAL_262 ? _EVAL_2267 : _EVAL_3864;
  assign _EVAL_727 = _EVAL_2535 ? _EVAL_2267 : _EVAL_821;
  assign _EVAL_2317 = _EVAL_4039 ? _EVAL_2267 : _EVAL_727;
  assign _EVAL_2106 = _EVAL_881 ? _EVAL_2267 : _EVAL_2317;
  assign _EVAL_1888 = _EVAL_3323 ? _EVAL_2267 : _EVAL_2106;
  assign _EVAL_592 = _EVAL_1416 ? _EVAL_2267 : _EVAL_1888;
  assign _EVAL_1148 = _EVAL_1873 ? _EVAL_2267 : _EVAL_592;
  assign _EVAL_1913 = _EVAL_590 ? _EVAL_2267 : _EVAL_1148;
  assign _EVAL_229 = _EVAL_1793 ? _EVAL_2267 : _EVAL_1913;
  assign _EVAL_525 = _EVAL_3895 & _EVAL_2267;
  assign _EVAL_3409 = _EVAL_525 & _EVAL_591;
  assign _EVAL_3510 = _EVAL_1635[78];
  assign _EVAL_2291 = _EVAL_3510 | LevelGateway_77__EVAL_3;
  assign _EVAL_375 = _EVAL_3510 == 1'h0;
  assign _EVAL_1432 = _EVAL_2999[93];
  assign _EVAL_1257 = _EVAL_3673 & _EVAL_1432;
  assign _EVAL_3476 = _EVAL_1257 & _EVAL_2267;
  assign _EVAL_3136 = _EVAL_3673 & _EVAL_3069;
  assign _EVAL_586 = _EVAL_1635[12];
  assign _EVAL_3269 = _EVAL_586 == 1'h0;
  assign _EVAL_3529 = _EVAL_1635[43];
  assign _EVAL_4032 = _EVAL_3529 | LevelGateway_42__EVAL_3;
  assign _EVAL_4041 = _EVAL_2999[88];
  assign _EVAL_4040 = _EVAL_2999[121];
  assign _EVAL_2731 = _EVAL_2999[75];
  assign _EVAL_2662 = _EVAL_1635[109];
  assign _EVAL_4043 = _EVAL_1635[32];
  assign _EVAL_3273 = _EVAL_4043 | LevelGateway_31__EVAL_3;
  assign _EVAL_3432 = Queue__EVAL[7:1];
  assign _EVAL_1064 = _EVAL_2999[125];
  assign _EVAL_3265 = _EVAL_3418 | LevelGateway_103__EVAL_3;
  assign _EVAL_3549 = _EVAL_514 | LevelGateway_95__EVAL_3;
  assign _EVAL_2565 = _EVAL_514 == 1'h0;
  assign _EVAL_1502 = _EVAL_2999[257];
  assign _EVAL_3981 = _EVAL_2999[3];
  assign _EVAL_3203 = _EVAL_1635[98];
  assign _EVAL_220 = _EVAL_3203 | LevelGateway_97__EVAL_3;
  assign _EVAL_1414 = _EVAL_3203 == 1'h0;
  assign _EVAL_3873 = _EVAL_2999[7];
  assign _EVAL_1922 = _EVAL_2999[99];
  assign _EVAL_3882 = _EVAL_2999[70];
  assign _EVAL_4062 = _EVAL_2999[78];
  assign _EVAL_3847 = _EVAL_2999[16];
  assign _EVAL_1764 = _EVAL_3673 & _EVAL_3847;
  assign _EVAL_2480 = _EVAL_1764 & _EVAL_2267;
  assign _EVAL_2697 = _EVAL_2480 & _EVAL_591;
  assign _EVAL_3707 = _EVAL_2999[40];
  assign _EVAL_2233 = _EVAL_2559 & _EVAL_2335;
  assign _EVAL_3588 = _EVAL_3673 & _EVAL_3884;
  assign _EVAL_710 = _EVAL_3588 & _EVAL_2267;
  assign _EVAL_2770 = _EVAL_710 & _EVAL_591;
  assign _EVAL_847 = _EVAL_2999[36];
  assign _EVAL_1202 = _EVAL_3673 & _EVAL_847;
  assign _EVAL_3429 = _EVAL_1202 & _EVAL_2267;
  assign _EVAL_2567 = _EVAL_2999[119];
  assign _EVAL_1069 = _EVAL_3673 & _EVAL_3882;
  assign _EVAL_2189 = _EVAL_2999[106];
  assign _EVAL_2388 = _EVAL_1635[28];
  assign _EVAL_2705 = _EVAL_2388 | LevelGateway_27__EVAL_3;
  assign _EVAL_2823 = _EVAL_2999[109];
  assign _EVAL_2503 = _EVAL_3673 & _EVAL_2823;
  assign _EVAL_1124 = _EVAL_1635[123];
  assign _EVAL_3011 = _EVAL_1124 == 1'h0;
  assign _EVAL_2320 = _EVAL_3673 & _EVAL_429;
  assign _EVAL_1100 = _EVAL_2320 & _EVAL_2267;
  assign _EVAL_927 = _EVAL_2999[123];
  assign _EVAL_3436 = _EVAL_3673 & _EVAL_927;
  assign _EVAL_2981 = _EVAL_3436 & _EVAL_2267;
  assign _EVAL_2467 = _EVAL_1635[102];
  assign _EVAL_3880 = _EVAL_2467 | LevelGateway_101__EVAL_3;
  assign _EVAL_2115 = {_EVAL_194,_EVAL_3283,_EVAL_912,_EVAL_3296,_EVAL_770,_EVAL_2838,_EVAL_730,_EVAL_1521};
  assign _EVAL_2629 = {_EVAL_715,_EVAL_1267,_EVAL_176,_EVAL_2942,_EVAL_3419,_EVAL_569,_EVAL_3199,_EVAL_3964,_EVAL_2115};
  assign _EVAL_1473 = {_EVAL_3713,_EVAL_3850,_EVAL_449,_EVAL_1471,_EVAL_1599,_EVAL_2938,_EVAL_741,_EVAL_2202,_EVAL_2288,_EVAL_2629};
  assign _EVAL_946 = {_EVAL_2688,_EVAL_2582,_EVAL_2803,_EVAL_2050,_EVAL_1313,_EVAL_3720,_EVAL_222,_EVAL_2485};
  assign _EVAL_2872 = {_EVAL_989,_EVAL_2684,_EVAL_427,_EVAL_1456,_EVAL_492,_EVAL_1315,_EVAL_462,_EVAL_2507};
  assign _EVAL_3380 = {_EVAL_1709,_EVAL_3715,_EVAL_3025,_EVAL_690,_EVAL_3899,_EVAL_2155,_EVAL_3407,_EVAL_1929,_EVAL_2872};
  assign _EVAL_1674 = {_EVAL_1073,_EVAL_2870,_EVAL_2341,_EVAL_2648,_EVAL_3137,_EVAL_1206,_EVAL_3527,_EVAL_2254,_EVAL_946,_EVAL_3380};
  assign _EVAL_594 = {_EVAL_2214,_EVAL_217,_EVAL_1708,_EVAL_3192,_EVAL_2666,_EVAL_269,_EVAL_2128,_EVAL_581};
  assign _EVAL_2883 = {_EVAL_1788,_EVAL_3759,_EVAL_163,_EVAL_2826,_EVAL_371,_EVAL_2209,_EVAL_2133};
  assign _EVAL_3972 = {_EVAL_1556,_EVAL_1121,_EVAL_3636,_EVAL_3750,_EVAL_1979,_EVAL_673,_EVAL_200,_EVAL_2807,_EVAL_2883};
  assign _EVAL_3999 = {_EVAL_3222,_EVAL_1597,_EVAL_3317,_EVAL_3505,_EVAL_448,_EVAL_387,_EVAL_306,_EVAL_614,_EVAL_594,_EVAL_3972};
  assign _EVAL_3572 = {_EVAL_1473,_EVAL_3239,_EVAL_1674,_EVAL_3999};
  assign _EVAL_1730 = _EVAL_1635[15];
  assign _EVAL_3334 = _EVAL_1730 | LevelGateway_14__EVAL_3;
  assign _EVAL_1439 = _EVAL_2999[54];
  assign _EVAL_732 = _EVAL_3282 & _EVAL_2267;
  assign _EVAL_308 = _EVAL_2999[110];
  assign _EVAL_2237 = _EVAL_3673 & _EVAL_308;
  assign _EVAL_1068 = _EVAL_2237 & _EVAL_2267;
  assign _EVAL_1948 = _EVAL_2999[71];
  assign _EVAL_987 = _EVAL_3673 & _EVAL_1948;
  assign _EVAL_3620 = _EVAL_987 & _EVAL_2267;
  assign _EVAL_1763 = _EVAL_3617 | LevelGateway_50__EVAL_3;
  assign _EVAL_1235 = _EVAL_2999[72];
  assign _EVAL_759 = _EVAL_3673 & _EVAL_1235;
  assign _EVAL_1297 = _EVAL_759 & _EVAL_2267;
  assign _EVAL_1650 = _EVAL_2999[32];
  assign _EVAL_219 = _EVAL_1635[22];
  assign _EVAL_1768 = _EVAL_2503 & _EVAL_2267;
  assign _EVAL_260 = _EVAL_2999[69];
  assign _EVAL_2743 = _EVAL_2999[35];
  assign _EVAL_1582 = _EVAL_1635[39];
  assign _EVAL_2627 = _EVAL_1582 | LevelGateway_38__EVAL_3;
  assign _EVAL_3682 = _EVAL_2999[66];
  assign _EVAL_1204 = _EVAL_3673 & _EVAL_3682;
  assign _EVAL_1837 = _EVAL_1204 & _EVAL_2267;
  assign _EVAL_335 = _EVAL_3705 == 1'h0;
  assign _EVAL_2449 = _EVAL_1635[82];
  assign _EVAL_1392 = _EVAL_2449 == 1'h0;
  assign _EVAL_1541 = _EVAL_1582 == 1'h0;
  assign _EVAL_2139 = _EVAL_4020 | LevelGateway_98__EVAL_3;
  assign _EVAL_2644 = _EVAL_2999[86];
  assign _EVAL_1237 = _EVAL_1805 == 1'h0;
  assign _EVAL_561 = _EVAL_3673 & _EVAL_3018;
  assign _EVAL_679 = _EVAL_561 & _EVAL_2267;
  assign _EVAL_3844 = _EVAL_2999[57];
  assign _EVAL_2545 = _EVAL_3673 & _EVAL_3844;
  assign _EVAL_2447 = _EVAL_2545 & _EVAL_2267;
  assign _EVAL_1957 = _EVAL_2447 & _EVAL_591;
  assign _EVAL_3287 = _EVAL_2999[55];
  assign _EVAL_326 = _EVAL_3673 & _EVAL_3287;
  assign _EVAL_4070 = _EVAL_326 & _EVAL_2267;
  assign _EVAL_954 = _EVAL_4070 & _EVAL_591;
  assign _EVAL_1213 = _EVAL_2999[13];
  assign _EVAL_1216 = _EVAL_2999[45];
  assign _EVAL_3615 = _EVAL_3673 & _EVAL_415;
  assign _EVAL_612 = _EVAL_679 & _EVAL_591;
  assign _EVAL_3101 = _EVAL_2999[9];
  assign _EVAL_896 = _EVAL_3156 & _EVAL_2267;
  assign _EVAL_412 = _EVAL_896 & _EVAL_591;
  assign _EVAL_3169 = _EVAL_1890 | LevelGateway_40__EVAL_3;
  assign _EVAL_1325 = _EVAL_2999[98];
  assign _EVAL_3350 = _EVAL_2999[27];
  assign _EVAL_2126 = _EVAL_1635[64];
  assign _EVAL_3185 = _EVAL_3476 & _EVAL_591;
  assign _EVAL_203 = _EVAL_1635[42];
  assign _EVAL_2325 = _EVAL_203 == 1'h0;
  assign _EVAL_315 = _EVAL_1956 & _EVAL_591;
  assign _EVAL_355 = _EVAL_3053 | LevelGateway_26__EVAL_3;
  assign _EVAL_3879 = _EVAL_3053 == 1'h0;
  assign _EVAL_2242 = _EVAL_3673 & _EVAL_2303;
  assign _EVAL_3041 = _EVAL_3673 & _EVAL_1502;
  assign _EVAL_2669 = _EVAL_3041 & _EVAL_2267;
  assign _EVAL_1564 = _EVAL_3459 == 1'h0;
  assign _EVAL_2455 = _EVAL_1635[9];
  assign _EVAL_1936 = _EVAL_2455 | LevelGateway_8__EVAL_3;
  assign _EVAL_2129 = _EVAL_2455 == 1'h0;
  assign _EVAL_1833 = _EVAL_2999[73];
  assign _EVAL_2468 = _EVAL_3673 & _EVAL_1648;
  assign _EVAL_1072 = _EVAL_2468 & _EVAL_2267;
  assign _EVAL_2097 = _EVAL_1072 & _EVAL_591;
  assign _EVAL_2023 = _EVAL_3673 & _EVAL_1922;
  assign _EVAL_1677 = _EVAL_3673 & _EVAL_3101;
  assign _EVAL_3991 = _EVAL_1635[2];
  assign _EVAL_1919 = _EVAL_3991 == 1'h0;
  assign _EVAL_1243 = _EVAL_1635[55];
  assign _EVAL_2144 = _EVAL_1635[53];
  assign _EVAL_3945 = _EVAL_2144 == 1'h0;
  assign _EVAL_2454 = _EVAL_1635[89];
  assign _EVAL_3784 = _EVAL_2454 == 1'h0;
  assign _EVAL_342 = _EVAL_1462 == 1'h0;
  assign _EVAL_3661 = _EVAL_3673 & _EVAL_2835;
  assign _EVAL_606 = _EVAL_3661 & _EVAL_2267;
  assign _EVAL_2690 = _EVAL_3594 & _EVAL_2354;
  assign _EVAL_2520 = _EVAL_2999[120];
  assign _EVAL_1013 = _EVAL_2999[113];
  assign _EVAL_3293 = _EVAL_3673 & _EVAL_1013;
  assign _EVAL_3659 = _EVAL_3293 & _EVAL_2267;
  assign _EVAL_3100 = _EVAL_3756 | LevelGateway_69__EVAL_3;
  assign _EVAL_3709 = _EVAL_3673 & _EVAL_2940;
  assign _EVAL_981 = _EVAL_3709 & _EVAL_2267;
  assign _EVAL_1182 = _EVAL_2999[15];
  assign _EVAL_2642 = _EVAL_3673 & _EVAL_1182;
  assign _EVAL_3853 = _EVAL_2642 & _EVAL_2267;
  assign _EVAL_3024 = _EVAL_3853 & _EVAL_591;
  assign _EVAL_994 = _EVAL_2415 & _EVAL_2267;
  assign _EVAL_2103 = _EVAL_1635[35];
  assign _EVAL_2682 = _EVAL_3673 & _EVAL_226;
  assign _EVAL_2229 = _EVAL_3615 & _EVAL_2267;
  assign _EVAL_4009 = _EVAL_2229 & _EVAL_809;
  assign _EVAL_3142 = _EVAL_3673 & _EVAL_3981;
  assign _EVAL_3266 = _EVAL_3142 & _EVAL_2267;
  assign _EVAL_1096 = _EVAL_2008 | LevelGateway_57__EVAL_3;
  assign _EVAL_1557 = _EVAL_3673 & _EVAL_1880;
  assign _EVAL_1492 = _EVAL_1557 & _EVAL_2267;
  assign _EVAL_691 = _EVAL_1492 & _EVAL_591;
  assign _EVAL_2167 = _EVAL_1635[66];
  assign _EVAL_3923 = _EVAL_3673 & _EVAL_3088;
  assign _EVAL_1211 = _EVAL_3923 & _EVAL_2267;
  assign _EVAL_2426 = _EVAL_1211 & _EVAL_591;
  assign _EVAL_2828 = _EVAL_3673 & _EVAL_2731;
  assign _EVAL_1200 = _EVAL_2828 & _EVAL_2267;
  assign _EVAL_3460 = _EVAL_3050 & _EVAL_591;
  assign _EVAL_2302 = _EVAL_2999[28];
  assign _EVAL_3903 = _EVAL_3673 & _EVAL_2302;
  assign _EVAL_1892 = _EVAL_3903 & _EVAL_2267;
  assign _EVAL_1841 = _EVAL_1892 & _EVAL_591;
  assign _EVAL_380 = _EVAL_2242 & _EVAL_2267;
  assign _EVAL_3832 = _EVAL_380 & _EVAL_591;
  assign _EVAL_3490 = _EVAL_1635[71];
  assign _EVAL_2788 = _EVAL_1853 == 1'h0;
  assign _EVAL_252 = _EVAL_3499 == 1'h0;
  assign _EVAL_720 = _EVAL_2103 | LevelGateway_34__EVAL_3;
  assign _EVAL_420 = _EVAL_1635[125];
  assign _EVAL_734 = _EVAL_420 | LevelGateway_124__EVAL_3;
  assign _EVAL_3868 = _EVAL_420 == 1'h0;
  assign _EVAL_3662 = _EVAL_1635[67];
  assign _EVAL_773 = _EVAL_3662 == 1'h0;
  assign _EVAL_1226 = _EVAL_2467 == 1'h0;
  assign _EVAL_2554 = _EVAL_1635[108];
  assign _EVAL_231 = _EVAL_1635[30];
  assign _EVAL_3667 = _EVAL_231 | LevelGateway_29__EVAL_3;
  assign _EVAL_1400 = _EVAL_2999[62];
  assign _EVAL_1602 = _EVAL_3673 & _EVAL_1400;
  assign _EVAL_3823 = _EVAL_1602 & _EVAL_2267;
  assign _EVAL_1338 = 10'h2 == _EVAL_1450;
  assign _EVAL_3244 = _EVAL_1873 ? {{29'd0}, _EVAL_251} : _EVAL_2728;
  assign _EVAL_2301 = _EVAL_590 ? {{29'd0}, _EVAL_285} : _EVAL_3244;
  assign _EVAL_1171 = _EVAL_1793 ? {{29'd0}, _EVAL_3102} : _EVAL_2301;
  assign _EVAL_1802 = _EVAL_1338 ? {{29'd0}, _EVAL_304} : _EVAL_1171;
  assign _EVAL_2011 = _EVAL_1635[73];
  assign _EVAL_2944 = _EVAL_2011 | LevelGateway_72__EVAL_3;
  assign _EVAL_3579 = _EVAL_2999[77];
  assign _EVAL_2886 = _EVAL_3673 & _EVAL_3579;
  assign _EVAL_1427 = _EVAL_2886 & _EVAL_2267;
  assign _EVAL_2143 = _EVAL_1427 & _EVAL_591;
  assign _EVAL_1671 = _EVAL_2449 | LevelGateway_81__EVAL_3;
  assign _EVAL_3687 = _EVAL_3673 & _EVAL_3707;
  assign _EVAL_1240 = _EVAL_2999[42];
  assign _EVAL_3012 = _EVAL_3673 & _EVAL_1240;
  assign _EVAL_1611 = _EVAL_3012 & _EVAL_2267;
  assign _EVAL_3618 = _EVAL_1611 & _EVAL_591;
  assign _EVAL_3625 = _EVAL_2011 == 1'h0;
  assign _EVAL_2539 = _EVAL_3673 & _EVAL_4054;
  assign _EVAL_2939 = _EVAL_2539 & _EVAL_2267;
  assign _EVAL_3337 = _EVAL_2939 & _EVAL_591;
  assign _EVAL_2187 = _EVAL_1635[8];
  assign _EVAL_2210 = _EVAL_2187 == 1'h0;
  assign _EVAL_925 = _EVAL_2999[92];
  assign _EVAL_3213 = _EVAL_2999[50];
  assign _EVAL_3887 = _EVAL_3673 & _EVAL_3213;
  assign _EVAL_345 = _EVAL_3887 & _EVAL_2267;
  assign _EVAL_667 = _EVAL_345 & _EVAL_591;
  assign _EVAL_2607 = _EVAL_3673 & _EVAL_3908;
  assign _EVAL_2304 = _EVAL_2607 & _EVAL_2267;
  assign _EVAL_1067 = _EVAL_2304 & _EVAL_591;
  assign _EVAL_3765 = _EVAL_2391 == 1'h0;
  assign _EVAL_3184 = _EVAL_1635[106];
  assign _EVAL_2910 = _EVAL_3184 | LevelGateway_105__EVAL_3;
  assign _EVAL_167 = _EVAL_3673 & _EVAL_3043;
  assign _EVAL_1370 = _EVAL_3673 & _EVAL_925;
  assign _EVAL_879 = _EVAL_1370 & _EVAL_2267;
  assign _EVAL_2557 = _EVAL_3673 & _EVAL_2644;
  assign _EVAL_1682 = _EVAL_3429 & _EVAL_591;
  assign _EVAL_2899 = _EVAL_3673 & _EVAL_3489;
  assign _EVAL_2494 = _EVAL_2899 & _EVAL_2267;
  assign _EVAL_3539 = _EVAL_2494 & _EVAL_591;
  assign _EVAL_1955 = _EVAL_1635[21];
  assign _EVAL_963 = _EVAL_1955 | LevelGateway_20__EVAL_3;
  assign _EVAL_3371 = _EVAL_1955 == 1'h0;
  assign _EVAL_3091 = _EVAL_3673 & _EVAL_3628;
  assign _EVAL_1617 = _EVAL_3091 & _EVAL_2267;
  assign _EVAL_3940 = _EVAL_1617 & _EVAL_591;
  assign _EVAL_316 = _EVAL_3594 & _EVAL_187;
  assign _EVAL_1357 = _EVAL_245 | LevelGateway_24__EVAL_3;
  assign _EVAL_310 = _EVAL_1635[19];
  assign _EVAL_2421 = _EVAL_310 == 1'h0;
  assign _EVAL_2378 = _EVAL_3490 | LevelGateway_70__EVAL_3;
  assign _EVAL_372 = _EVAL_3490 == 1'h0;
  assign _EVAL_3006 = _EVAL_2746 | LevelGateway_46__EVAL_3;
  assign _EVAL_865 = _EVAL_2183 | LevelGateway_89__EVAL_3;
  assign _EVAL_1751 = _EVAL_2183 == 1'h0;
  assign _EVAL_812 = _EVAL_3673 & _EVAL_1475;
  assign _EVAL_3822 = _EVAL_812 & _EVAL_2267;
  assign _EVAL_2533 = _EVAL_3822 & _EVAL_591;
  assign _EVAL_2952 = _EVAL_3662 | LevelGateway_66__EVAL_3;
  assign _EVAL_2416 = _EVAL_3673 & _EVAL_1907;
  assign _EVAL_2579 = _EVAL_2416 & _EVAL_2267;
  assign _EVAL_3825 = _EVAL_2662 | LevelGateway_108__EVAL_3;
  assign _EVAL_1424 = _EVAL_2662 == 1'h0;
  assign _EVAL_2818 = _EVAL_1635[119];
  assign _EVAL_1614 = _EVAL_2818 | LevelGateway_118__EVAL_3;
  assign _EVAL_1858 = _EVAL_2818 == 1'h0;
  assign _EVAL_2971 = _EVAL_3673 & _EVAL_3350;
  assign _EVAL_2137 = _EVAL_2971 & _EVAL_2267;
  assign _EVAL_313 = _EVAL_2137 & _EVAL_591;
  assign _EVAL_3107 = _EVAL_2023 & _EVAL_2267;
  assign _EVAL_1225 = _EVAL_3107 & _EVAL_591;
  assign _EVAL_295 = _EVAL_2999[114];
  assign _EVAL_3384 = _EVAL_3673 & _EVAL_295;
  assign _EVAL_830 = _EVAL_3384 & _EVAL_2267;
  assign _EVAL_3157 = _EVAL_3961 & _EVAL_2267;
  assign _EVAL_1027 = _EVAL_3157 & _EVAL_591;
  assign _EVAL_1131 = _EVAL_3673 & _EVAL_1213;
  assign _EVAL_832 = _EVAL_1131 & _EVAL_2267;
  assign _EVAL_1558 = _EVAL_832 & _EVAL_591;
  assign _EVAL_557 = _EVAL_2782 == 1'h0;
  assign _EVAL_2686 = _EVAL_3673 & _EVAL_1650;
  assign _EVAL_2854 = _EVAL_1635[95];
  assign _EVAL_1816 = _EVAL_2854 | LevelGateway_94__EVAL_3;
  assign _EVAL_3547 = _EVAL_3673 & _EVAL_985;
  assign _EVAL_3589 = _EVAL_3673 & _EVAL_265;
  assign _EVAL_1210 = _EVAL_3589 & _EVAL_2267;
  assign _EVAL_3064 = _EVAL_1210 & _EVAL_591;
  assign _EVAL_1835 = _EVAL_1635[54];
  assign _EVAL_360 = _EVAL_1835 | LevelGateway_53__EVAL_3;
  assign _EVAL_1723 = _EVAL_4020 == 1'h0;
  assign _EVAL_4064 = _EVAL_1635[62];
  assign _EVAL_221 = _EVAL_4064 | LevelGateway_61__EVAL_3;
  assign _EVAL_3946 = _EVAL_4064 == 1'h0;
  assign _EVAL_712 = _EVAL_1635[26];
  assign _EVAL_971 = _EVAL_712 == 1'h0;
  assign _EVAL_1161 = _EVAL_1100 & _EVAL_591;
  assign _EVAL_723 = _EVAL_1635[1];
  assign _EVAL_956 = _EVAL_723 | LevelGateway__EVAL_3;
  assign _EVAL_731 = _EVAL_723 == 1'h0;
  assign _EVAL_539 = _EVAL_3673 & _EVAL_1613;
  assign _EVAL_505 = _EVAL_539 & _EVAL_2267;
  assign _EVAL_1633 = _EVAL_1635[4];
  assign _EVAL_875 = _EVAL_3673 & _EVAL_824;
  assign _EVAL_1019 = _EVAL_875 & _EVAL_2267;
  assign _EVAL_3374 = _EVAL_3673 & _EVAL_873;
  assign _EVAL_1527 = _EVAL_3374 & _EVAL_2267;
  assign _EVAL_1120 = _EVAL_3620 & _EVAL_591;
  assign _EVAL_2608 = _EVAL_2999[82];
  assign _EVAL_1555 = _EVAL_3673 & _EVAL_2608;
  assign _EVAL_1784 = _EVAL_1164 & _EVAL_591;
  assign _EVAL_381 = _EVAL_3673 & _EVAL_845;
  assign _EVAL_1454 = _EVAL_381 & _EVAL_2267;
  assign _EVAL_1113 = _EVAL_2999[46];
  assign _EVAL_3952 = _EVAL_1635[33];
  assign _EVAL_1848 = _EVAL_2631 & _EVAL_2267;
  assign _EVAL_190 = _EVAL_3266 & _EVAL_591;
  assign _EVAL_2893 = _EVAL_3509 | LevelGateway_5__EVAL_3;
  assign _EVAL_2225 = _EVAL_586 | LevelGateway_11__EVAL_3;
  assign _EVAL_1509 = _EVAL_3673 & _EVAL_1886;
  assign _EVAL_820 = _EVAL_1635[13];
  assign _EVAL_242 = _EVAL_820 | LevelGateway_12__EVAL_3;
  assign _EVAL_571 = _EVAL_1454 & _EVAL_591;
  assign _EVAL_2169 = _EVAL_1124 | LevelGateway_122__EVAL_3;
  assign _EVAL_199 = _EVAL_3240 | LevelGateway_104__EVAL_3;
  assign _EVAL_2131 = _EVAL_167 & _EVAL_2267;
  assign _EVAL_2365 = _EVAL_245 == 1'h0;
  assign _EVAL_2482 = _EVAL_1785 | LevelGateway_9__EVAL_3;
  assign _EVAL_2651 = _EVAL_3673 & _EVAL_926;
  assign _EVAL_3338 = _EVAL_2651 & _EVAL_2267;
  assign _EVAL_1655 = _EVAL_3338 & _EVAL_591;
  assign _EVAL_2889 = _EVAL_1635[103];
  assign _EVAL_1350 = _EVAL_2889 | LevelGateway_102__EVAL_3;
  assign _EVAL_1740 = _EVAL_2889 == 1'h0;
  assign _EVAL_815 = Queue__EVAL_13;
  assign _EVAL_788 = _EVAL_3991 | LevelGateway_1__EVAL_3;
  assign _EVAL_1070 = _EVAL_1635[97];
  assign _EVAL_1771 = _EVAL_1070 | LevelGateway_96__EVAL_3;
  assign _EVAL_346 = _EVAL_3673 & _EVAL_2567;
  assign _EVAL_1076 = _EVAL_346 & _EVAL_2267;
  assign _EVAL_476 = _EVAL_1635[112];
  assign _EVAL_2698 = _EVAL_476 | LevelGateway_111__EVAL_3;
  assign _EVAL_1386 = _EVAL_1837 & _EVAL_591;
  assign _EVAL_363 = _EVAL_3673 & _EVAL_4040;
  assign _EVAL_2382 = _EVAL_476 == 1'h0;
  assign _EVAL_268 = _EVAL_2999[115];
  assign _EVAL_2827 = _EVAL_231 == 1'h0;
  assign _EVAL_3047 = _EVAL_712 | LevelGateway_25__EVAL_3;
  assign _EVAL_2005 = _EVAL_3687 & _EVAL_2267;
  assign _EVAL_866 = _EVAL_2005 & _EVAL_591;
  assign _EVAL_793 = _EVAL_1635[72];
  assign _EVAL_3553 = _EVAL_1635[115];
  assign _EVAL_3469 = 128'h1 << _EVAL_666;
  assign _EVAL_3491 = _EVAL_1990 ? _EVAL_3469 : 128'h0;
  assign _EVAL_3263 = _EVAL_2144 | LevelGateway_52__EVAL_3;
  assign _EVAL_2430 = _EVAL_1835 == 1'h0;
  assign _EVAL_631 = _EVAL_1549 == 1'h0;
  assign _EVAL_2963 = _EVAL_189 == 1'h0;
  assign _EVAL_1081 = _EVAL_3673 & _EVAL_1325;
  assign _EVAL_1756 = _EVAL_1243 | LevelGateway_54__EVAL_3;
  assign _EVAL_3896 = _EVAL_2126 == 1'h0;
  assign _EVAL_3769 = _EVAL_795 == 1'h0;
  assign _EVAL_3150 = _EVAL_1635[3];
  assign _EVAL_3065 = _EVAL_3150 | LevelGateway_2__EVAL_3;
  assign _EVAL_2017 = _EVAL_3150 == 1'h0;
  assign _EVAL_2058 = _EVAL_879 & _EVAL_591;
  assign _EVAL_1062 = _EVAL_1635[107];
  assign _EVAL_1690 = _EVAL_820 == 1'h0;
  assign _EVAL_780 = _EVAL_1635[40];
  assign _EVAL_395 = _EVAL_3673 & _EVAL_3873;
  assign _EVAL_1175 = _EVAL_1635[45];
  assign _EVAL_3099 = _EVAL_1175 | LevelGateway_44__EVAL_3;
  assign _EVAL_2601 = _EVAL_1175 == 1'h0;
  assign _EVAL_1999 = _EVAL_1070 == 1'h0;
  assign _EVAL_2911 = _EVAL_2686 & _EVAL_2267;
  assign _EVAL_3632 = _EVAL_3959 & _EVAL_2267;
  assign _EVAL_3388 = _EVAL_3673 & _EVAL_2122;
  assign _EVAL_2527 = {_EVAL_3623,_EVAL_1697,_EVAL_2188,_EVAL_2018,_EVAL_1776,_EVAL_2754,_EVAL_2073,_EVAL_1162,_EVAL_3497};
  assign _EVAL_3799 = _EVAL_310 | LevelGateway_18__EVAL_3;
  assign _EVAL_3921 = _EVAL_2125 & _EVAL_2267;
  assign _EVAL_3198 = _EVAL_3921 & _EVAL_591;
  assign _EVAL_2438 = _EVAL_3673 & _EVAL_1531;
  assign _EVAL_1506 = _EVAL_219 == 1'h0;
  assign _EVAL_1550 = _EVAL_1635[111];
  assign _EVAL_2589 = _EVAL_1635[77];
  assign _EVAL_1242 = _EVAL_2589 | LevelGateway_76__EVAL_3;
  assign _EVAL_807 = _EVAL_2229 & _EVAL_2335;
  assign _EVAL_1773 = _EVAL_2229 & _EVAL_187;
  assign _EVAL_2059 = _EVAL_3673 & _EVAL_1216;
  assign _EVAL_3112 = _EVAL_2059 & _EVAL_2267;
  assign _EVAL_2330 = _EVAL_1555 & _EVAL_2267;
  assign _EVAL_796 = _EVAL_2330 & _EVAL_591;
  assign _EVAL_1066 = _EVAL_3673 & _EVAL_1064;
  assign _EVAL_2715 = _EVAL_1066 & _EVAL_2267;
  assign _EVAL_1205 = _EVAL_2715 & _EVAL_591;
  assign _EVAL_3353 = _EVAL_3632 & _EVAL_591;
  assign _EVAL_3314 = _EVAL_3673 & _EVAL_353;
  assign _EVAL_1477 = _EVAL_3673 & _EVAL_1230;
  assign _EVAL_1485 = _EVAL_1477 & _EVAL_2267;
  assign _EVAL_3566 = _EVAL_2279 | LevelGateway_68__EVAL_3;
  assign _EVAL_1769 = _EVAL_3673 & _EVAL_2520;
  assign _EVAL_1899 = _EVAL_1769 & _EVAL_2267;
  assign _EVAL_1571 = _EVAL_2103 == 1'h0;
  assign _EVAL_4028 = _EVAL_2589 == 1'h0;
  assign _EVAL_2739 = _EVAL_263 | LevelGateway_19__EVAL_3;
  assign _EVAL_1815 = _EVAL_2136 == 1'h0;
  assign _EVAL_1737 = _EVAL_3673 & _EVAL_4062;
  assign _EVAL_3433 = _EVAL_1737 & _EVAL_2267;
  assign _EVAL_2511 = _EVAL_3433 & _EVAL_591;
  assign _EVAL_1291 = _EVAL_395 & _EVAL_2267;
  assign _EVAL_682 = _EVAL_1550 | LevelGateway_110__EVAL_3;
  assign _EVAL_3515 = _EVAL_3673 & _EVAL_1439;
  assign _EVAL_3629 = _EVAL_3515 & _EVAL_2267;
  assign _EVAL_2309 = _EVAL_3547 & _EVAL_2267;
  assign _EVAL_2903 = _EVAL_2669 & _EVAL_809;
  assign _EVAL_3890 = _EVAL_2554 | LevelGateway_107__EVAL_3;
  assign _EVAL_3329 = _EVAL_1635[57];
  assign _EVAL_2142 = _EVAL_2187 | LevelGateway_7__EVAL_3;
  assign _EVAL_1094 = _EVAL_3553 | LevelGateway_114__EVAL_3;
  assign _EVAL_2358 = _EVAL_3553 == 1'h0;
  assign _EVAL_1287 = _EVAL_3673 & _EVAL_1833;
  assign _EVAL_1135 = _EVAL_3673 & _EVAL_4041;
  assign _EVAL_867 = _EVAL_1135 & _EVAL_2267;
  assign _EVAL_2150 = _EVAL_3673 & _EVAL_822;
  assign _EVAL_3683 = _EVAL_1289 & _EVAL_591;
  assign _EVAL_1927 = _EVAL_1062 == 1'h0;
  assign _EVAL_3486 = _EVAL_1635[122];
  assign _EVAL_2206 = _EVAL_3486 == 1'h0;
  assign _EVAL_1109 = _EVAL_3673 & _EVAL_260;
  assign _EVAL_3028 = _EVAL_1109 & _EVAL_2267;
  assign _EVAL_3681 = _EVAL_3028 & _EVAL_591;
  assign _EVAL_1725 = _EVAL_1635[92];
  assign _EVAL_2084 = _EVAL_1725 == 1'h0;
  assign _EVAL_3135 = _EVAL_3314 & _EVAL_2267;
  assign _EVAL_1015 = _EVAL_3135 & _EVAL_591;
  assign _EVAL_3045 = _EVAL_1635[116];
  assign _EVAL_2791 = _EVAL_3045 == 1'h0;
  assign _EVAL_3993 = _EVAL_1633 | LevelGateway_3__EVAL_3;
  assign _EVAL_2120 = _EVAL_1635[79];
  assign _EVAL_1540 = _EVAL_2120 | LevelGateway_78__EVAL_3;
  assign _EVAL_1585 = _EVAL_780 | LevelGateway_39__EVAL_3;
  assign _EVAL_3663 = _EVAL_780 == 1'h0;
  assign _EVAL_1966 = _EVAL_2366 & _EVAL_591;
  assign _EVAL_3519 = _EVAL_3329 | LevelGateway_56__EVAL_3;
  assign _EVAL_1596 = _EVAL_2854 == 1'h0;
  assign _EVAL_1434 = _EVAL_585 == 1'h0;
  assign _EVAL_2257 = _EVAL_1677 & _EVAL_2267;
  assign _EVAL_447 = _EVAL_1635[83];
  assign _EVAL_1758 = _EVAL_447 | LevelGateway_82__EVAL_3;
  assign _EVAL_3410 = _EVAL_363 & _EVAL_2267;
  assign _EVAL_1063 = _EVAL_1635[100];
  assign _EVAL_1144 = _EVAL_1063 | LevelGateway_99__EVAL_3;
  assign _EVAL_2885 = _EVAL_1063 == 1'h0;
  assign _EVAL_2117 = _EVAL_1635[34];
  assign _EVAL_1333 = _EVAL_2117 | LevelGateway_33__EVAL_3;
  assign _EVAL_2786 = _EVAL_2117 == 1'h0;
  assign _EVAL_2163 = _EVAL_1550 == 1'h0;
  assign _EVAL_1827 = _EVAL_1635[80];
  assign _EVAL_473 = _EVAL_1827 == 1'h0;
  assign _EVAL_2767 = _EVAL_1635[124];
  assign _EVAL_2704 = _EVAL_2767 | LevelGateway_123__EVAL_3;
  assign _EVAL_968 = _EVAL_2767 == 1'h0;
  assign _EVAL_479 = _EVAL_3112 & _EVAL_591;
  assign _EVAL_2764 = _EVAL_1635[61];
  assign _EVAL_864 = _EVAL_2764 | LevelGateway_60__EVAL_3;
  assign _EVAL_3013 = _EVAL_2764 == 1'h0;
  assign _EVAL_1640 = 10'h1 == _EVAL_1450;
  assign _EVAL_3710 = _EVAL_1338 ? _EVAL_2267 : _EVAL_229;
  assign _EVAL_1190 = _EVAL_1640 ? _EVAL_2267 : _EVAL_3710;
  assign _EVAL_2639 = _EVAL_2669 & _EVAL_187;
  assign _EVAL_3186 = _EVAL_1635[50];
  assign _EVAL_171 = _EVAL_3186 | LevelGateway_49__EVAL_3;
  assign _EVAL_3677 = _EVAL_3186 == 1'h0;
  assign _EVAL_2588 = _EVAL_3673 & _EVAL_1533;
  assign _EVAL_718 = _EVAL_2588 & _EVAL_2267;
  assign _EVAL_1472 = _EVAL_1408 & _EVAL_591;
  assign _EVAL_2913 = _EVAL_3045 | LevelGateway_115__EVAL_3;
  assign _EVAL_797 = _EVAL_1635[16];
  assign _EVAL_3749 = _EVAL_797 | LevelGateway_15__EVAL_3;
  assign _EVAL_2593 = _EVAL_797 == 1'h0;
  assign _EVAL_2425 = _EVAL_1704 == 1'h0;
  assign _EVAL_3351 = _EVAL_3673 & _EVAL_2189;
  assign _EVAL_450 = _EVAL_3351 & _EVAL_2267;
  assign _EVAL_1799 = _EVAL_2126 | LevelGateway_63__EVAL_3;
  assign _EVAL_2316 = _EVAL_447 == 1'h0;
  assign _EVAL_3139 = _EVAL_1635[91];
  assign _EVAL_3426 = _EVAL_3139 | LevelGateway_90__EVAL_3;
  assign _EVAL_2064 = _EVAL_3139 == 1'h0;
  assign _EVAL_2404 = _EVAL_3756 == 1'h0;
  assign _EVAL_2597 = _EVAL_4043 == 1'h0;
  assign _EVAL_986 = _EVAL_1992 | LevelGateway_74__EVAL_3;
  assign _EVAL_3719 = _EVAL_3673 & _EVAL_1113;
  assign _EVAL_4010 = _EVAL_3719 & _EVAL_2267;
  assign _EVAL_3997 = _EVAL_4010 & _EVAL_591;
  assign _EVAL_2408 = _EVAL_3220 & _EVAL_591;
  assign _EVAL_1178 = _EVAL_1068 & _EVAL_591;
  assign _EVAL_1465 = _EVAL_203 | LevelGateway_41__EVAL_3;
  assign _EVAL_1845 = _EVAL_1243 == 1'h0;
  assign _EVAL_299 = _EVAL_1725 | LevelGateway_91__EVAL_3;
  assign _EVAL_2109 = _EVAL_3930 & _EVAL_591;
  assign _EVAL_2037 = _EVAL_1287 & _EVAL_2267;
  assign _EVAL_391 = _EVAL_2037 & _EVAL_591;
  assign _EVAL_1449 = _EVAL_3584 & _EVAL_2267;
  assign _EVAL_3774 = _EVAL_1449 & _EVAL_591;
  assign _EVAL_341 = _EVAL_3329 == 1'h0;
  assign _EVAL_2581 = _EVAL_1069 & _EVAL_2267;
  assign _EVAL_1311 = _EVAL_2581 & _EVAL_591;
  assign _EVAL_3796 = _EVAL_2454 | LevelGateway_88__EVAL_3;
  assign _EVAL_1093 = _EVAL_219 | LevelGateway_21__EVAL_3;
  assign _EVAL_2654 = _EVAL_1291 & _EVAL_591;
  assign _EVAL_3456 = _EVAL_3629 & _EVAL_591;
  assign _EVAL_3842 = _EVAL_1503 & _EVAL_591;
  assign _EVAL_1728 = _EVAL_2309 & _EVAL_591;
  assign _EVAL_2411 = _EVAL_2131 & _EVAL_591;
  assign _EVAL_2015 = _EVAL_1076 & _EVAL_591;
  assign _EVAL_2563 = _EVAL_2669 & _EVAL_2354;
  assign _EVAL_1559 = _EVAL_3529 == 1'h0;
  assign _EVAL_1246 = _EVAL_2782 | LevelGateway_93__EVAL_3;
  assign _EVAL_1244 = _EVAL_2333 == 1'h0;
  assign _EVAL_1042 = _EVAL_2579 & _EVAL_591;
  assign _EVAL_3751 = _EVAL_1890 == 1'h0;
  assign _EVAL_3650 = _EVAL_1527 & _EVAL_591;
  assign _EVAL_2070 = _EVAL_3673 & _EVAL_2743;
  assign _EVAL_2806 = _EVAL_2070 & _EVAL_2267;
  assign _EVAL_3020 = Queue__EVAL[23:16];
  assign _EVAL_3724 = _EVAL_1635[23];
  assign _EVAL_2590 = _EVAL_3724 | LevelGateway_22__EVAL_3;
  assign _EVAL_3284 = _EVAL_1297 & _EVAL_591;
  assign _EVAL_1378 = _EVAL_2229 & _EVAL_2354;
  assign _EVAL_3214 = _EVAL_606 & _EVAL_591;
  assign _EVAL_570 = _EVAL_793 == 1'h0;
  assign _EVAL_3998 = _EVAL_1085 & _EVAL_591;
  assign _EVAL_2218 = _EVAL_2532 & _EVAL_591;
  assign _EVAL_706 = _EVAL_3823 & _EVAL_591;
  assign _EVAL_4027 = _EVAL_1640 ? {{29'd0}, _EVAL_1156} : _EVAL_1802;
  assign _EVAL_688 = Queue__EVAL[7:0];
  assign _EVAL_2099 = _EVAL_718 & _EVAL_591;
  assign _EVAL_541 = _EVAL_899 & _EVAL_591;
  assign _EVAL_1139 = _EVAL_830 & _EVAL_591;
  assign _EVAL_1157 = _EVAL_2806 & _EVAL_591;
  assign _EVAL_2909 = _EVAL_3388 & _EVAL_2267;
  assign _EVAL_1218 = _EVAL_3504 & _EVAL_2267;
  assign _EVAL_4061 = _EVAL_1218 & _EVAL_591;
  assign _EVAL_3191 = _EVAL_207 & _EVAL_591;
  assign _EVAL_3281 = _EVAL_3434 == 1'h0;
  assign _EVAL_1251 = _EVAL_1633 == 1'h0;
  assign _EVAL_2278 = _EVAL_1915 | LevelGateway_6__EVAL_3;
  assign _EVAL_214 = _EVAL_2167 | LevelGateway_65__EVAL_3;
  assign _EVAL_3892 = _EVAL_2554 == 1'h0;
  assign _EVAL_3005 = _EVAL_505 & _EVAL_591;
  assign _EVAL_2898 = _EVAL_3184 == 1'h0;
  assign _EVAL_1461 = _EVAL_994 & _EVAL_591;
  assign _EVAL_3543 = _EVAL_2682 & _EVAL_2267;
  assign _EVAL_3275 = _EVAL_3952 | LevelGateway_32__EVAL_3;
  assign _EVAL_1998 = _EVAL_1019 & _EVAL_591;
  assign _EVAL_2751 = _EVAL_2120 == 1'h0;
  assign _EVAL_2785 = _EVAL_450 & _EVAL_591;
  assign _EVAL_3649 = _EVAL_540 == 1'h0;
  assign _EVAL_1632 = _EVAL_1827 | LevelGateway_79__EVAL_3;
  assign _EVAL_3669 = _EVAL_2438 & _EVAL_2267;
  assign _EVAL_1874 = _EVAL_2557 & _EVAL_2267;
  assign _EVAL_1082 = _EVAL_1874 & _EVAL_591;
  assign _EVAL_3766 = _EVAL_3724 == 1'h0;
  assign _EVAL_3070 = _EVAL_1856 == 1'h0;
  assign _EVAL_1479 = _EVAL_2167 == 1'h0;
  assign _EVAL_2737 = _EVAL_1002 | LevelGateway_100__EVAL_3;
  assign _EVAL_457 = _EVAL_1062 | LevelGateway_106__EVAL_3;
  assign _EVAL_1134 = _EVAL_1509 & _EVAL_2267;
  assign _EVAL_3738 = _EVAL_1134 & _EVAL_591;
  assign _EVAL_3356 = _EVAL_3509 == 1'h0;
  assign _EVAL_2603 = _EVAL_3410 & _EVAL_591;
  assign _EVAL_3495 = _EVAL_3136 & _EVAL_2267;
  assign _EVAL_1403 = _EVAL_3495 & _EVAL_591;
  assign _EVAL_1591 = _EVAL_2909 & _EVAL_591;
  assign _EVAL_1510 = _EVAL_2514 & _EVAL_591;
  assign _EVAL_3583 = _EVAL_732 & _EVAL_591;
  assign _EVAL_298 = _EVAL_3669 & _EVAL_591;
  assign _EVAL_2160 = _EVAL_1899 & _EVAL_591;
  assign _EVAL_2261 = _EVAL_2388 == 1'h0;
  assign _EVAL_1453 = _EVAL_3952 == 1'h0;
  assign _EVAL_1197 = _EVAL_3166 & _EVAL_2267;
  assign _EVAL_1863 = _EVAL_3673 & _EVAL_268;
  assign _EVAL_2198 = _EVAL_1863 & _EVAL_2267;
  assign _EVAL_2844 = _EVAL_1730 == 1'h0;
  assign _EVAL_1187 = _EVAL_2257 & _EVAL_591;
  assign _EVAL_608 = _EVAL_793 | LevelGateway_71__EVAL_3;
  assign _EVAL_816 = _EVAL_2150 & _EVAL_2267;
  assign _EVAL_3103 = _EVAL_816 & _EVAL_591;
  assign _EVAL_359 = _EVAL_2198 & _EVAL_591;
  assign _EVAL_182 = _EVAL_1768 & _EVAL_591;
  assign _EVAL_1918 = _EVAL_1081 & _EVAL_2267;
  assign _EVAL_651 = _EVAL_1918 & _EVAL_591;
  assign _EVAL_3939 = _EVAL_2911 & _EVAL_591;
  assign _EVAL_1663 = _EVAL_2669 & _EVAL_2335;
  assign _EVAL_3764 = _EVAL_1839 & _EVAL_591;
  assign _EVAL_2776 = _EVAL_2559 & _EVAL_187;
  assign _EVAL_1446 = _EVAL_1200 & _EVAL_591;
  assign _EVAL_1025 = _EVAL_1485 & _EVAL_591;
  assign _EVAL_2729 = _EVAL_867 & _EVAL_591;
  assign _EVAL_1159 = _EVAL_3688 | LevelGateway_87__EVAL_3;
  assign _EVAL_3581 = _EVAL_3486 | LevelGateway_121__EVAL_3;
  assign _EVAL_1861 = Queue__EVAL[15:8];
  assign _EVAL_975 = _EVAL_3543 & _EVAL_591;
  assign _EVAL_2439 = _EVAL_632 & _EVAL_591;
  assign _EVAL_2663 = _EVAL_3659 & _EVAL_591;
  assign _EVAL_576 = _EVAL_981 & _EVAL_591;
  assign _EVAL_1271 = _EVAL_1197 & _EVAL_591;
  assign _EVAL_1842 = _EVAL_1848 & _EVAL_591;
  assign _EVAL_2744 = _EVAL_2981 & _EVAL_591;
  assign _EVAL_3965 = Queue__EVAL[2:0];
  assign LevelGateway_32__EVAL_2 = _EVAL_105;
  assign LevelGateway_102__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_62 = _EVAL_2536;
  assign PLICFanIn__EVAL_49 = _EVAL_1819;
  assign LevelGateway_104__EVAL_0 = _EVAL_3199 == 1'h0;
  assign LevelGateway_40__EVAL = _EVAL_3491[41];
  assign LevelGateway_6__EVAL_1 = _EVAL_71;
  assign LevelGateway_99__EVAL_0 = _EVAL_3296 == 1'h0;
  assign LevelGateway_25__EVAL_1 = _EVAL_29;
  assign LevelGateway_119__EVAL = _EVAL_3491[120];
  assign LevelGateway_97__EVAL_2 = _EVAL_105;
  assign LevelGateway_17__EVAL_1 = _EVAL_96;
  assign LevelGateway_68__EVAL = _EVAL_3491[69];
  assign PLICFanIn__EVAL_109 = _EVAL_2677;
  assign LevelGateway_80__EVAL_4 = _EVAL_142;
  assign LevelGateway_49__EVAL_1 = _EVAL_22;
  assign LevelGateway_108__EVAL = _EVAL_3491[109];
  assign LevelGateway_56__EVAL_1 = _EVAL_90;
  assign LevelGateway_18__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_29 = _EVAL_1088;
  assign LevelGateway_11__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_40 = _EVAL_1870;
  assign LevelGateway_78__EVAL = _EVAL_3491[79];
  assign LevelGateway_5__EVAL_2 = _EVAL_105;
  assign LevelGateway_16__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_127 = _EVAL_3118;
  assign LevelGateway_87__EVAL = _EVAL_3491[88];
  assign LevelGateway_22__EVAL_2 = _EVAL_105;
  assign LevelGateway_48__EVAL_0 = _EVAL_222 == 1'h0;
  assign LevelGateway_121__EVAL_2 = _EVAL_105;
  assign LevelGateway_32__EVAL_1 = _EVAL_133;
  assign LevelGateway_117__EVAL_1 = _EVAL_45;
  assign LevelGateway_97__EVAL_4 = _EVAL_142;
  assign LevelGateway_109__EVAL_1 = _EVAL_81;
  assign LevelGateway_57__EVAL_0 = _EVAL_1206 == 1'h0;
  assign LevelGateway_58__EVAL_1 = _EVAL_123;
  assign LevelGateway_94__EVAL = _EVAL_3491[95];
  assign LevelGateway_114__EVAL_2 = _EVAL_105;
  assign LevelGateway_42__EVAL_0 = _EVAL_3899 == 1'h0;
  assign LevelGateway_71__EVAL_0 = _EVAL_3039 == 1'h0;
  assign PLICFanIn__EVAL_108 = _EVAL_251;
  assign LevelGateway_60__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_103 = _EVAL_285;
  assign LevelGateway_70__EVAL_0 = _EVAL_552 == 1'h0;
  assign PLICFanIn__EVAL_34 = _EVAL_1680;
  assign LevelGateway_32__EVAL_0 = _EVAL_462 == 1'h0;
  assign LevelGateway_89__EVAL_4 = _EVAL_142;
  assign LevelGateway_113__EVAL_1 = _EVAL_41;
  assign LevelGateway_12__EVAL_0 = _EVAL_3636 == 1'h0;
  assign LevelGateway_10__EVAL_4 = _EVAL_142;
  assign LevelGateway_43__EVAL = _EVAL_3491[44];
  assign PLICFanIn__EVAL_69 = _EVAL_1239;
  assign LevelGateway_52__EVAL_1 = _EVAL_23;
  assign LevelGateway_35__EVAL_4 = _EVAL_142;
  assign LevelGateway_2__EVAL_0 = _EVAL_371 == 1'h0;
  assign LevelGateway_106__EVAL_1 = _EVAL_82;
  assign LevelGateway_11__EVAL_2 = _EVAL_105;
  assign LevelGateway_75__EVAL_0 = _EVAL_1930 == 1'h0;
  assign LevelGateway_90__EVAL = _EVAL_3491[91];
  assign LevelGateway_31__EVAL_1 = _EVAL_113;
  assign LevelGateway_6__EVAL = _EVAL_3491[7];
  assign LevelGateway_120__EVAL_4 = _EVAL_142;
  assign LevelGateway_49__EVAL_0 = _EVAL_3720 == 1'h0;
  assign LevelGateway_94__EVAL_1 = _EVAL_122;
  assign PLICFanIn__EVAL_51 = _EVAL_3336;
  assign PLICFanIn__EVAL_39 = _EVAL_331;
  assign LevelGateway_71__EVAL_1 = _EVAL_24;
  assign PLICFanIn__EVAL_98 = _EVAL_444;
  assign LevelGateway_50__EVAL_2 = _EVAL_105;
  assign LevelGateway_100__EVAL_2 = _EVAL_105;
  assign LevelGateway_35__EVAL_1 = _EVAL_2;
  assign _EVAL_130 = _EVAL_1190 ? _EVAL_4027 : 32'h0;
  assign LevelGateway_101__EVAL_1 = _EVAL_85;
  assign LevelGateway_59__EVAL_0 = _EVAL_2648 == 1'h0;
  assign LevelGateway_76__EVAL_0 = _EVAL_212 == 1'h0;
  assign LevelGateway_8__EVAL_4 = _EVAL_142;
  assign LevelGateway_67__EVAL_0 = _EVAL_421 == 1'h0;
  assign LevelGateway_103__EVAL_4 = _EVAL_142;
  assign LevelGateway_81__EVAL = _EVAL_3491[82];
  assign LevelGateway_94__EVAL_2 = _EVAL_105;
  assign LevelGateway_41__EVAL_0 = _EVAL_2155 == 1'h0;
  assign LevelGateway_55__EVAL = _EVAL_3491[56];
  assign LevelGateway_48__EVAL_4 = _EVAL_142;
  assign LevelGateway_22__EVAL_4 = _EVAL_142;
  assign LevelGateway_27__EVAL_0 = _EVAL_3505 == 1'h0;
  assign LevelGateway__EVAL_0 = _EVAL_2133 == 1'h0;
  assign LevelGateway_116__EVAL_2 = _EVAL_105;
  assign LevelGateway_91__EVAL_2 = _EVAL_105;
  assign LevelGateway_126__EVAL_2 = _EVAL_105;
  assign LevelGateway_64__EVAL_4 = _EVAL_142;
  assign LevelGateway_123__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_104 = _EVAL_2110;
  assign LevelGateway_64__EVAL_1 = _EVAL_53;
  assign LevelGateway_85__EVAL_0 = _EVAL_3245 == 1'h0;
  assign LevelGateway_91__EVAL_0 = _EVAL_3279 == 1'h0;
  assign LevelGateway_116__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_20 = _EVAL_2035;
  assign LevelGateway_28__EVAL_4 = _EVAL_142;
  assign LevelGateway_36__EVAL_4 = _EVAL_142;
  assign LevelGateway_111__EVAL_1 = _EVAL_110;
  assign LevelGateway_57__EVAL = _EVAL_3491[58];
  assign PLICFanIn__EVAL_74 = _EVAL_3645;
  assign LevelGateway_91__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_118 = _EVAL_2965;
  assign LevelGateway_59__EVAL = _EVAL_3491[60];
  assign LevelGateway_22__EVAL = _EVAL_3491[23];
  assign LevelGateway_12__EVAL_1 = _EVAL_139;
  assign LevelGateway_2__EVAL_4 = _EVAL_142;
  assign LevelGateway_101__EVAL = _EVAL_3491[102];
  assign LevelGateway_47__EVAL_4 = _EVAL_142;
  assign LevelGateway_44__EVAL_1 = _EVAL_64;
  assign LevelGateway_1__EVAL_0 = _EVAL_2209 == 1'h0;
  assign PLICFanIn__EVAL_17 = _EVAL_3731;
  assign LevelGateway_40__EVAL_4 = _EVAL_142;
  assign LevelGateway_101__EVAL_0 = _EVAL_3283 == 1'h0;
  assign PLICFanIn__EVAL_0 = _EVAL_648;
  assign LevelGateway_102__EVAL_0 = _EVAL_194 == 1'h0;
  assign LevelGateway_110__EVAL = _EVAL_3491[111];
  assign LevelGateway_77__EVAL_1 = _EVAL_141;
  assign LevelGateway_73__EVAL_0 = _EVAL_2159 == 1'h0;
  assign LevelGateway_39__EVAL = _EVAL_3491[40];
  assign LevelGateway_83__EVAL = _EVAL_3491[84];
  assign LevelGateway_48__EVAL_1 = _EVAL_30;
  assign PLICFanIn__EVAL_48 = _EVAL_4066;
  assign PLICFanIn__EVAL_122 = _EVAL_2484;
  assign LevelGateway_81__EVAL_0 = _EVAL_3299 == 1'h0;
  assign LevelGateway_109__EVAL_2 = _EVAL_105;
  assign LevelGateway_31__EVAL_4 = _EVAL_142;
  assign LevelGateway_6__EVAL_2 = _EVAL_105;
  assign LevelGateway_84__EVAL_1 = _EVAL_21;
  assign LevelGateway_122__EVAL_4 = _EVAL_142;
  assign LevelGateway_9__EVAL_0 = _EVAL_673 == 1'h0;
  assign _EVAL_138 = _EVAL_1444 > _EVAL_663;
  assign LevelGateway_6__EVAL_4 = _EVAL_142;
  assign LevelGateway_60__EVAL_4 = _EVAL_142;
  assign LevelGateway_106__EVAL_2 = _EVAL_105;
  assign LevelGateway_51__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_45 = _EVAL_1980;
  assign LevelGateway_23__EVAL_2 = _EVAL_105;
  assign LevelGateway_54__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_81 = _EVAL_3571;
  assign LevelGateway_5__EVAL_4 = _EVAL_142;
  assign LevelGateway_17__EVAL = _EVAL_3491[18];
  assign PLICFanIn__EVAL_67 = _EVAL_1786;
  assign LevelGateway_39__EVAL_1 = _EVAL_124;
  assign LevelGateway_49__EVAL_4 = _EVAL_142;
  assign LevelGateway_100__EVAL = _EVAL_3491[101];
  assign LevelGateway_98__EVAL_0 = _EVAL_770 == 1'h0;
  assign LevelGateway_63__EVAL_2 = _EVAL_105;
  assign LevelGateway_103__EVAL_0 = _EVAL_3964 == 1'h0;
  assign LevelGateway_102__EVAL_4 = _EVAL_142;
  assign LevelGateway_80__EVAL = _EVAL_3491[81];
  assign LevelGateway_99__EVAL = _EVAL_3491[100];
  assign LevelGateway_85__EVAL_1 = _EVAL_31;
  assign PLICFanIn__EVAL_30 = _EVAL_675;
  assign LevelGateway_32__EVAL_4 = _EVAL_142;
  assign LevelGateway_99__EVAL_1 = _EVAL_18;
  assign LevelGateway_107__EVAL = _EVAL_3491[108];
  assign LevelGateway_17__EVAL_4 = _EVAL_142;
  assign LevelGateway_98__EVAL = _EVAL_3491[99];
  assign LevelGateway_88__EVAL_1 = _EVAL_42;
  assign LevelGateway_95__EVAL_2 = _EVAL_105;
  assign LevelGateway_47__EVAL_1 = _EVAL_87;
  assign LevelGateway_117__EVAL_4 = _EVAL_142;
  assign LevelGateway_40__EVAL_0 = _EVAL_3407 == 1'h0;
  assign LevelGateway_55__EVAL_2 = _EVAL_105;
  assign LevelGateway_114__EVAL_0 = _EVAL_1753 == 1'h0;
  assign PLICFanIn__EVAL_107 = _EVAL_2481;
  assign LevelGateway_69__EVAL_1 = _EVAL_25;
  assign LevelGateway_3__EVAL_2 = _EVAL_105;
  assign LevelGateway_31__EVAL = _EVAL_3491[32];
  assign PLICFanIn__EVAL_9 = _EVAL_2491;
  assign LevelGateway_8__EVAL_0 = _EVAL_200 == 1'h0;
  assign LevelGateway_98__EVAL_4 = _EVAL_142;
  assign LevelGateway_35__EVAL = _EVAL_3491[36];
  assign LevelGateway_83__EVAL_2 = _EVAL_105;
  assign LevelGateway_16__EVAL_0 = _EVAL_2128 == 1'h0;
  assign LevelGateway_93__EVAL_0 = _EVAL_3788 == 1'h0;
  assign LevelGateway_87__EVAL_0 = _EVAL_2972 == 1'h0;
  assign LevelGateway_33__EVAL_1 = _EVAL_70;
  assign LevelGateway_54__EVAL_0 = _EVAL_2688 == 1'h0;
  assign LevelGateway_117__EVAL_0 = _EVAL_519 == 1'h0;
  assign LevelGateway_111__EVAL_0 = _EVAL_1496 == 1'h0;
  assign PLICFanIn__EVAL_31 = _EVAL_3056;
  assign LevelGateway_118__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL = _EVAL_2290;
  assign LevelGateway_81__EVAL_1 = _EVAL_118;
  assign LevelGateway_120__EVAL_0 = _EVAL_741 == 1'h0;
  assign PLICFanIn__EVAL_82 = _EVAL_155;
  assign LevelGateway_61__EVAL_1 = _EVAL_78;
  assign LevelGateway_6__EVAL_0 = _EVAL_1788 == 1'h0;
  assign LevelGateway_63__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_25 = _EVAL_1127;
  assign LevelGateway_16__EVAL_2 = _EVAL_105;
  assign LevelGateway_97__EVAL_0 = _EVAL_2838 == 1'h0;
  assign PLICFanIn__EVAL_88 = _EVAL_1962;
  assign PLICFanIn__EVAL_4 = _EVAL_354;
  assign LevelGateway_7__EVAL_0 = _EVAL_2807 == 1'h0;
  assign LevelGateway_88__EVAL_0 = _EVAL_1270 == 1'h0;
  assign PLICFanIn__EVAL_72 = _EVAL_3909;
  assign PLICFanIn__EVAL_113 = _EVAL_2527 & _EVAL_3572;
  assign LevelGateway_1__EVAL_1 = _EVAL_116;
  assign PLICFanIn__EVAL_42 = _EVAL_3721;
  assign LevelGateway_34__EVAL = _EVAL_3491[35];
  assign LevelGateway_120__EVAL_2 = _EVAL_105;
  assign LevelGateway__EVAL = _EVAL_3491[1];
  assign LevelGateway_24__EVAL_1 = _EVAL_80;
  assign LevelGateway_113__EVAL_4 = _EVAL_142;
  assign LevelGateway_108__EVAL_0 = _EVAL_176 == 1'h0;
  assign PLICFanIn__EVAL_128 = _EVAL_548;
  assign LevelGateway_46__EVAL_4 = _EVAL_142;
  assign LevelGateway_47__EVAL = _EVAL_3491[48];
  assign LevelGateway_104__EVAL_2 = _EVAL_105;
  assign LevelGateway_100__EVAL_0 = _EVAL_912 == 1'h0;
  assign LevelGateway_107__EVAL_0 = _EVAL_2942 == 1'h0;
  assign LevelGateway_21__EVAL_4 = _EVAL_142;
  assign LevelGateway_50__EVAL = _EVAL_3491[51];
  assign LevelGateway_45__EVAL_0 = _EVAL_3715 == 1'h0;
  assign LevelGateway_44__EVAL_2 = _EVAL_105;
  assign LevelGateway_86__EVAL_1 = _EVAL_83;
  assign LevelGateway_36__EVAL_2 = _EVAL_105;
  assign LevelGateway_108__EVAL_2 = _EVAL_105;
  assign LevelGateway_79__EVAL_0 = _EVAL_1580 == 1'h0;
  assign LevelGateway_73__EVAL_1 = _EVAL_65;
  assign LevelGateway_72__EVAL_1 = _EVAL_92;
  assign PLICFanIn__EVAL_60 = _EVAL_762;
  assign PLICFanIn__EVAL_47 = _EVAL_2937;
  assign LevelGateway_84__EVAL_2 = _EVAL_105;
  assign LevelGateway_23__EVAL_0 = _EVAL_614 == 1'h0;
  assign PLICFanIn__EVAL_15 = _EVAL_2760;
  assign LevelGateway_105__EVAL = _EVAL_3491[106];
  assign LevelGateway__EVAL_1 = _EVAL_127;
  assign LevelGateway_48__EVAL_2 = _EVAL_105;
  assign LevelGateway_25__EVAL_0 = _EVAL_387 == 1'h0;
  assign LevelGateway_46__EVAL_2 = _EVAL_105;
  assign LevelGateway_74__EVAL_1 = _EVAL_50;
  assign LevelGateway_30__EVAL_2 = _EVAL_105;
  assign LevelGateway_53__EVAL_2 = _EVAL_105;
  assign LevelGateway_122__EVAL = _EVAL_3491[123];
  assign LevelGateway_56__EVAL_4 = _EVAL_142;
  assign LevelGateway_74__EVAL = _EVAL_3491[75];
  assign LevelGateway_111__EVAL = _EVAL_3491[112];
  assign LevelGateway_23__EVAL_1 = _EVAL_4;
  assign LevelGateway_59__EVAL_1 = _EVAL_93;
  assign LevelGateway_80__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_28 = _EVAL_2111;
  assign LevelGateway_73__EVAL = _EVAL_3491[74];
  assign LevelGateway_41__EVAL_2 = _EVAL_105;
  assign LevelGateway_68__EVAL_2 = _EVAL_105;
  assign LevelGateway_67__EVAL_2 = _EVAL_105;
  assign LevelGateway_67__EVAL_1 = _EVAL_88;
  assign LevelGateway_96__EVAL = _EVAL_3491[97];
  assign LevelGateway_14__EVAL_2 = _EVAL_105;
  assign LevelGateway_33__EVAL_0 = _EVAL_1315 == 1'h0;
  assign LevelGateway_19__EVAL = _EVAL_3491[20];
  assign LevelGateway_82__EVAL_4 = _EVAL_142;
  assign LevelGateway_65__EVAL_0 = _EVAL_4034 == 1'h0;
  assign LevelGateway_58__EVAL = _EVAL_3491[59];
  assign LevelGateway_29__EVAL = _EVAL_3491[30];
  assign Queue__EVAL_11 = _EVAL_105;
  assign LevelGateway_69__EVAL_0 = _EVAL_3023 == 1'h0;
  assign LevelGateway_125__EVAL_1 = _EVAL_95;
  assign LevelGateway_53__EVAL_4 = _EVAL_142;
  assign LevelGateway_10__EVAL_0 = _EVAL_1979 == 1'h0;
  assign LevelGateway_7__EVAL_1 = _EVAL_46;
  assign LevelGateway_75__EVAL_1 = _EVAL_100;
  assign LevelGateway_44__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_93 = _EVAL_4013;
  assign LevelGateway_103__EVAL_1 = _EVAL_106;
  assign LevelGateway_86__EVAL = _EVAL_3491[87];
  assign LevelGateway_19__EVAL_1 = _EVAL_97;
  assign LevelGateway_122__EVAL_1 = _EVAL_27;
  assign LevelGateway_12__EVAL_2 = _EVAL_105;
  assign LevelGateway_46__EVAL_1 = _EVAL_48;
  assign LevelGateway_118__EVAL = _EVAL_3491[119];
  assign PLICFanIn__EVAL_77 = _EVAL_3216;
  assign LevelGateway_50__EVAL_0 = _EVAL_1313 == 1'h0;
  assign PLICFanIn__EVAL_54 = _EVAL_2306;
  assign LevelGateway_100__EVAL_1 = _EVAL_10;
  assign LevelGateway_103__EVAL = _EVAL_3491[104];
  assign LevelGateway_11__EVAL_1 = _EVAL_44;
  assign PLICFanIn__EVAL_75 = _EVAL_2055;
  assign LevelGateway_117__EVAL_2 = _EVAL_105;
  assign LevelGateway_21__EVAL_0 = _EVAL_217 == 1'h0;
  assign LevelGateway_53__EVAL_0 = _EVAL_2582 == 1'h0;
  assign LevelGateway_78__EVAL_0 = _EVAL_2850 == 1'h0;
  assign LevelGateway_58__EVAL_4 = _EVAL_142;
  assign LevelGateway_21__EVAL = _EVAL_3491[22];
  assign LevelGateway_31__EVAL_2 = _EVAL_105;
  assign LevelGateway_111__EVAL_2 = _EVAL_105;
  assign LevelGateway_4__EVAL_4 = _EVAL_142;
  assign LevelGateway_49__EVAL = _EVAL_3491[50];
  assign LevelGateway_112__EVAL_4 = _EVAL_142;
  assign LevelGateway_8__EVAL = _EVAL_3491[9];
  assign LevelGateway_37__EVAL_0 = _EVAL_2684 == 1'h0;
  assign LevelGateway_11__EVAL_0 = _EVAL_3750 == 1'h0;
  assign LevelGateway_52__EVAL = _EVAL_3491[53];
  assign PLICFanIn__EVAL_70 = _EVAL_2334;
  assign LevelGateway_61__EVAL = _EVAL_3491[62];
  assign LevelGateway_39__EVAL_0 = _EVAL_1929 == 1'h0;
  assign PLICFanIn__EVAL_52 = _EVAL_3843;
  assign LevelGateway_60__EVAL_1 = _EVAL_7;
  assign LevelGateway_29__EVAL_0 = _EVAL_1597 == 1'h0;
  assign LevelGateway_13__EVAL_4 = _EVAL_142;
  assign LevelGateway_24__EVAL_4 = _EVAL_142;
  assign LevelGateway_105__EVAL_0 = _EVAL_569 == 1'h0;
  assign LevelGateway_13__EVAL_1 = _EVAL_76;
  assign LevelGateway_56__EVAL_0 = _EVAL_3527 == 1'h0;
  assign LevelGateway_15__EVAL = _EVAL_3491[16];
  assign LevelGateway_39__EVAL_4 = _EVAL_142;
  assign LevelGateway_24__EVAL_0 = _EVAL_306 == 1'h0;
  assign PLICFanIn__EVAL_26 = _EVAL_247;
  assign LevelGateway_26__EVAL_2 = _EVAL_105;
  assign LevelGateway_54__EVAL_2 = _EVAL_105;
  assign LevelGateway_107__EVAL_2 = _EVAL_105;
  assign LevelGateway_78__EVAL_4 = _EVAL_142;
  assign LevelGateway_49__EVAL_2 = _EVAL_105;
  assign LevelGateway_119__EVAL_2 = _EVAL_105;
  assign LevelGateway_18__EVAL_2 = _EVAL_105;
  assign LevelGateway_77__EVAL_0 = _EVAL_880 == 1'h0;
  assign PLICFanIn__EVAL_73 = _EVAL_3267;
  assign LevelGateway_3__EVAL = _EVAL_3491[4];
  assign LevelGateway_66__EVAL_1 = _EVAL_89;
  assign LevelGateway_15__EVAL_0 = _EVAL_581 == 1'h0;
  assign LevelGateway_50__EVAL_1 = _EVAL_54;
  assign LevelGateway_92__EVAL_2 = _EVAL_105;
  assign LevelGateway_9__EVAL_4 = _EVAL_142;
  assign LevelGateway_30__EVAL_0 = _EVAL_3222 == 1'h0;
  assign LevelGateway_118__EVAL_2 = _EVAL_105;
  assign LevelGateway_115__EVAL_1 = _EVAL_40;
  assign PLICFanIn__EVAL_10 = _EVAL_3195;
  assign PLICFanIn__EVAL_64 = _EVAL_3331;
  assign LevelGateway_9__EVAL = _EVAL_3491[10];
  assign LevelGateway_1__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_97 = _EVAL_1142;
  assign LevelGateway_46__EVAL_0 = _EVAL_1709 == 1'h0;
  assign LevelGateway_82__EVAL_0 = _EVAL_1261 == 1'h0;
  assign LevelGateway_82__EVAL_1 = _EVAL_8;
  assign LevelGateway_28__EVAL_2 = _EVAL_105;
  assign LevelGateway_18__EVAL_0 = _EVAL_2666 == 1'h0;
  assign PLICFanIn__EVAL_63 = _EVAL_3552;
  assign _EVAL_15 = Queue__EVAL_12;
  assign LevelGateway_92__EVAL_0 = _EVAL_3783 == 1'h0;
  assign LevelGateway_123__EVAL_4 = _EVAL_142;
  assign LevelGateway_53__EVAL = _EVAL_3491[54];
  assign LevelGateway_90__EVAL_1 = _EVAL_140;
  assign LevelGateway_68__EVAL_4 = _EVAL_142;
  assign LevelGateway_106__EVAL_4 = _EVAL_142;
  assign LevelGateway_93__EVAL = _EVAL_3491[94];
  assign LevelGateway_91__EVAL = _EVAL_3491[92];
  assign PLICFanIn__EVAL_119 = _EVAL_3014;
  assign LevelGateway_58__EVAL_0 = _EVAL_3137 == 1'h0;
  assign LevelGateway_109__EVAL = _EVAL_3491[110];
  assign PLICFanIn__EVAL_94 = _EVAL_4050;
  assign LevelGateway_42__EVAL_1 = _EVAL_115;
  assign LevelGateway_14__EVAL_1 = _EVAL_35;
  assign LevelGateway_108__EVAL_4 = _EVAL_142;
  assign LevelGateway_61__EVAL_2 = _EVAL_105;
  assign LevelGateway_55__EVAL_0 = _EVAL_2254 == 1'h0;
  assign LevelGateway_115__EVAL_0 = _EVAL_3167 == 1'h0;
  assign LevelGateway_99__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_80 = _EVAL_3204;
  assign LevelGateway_126__EVAL_4 = _EVAL_142;
  assign LevelGateway_77__EVAL_4 = _EVAL_142;
  assign LevelGateway_35__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_57 = _EVAL_3768;
  assign LevelGateway_119__EVAL_0 = _EVAL_2202 == 1'h0;
  assign LevelGateway_98__EVAL_2 = _EVAL_105;
  assign LevelGateway_70__EVAL_1 = _EVAL_103;
  assign LevelGateway_124__EVAL = _EVAL_3491[125];
  assign Queue__EVAL_9 = _EVAL_131;
  assign LevelGateway_64__EVAL_2 = _EVAL_105;
  assign LevelGateway_11__EVAL = _EVAL_3491[12];
  assign LevelGateway_120__EVAL_1 = _EVAL_120;
  assign LevelGateway_25__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_100 = _EVAL_3113;
  assign LevelGateway_33__EVAL_2 = _EVAL_105;
  assign LevelGateway_36__EVAL = _EVAL_3491[37];
  assign LevelGateway_22__EVAL_1 = _EVAL_11;
  assign LevelGateway_83__EVAL_4 = _EVAL_142;
  assign LevelGateway_26__EVAL = _EVAL_3491[27];
  assign LevelGateway_89__EVAL_2 = _EVAL_105;
  assign LevelGateway_70__EVAL = _EVAL_3491[71];
  assign LevelGateway_56__EVAL = _EVAL_3491[57];
  assign LevelGateway_89__EVAL_1 = _EVAL_114;
  assign PLICFanIn__EVAL_46 = _EVAL_3591;
  assign LevelGateway_9__EVAL_1 = _EVAL_49;
  assign PLICFanIn__EVAL_2 = _EVAL_3573;
  assign LevelGateway_86__EVAL_4 = _EVAL_142;
  assign LevelGateway_3__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_87 = _EVAL_757;
  assign LevelGateway_106__EVAL_0 = _EVAL_3419 == 1'h0;
  assign LevelGateway_45__EVAL_2 = _EVAL_105;
  assign LevelGateway__EVAL_2 = _EVAL_105;
  assign LevelGateway_5__EVAL_1 = _EVAL_129;
  assign LevelGateway_17__EVAL_2 = _EVAL_105;
  assign LevelGateway_121__EVAL_1 = _EVAL_43;
  assign LevelGateway_114__EVAL_4 = _EVAL_142;
  assign LevelGateway_41__EVAL = _EVAL_3491[42];
  assign PLICFanIn__EVAL_43 = _EVAL_3242;
  assign LevelGateway_71__EVAL = _EVAL_3491[72];
  assign LevelGateway_95__EVAL_4 = _EVAL_142;
  assign LevelGateway_24__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_3 = _EVAL_3563;
  assign LevelGateway_87__EVAL_1 = _EVAL_125;
  assign PLICFanIn__EVAL_86 = _EVAL_3943;
  assign LevelGateway_51__EVAL_0 = _EVAL_2050 == 1'h0;
  assign LevelGateway_75__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_21 = _EVAL_304;
  assign PLICFanIn__EVAL_89 = _EVAL_3312;
  assign PLICFanIn__EVAL_12 = _EVAL_1801;
  assign LevelGateway_124__EVAL_2 = _EVAL_105;
  assign LevelGateway_57__EVAL_1 = _EVAL_108;
  assign LevelGateway_118__EVAL_1 = _EVAL_94;
  assign LevelGateway_8__EVAL_1 = _EVAL_52;
  assign LevelGateway_125__EVAL_4 = _EVAL_142;
  assign LevelGateway_57__EVAL_2 = _EVAL_105;
  assign Queue__EVAL_4 = _EVAL_59;
  assign LevelGateway_97__EVAL_1 = _EVAL_47;
  assign LevelGateway_73__EVAL_2 = _EVAL_105;
  assign LevelGateway_18__EVAL = _EVAL_3491[19];
  assign LevelGateway_1__EVAL_2 = _EVAL_105;
  assign LevelGateway_20__EVAL_4 = _EVAL_142;
  assign LevelGateway_64__EVAL = _EVAL_3491[65];
  assign LevelGateway_126__EVAL_0 = _EVAL_3713 == 1'h0;
  assign PLICFanIn__EVAL_92 = _EVAL_2646;
  assign LevelGateway_69__EVAL = _EVAL_3491[70];
  assign PLICFanIn__EVAL_1 = _EVAL_1212;
  assign LevelGateway_92__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_101 = _EVAL_481;
  assign LevelGateway_2__EVAL_1 = _EVAL_68;
  assign LevelGateway_86__EVAL_2 = _EVAL_105;
  assign LevelGateway_89__EVAL_0 = _EVAL_3996 == 1'h0;
  assign LevelGateway_36__EVAL_1 = _EVAL_17;
  assign LevelGateway_122__EVAL_2 = _EVAL_105;
  assign LevelGateway_66__EVAL_2 = _EVAL_105;
  assign LevelGateway_5__EVAL = _EVAL_3491[6];
  assign LevelGateway_63__EVAL_1 = _EVAL_61;
  assign LevelGateway_51__EVAL = _EVAL_3491[52];
  assign LevelGateway_80__EVAL_1 = _EVAL_57;
  assign LevelGateway_71__EVAL_4 = _EVAL_142;
  assign LevelGateway_106__EVAL = _EVAL_3491[107];
  assign PLICFanIn__EVAL_126 = _EVAL_188;
  assign LevelGateway_52__EVAL_2 = _EVAL_105;
  assign LevelGateway_2__EVAL = _EVAL_3491[3];
  assign LevelGateway_19__EVAL_4 = _EVAL_142;
  assign LevelGateway_80__EVAL_0 = _EVAL_1536 == 1'h0;
  assign Queue__EVAL_7 = _EVAL_84;
  assign LevelGateway_60__EVAL_0 = _EVAL_2341 == 1'h0;
  assign LevelGateway_60__EVAL = _EVAL_3491[61];
  assign PLICFanIn__EVAL_66 = _EVAL_485;
  assign LevelGateway_3__EVAL_1 = _EVAL_55;
  assign LevelGateway_69__EVAL_2 = _EVAL_105;
  assign LevelGateway_10__EVAL_1 = _EVAL_37;
  assign LevelGateway_62__EVAL_2 = _EVAL_105;
  assign LevelGateway_17__EVAL_0 = _EVAL_269 == 1'h0;
  assign LevelGateway_31__EVAL_0 = _EVAL_2507 == 1'h0;
  assign Queue__EVAL_2 = _EVAL_142;
  assign PLICFanIn__EVAL_61 = _EVAL_750;
  assign LevelGateway_24__EVAL = _EVAL_3491[25];
  assign LevelGateway_67__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_105 = _EVAL_2231;
  assign _EVAL_38 = {{2'd0}, _EVAL_815};
  assign LevelGateway_120__EVAL = _EVAL_3491[121];
  assign LevelGateway_38__EVAL_2 = _EVAL_105;
  assign LevelGateway_10__EVAL = _EVAL_3491[11];
  assign LevelGateway_8__EVAL_2 = _EVAL_105;
  assign LevelGateway_23__EVAL = _EVAL_3491[24];
  assign LevelGateway_121__EVAL_4 = _EVAL_142;
  assign LevelGateway_4__EVAL_1 = _EVAL_34;
  assign LevelGateway_59__EVAL_4 = _EVAL_142;
  assign LevelGateway_67__EVAL = _EVAL_3491[68];
  assign LevelGateway_32__EVAL = _EVAL_3491[33];
  assign LevelGateway_14__EVAL_0 = _EVAL_1556 == 1'h0;
  assign LevelGateway_39__EVAL_2 = _EVAL_105;
  assign LevelGateway_105__EVAL_1 = _EVAL_137;
  assign PLICFanIn__EVAL_106 = _EVAL_2881;
  assign LevelGateway_13__EVAL_0 = _EVAL_1121 == 1'h0;
  assign PLICFanIn__EVAL_125 = _EVAL_2851;
  assign LevelGateway_47__EVAL_0 = _EVAL_2485 == 1'h0;
  assign LevelGateway_95__EVAL_0 = _EVAL_1521 == 1'h0;
  assign Queue__EVAL_0 = {_EVAL_20,_EVAL_79};
  assign LevelGateway_34__EVAL_4 = _EVAL_142;
  assign LevelGateway_4__EVAL = _EVAL_3491[5];
  assign LevelGateway_45__EVAL = _EVAL_3491[46];
  assign LevelGateway_108__EVAL_1 = _EVAL_134;
  assign LevelGateway_88__EVAL_4 = _EVAL_142;
  assign LevelGateway_7__EVAL = _EVAL_3491[8];
  assign LevelGateway_29__EVAL_1 = _EVAL_28;
  assign PLICFanIn__EVAL_78 = _EVAL_2584;
  assign PLICFanIn__EVAL_23 = _EVAL_1151;
  assign LevelGateway_38__EVAL_4 = _EVAL_142;
  assign LevelGateway_72__EVAL = _EVAL_3491[73];
  assign LevelGateway_102__EVAL_1 = _EVAL_109;
  assign LevelGateway_83__EVAL_1 = _EVAL_33;
  assign PLICFanIn__EVAL_53 = _EVAL_768;
  assign LevelGateway_34__EVAL_0 = _EVAL_492 == 1'h0;
  assign LevelGateway_15__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_24 = _EVAL_2958;
  assign LevelGateway_29__EVAL_2 = _EVAL_105;
  assign LevelGateway_76__EVAL = _EVAL_3491[77];
  assign LevelGateway_37__EVAL_1 = _EVAL_56;
  assign LevelGateway_104__EVAL_1 = _EVAL_74;
  assign PLICFanIn__EVAL_120 = _EVAL_1660;
  assign LevelGateway_90__EVAL_0 = _EVAL_3757 == 1'h0;
  assign PLICFanIn__EVAL_7 = _EVAL_2256;
  assign LevelGateway_125__EVAL_2 = _EVAL_105;
  assign LevelGateway_13__EVAL_2 = _EVAL_105;
  assign LevelGateway_38__EVAL_0 = _EVAL_989 == 1'h0;
  assign LevelGateway_79__EVAL_2 = _EVAL_105;
  assign LevelGateway_27__EVAL = _EVAL_3491[28];
  assign LevelGateway_116__EVAL_1 = _EVAL_102;
  assign LevelGateway_107__EVAL_4 = _EVAL_142;
  assign LevelGateway_62__EVAL = _EVAL_3491[63];
  assign LevelGateway_91__EVAL_1 = _EVAL_63;
  assign PLICFanIn__EVAL_124 = _EVAL_512;
  assign LevelGateway_10__EVAL_2 = _EVAL_105;
  assign LevelGateway_51__EVAL_2 = _EVAL_105;
  assign LevelGateway_115__EVAL = _EVAL_3491[116];
  assign PLICFanIn__EVAL_56 = _EVAL_835;
  assign LevelGateway_84__EVAL_0 = _EVAL_3551 == 1'h0;
  assign LevelGateway_41__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_84 = _EVAL_1280;
  assign LevelGateway_43__EVAL_4 = _EVAL_142;
  assign LevelGateway_21__EVAL_1 = _EVAL_77;
  assign PLICFanIn__EVAL_37 = _EVAL_3008;
  assign Queue__EVAL_8 = _EVAL_910[23:0];
  assign PLICFanIn__EVAL_116 = _EVAL_1783;
  assign LevelGateway_93__EVAL_1 = _EVAL_136;
  assign LevelGateway_88__EVAL_2 = _EVAL_105;
  assign LevelGateway_64__EVAL_0 = _EVAL_947 == 1'h0;
  assign LevelGateway_66__EVAL_4 = _EVAL_142;
  assign LevelGateway_96__EVAL_0 = _EVAL_730 == 1'h0;
  assign LevelGateway_110__EVAL_0 = _EVAL_715 == 1'h0;
  assign LevelGateway_57__EVAL_4 = _EVAL_142;
  assign LevelGateway_124__EVAL_4 = _EVAL_142;
  assign LevelGateway_92__EVAL = _EVAL_3491[93];
  assign Queue__EVAL_14 = _EVAL_69;
  assign PLICFanIn__EVAL_6 = _EVAL_3740;
  assign LevelGateway_89__EVAL = _EVAL_3491[90];
  assign LevelGateway_94__EVAL_4 = _EVAL_142;
  assign LevelGateway_63__EVAL = _EVAL_3491[64];
  assign LevelGateway_82__EVAL_2 = _EVAL_105;
  assign LevelGateway_61__EVAL_4 = _EVAL_142;
  assign LevelGateway_68__EVAL_0 = _EVAL_2701 == 1'h0;
  assign LevelGateway_103__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_123 = _EVAL_286;
  assign LevelGateway_27__EVAL_2 = _EVAL_105;
  assign LevelGateway_15__EVAL_1 = _EVAL_26;
  assign LevelGateway_81__EVAL_4 = _EVAL_142;
  assign LevelGateway_48__EVAL = _EVAL_3491[49];
  assign LevelGateway_79__EVAL_1 = _EVAL_16;
  assign LevelGateway_77__EVAL_2 = _EVAL_105;
  assign LevelGateway_33__EVAL = _EVAL_3491[34];
  assign LevelGateway_83__EVAL_0 = _EVAL_3728 == 1'h0;
  assign LevelGateway_119__EVAL_1 = _EVAL_1;
  assign LevelGateway_90__EVAL_4 = _EVAL_142;
  assign LevelGateway_58__EVAL_2 = _EVAL_105;
  assign LevelGateway_92__EVAL_1 = _EVAL_9;
  assign LevelGateway_76__EVAL_1 = _EVAL_126;
  assign LevelGateway_1__EVAL = _EVAL_3491[2];
  assign LevelGateway_62__EVAL_0 = _EVAL_1073 == 1'h0;
  assign LevelGateway_62__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_96 = _EVAL_1122;
  assign LevelGateway_75__EVAL_2 = _EVAL_105;
  assign LevelGateway_88__EVAL = _EVAL_3491[89];
  assign LevelGateway_90__EVAL_2 = _EVAL_105;
  assign LevelGateway_20__EVAL_0 = _EVAL_1708 == 1'h0;
  assign LevelGateway_109__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_16 = _EVAL_3608;
  assign LevelGateway_69__EVAL_4 = _EVAL_142;
  assign LevelGateway_42__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_41 = _EVAL_1351;
  assign LevelGateway_71__EVAL_2 = _EVAL_105;
  assign LevelGateway_53__EVAL_1 = _EVAL_66;
  assign LevelGateway_43__EVAL_0 = _EVAL_690 == 1'h0;
  assign LevelGateway_113__EVAL = _EVAL_3491[114];
  assign LevelGateway_105__EVAL_2 = _EVAL_105;
  assign LevelGateway_45__EVAL_1 = _EVAL_5;
  assign LevelGateway_72__EVAL_0 = _EVAL_497 == 1'h0;
  assign LevelGateway_37__EVAL_2 = _EVAL_105;
  assign LevelGateway_115__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_5 = _EVAL_1365;
  assign LevelGateway_34__EVAL_1 = _EVAL_119;
  assign LevelGateway_118__EVAL_0 = _EVAL_4063 == 1'h0;
  assign LevelGateway_122__EVAL_0 = _EVAL_1599 == 1'h0;
  assign PLICFanIn__EVAL_83 = _EVAL_902;
  assign LevelGateway_65__EVAL_4 = _EVAL_142;
  assign LevelGateway_25__EVAL_4 = _EVAL_142;
  assign LevelGateway_66__EVAL = _EVAL_3491[67];
  assign LevelGateway_87__EVAL_4 = _EVAL_142;
  assign Queue__EVAL_1 = _EVAL_86 == 3'h4;
  assign PLICFanIn__EVAL_102 = _EVAL_1390;
  assign LevelGateway_20__EVAL_1 = _EVAL_128;
  assign LevelGateway_40__EVAL_2 = _EVAL_105;
  assign LevelGateway_78__EVAL_2 = _EVAL_105;
  assign LevelGateway_30__EVAL_1 = _EVAL_72;
  assign LevelGateway_18__EVAL_1 = _EVAL_99;
  assign LevelGateway_74__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_117 = _EVAL_1562;
  assign LevelGateway_113__EVAL_0 = _EVAL_1917 == 1'h0;
  assign LevelGateway_75__EVAL = _EVAL_3491[76];
  assign LevelGateway_62__EVAL_1 = _EVAL_36;
  assign LevelGateway_68__EVAL_1 = _EVAL_73;
  assign LevelGateway_26__EVAL_0 = _EVAL_448 == 1'h0;
  assign LevelGateway_12__EVAL_4 = _EVAL_142;
  assign LevelGateway_54__EVAL = _EVAL_3491[55];
  assign PLICFanIn__EVAL_121 = _EVAL_3274;
  assign LevelGateway_107__EVAL_1 = _EVAL_0;
  assign LevelGateway_95__EVAL_1 = _EVAL_144;
  assign LevelGateway_101__EVAL_2 = _EVAL_105;
  assign LevelGateway_45__EVAL_4 = _EVAL_142;
  assign LevelGateway_25__EVAL = _EVAL_3491[26];
  assign PLICFanIn__EVAL_95 = _EVAL_1156;
  assign LevelGateway_43__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_27 = _EVAL_1738;
  assign LevelGateway_86__EVAL_0 = _EVAL_2809 == 1'h0;
  assign LevelGateway_7__EVAL_4 = _EVAL_142;
  assign LevelGateway_7__EVAL_2 = _EVAL_105;
  assign LevelGateway_93__EVAL_2 = _EVAL_105;
  assign LevelGateway_12__EVAL = _EVAL_3491[13];
  assign LevelGateway_110__EVAL_4 = _EVAL_142;
  assign LevelGateway_42__EVAL_2 = _EVAL_105;
  assign LevelGateway_101__EVAL_4 = _EVAL_142;
  assign LevelGateway_121__EVAL = _EVAL_3491[122];
  assign LevelGateway_114__EVAL_1 = _EVAL_121;
  assign PLICFanIn__EVAL_14 = _EVAL_1253;
  assign LevelGateway_98__EVAL_1 = _EVAL_111;
  assign LevelGateway_26__EVAL_1 = _EVAL_19;
  assign LevelGateway_85__EVAL = _EVAL_3491[86];
  assign LevelGateway_100__EVAL_4 = _EVAL_142;
  assign LevelGateway_27__EVAL_4 = _EVAL_142;
  assign LevelGateway_84__EVAL = _EVAL_3491[85];
  assign LevelGateway_119__EVAL_4 = _EVAL_142;
  assign LevelGateway_41__EVAL_1 = _EVAL_135;
  assign PLICFanIn__EVAL_76 = _EVAL_2311;
  assign LevelGateway_111__EVAL_4 = _EVAL_142;
  assign LevelGateway_13__EVAL = _EVAL_3491[14];
  assign LevelGateway_113__EVAL_2 = _EVAL_105;
  assign LevelGateway_19__EVAL_0 = _EVAL_3192 == 1'h0;
  assign LevelGateway_77__EVAL = _EVAL_3491[78];
  assign LevelGateway_56__EVAL_2 = _EVAL_105;
  assign LevelGateway_26__EVAL_4 = _EVAL_142;
  assign LevelGateway_14__EVAL_4 = _EVAL_142;
  assign LevelGateway_87__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_58 = _EVAL_2810;
  assign LevelGateway_124__EVAL_1 = _EVAL_32;
  assign LevelGateway_21__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_99 = _EVAL_2653;
  assign LevelGateway_65__EVAL_1 = _EVAL_112;
  assign LevelGateway_76__EVAL_2 = _EVAL_105;
  assign LevelGateway_97__EVAL = _EVAL_3491[98];
  assign LevelGateway_112__EVAL_1 = _EVAL_6;
  assign LevelGateway_16__EVAL_1 = _EVAL_39;
  assign LevelGateway_126__EVAL_1 = _EVAL_91;
  assign PLICFanIn__EVAL_55 = _EVAL_3102;
  assign LevelGateway_38__EVAL = _EVAL_3491[39];
  assign LevelGateway_114__EVAL = _EVAL_3491[115];
  assign LevelGateway_110__EVAL_1 = _EVAL_107;
  assign _EVAL_62 = _EVAL_291[1:0];
  assign LevelGateway_94__EVAL_0 = _EVAL_2953 == 1'h0;
  assign PLICFanIn__EVAL_33 = _EVAL_1176;
  assign LevelGateway_123__EVAL_0 = _EVAL_1471 == 1'h0;
  assign LevelGateway_104__EVAL_4 = _EVAL_142;
  assign LevelGateway_28__EVAL_1 = _EVAL_14;
  assign LevelGateway_112__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_59 = _EVAL_2720;
  assign LevelGateway_99__EVAL_2 = _EVAL_105;
  assign LevelGateway_61__EVAL_0 = _EVAL_2870 == 1'h0;
  assign LevelGateway_85__EVAL_2 = _EVAL_105;
  assign LevelGateway_52__EVAL_0 = _EVAL_2803 == 1'h0;
  assign LevelGateway_124__EVAL_0 = _EVAL_449 == 1'h0;
  assign LevelGateway_9__EVAL_2 = _EVAL_105;
  assign LevelGateway_65__EVAL_2 = _EVAL_105;
  assign LevelGateway_50__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_65 = _EVAL_765;
  assign LevelGateway_65__EVAL = _EVAL_3491[66];
  assign LevelGateway_78__EVAL_1 = _EVAL_12;
  assign LevelGateway_96__EVAL_1 = _EVAL_104;
  assign LevelGateway_55__EVAL_4 = _EVAL_142;
  assign LevelGateway_14__EVAL = _EVAL_3491[15];
  assign PLICFanIn__EVAL_114 = _EVAL_2336;
  assign LevelGateway_126__EVAL = _EVAL_3491[127];
  assign LevelGateway_20__EVAL = _EVAL_3491[21];
  assign LevelGateway_36__EVAL_0 = _EVAL_427 == 1'h0;
  assign LevelGateway_123__EVAL = _EVAL_3491[124];
  assign LevelGateway_110__EVAL_2 = _EVAL_105;
  assign LevelGateway__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_110 = _EVAL_1526;
  assign PLICFanIn__EVAL_71 = _EVAL_3644;
  assign LevelGateway_116__EVAL = _EVAL_3491[117];
  assign LevelGateway_28__EVAL = _EVAL_3491[29];
  assign LevelGateway_105__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_11 = _EVAL_1438;
  assign LevelGateway_76__EVAL_4 = _EVAL_142;
  assign LevelGateway_34__EVAL_2 = _EVAL_105;
  assign LevelGateway_96__EVAL_4 = _EVAL_142;
  assign LevelGateway_72__EVAL_4 = _EVAL_142;
  assign LevelGateway_28__EVAL_0 = _EVAL_3317 == 1'h0;
  assign LevelGateway_4__EVAL_2 = _EVAL_105;
  assign LevelGateway_125__EVAL = _EVAL_3491[126];
  assign LevelGateway_79__EVAL = _EVAL_3491[80];
  assign LevelGateway_112__EVAL_0 = _EVAL_480 == 1'h0;
  assign PLICFanIn__EVAL_115 = _EVAL_1433;
  assign LevelGateway_44__EVAL = _EVAL_3491[45];
  assign LevelGateway_30__EVAL_4 = _EVAL_142;
  assign LevelGateway_112__EVAL = _EVAL_3491[113];
  assign LevelGateway_46__EVAL = _EVAL_3491[47];
  assign PLICFanIn__EVAL_90 = _EVAL_3554;
  assign LevelGateway_22__EVAL_0 = _EVAL_2214 == 1'h0;
  assign LevelGateway_74__EVAL_0 = _EVAL_3361 == 1'h0;
  assign LevelGateway_2__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_111 = _EVAL_1035;
  assign PLICFanIn__EVAL_50 = _EVAL_2121;
  assign LevelGateway_42__EVAL = _EVAL_3491[43];
  assign LevelGateway_27__EVAL_1 = _EVAL_132;
  assign LevelGateway_20__EVAL_2 = _EVAL_105;
  assign LevelGateway_70__EVAL_4 = _EVAL_142;
  assign LevelGateway_73__EVAL_4 = _EVAL_142;
  assign LevelGateway_52__EVAL_4 = _EVAL_142;
  assign LevelGateway_72__EVAL_2 = _EVAL_105;
  assign LevelGateway_109__EVAL_0 = _EVAL_1267 == 1'h0;
  assign LevelGateway_23__EVAL_4 = _EVAL_142;
  assign LevelGateway_115__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_112 = _EVAL_147;
  assign LevelGateway_38__EVAL_1 = _EVAL_75;
  assign LevelGateway_102__EVAL = _EVAL_3491[103];
  assign LevelGateway_51__EVAL_1 = _EVAL_67;
  assign LevelGateway_74__EVAL_2 = _EVAL_105;
  assign LevelGateway_35__EVAL_0 = _EVAL_1456 == 1'h0;
  assign LevelGateway_81__EVAL_2 = _EVAL_105;
  assign LevelGateway_44__EVAL_0 = _EVAL_3025 == 1'h0;
  assign PLICFanIn__EVAL_79 = _EVAL_293;
  assign LevelGateway_5__EVAL_0 = _EVAL_3759 == 1'h0;
  assign LevelGateway_96__EVAL_2 = _EVAL_105;
  assign PLICFanIn__EVAL_38 = _EVAL_3804;
  assign LevelGateway_79__EVAL_4 = _EVAL_142;
  assign _EVAL_3 = Queue__EVAL_5;
  assign LevelGateway_3__EVAL_0 = _EVAL_2826 == 1'h0;
  assign PLICFanIn__EVAL_35 = _EVAL_739;
  assign PLICFanIn__EVAL_22 = _EVAL_3801;
  assign LevelGateway_37__EVAL_4 = _EVAL_142;
  assign LevelGateway_43__EVAL_1 = _EVAL_101;
  assign LevelGateway_117__EVAL = _EVAL_3491[118];
  assign LevelGateway_4__EVAL_0 = _EVAL_163 == 1'h0;
  assign LevelGateway_54__EVAL_1 = _EVAL_60;
  assign LevelGateway_104__EVAL = _EVAL_3491[105];
  assign LevelGateway_125__EVAL_0 = _EVAL_3850 == 1'h0;
  assign PLICFanIn__EVAL_91 = _EVAL_410;
  assign LevelGateway_47__EVAL_2 = _EVAL_105;
  assign LevelGateway_93__EVAL_4 = _EVAL_142;
  assign LevelGateway_40__EVAL_1 = _EVAL_13;
  assign PLICFanIn__EVAL_18 = _EVAL_1168;
  assign PLICFanIn__EVAL_68 = _EVAL_3733;
  assign LevelGateway_66__EVAL_0 = _EVAL_3359 == 1'h0;
  assign LevelGateway_116__EVAL_0 = _EVAL_1938 == 1'h0;
  assign LevelGateway_63__EVAL_0 = _EVAL_1587 == 1'h0;
  assign LevelGateway_84__EVAL_4 = _EVAL_142;
  assign LevelGateway_29__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_44 = _EVAL_2356;
  assign LevelGateway_15__EVAL_2 = _EVAL_105;
  assign LevelGateway_55__EVAL_1 = _EVAL_98;
  assign PLICFanIn__EVAL_85 = _EVAL_1266;
  assign LevelGateway_37__EVAL = _EVAL_3491[38];
  assign LevelGateway_82__EVAL = _EVAL_3491[83];
  assign LevelGateway_30__EVAL = _EVAL_3491[31];
  assign LevelGateway_33__EVAL_4 = _EVAL_142;
  assign LevelGateway_16__EVAL = _EVAL_3491[17];
  assign LevelGateway_85__EVAL_4 = _EVAL_142;
  assign PLICFanIn__EVAL_19 = _EVAL_3383;
  assign LevelGateway_123__EVAL_1 = _EVAL_117;
  assign LevelGateway_121__EVAL_0 = _EVAL_2938 == 1'h0;
  assign _EVAL = _EVAL_291[13:2];
  assign LevelGateway_70__EVAL_2 = _EVAL_105;
  assign LevelGateway_95__EVAL = _EVAL_3491[96];
  assign PLICFanIn__EVAL_8 = _EVAL_2500;
  assign PLICFanIn__EVAL_13 = _EVAL_3315;
  assign LevelGateway_59__EVAL_2 = _EVAL_105;
  assign LevelGateway_19__EVAL_2 = _EVAL_105;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_147 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_155 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_163 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_176 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_188 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_194 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_200 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_212 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_217 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_222 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_247 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_251 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_269 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_285 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_286 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_293 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_304 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_306 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_331 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_354 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_366 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_371 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_387 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_410 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_421 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_427 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_444 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_448 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_449 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_462 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_480 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_481 = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_485 = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_492 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_497 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_512 = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_519 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_548 = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_552 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_569 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_581 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_614 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_648 = _RAND_42[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_663 = _RAND_43[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_673 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_675 = _RAND_45[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_690 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_715 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_730 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_739 = _RAND_49[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_741 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_750 = _RAND_51[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_757 = _RAND_52[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_762 = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_765 = _RAND_54[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_768 = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_770 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_835 = _RAND_57[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_880 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_902 = _RAND_59[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_912 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_947 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_989 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1035 = _RAND_63[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1073 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1088 = _RAND_65[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1121 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1122 = _RAND_67[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1127 = _RAND_68[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1142 = _RAND_69[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1151 = _RAND_70[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1156 = _RAND_71[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1162 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1168 = _RAND_73[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1176 = _RAND_74[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1206 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1212 = _RAND_76[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1239 = _RAND_77[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1253 = _RAND_78[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1261 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1266 = _RAND_80[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1267 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1270 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1280 = _RAND_83[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1313 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1315 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1351 = _RAND_86[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1365 = _RAND_87[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1390 = _RAND_88[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1433 = _RAND_89[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1438 = _RAND_90[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1444 = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1456 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1471 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1496 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1521 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1526 = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1536 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1556 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1562 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1580 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1587 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1597 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1599 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1639 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1660 = _RAND_105[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1680 = _RAND_106[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_1697 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1698 = _RAND_108[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_1708 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1709 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1738 = _RAND_111[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1753 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1776 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _EVAL_1783 = _RAND_114[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_1786 = _RAND_115[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1788 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1801 = _RAND_117[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1819 = _RAND_118[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_1870 = _RAND_119[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1917 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1929 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1930 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1938 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_1962 = _RAND_124[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_1979 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_1980 = _RAND_126[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_2018 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_2035 = _RAND_128[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_2050 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_2055 = _RAND_130[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_2073 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_2110 = _RAND_132[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_2111 = _RAND_133[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_2121 = _RAND_134[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_2128 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_2133 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_2155 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_2159 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_2188 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_2202 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_2209 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _EVAL_2214 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2231 = _RAND_143[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _EVAL_2254 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _EVAL_2256 = _RAND_145[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2290 = _RAND_146[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _EVAL_2306 = _RAND_147[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _EVAL_2311 = _RAND_148[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _EVAL_2334 = _RAND_149[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _EVAL_2336 = _RAND_150[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _EVAL_2341 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _EVAL_2356 = _RAND_152[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _EVAL_2481 = _RAND_153[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _EVAL_2484 = _RAND_154[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _EVAL_2485 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _EVAL_2491 = _RAND_156[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _EVAL_2500 = _RAND_157[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _EVAL_2507 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _EVAL_2536 = _RAND_159[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _EVAL_2582 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _EVAL_2584 = _RAND_161[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _EVAL_2646 = _RAND_162[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _EVAL_2648 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _EVAL_2653 = _RAND_164[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _EVAL_2666 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _EVAL_2677 = _RAND_166[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _EVAL_2684 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _EVAL_2688 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _EVAL_2701 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _EVAL_2720 = _RAND_170[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _EVAL_2754 = _RAND_171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _EVAL_2760 = _RAND_172[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _EVAL_2803 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _EVAL_2807 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _EVAL_2809 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _EVAL_2810 = _RAND_176[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _EVAL_2826 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _EVAL_2838 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _EVAL_2850 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _EVAL_2851 = _RAND_180[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _EVAL_2870 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _EVAL_2881 = _RAND_182[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _EVAL_2937 = _RAND_183[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _EVAL_2938 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _EVAL_2942 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _EVAL_2953 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _EVAL_2958 = _RAND_187[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _EVAL_2965 = _RAND_188[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _EVAL_2972 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _EVAL_3008 = _RAND_190[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _EVAL_3014 = _RAND_191[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _EVAL_3023 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _EVAL_3025 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _EVAL_3039 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _EVAL_3056 = _RAND_195[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _EVAL_3102 = _RAND_196[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _EVAL_3113 = _RAND_197[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _EVAL_3118 = _RAND_198[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _EVAL_3137 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _EVAL_3167 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _EVAL_3192 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _EVAL_3195 = _RAND_202[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _EVAL_3199 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _EVAL_3204 = _RAND_204[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _EVAL_3216 = _RAND_205[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _EVAL_3222 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _EVAL_3235 = _RAND_207[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _EVAL_3242 = _RAND_208[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _EVAL_3245 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _EVAL_3267 = _RAND_210[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _EVAL_3274 = _RAND_211[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _EVAL_3279 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _EVAL_3283 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _EVAL_3296 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _EVAL_3299 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _EVAL_3312 = _RAND_216[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _EVAL_3315 = _RAND_217[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _EVAL_3317 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _EVAL_3331 = _RAND_219[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _EVAL_3336 = _RAND_220[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _EVAL_3359 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _EVAL_3361 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _EVAL_3383 = _RAND_223[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _EVAL_3407 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _EVAL_3419 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _EVAL_3421 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _EVAL_3488 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _EVAL_3505 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _EVAL_3527 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _EVAL_3551 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _EVAL_3552 = _RAND_231[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _EVAL_3554 = _RAND_232[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _EVAL_3563 = _RAND_233[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _EVAL_3571 = _RAND_234[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _EVAL_3573 = _RAND_235[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _EVAL_3591 = _RAND_236[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _EVAL_3608 = _RAND_237[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _EVAL_3623 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _EVAL_3636 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _EVAL_3644 = _RAND_240[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _EVAL_3645 = _RAND_241[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _EVAL_3713 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _EVAL_3715 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _EVAL_3720 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _EVAL_3721 = _RAND_245[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _EVAL_3728 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _EVAL_3731 = _RAND_247[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _EVAL_3733 = _RAND_248[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _EVAL_3740 = _RAND_249[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _EVAL_3743 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _EVAL_3750 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _EVAL_3757 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _EVAL_3759 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _EVAL_3768 = _RAND_254[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _EVAL_3783 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _EVAL_3788 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _EVAL_3801 = _RAND_257[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _EVAL_3804 = _RAND_258[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _EVAL_3843 = _RAND_259[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _EVAL_3850 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _EVAL_3870 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _EVAL_3899 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _EVAL_3909 = _RAND_263[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _EVAL_3913 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _EVAL_3943 = _RAND_265[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _EVAL_3964 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _EVAL_3996 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _EVAL_4013 = _RAND_268[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _EVAL_4034 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _EVAL_4050 = _RAND_270[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _EVAL_4063 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _EVAL_4066 = _RAND_272[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_142) begin
    if (_EVAL_1139) begin
      _EVAL_147 <= _EVAL_3965;
    end
    if (_EVAL_1841) begin
      _EVAL_155 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_163 <= 1'h0;
    end else begin
      if (_EVAL_622) begin
        _EVAL_163 <= _EVAL_3281;
      end
    end
    if (_EVAL_105) begin
      _EVAL_176 <= 1'h0;
    end else begin
      if (_EVAL_3825) begin
        _EVAL_176 <= _EVAL_1424;
      end
    end
    if (_EVAL_3103) begin
      _EVAL_188 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_194 <= 1'h0;
    end else begin
      if (_EVAL_1350) begin
        _EVAL_194 <= _EVAL_1740;
      end
    end
    if (_EVAL_105) begin
      _EVAL_200 <= 1'h0;
    end else begin
      if (_EVAL_1936) begin
        _EVAL_200 <= _EVAL_2129;
      end
    end
    if (_EVAL_105) begin
      _EVAL_212 <= 1'h0;
    end else begin
      if (_EVAL_1242) begin
        _EVAL_212 <= _EVAL_4028;
      end
    end
    if (_EVAL_105) begin
      _EVAL_217 <= 1'h0;
    end else begin
      if (_EVAL_1093) begin
        _EVAL_217 <= _EVAL_1506;
      end
    end
    if (_EVAL_105) begin
      _EVAL_222 <= 1'h0;
    end else begin
      if (_EVAL_2578) begin
        _EVAL_222 <= _EVAL_2956;
      end
    end
    if (_EVAL_3337) begin
      _EVAL_247 <= _EVAL_3965;
    end
    if (_EVAL_3064) begin
      _EVAL_251 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_269 <= 1'h0;
    end else begin
      if (_EVAL_2852) begin
        _EVAL_269 <= _EVAL_4026;
      end
    end
    if (_EVAL_3842) begin
      _EVAL_285 <= _EVAL_3965;
    end
    if (_EVAL_2001) begin
      _EVAL_286 <= _EVAL_3965;
    end
    if (_EVAL_3191) begin
      _EVAL_293 <= _EVAL_3965;
    end
    if (_EVAL_612) begin
      _EVAL_304 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_306 <= 1'h0;
    end else begin
      if (_EVAL_1357) begin
        _EVAL_306 <= _EVAL_2365;
      end
    end
    if (_EVAL_2729) begin
      _EVAL_331 <= _EVAL_3965;
    end
    if (_EVAL_3005) begin
      _EVAL_354 <= _EVAL_3965;
    end
    if (_EVAL_2639) begin
      _EVAL_366 <= _EVAL_2047;
    end
    if (_EVAL_105) begin
      _EVAL_371 <= 1'h0;
    end else begin
      if (_EVAL_3065) begin
        _EVAL_371 <= _EVAL_2017;
      end
    end
    if (_EVAL_105) begin
      _EVAL_387 <= 1'h0;
    end else begin
      if (_EVAL_3047) begin
        _EVAL_387 <= _EVAL_971;
      end
    end
    if (_EVAL_3185) begin
      _EVAL_410 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_421 <= 1'h0;
    end else begin
      if (_EVAL_2208) begin
        _EVAL_421 <= _EVAL_3070;
      end
    end
    if (_EVAL_105) begin
      _EVAL_427 <= 1'h0;
    end else begin
      if (_EVAL_509) begin
        _EVAL_427 <= _EVAL_3765;
      end
    end
    if (_EVAL_2660) begin
      _EVAL_444 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_448 <= 1'h0;
    end else begin
      if (_EVAL_355) begin
        _EVAL_448 <= _EVAL_3879;
      end
    end
    if (_EVAL_105) begin
      _EVAL_449 <= 1'h0;
    end else begin
      if (_EVAL_734) begin
        _EVAL_449 <= _EVAL_3868;
      end
    end
    if (_EVAL_105) begin
      _EVAL_462 <= 1'h0;
    end else begin
      if (_EVAL_3275) begin
        _EVAL_462 <= _EVAL_1453;
      end
    end
    if (_EVAL_105) begin
      _EVAL_480 <= 1'h0;
    end else begin
      if (_EVAL_1264) begin
        _EVAL_480 <= _EVAL_3649;
      end
    end
    if (_EVAL_2654) begin
      _EVAL_481 <= _EVAL_3965;
    end
    if (_EVAL_576) begin
      _EVAL_485 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_492 <= 1'h0;
    end else begin
      if (_EVAL_720) begin
        _EVAL_492 <= _EVAL_1571;
      end
    end
    if (_EVAL_105) begin
      _EVAL_497 <= 1'h0;
    end else begin
      if (_EVAL_2944) begin
        _EVAL_497 <= _EVAL_3625;
      end
    end
    if (_EVAL_866) begin
      _EVAL_512 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_519 <= 1'h0;
    end else begin
      if (_EVAL_3424) begin
        _EVAL_519 <= _EVAL_3755;
      end
    end
    if (_EVAL_1120) begin
      _EVAL_548 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_552 <= 1'h0;
    end else begin
      if (_EVAL_2378) begin
        _EVAL_552 <= _EVAL_372;
      end
    end
    if (_EVAL_105) begin
      _EVAL_569 <= 1'h0;
    end else begin
      if (_EVAL_2910) begin
        _EVAL_569 <= _EVAL_2898;
      end
    end
    if (_EVAL_105) begin
      _EVAL_581 <= 1'h0;
    end else begin
      if (_EVAL_3749) begin
        _EVAL_581 <= _EVAL_2593;
      end
    end
    if (_EVAL_105) begin
      _EVAL_614 <= 1'h0;
    end else begin
      if (_EVAL_1486) begin
        _EVAL_614 <= _EVAL_2907;
      end
    end
    if (_EVAL_2160) begin
      _EVAL_648 <= _EVAL_3965;
    end
    if (_EVAL_298) begin
      _EVAL_663 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_673 <= 1'h0;
    end else begin
      if (_EVAL_2482) begin
        _EVAL_673 <= _EVAL_1452;
      end
    end
    if (_EVAL_3539) begin
      _EVAL_675 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_690 <= 1'h0;
    end else begin
      if (_EVAL_917) begin
        _EVAL_690 <= _EVAL_2573;
      end
    end
    if (_EVAL_105) begin
      _EVAL_715 <= 1'h0;
    end else begin
      if (_EVAL_682) begin
        _EVAL_715 <= _EVAL_2163;
      end
    end
    if (_EVAL_105) begin
      _EVAL_730 <= 1'h0;
    end else begin
      if (_EVAL_1771) begin
        _EVAL_730 <= _EVAL_1999;
      end
    end
    if (_EVAL_2869) begin
      _EVAL_739 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_741 <= 1'h0;
    end else begin
      if (_EVAL_1265) begin
        _EVAL_741 <= _EVAL_428;
      end
    end
    if (_EVAL_1161) begin
      _EVAL_750 <= _EVAL_3965;
    end
    if (_EVAL_4061) begin
      _EVAL_757 <= _EVAL_3965;
    end
    if (_EVAL_1998) begin
      _EVAL_762 <= _EVAL_3965;
    end
    if (_EVAL_1461) begin
      _EVAL_765 <= _EVAL_3965;
    end
    if (_EVAL_2099) begin
      _EVAL_768 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_770 <= 1'h0;
    end else begin
      if (_EVAL_2139) begin
        _EVAL_770 <= _EVAL_1723;
      end
    end
    if (_EVAL_1386) begin
      _EVAL_835 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_880 <= 1'h0;
    end else begin
      if (_EVAL_2291) begin
        _EVAL_880 <= _EVAL_375;
      end
    end
    if (_EVAL_3650) begin
      _EVAL_902 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_912 <= 1'h0;
    end else begin
      if (_EVAL_2737) begin
        _EVAL_912 <= _EVAL_565;
      end
    end
    if (_EVAL_105) begin
      _EVAL_947 <= 1'h0;
    end else begin
      if (_EVAL_2277) begin
        _EVAL_947 <= _EVAL_1815;
      end
    end
    if (_EVAL_105) begin
      _EVAL_989 <= 1'h0;
    end else begin
      if (_EVAL_2627) begin
        _EVAL_989 <= _EVAL_1541;
      end
    end
    if (_EVAL_2048) begin
      _EVAL_1035 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1073 <= 1'h0;
    end else begin
      if (_EVAL_1887) begin
        _EVAL_1073 <= _EVAL_335;
      end
    end
    if (_EVAL_2663) begin
      _EVAL_1088 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1121 <= 1'h0;
    end else begin
      if (_EVAL_1914) begin
        _EVAL_1121 <= _EVAL_631;
      end
    end
    if (_EVAL_532) begin
      _EVAL_1122 <= _EVAL_3965;
    end
    if (_EVAL_1082) begin
      _EVAL_1127 <= _EVAL_3965;
    end
    if (_EVAL_1966) begin
      _EVAL_1142 <= _EVAL_3965;
    end
    if (_EVAL_3152) begin
      _EVAL_1151 <= _EVAL_3965;
    end
    if (_EVAL_1784) begin
      _EVAL_1156 <= _EVAL_3965;
    end
    if (_EVAL_4009) begin
      _EVAL_1162 <= _EVAL_688;
    end
    if (_EVAL_651) begin
      _EVAL_1168 <= _EVAL_3965;
    end
    if (_EVAL_1215) begin
      _EVAL_1176 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1206 <= 1'h0;
    end else begin
      if (_EVAL_1096) begin
        _EVAL_1206 <= _EVAL_3680;
      end
    end
    if (_EVAL_2511) begin
      _EVAL_1212 <= _EVAL_3965;
    end
    if (_EVAL_2785) begin
      _EVAL_1239 <= _EVAL_3965;
    end
    if (_EVAL_660) begin
      _EVAL_1253 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1261 <= 1'h0;
    end else begin
      if (_EVAL_1758) begin
        _EVAL_1261 <= _EVAL_2316;
      end
    end
    if (_EVAL_3409) begin
      _EVAL_1266 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1267 <= 1'h0;
    end else begin
      if (_EVAL_3390) begin
        _EVAL_1267 <= _EVAL_342;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1270 <= 1'h0;
    end else begin
      if (_EVAL_3796) begin
        _EVAL_1270 <= _EVAL_3784;
      end
    end
    if (_EVAL_1548) begin
      _EVAL_1280 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1313 <= 1'h0;
    end else begin
      if (_EVAL_1763) begin
        _EVAL_1313 <= _EVAL_2140;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1315 <= 1'h0;
    end else begin
      if (_EVAL_1333) begin
        _EVAL_1315 <= _EVAL_2786;
      end
    end
    if (_EVAL_2603) begin
      _EVAL_1351 <= _EVAL_3965;
    end
    if (_EVAL_1591) begin
      _EVAL_1365 <= _EVAL_3965;
    end
    if (_EVAL_391) begin
      _EVAL_1390 <= _EVAL_3965;
    end
    if (_EVAL_3997) begin
      _EVAL_1433 <= _EVAL_3965;
    end
    if (_EVAL_3456) begin
      _EVAL_1438 <= _EVAL_3965;
    end
    _EVAL_1444 <= PLICFanIn__EVAL_32;
    if (_EVAL_105) begin
      _EVAL_1456 <= 1'h0;
    end else begin
      if (_EVAL_2463) begin
        _EVAL_1456 <= _EVAL_2425;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1471 <= 1'h0;
    end else begin
      if (_EVAL_2704) begin
        _EVAL_1471 <= _EVAL_968;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1496 <= 1'h0;
    end else begin
      if (_EVAL_2698) begin
        _EVAL_1496 <= _EVAL_2382;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1521 <= 1'h0;
    end else begin
      if (_EVAL_3549) begin
        _EVAL_1521 <= _EVAL_2565;
      end
    end
    if (_EVAL_541) begin
      _EVAL_1526 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1536 <= 1'h0;
    end else begin
      if (_EVAL_1229) begin
        _EVAL_1536 <= _EVAL_1397;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1556 <= 1'h0;
    end else begin
      if (_EVAL_3334) begin
        _EVAL_1556 <= _EVAL_2844;
      end
    end
    if (_EVAL_3939) begin
      _EVAL_1562 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1580 <= 1'h0;
    end else begin
      if (_EVAL_1632) begin
        _EVAL_1580 <= _EVAL_473;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1587 <= 1'h0;
    end else begin
      if (_EVAL_1799) begin
        _EVAL_1587 <= _EVAL_3896;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1597 <= 1'h0;
    end else begin
      if (_EVAL_3667) begin
        _EVAL_1597 <= _EVAL_2827;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1599 <= 1'h0;
    end else begin
      if (_EVAL_2169) begin
        _EVAL_1599 <= _EVAL_3011;
      end
    end
    if (_EVAL_2865) begin
      _EVAL_1639 <= _EVAL_1861;
    end
    if (_EVAL_1728) begin
      _EVAL_1660 <= _EVAL_3965;
    end
    if (_EVAL_1311) begin
      _EVAL_1680 <= _EVAL_3965;
    end
    if (_EVAL_2515) begin
      _EVAL_1697 <= _EVAL_3020;
    end
    if (_EVAL_2696) begin
      _EVAL_1698 <= _EVAL_3432;
    end
    if (_EVAL_105) begin
      _EVAL_1708 <= 1'h0;
    end else begin
      if (_EVAL_963) begin
        _EVAL_1708 <= _EVAL_3371;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1709 <= 1'h0;
    end else begin
      if (_EVAL_3006) begin
        _EVAL_1709 <= _EVAL_3078;
      end
    end
    if (_EVAL_2058) begin
      _EVAL_1738 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1753 <= 1'h0;
    end else begin
      if (_EVAL_1094) begin
        _EVAL_1753 <= _EVAL_2358;
      end
    end
    if (_EVAL_1773) begin
      _EVAL_1776 <= _EVAL_2047;
    end
    if (_EVAL_3832) begin
      _EVAL_1783 <= _EVAL_3965;
    end
    if (_EVAL_2057) begin
      _EVAL_1786 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1788 <= 1'h0;
    end else begin
      if (_EVAL_2278) begin
        _EVAL_1788 <= _EVAL_1958;
      end
    end
    if (_EVAL_1558) begin
      _EVAL_1801 <= _EVAL_3965;
    end
    if (_EVAL_3683) begin
      _EVAL_1819 <= _EVAL_3965;
    end
    if (_EVAL_3024) begin
      _EVAL_1870 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1917 <= 1'h0;
    end else begin
      if (_EVAL_1500) begin
        _EVAL_1917 <= _EVAL_2443;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1929 <= 1'h0;
    end else begin
      if (_EVAL_1585) begin
        _EVAL_1929 <= _EVAL_3663;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1930 <= 1'h0;
    end else begin
      if (_EVAL_303) begin
        _EVAL_1930 <= _EVAL_3443;
      end
    end
    if (_EVAL_105) begin
      _EVAL_1938 <= 1'h0;
    end else begin
      if (_EVAL_2346) begin
        _EVAL_1938 <= _EVAL_2788;
      end
    end
    if (_EVAL_3764) begin
      _EVAL_1962 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_1979 <= 1'h0;
    end else begin
      if (_EVAL_3292) begin
        _EVAL_1979 <= _EVAL_3256;
      end
    end
    if (_EVAL_2744) begin
      _EVAL_1980 <= _EVAL_3965;
    end
    if (_EVAL_2825) begin
      _EVAL_2018 <= _EVAL_688;
    end
    if (_EVAL_1472) begin
      _EVAL_2035 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2050 <= 1'h0;
    end else begin
      if (_EVAL_3595) begin
        _EVAL_2050 <= _EVAL_3534;
      end
    end
    if (_EVAL_1655) begin
      _EVAL_2055 <= _EVAL_3965;
    end
    if (_EVAL_807) begin
      _EVAL_2073 <= _EVAL_1861;
    end
    if (_EVAL_1187) begin
      _EVAL_2110 <= _EVAL_3965;
    end
    if (_EVAL_1510) begin
      _EVAL_2111 <= _EVAL_3965;
    end
    if (_EVAL_2408) begin
      _EVAL_2121 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2128 <= 1'h0;
    end else begin
      if (_EVAL_1294) begin
        _EVAL_2128 <= _EVAL_2963;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2133 <= 1'h0;
    end else begin
      if (_EVAL_956) begin
        _EVAL_2133 <= _EVAL_731;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2155 <= 1'h0;
    end else begin
      if (_EVAL_1465) begin
        _EVAL_2155 <= _EVAL_2325;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2159 <= 1'h0;
    end else begin
      if (_EVAL_4068) begin
        _EVAL_2159 <= _EVAL_2969;
      end
    end
    if (_EVAL_2233) begin
      _EVAL_2188 <= _EVAL_1861;
    end
    if (_EVAL_105) begin
      _EVAL_2202 <= 1'h0;
    end else begin
      if (_EVAL_3675) begin
        _EVAL_2202 <= _EVAL_3769;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2209 <= 1'h0;
    end else begin
      if (_EVAL_788) begin
        _EVAL_2209 <= _EVAL_1919;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2214 <= 1'h0;
    end else begin
      if (_EVAL_2590) begin
        _EVAL_2214 <= _EVAL_3766;
      end
    end
    if (_EVAL_706) begin
      _EVAL_2231 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2254 <= 1'h0;
    end else begin
      if (_EVAL_274) begin
        _EVAL_2254 <= _EVAL_1136;
      end
    end
    if (_EVAL_2533) begin
      _EVAL_2256 <= _EVAL_3965;
    end
    if (_EVAL_2015) begin
      _EVAL_2290 <= _EVAL_3965;
    end
    if (_EVAL_359) begin
      _EVAL_2306 <= _EVAL_3965;
    end
    if (_EVAL_1403) begin
      _EVAL_2311 <= _EVAL_3965;
    end
    if (_EVAL_2439) begin
      _EVAL_2334 <= _EVAL_3965;
    end
    if (_EVAL_1355) begin
      _EVAL_2336 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2341 <= 1'h0;
    end else begin
      if (_EVAL_864) begin
        _EVAL_2341 <= _EVAL_3013;
      end
    end
    if (_EVAL_3214) begin
      _EVAL_2356 <= _EVAL_3965;
    end
    if (_EVAL_1271) begin
      _EVAL_2481 <= _EVAL_3965;
    end
    if (_EVAL_667) begin
      _EVAL_2484 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2485 <= 1'h0;
    end else begin
      if (_EVAL_2624) begin
        _EVAL_2485 <= _EVAL_401;
      end
    end
    if (_EVAL_2426) begin
      _EVAL_2491 <= _EVAL_3965;
    end
    if (_EVAL_2218) begin
      _EVAL_2500 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2507 <= 1'h0;
    end else begin
      if (_EVAL_3273) begin
        _EVAL_2507 <= _EVAL_2597;
      end
    end
    if (_EVAL_1232) begin
      _EVAL_2536 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2582 <= 1'h0;
    end else begin
      if (_EVAL_360) begin
        _EVAL_2582 <= _EVAL_2430;
      end
    end
    if (_EVAL_3353) begin
      _EVAL_2584 <= _EVAL_3965;
    end
    if (_EVAL_1027) begin
      _EVAL_2646 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2648 <= 1'h0;
    end else begin
      if (_EVAL_574) begin
        _EVAL_2648 <= _EVAL_2750;
      end
    end
    if (_EVAL_3744) begin
      _EVAL_2653 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2666 <= 1'h0;
    end else begin
      if (_EVAL_3799) begin
        _EVAL_2666 <= _EVAL_2421;
      end
    end
    if (_EVAL_3198) begin
      _EVAL_2677 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2684 <= 1'h0;
    end else begin
      if (_EVAL_248) begin
        _EVAL_2684 <= _EVAL_1564;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2688 <= 1'h0;
    end else begin
      if (_EVAL_1756) begin
        _EVAL_2688 <= _EVAL_1845;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2701 <= 1'h0;
    end else begin
      if (_EVAL_3566) begin
        _EVAL_2701 <= _EVAL_2574;
      end
    end
    if (_EVAL_3583) begin
      _EVAL_2720 <= _EVAL_3965;
    end
    if (_EVAL_1378) begin
      _EVAL_2754 <= _EVAL_3020;
    end
    if (_EVAL_571) begin
      _EVAL_2760 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2803 <= 1'h0;
    end else begin
      if (_EVAL_3263) begin
        _EVAL_2803 <= _EVAL_3945;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2807 <= 1'h0;
    end else begin
      if (_EVAL_2142) begin
        _EVAL_2807 <= _EVAL_2210;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2809 <= 1'h0;
    end else begin
      if (_EVAL_320) begin
        _EVAL_2809 <= _EVAL_2555;
      end
    end
    if (_EVAL_1682) begin
      _EVAL_2810 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2826 <= 1'h0;
    end else begin
      if (_EVAL_3993) begin
        _EVAL_2826 <= _EVAL_1251;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2838 <= 1'h0;
    end else begin
      if (_EVAL_220) begin
        _EVAL_2838 <= _EVAL_1414;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2850 <= 1'h0;
    end else begin
      if (_EVAL_1540) begin
        _EVAL_2850 <= _EVAL_2751;
      end
    end
    if (_EVAL_3774) begin
      _EVAL_2851 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2870 <= 1'h0;
    end else begin
      if (_EVAL_221) begin
        _EVAL_2870 <= _EVAL_3946;
      end
    end
    if (_EVAL_2097) begin
      _EVAL_2881 <= _EVAL_3965;
    end
    if (_EVAL_2697) begin
      _EVAL_2937 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2938 <= 1'h0;
    end else begin
      if (_EVAL_3581) begin
        _EVAL_2938 <= _EVAL_2206;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2942 <= 1'h0;
    end else begin
      if (_EVAL_3890) begin
        _EVAL_2942 <= _EVAL_3892;
      end
    end
    if (_EVAL_105) begin
      _EVAL_2953 <= 1'h0;
    end else begin
      if (_EVAL_1816) begin
        _EVAL_2953 <= _EVAL_1596;
      end
    end
    if (_EVAL_954) begin
      _EVAL_2958 <= _EVAL_3965;
    end
    if (_EVAL_1707) begin
      _EVAL_2965 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_2972 <= 1'h0;
    end else begin
      if (_EVAL_1159) begin
        _EVAL_2972 <= _EVAL_2917;
      end
    end
    if (_EVAL_313) begin
      _EVAL_3008 <= _EVAL_3965;
    end
    if (_EVAL_4001) begin
      _EVAL_3014 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3023 <= 1'h0;
    end else begin
      if (_EVAL_3100) begin
        _EVAL_3023 <= _EVAL_2404;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3025 <= 1'h0;
    end else begin
      if (_EVAL_3099) begin
        _EVAL_3025 <= _EVAL_2601;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3039 <= 1'h0;
    end else begin
      if (_EVAL_608) begin
        _EVAL_3039 <= _EVAL_570;
      end
    end
    if (_EVAL_2109) begin
      _EVAL_3056 <= _EVAL_3965;
    end
    if (_EVAL_190) begin
      _EVAL_3102 <= _EVAL_3965;
    end
    if (_EVAL_2845) begin
      _EVAL_3113 <= _EVAL_3965;
    end
    if (_EVAL_2770) begin
      _EVAL_3118 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3137 <= 1'h0;
    end else begin
      if (_EVAL_195) begin
        _EVAL_3137 <= _EVAL_252;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3167 <= 1'h0;
    end else begin
      if (_EVAL_2913) begin
        _EVAL_3167 <= _EVAL_2791;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3192 <= 1'h0;
    end else begin
      if (_EVAL_2739) begin
        _EVAL_3192 <= _EVAL_3641;
      end
    end
    if (_EVAL_2411) begin
      _EVAL_3195 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3199 <= 1'h0;
    end else begin
      if (_EVAL_199) begin
        _EVAL_3199 <= _EVAL_2156;
      end
    end
    if (_EVAL_975) begin
      _EVAL_3204 <= _EVAL_3965;
    end
    if (_EVAL_466) begin
      _EVAL_3216 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3222 <= 1'h0;
    end else begin
      if (_EVAL_3546) begin
        _EVAL_3222 <= _EVAL_1855;
      end
    end
    _EVAL_3235 <= PLICFanIn__EVAL_36;
    if (_EVAL_3460) begin
      _EVAL_3242 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3245 <= 1'h0;
    end else begin
      if (_EVAL_2902) begin
        _EVAL_3245 <= _EVAL_488;
      end
    end
    if (_EVAL_412) begin
      _EVAL_3267 <= _EVAL_3965;
    end
    if (_EVAL_3940) begin
      _EVAL_3274 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3279 <= 1'h0;
    end else begin
      if (_EVAL_299) begin
        _EVAL_3279 <= _EVAL_2084;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3283 <= 1'h0;
    end else begin
      if (_EVAL_3880) begin
        _EVAL_3283 <= _EVAL_1226;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3296 <= 1'h0;
    end else begin
      if (_EVAL_1144) begin
        _EVAL_3296 <= _EVAL_2885;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3299 <= 1'h0;
    end else begin
      if (_EVAL_1671) begin
        _EVAL_3299 <= _EVAL_1392;
      end
    end
    if (_EVAL_3284) begin
      _EVAL_3312 <= _EVAL_3965;
    end
    if (_EVAL_1309) begin
      _EVAL_3315 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3317 <= 1'h0;
    end else begin
      if (_EVAL_3586) begin
        _EVAL_3317 <= _EVAL_1434;
      end
    end
    if (_EVAL_2143) begin
      _EVAL_3331 <= _EVAL_3965;
    end
    if (_EVAL_1446) begin
      _EVAL_3336 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3359 <= 1'h0;
    end else begin
      if (_EVAL_2952) begin
        _EVAL_3359 <= _EVAL_773;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3361 <= 1'h0;
    end else begin
      if (_EVAL_986) begin
        _EVAL_3361 <= _EVAL_846;
      end
    end
    if (_EVAL_1025) begin
      _EVAL_3383 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3407 <= 1'h0;
    end else begin
      if (_EVAL_3169) begin
        _EVAL_3407 <= _EVAL_3751;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3419 <= 1'h0;
    end else begin
      if (_EVAL_457) begin
        _EVAL_3419 <= _EVAL_1927;
      end
    end
    if (_EVAL_2690) begin
      _EVAL_3421 <= _EVAL_3020;
    end
    if (_EVAL_2903) begin
      _EVAL_3488 <= _EVAL_688;
    end
    if (_EVAL_105) begin
      _EVAL_3505 <= 1'h0;
    end else begin
      if (_EVAL_2705) begin
        _EVAL_3505 <= _EVAL_2261;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3527 <= 1'h0;
    end else begin
      if (_EVAL_3519) begin
        _EVAL_3527 <= _EVAL_341;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3551 <= 1'h0;
    end else begin
      if (_EVAL_1259) begin
        _EVAL_3551 <= _EVAL_2628;
      end
    end
    if (_EVAL_1067) begin
      _EVAL_3552 <= _EVAL_3965;
    end
    if (_EVAL_1157) begin
      _EVAL_3554 <= _EVAL_3965;
    end
    if (_EVAL_3681) begin
      _EVAL_3563 <= _EVAL_3965;
    end
    if (_EVAL_3726) begin
      _EVAL_3571 <= _EVAL_3965;
    end
    if (_EVAL_3998) begin
      _EVAL_3573 <= _EVAL_3965;
    end
    if (_EVAL_1205) begin
      _EVAL_3591 <= _EVAL_3965;
    end
    if (_EVAL_1842) begin
      _EVAL_3608 <= _EVAL_3965;
    end
    if (_EVAL_2776) begin
      _EVAL_3623 <= _EVAL_2047;
    end
    if (_EVAL_105) begin
      _EVAL_3636 <= 1'h0;
    end else begin
      if (_EVAL_242) begin
        _EVAL_3636 <= _EVAL_1690;
      end
    end
    if (_EVAL_1957) begin
      _EVAL_3644 <= _EVAL_3965;
    end
    if (_EVAL_3738) begin
      _EVAL_3645 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3713 <= 1'h0;
    end else begin
      if (_EVAL_3852) begin
        _EVAL_3713 <= _EVAL_1843;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3715 <= 1'h0;
    end else begin
      if (_EVAL_1077) begin
        _EVAL_3715 <= _EVAL_1237;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3720 <= 1'h0;
    end else begin
      if (_EVAL_171) begin
        _EVAL_3720 <= _EVAL_3677;
      end
    end
    if (_EVAL_3618) begin
      _EVAL_3721 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3728 <= 1'h0;
    end else begin
      if (_EVAL_1021) begin
        _EVAL_3728 <= _EVAL_1244;
      end
    end
    if (_EVAL_2130) begin
      _EVAL_3731 <= _EVAL_3965;
    end
    if (_EVAL_1225) begin
      _EVAL_3733 <= _EVAL_3965;
    end
    if (_EVAL_1015) begin
      _EVAL_3740 <= _EVAL_3965;
    end
    if (_EVAL_316) begin
      _EVAL_3743 <= _EVAL_2047;
    end
    if (_EVAL_105) begin
      _EVAL_3750 <= 1'h0;
    end else begin
      if (_EVAL_2225) begin
        _EVAL_3750 <= _EVAL_3269;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3757 <= 1'h0;
    end else begin
      if (_EVAL_3426) begin
        _EVAL_3757 <= _EVAL_2064;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3759 <= 1'h0;
    end else begin
      if (_EVAL_2893) begin
        _EVAL_3759 <= _EVAL_3356;
      end
    end
    if (_EVAL_796) begin
      _EVAL_3768 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3783 <= 1'h0;
    end else begin
      if (_EVAL_2548) begin
        _EVAL_3783 <= _EVAL_3252;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3788 <= 1'h0;
    end else begin
      if (_EVAL_1246) begin
        _EVAL_3788 <= _EVAL_557;
      end
    end
    if (_EVAL_3234) begin
      _EVAL_3801 <= _EVAL_3965;
    end
    if (_EVAL_1178) begin
      _EVAL_3804 <= _EVAL_3965;
    end
    if (_EVAL_315) begin
      _EVAL_3843 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3850 <= 1'h0;
    end else begin
      if (_EVAL_3431) begin
        _EVAL_3850 <= _EVAL_1986;
      end
    end
    if (_EVAL_2563) begin
      _EVAL_3870 <= _EVAL_3020;
    end
    if (_EVAL_105) begin
      _EVAL_3899 <= 1'h0;
    end else begin
      if (_EVAL_4032) begin
        _EVAL_3899 <= _EVAL_1559;
      end
    end
    if (_EVAL_1042) begin
      _EVAL_3909 <= _EVAL_3965;
    end
    if (_EVAL_1663) begin
      _EVAL_3913 <= _EVAL_1861;
    end
    if (_EVAL_182) begin
      _EVAL_3943 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_3964 <= 1'h0;
    end else begin
      if (_EVAL_3265) begin
        _EVAL_3964 <= _EVAL_4056;
      end
    end
    if (_EVAL_105) begin
      _EVAL_3996 <= 1'h0;
    end else begin
      if (_EVAL_865) begin
        _EVAL_3996 <= _EVAL_1751;
      end
    end
    if (_EVAL_479) begin
      _EVAL_4013 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_4034 <= 1'h0;
    end else begin
      if (_EVAL_214) begin
        _EVAL_4034 <= _EVAL_1479;
      end
    end
    if (_EVAL_691) begin
      _EVAL_4050 <= _EVAL_3965;
    end
    if (_EVAL_105) begin
      _EVAL_4063 <= 1'h0;
    end else begin
      if (_EVAL_1614) begin
        _EVAL_4063 <= _EVAL_1858;
      end
    end
    if (_EVAL_1337) begin
      _EVAL_4066 <= _EVAL_3965;
    end
  end
endmodule
