//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_123_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [6:0]  _EVAL_7,
  input  [13:0] _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input  [6:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_38;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_42;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_127;
  reg [31:0] _RAND_2;
  reg [5:0] _EVAL_142;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_170;
  reg [31:0] _RAND_4;
  reg [72:0] _EVAL_173;
  reg [95:0] _RAND_5;
  reg [3:0] _EVAL_207;
  reg [31:0] _RAND_6;
  reg [6:0] _EVAL_217;
  reg [31:0] _RAND_7;
  reg [5:0] _EVAL_237;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_243;
  reg [31:0] _RAND_9;
  reg [13:0] _EVAL_251;
  reg [31:0] _RAND_10;
  reg [5:0] _EVAL_254;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_273;
  reg [31:0] _RAND_12;
  reg [6:0] _EVAL_295;
  reg [31:0] _RAND_13;
  wire  _EVAL_192;
  wire [1:0] _EVAL_77;
  wire [1:0] _EVAL_167;
  wire  _EVAL_265;
  wire  _EVAL_246;
  wire  _EVAL_122;
  wire  _EVAL_232;
  wire  _EVAL_40;
  wire  _EVAL_163;
  wire  _EVAL_298;
  wire  _EVAL_97;
  wire [127:0] _EVAL_125;
  wire [127:0] _EVAL_226;
  wire [72:0] _EVAL_143;
  wire [72:0] _EVAL_116;
  wire [72:0] _EVAL_35;
  wire  _EVAL_105;
  wire  _EVAL_140;
  wire  _EVAL_21;
  wire [2:0] _EVAL_294;
  wire  _EVAL_101;
  wire  _EVAL_137;
  wire  _EVAL_196;
  wire  _EVAL_227;
  wire  _EVAL_138;
  wire [22:0] _EVAL_181;
  wire [7:0] _EVAL_156;
  wire [7:0] _EVAL_281;
  wire [5:0] _EVAL_81;
  wire [5:0] _EVAL_212;
  wire  _EVAL_128;
  wire  _EVAL_58;
  wire  _EVAL_60;
  wire [3:0] _EVAL_49;
  wire  _EVAL_255;
  wire [2:0] _EVAL_183;
  wire  _EVAL_56;
  wire  _EVAL_98;
  wire  _EVAL_111;
  wire  _EVAL_287;
  wire  _EVAL_65;
  wire  _EVAL_57;
  wire  _EVAL_147;
  wire  _EVAL_130;
  wire  _EVAL_70;
  wire  _EVAL_19;
  wire  _EVAL_126;
  wire  _EVAL_83;
  wire  _EVAL_28;
  wire  _EVAL_61;
  wire  _EVAL_200;
  wire  _EVAL_110;
  wire  _EVAL_230;
  wire  _EVAL_145;
  wire  _EVAL_53;
  wire  _EVAL_129;
  wire  _EVAL_191;
  wire  _EVAL_34;
  wire  _EVAL_228;
  wire  _EVAL_185;
  wire  _EVAL_283;
  wire  _EVAL_271;
  wire  _EVAL_219;
  wire  _EVAL_204;
  wire  _EVAL_155;
  wire  _EVAL_288;
  wire  _EVAL_29;
  wire  _EVAL_233;
  wire  _EVAL_115;
  wire  _EVAL_258;
  wire  _EVAL_133;
  wire  _EVAL_73;
  wire [3:0] _EVAL_221;
  wire  _EVAL_260;
  wire  _EVAL_248;
  wire [22:0] _EVAL_88;
  wire [7:0] _EVAL_31;
  wire [7:0] _EVAL_44;
  wire [5:0] _EVAL_36;
  wire  _EVAL_266;
  wire  _EVAL_199;
  wire  _EVAL_102;
  wire  _EVAL_108;
  wire  _EVAL_247;
  wire  _EVAL_250;
  wire  _EVAL_162;
  wire  _EVAL_93;
  wire  _EVAL_176;
  wire  _EVAL_20;
  wire [3:0] _EVAL_54;
  wire  _EVAL_112;
  wire [13:0] _EVAL_187;
  wire [14:0] _EVAL_291;
  wire  _EVAL_141;
  wire  _EVAL_244;
  wire  _EVAL_236;
  wire  _EVAL_180;
  wire  _EVAL_68;
  wire  _EVAL_104;
  wire  _EVAL_94;
  wire [127:0] _EVAL_166;
  wire [127:0] _EVAL_85;
  wire [72:0] _EVAL_120;
  wire [72:0] _EVAL_67;
  wire [3:0] _EVAL_30;
  wire [3:0] _EVAL_134;
  wire [3:0] _EVAL_62;
  wire  _EVAL_252;
  wire  _EVAL_216;
  wire  _EVAL_69;
  wire  _EVAL_229;
  wire  _EVAL_178;
  wire  _EVAL_75;
  wire  _EVAL_205;
  wire  _EVAL_224;
  wire  _EVAL_24;
  wire  _EVAL_272;
  wire  _EVAL_285;
  wire  _EVAL_293;
  wire  _EVAL_76;
  wire  _EVAL_165;
  wire  _EVAL_179;
  wire  _EVAL_231;
  wire  _EVAL_106;
  wire  _EVAL_113;
  wire  _EVAL_189;
  wire  _EVAL_84;
  wire  _EVAL_282;
  wire  _EVAL_259;
  wire  _EVAL_239;
  wire  _EVAL_18;
  wire  _EVAL_203;
  wire  _EVAL_245;
  wire  _EVAL_161;
  wire [72:0] _EVAL_171;
  wire [72:0] _EVAL_209;
  wire [72:0] _EVAL_121;
  wire  _EVAL_214;
  wire  _EVAL_89;
  wire  _EVAL_74;
  wire  _EVAL_17;
  wire  _EVAL_175;
  wire [5:0] _EVAL_268;
  wire  _EVAL_249;
  wire  _EVAL_146;
  wire  _EVAL_131;
  wire  _EVAL_264;
  wire  _EVAL_208;
  wire  _EVAL_132;
  wire  _EVAL_160;
  wire  _EVAL_186;
  wire  _EVAL_284;
  wire  _EVAL_276;
  wire  _EVAL_218;
  wire  _EVAL_151;
  wire  _EVAL_159;
  wire  _EVAL_280;
  wire [5:0] _EVAL_234;
  wire [14:0] _EVAL_52;
  wire  _EVAL_72;
  wire  _EVAL_241;
  wire  _EVAL_198;
  wire  _EVAL_124;
  wire  _EVAL_222;
  wire  _EVAL_193;
  wire  _EVAL_242;
  wire  _EVAL_211;
  wire  _EVAL_292;
  wire  _EVAL_262;
  wire  _EVAL_257;
  wire  _EVAL_174;
  wire [14:0] _EVAL_261;
  wire  _EVAL_87;
  wire  _EVAL_99;
  wire  _EVAL_26;
  wire  _EVAL_263;
  wire  _EVAL_107;
  wire  _EVAL_22;
  wire  _EVAL_190;
  wire  _EVAL_103;
  wire  _EVAL_210;
  wire  _EVAL_33;
  wire  _EVAL_289;
  wire  _EVAL_150;
  wire  _EVAL_201;
  wire  _EVAL_71;
  wire  _EVAL_48;
  wire  _EVAL_80;
  wire  _EVAL_154;
  wire  _EVAL_96;
  wire  _EVAL_275;
  wire  _EVAL_296;
  wire  _EVAL_153;
  wire  _EVAL_256;
  wire  _EVAL_144;
  wire  _EVAL_297;
  wire  _EVAL_135;
  wire  _EVAL_177;
  wire  _EVAL_123;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_37;
  wire  _EVAL_136;
  wire  _EVAL_100;
  wire  _EVAL_157;
  wire  _EVAL_119;
  wire [13:0] _EVAL_91;
  wire [13:0] _EVAL_182;
  wire  _EVAL_39;
  wire  _EVAL_23;
  wire  _EVAL_172;
  wire  _EVAL_109;
  wire  _EVAL_51;
  wire  _EVAL_45;
  wire  _EVAL_43;
  wire  _EVAL_92;
  wire  _EVAL_90;
  wire  _EVAL_206;
  wire  _EVAL_253;
  wire  _EVAL_269;
  wire  _EVAL_41;
  wire  _EVAL_290;
  wire  _EVAL_240;
  wire  _EVAL_202;
  wire  _EVAL_63;
  wire  _EVAL_235;
  wire  _EVAL_139;
  wire [5:0] _EVAL_164;
  wire  _EVAL_184;
  wire  _EVAL_95;
  wire  _EVAL_47;
  wire  _EVAL_238;
  wire  _EVAL_168;
  wire  _EVAL_79;
  wire  _EVAL_59;
  wire  _EVAL_117;
  wire  _EVAL_195;
  wire [31:0] _EVAL_152;
  wire  _EVAL_50;
  wire  _EVAL_223;
  wire  _EVAL_194;
  wire  _EVAL_286;
  wire  _EVAL_78;
  wire  _EVAL_82;
  wire  _EVAL_267;
  wire  _EVAL_277;
  wire  _EVAL_158;
  wire  _EVAL_64;
  wire  _EVAL_118;
  wire  _EVAL_220;
  wire  _EVAL_46;
  wire  _EVAL_25;
  wire  _EVAL_27;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_192 = _EVAL_9[0];
  assign _EVAL_77 = 2'h1 << _EVAL_192;
  assign _EVAL_167 = _EVAL_77 | 2'h1;
  assign _EVAL_265 = _EVAL_167[0];
  assign _EVAL_246 = _EVAL_8[1];
  assign _EVAL_122 = _EVAL_8[0];
  assign _EVAL_232 = _EVAL_246 & _EVAL_122;
  assign _EVAL_40 = _EVAL_265 & _EVAL_232;
  assign _EVAL_163 = _EVAL_6 & _EVAL_10;
  assign _EVAL_298 = _EVAL_254 == 6'h0;
  assign _EVAL_97 = _EVAL_163 & _EVAL_298;
  assign _EVAL_125 = 128'h1 << _EVAL_11;
  assign _EVAL_226 = _EVAL_97 ? _EVAL_125 : 128'h0;
  assign _EVAL_143 = _EVAL_226[72:0];
  assign _EVAL_116 = _EVAL_143 | _EVAL_173;
  assign _EVAL_35 = _EVAL_116 >> _EVAL_7;
  assign _EVAL_105 = _EVAL_35[0];
  assign _EVAL_140 = _EVAL_3 == 3'h1;
  assign _EVAL_21 = _EVAL_10 & _EVAL_140;
  assign _EVAL_294 = _EVAL_11[2:0];
  assign _EVAL_101 = 3'h1 <= _EVAL_294;
  assign _EVAL_137 = _EVAL_5 <= 3'h2;
  assign _EVAL_196 = _EVAL_137 | _EVAL_13;
  assign _EVAL_227 = _EVAL_3[2];
  assign _EVAL_138 = _EVAL_227 == 1'h0;
  assign _EVAL_181 = 23'hff << _EVAL_9;
  assign _EVAL_156 = _EVAL_181[7:0];
  assign _EVAL_281 = ~ _EVAL_156;
  assign _EVAL_81 = _EVAL_281[7:2];
  assign _EVAL_212 = _EVAL_254 - 6'h1;
  assign _EVAL_128 = _EVAL & _EVAL_15;
  assign _EVAL_58 = _EVAL_237 == 6'h0;
  assign _EVAL_60 = _EVAL_128 & _EVAL_58;
  assign _EVAL_49 = _EVAL_7[6:3];
  assign _EVAL_255 = _EVAL_49 == 4'h8;
  assign _EVAL_183 = _EVAL_7[2:0];
  assign _EVAL_56 = 3'h1 <= _EVAL_183;
  assign _EVAL_98 = _EVAL_255 & _EVAL_56;
  assign _EVAL_111 = _EVAL_0 == _EVAL_38;
  assign _EVAL_287 = _EVAL_111 | _EVAL_13;
  assign _EVAL_65 = _EVAL_287 == 1'h0;
  assign _EVAL_57 = _EVAL_8 == _EVAL_251;
  assign _EVAL_147 = _EVAL_57 | _EVAL_13;
  assign _EVAL_130 = _EVAL_147 == 1'h0;
  assign _EVAL_70 = _EVAL_5 == _EVAL_127;
  assign _EVAL_19 = _EVAL_70 | _EVAL_13;
  assign _EVAL_126 = _EVAL_19 == 1'h0;
  assign _EVAL_83 = _EVAL_7 == 7'h48;
  assign _EVAL_28 = _EVAL_7 == 7'h40;
  assign _EVAL_61 = _EVAL_83 | _EVAL_28;
  assign _EVAL_200 = _EVAL_61 | _EVAL_98;
  assign _EVAL_110 = _EVAL_7 == 7'h20;
  assign _EVAL_230 = _EVAL_200 | _EVAL_110;
  assign _EVAL_145 = _EVAL_173 != 73'h0;
  assign _EVAL_53 = _EVAL_145 == 1'h0;
  assign _EVAL_129 = plusarg_reader_out == 32'h0;
  assign _EVAL_191 = _EVAL_53 | _EVAL_129;
  assign _EVAL_34 = _EVAL_273 < plusarg_reader_out;
  assign _EVAL_228 = _EVAL_191 | _EVAL_34;
  assign _EVAL_185 = _EVAL_228 | _EVAL_13;
  assign _EVAL_283 = _EVAL_9 >= 4'h2;
  assign _EVAL_271 = _EVAL_167[1];
  assign _EVAL_219 = _EVAL_246 == 1'h0;
  assign _EVAL_204 = _EVAL_271 & _EVAL_219;
  assign _EVAL_155 = _EVAL_283 | _EVAL_204;
  assign _EVAL_288 = _EVAL_122 == 1'h0;
  assign _EVAL_29 = _EVAL_219 & _EVAL_288;
  assign _EVAL_233 = _EVAL_265 & _EVAL_29;
  assign _EVAL_115 = _EVAL_155 | _EVAL_233;
  assign _EVAL_258 = _EVAL_185 == 1'h0;
  assign _EVAL_133 = _EVAL_0 == 3'h2;
  assign _EVAL_73 = _EVAL_15 & _EVAL_133;
  assign _EVAL_221 = _EVAL_11[6:3];
  assign _EVAL_260 = _EVAL_221 == 4'h8;
  assign _EVAL_248 = _EVAL_5 != 3'h0;
  assign _EVAL_88 = 23'hff << _EVAL_12;
  assign _EVAL_31 = _EVAL_88[7:0];
  assign _EVAL_44 = ~ _EVAL_31;
  assign _EVAL_36 = _EVAL_44[7:2];
  assign _EVAL_266 = _EVAL_11 == 7'h48;
  assign _EVAL_199 = _EVAL_271 & _EVAL_246;
  assign _EVAL_102 = _EVAL_283 | _EVAL_199;
  assign _EVAL_108 = _EVAL_102 | _EVAL_40;
  assign _EVAL_247 = _EVAL_246 & _EVAL_288;
  assign _EVAL_250 = _EVAL_265 & _EVAL_247;
  assign _EVAL_162 = _EVAL_102 | _EVAL_250;
  assign _EVAL_93 = _EVAL_219 & _EVAL_122;
  assign _EVAL_176 = _EVAL_265 & _EVAL_93;
  assign _EVAL_20 = _EVAL_155 | _EVAL_176;
  assign _EVAL_54 = {_EVAL_108,_EVAL_162,_EVAL_20,_EVAL_115};
  assign _EVAL_112 = _EVAL_1 == _EVAL_54;
  assign _EVAL_187 = _EVAL_8 ^ 14'h3000;
  assign _EVAL_291 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_141 = _EVAL_0 <= 3'h6;
  assign _EVAL_244 = _EVAL_141 | _EVAL_13;
  assign _EVAL_236 = _EVAL_244 == 1'h0;
  assign _EVAL_180 = _EVAL_3 == 3'h3;
  assign _EVAL_68 = _EVAL_0 == 3'h6;
  assign _EVAL_104 = _EVAL_68 == 1'h0;
  assign _EVAL_94 = _EVAL_60 & _EVAL_104;
  assign _EVAL_166 = 128'h1 << _EVAL_7;
  assign _EVAL_85 = _EVAL_94 ? _EVAL_166 : 128'h0;
  assign _EVAL_120 = _EVAL_85[72:0];
  assign _EVAL_67 = ~ _EVAL_120;
  assign _EVAL_30 = ~ _EVAL_1;
  assign _EVAL_134 = ~ _EVAL_54;
  assign _EVAL_62 = _EVAL_1 & _EVAL_134;
  assign _EVAL_252 = _EVAL_62 == 4'h0;
  assign _EVAL_216 = _EVAL_252 | _EVAL_13;
  assign _EVAL_69 = _EVAL_12 == _EVAL_207;
  assign _EVAL_229 = _EVAL_69 | _EVAL_13;
  assign _EVAL_178 = _EVAL_49 == 4'h0;
  assign _EVAL_75 = _EVAL_230 | _EVAL_178;
  assign _EVAL_205 = _EVAL_49 == 4'h1;
  assign _EVAL_224 = _EVAL_75 | _EVAL_205;
  assign _EVAL_24 = _EVAL_49 == 4'h2;
  assign _EVAL_272 = _EVAL_224 | _EVAL_24;
  assign _EVAL_285 = _EVAL_49 == 4'h3;
  assign _EVAL_293 = _EVAL_272 | _EVAL_285;
  assign _EVAL_76 = _EVAL_3 == 3'h7;
  assign _EVAL_165 = _EVAL_10 & _EVAL_76;
  assign _EVAL_179 = _EVAL_11 == 7'h40;
  assign _EVAL_231 = _EVAL_266 | _EVAL_179;
  assign _EVAL_106 = _EVAL_260 & _EVAL_101;
  assign _EVAL_113 = _EVAL_231 | _EVAL_106;
  assign _EVAL_189 = _EVAL_0 == 3'h0;
  assign _EVAL_84 = _EVAL_15 & _EVAL_189;
  assign _EVAL_282 = _EVAL_11 == _EVAL_295;
  assign _EVAL_259 = _EVAL_282 | _EVAL_13;
  assign _EVAL_239 = _EVAL_9 == _EVAL_170;
  assign _EVAL_18 = _EVAL_239 | _EVAL_13;
  assign _EVAL_203 = _EVAL_18 == 1'h0;
  assign _EVAL_245 = _EVAL_3 == 3'h2;
  assign _EVAL_161 = _EVAL_10 & _EVAL_245;
  assign _EVAL_171 = _EVAL_173 | _EVAL_143;
  assign _EVAL_209 = _EVAL_171 & _EVAL_67;
  assign _EVAL_121 = _EVAL_173 >> _EVAL_11;
  assign _EVAL_214 = _EVAL_143 != 73'h0;
  assign _EVAL_89 = _EVAL_214 == 1'h0;
  assign _EVAL_74 = _EVAL_10 & _EVAL_180;
  assign _EVAL_17 = _EVAL_142 == 6'h0;
  assign _EVAL_175 = _EVAL_0[0];
  assign _EVAL_268 = _EVAL_142 - 6'h1;
  assign _EVAL_249 = _EVAL_11 == 7'h20;
  assign _EVAL_146 = _EVAL_113 | _EVAL_249;
  assign _EVAL_131 = _EVAL_221 == 4'h0;
  assign _EVAL_264 = _EVAL_146 | _EVAL_131;
  assign _EVAL_208 = _EVAL_221 == 4'h1;
  assign _EVAL_132 = _EVAL_264 | _EVAL_208;
  assign _EVAL_160 = _EVAL_221 == 4'h2;
  assign _EVAL_186 = _EVAL_132 | _EVAL_160;
  assign _EVAL_284 = _EVAL_128 & _EVAL_17;
  assign _EVAL_276 = _EVAL_143 != _EVAL_120;
  assign _EVAL_218 = _EVAL_276 | _EVAL_89;
  assign _EVAL_151 = _EVAL_218 | _EVAL_13;
  assign _EVAL_159 = _EVAL_151 == 1'h0;
  assign _EVAL_280 = _EVAL_243 == 6'h0;
  assign _EVAL_234 = _EVAL_243 - 6'h1;
  assign _EVAL_52 = $signed(_EVAL_291) & $signed(-15'sh1000);
  assign _EVAL_72 = _EVAL_17 == 1'h0;
  assign _EVAL_241 = _EVAL_9 <= 4'h8;
  assign _EVAL_198 = _EVAL_283 | _EVAL_13;
  assign _EVAL_124 = _EVAL_198 == 1'h0;
  assign _EVAL_222 = _EVAL_112 | _EVAL_13;
  assign _EVAL_193 = _EVAL_222 == 1'h0;
  assign _EVAL_242 = _EVAL_9 <= 4'h2;
  assign _EVAL_211 = _EVAL_12 >= 4'h2;
  assign _EVAL_292 = _EVAL_211 | _EVAL_13;
  assign _EVAL_262 = _EVAL_292 == 1'h0;
  assign _EVAL_257 = _EVAL_5 == 3'h0;
  assign _EVAL_174 = _EVAL_257 | _EVAL_13;
  assign _EVAL_261 = $signed(_EVAL_52);
  assign _EVAL_87 = $signed(_EVAL_261) == $signed(15'sh0);
  assign _EVAL_99 = _EVAL_242 & _EVAL_87;
  assign _EVAL_26 = _EVAL_105 | _EVAL_13;
  assign _EVAL_263 = _EVAL_26 == 1'h0;
  assign _EVAL_107 = _EVAL_3 == _EVAL_42;
  assign _EVAL_22 = _EVAL_107 | _EVAL_13;
  assign _EVAL_190 = _EVAL_22 == 1'h0;
  assign _EVAL_103 = _EVAL_5 <= 3'h3;
  assign _EVAL_210 = _EVAL_103 | _EVAL_13;
  assign _EVAL_33 = _EVAL_210 == 1'h0;
  assign _EVAL_289 = _EVAL_3 == 3'h4;
  assign _EVAL_150 = _EVAL_10 & _EVAL_289;
  assign _EVAL_201 = _EVAL_3 == 3'h5;
  assign _EVAL_71 = _EVAL_10 & _EVAL_201;
  assign _EVAL_48 = _EVAL_241 & _EVAL_87;
  assign _EVAL_80 = _EVAL_48 | _EVAL_13;
  assign _EVAL_154 = _EVAL_80 == 1'h0;
  assign _EVAL_96 = _EVAL_2 == 1'h0;
  assign _EVAL_275 = _EVAL_96 | _EVAL_13;
  assign _EVAL_296 = _EVAL_275 == 1'h0;
  assign _EVAL_153 = 4'h6 == _EVAL_9;
  assign _EVAL_256 = _EVAL_3 == 3'h0;
  assign _EVAL_144 = _EVAL_163 & _EVAL_280;
  assign _EVAL_297 = _EVAL_221 == 4'h3;
  assign _EVAL_135 = _EVAL_186 | _EVAL_297;
  assign _EVAL_177 = _EVAL_248 | _EVAL_13;
  assign _EVAL_123 = _EVAL_177 == 1'h0;
  assign _EVAL_148 = _EVAL_30 == 4'h0;
  assign _EVAL_149 = _EVAL_148 | _EVAL_13;
  assign _EVAL_37 = _EVAL_0 == 3'h4;
  assign _EVAL_136 = _EVAL_15 & _EVAL_37;
  assign _EVAL_100 = _EVAL_135 | _EVAL_13;
  assign _EVAL_157 = _EVAL_100 == 1'h0;
  assign _EVAL_119 = _EVAL_293 | _EVAL_13;
  assign _EVAL_91 = {{6'd0}, _EVAL_281};
  assign _EVAL_182 = _EVAL_8 & _EVAL_91;
  assign _EVAL_39 = _EVAL_3 == 3'h6;
  assign _EVAL_23 = _EVAL_14 | _EVAL_13;
  assign _EVAL_172 = _EVAL_196 == 1'h0;
  assign _EVAL_109 = _EVAL_0 == 3'h1;
  assign _EVAL_51 = _EVAL_14 == 1'h0;
  assign _EVAL_45 = _EVAL_51 | _EVAL_13;
  assign _EVAL_43 = _EVAL_45 == 1'h0;
  assign _EVAL_92 = _EVAL_182 == 14'h0;
  assign _EVAL_90 = _EVAL_92 | _EVAL_13;
  assign _EVAL_206 = _EVAL_90 == 1'h0;
  assign _EVAL_253 = _EVAL_121[0];
  assign _EVAL_269 = _EVAL_253 == 1'h0;
  assign _EVAL_41 = _EVAL_13 == 1'h0;
  assign _EVAL_290 = _EVAL_119 == 1'h0;
  assign _EVAL_240 = _EVAL_179 ? _EVAL_153 : 1'h0;
  assign _EVAL_202 = _EVAL_240 | _EVAL_13;
  assign _EVAL_63 = _EVAL_202 == 1'h0;
  assign _EVAL_235 = _EVAL_23 == 1'h0;
  assign _EVAL_139 = _EVAL_15 & _EVAL_109;
  assign _EVAL_164 = _EVAL_237 - 6'h1;
  assign _EVAL_184 = _EVAL_10 & _EVAL_39;
  assign _EVAL_95 = _EVAL_7 == _EVAL_217;
  assign _EVAL_47 = _EVAL_95 | _EVAL_13;
  assign _EVAL_238 = _EVAL_47 == 1'h0;
  assign _EVAL_168 = _EVAL_15 & _EVAL_72;
  assign _EVAL_79 = _EVAL_174 == 1'h0;
  assign _EVAL_59 = _EVAL_269 | _EVAL_13;
  assign _EVAL_117 = _EVAL_0 == 3'h5;
  assign _EVAL_195 = _EVAL_15 & _EVAL_117;
  assign _EVAL_152 = _EVAL_273 + 32'h1;
  assign _EVAL_50 = _EVAL_229 == 1'h0;
  assign _EVAL_223 = _EVAL_259 == 1'h0;
  assign _EVAL_194 = _EVAL_5 <= 3'h4;
  assign _EVAL_286 = _EVAL_194 | _EVAL_13;
  assign _EVAL_78 = _EVAL_286 == 1'h0;
  assign _EVAL_82 = _EVAL_99 | _EVAL_13;
  assign _EVAL_267 = _EVAL_82 == 1'h0;
  assign _EVAL_277 = _EVAL_216 == 1'h0;
  assign _EVAL_158 = _EVAL_280 == 1'h0;
  assign _EVAL_64 = _EVAL_10 & _EVAL_158;
  assign _EVAL_118 = _EVAL_10 & _EVAL_256;
  assign _EVAL_220 = _EVAL_163 | _EVAL_128;
  assign _EVAL_46 = _EVAL_15 & _EVAL_68;
  assign _EVAL_25 = _EVAL_149 == 1'h0;
  assign _EVAL_27 = _EVAL_59 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_38 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_42 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_127 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_142 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_170 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  _EVAL_173 = _RAND_5[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_207 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_217 = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_237 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_243 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_251 = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_254 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_273 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_295 = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_284) begin
      _EVAL_38 <= _EVAL_0;
    end
    if (_EVAL_144) begin
      _EVAL_42 <= _EVAL_3;
    end
    if (_EVAL_144) begin
      _EVAL_127 <= _EVAL_5;
    end
    if (_EVAL_13) begin
      _EVAL_142 <= 6'h0;
    end else begin
      if (_EVAL_128) begin
        if (_EVAL_17) begin
          if (_EVAL_175) begin
            _EVAL_142 <= _EVAL_36;
          end else begin
            _EVAL_142 <= 6'h0;
          end
        end else begin
          _EVAL_142 <= _EVAL_268;
        end
      end
    end
    if (_EVAL_144) begin
      _EVAL_170 <= _EVAL_9;
    end
    if (_EVAL_13) begin
      _EVAL_173 <= 73'h0;
    end else begin
      _EVAL_173 <= _EVAL_209;
    end
    if (_EVAL_284) begin
      _EVAL_207 <= _EVAL_12;
    end
    if (_EVAL_284) begin
      _EVAL_217 <= _EVAL_7;
    end
    if (_EVAL_13) begin
      _EVAL_237 <= 6'h0;
    end else begin
      if (_EVAL_128) begin
        if (_EVAL_58) begin
          if (_EVAL_175) begin
            _EVAL_237 <= _EVAL_36;
          end else begin
            _EVAL_237 <= 6'h0;
          end
        end else begin
          _EVAL_237 <= _EVAL_164;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_243 <= 6'h0;
    end else begin
      if (_EVAL_163) begin
        if (_EVAL_280) begin
          if (_EVAL_138) begin
            _EVAL_243 <= _EVAL_81;
          end else begin
            _EVAL_243 <= 6'h0;
          end
        end else begin
          _EVAL_243 <= _EVAL_234;
        end
      end
    end
    if (_EVAL_144) begin
      _EVAL_251 <= _EVAL_8;
    end
    if (_EVAL_13) begin
      _EVAL_254 <= 6'h0;
    end else begin
      if (_EVAL_163) begin
        if (_EVAL_298) begin
          if (_EVAL_138) begin
            _EVAL_254 <= _EVAL_81;
          end else begin
            _EVAL_254 <= 6'h0;
          end
        end else begin
          _EVAL_254 <= _EVAL_212;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_273 <= 32'h0;
    end else begin
      if (_EVAL_220) begin
        _EVAL_273 <= 32'h0;
      end else begin
        _EVAL_273 <= _EVAL_152;
      end
    end
    if (_EVAL_144) begin
      _EVAL_295 <= _EVAL_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e1702be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7ab2b43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf87cd8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8c54842)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2ca273e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22f18dd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4df809a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e58ab7a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b42c1963)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f500673)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb75be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb434cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89d0c247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd5c382d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a44afbd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(285f7329)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73fb9d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8241cd68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1766f8b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6638bbe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b2834f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7badc8e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbaef6f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fa1294d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f947cd44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c5d1efa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8123e1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfb3b714)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(312205f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0660086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d452264f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(867057fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69738b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bafb24fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b729448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea40719e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f989a5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(584769d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2801f87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a850d32d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba2de6fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c468a740)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81cf64f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da185ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(837578dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2ae0420)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3de3677)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc00f87d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e63c44c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(987c7e87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14eba7af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcad3178)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a9c7882)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ec765ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e701518)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53b313ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bf53f59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c40a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e0e751d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(457f3987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ef0534c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60484da7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42158045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb5e3677)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6086441a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8052c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74c0c8b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(759d50a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd29ff56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(352128a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1be2857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdf83612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c17f23c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78fb97f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12952b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ff738e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffc70349)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c324123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce0d3a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
