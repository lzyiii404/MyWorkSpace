//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_153_assert(
  input  [2:0]  _EVAL,
  input  [6:0]  _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [14:0] _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [6:0]  _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_83;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_115;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_129;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_140;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_149;
  reg [31:0] _RAND_4;
  reg [6:0] _EVAL_152;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_153;
  reg [31:0] _RAND_6;
  reg [6:0] _EVAL_161;
  reg [31:0] _RAND_7;
  reg [72:0] _EVAL_184;
  reg [95:0] _RAND_8;
  reg [3:0] _EVAL_191;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_200;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_208;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_278;
  reg [31:0] _RAND_12;
  reg [14:0] _EVAL_284;
  reg [31:0] _RAND_13;
  wire [12:0] _EVAL_39;
  wire [5:0] _EVAL_233;
  wire [5:0] _EVAL_175;
  wire [14:0] _EVAL_22;
  wire [14:0] _EVAL_276;
  wire  _EVAL_282;
  wire  _EVAL_92;
  wire  _EVAL_195;
  wire  _EVAL_183;
  wire  _EVAL_41;
  wire  _EVAL_135;
  wire  _EVAL_48;
  wire  _EVAL_221;
  wire  _EVAL_75;
  wire  _EVAL_265;
  wire [3:0] _EVAL_43;
  wire  _EVAL_146;
  wire [2:0] _EVAL_68;
  wire  _EVAL_24;
  wire  _EVAL_180;
  wire  _EVAL_269;
  wire  _EVAL_263;
  wire  _EVAL_193;
  wire [3:0] _EVAL_279;
  wire  _EVAL_216;
  wire  _EVAL_262;
  wire [1:0] _EVAL_80;
  wire [1:0] _EVAL_203;
  wire  _EVAL_72;
  wire  _EVAL_272;
  wire  _EVAL_242;
  wire  _EVAL_34;
  wire  _EVAL_81;
  wire  _EVAL_170;
  wire  _EVAL_125;
  wire  _EVAL_209;
  wire  _EVAL_53;
  wire [127:0] _EVAL_266;
  wire [127:0] _EVAL_160;
  wire [72:0] _EVAL_95;
  wire  _EVAL_245;
  wire  _EVAL_229;
  wire  _EVAL_204;
  wire  _EVAL_267;
  wire  _EVAL_164;
  wire  _EVAL_90;
  wire [127:0] _EVAL_220;
  wire [127:0] _EVAL_287;
  wire [72:0] _EVAL_89;
  wire  _EVAL_154;
  wire  _EVAL_118;
  wire  _EVAL_35;
  wire  _EVAL_222;
  wire  _EVAL_162;
  wire [3:0] _EVAL_138;
  wire  _EVAL_261;
  wire [72:0] _EVAL_70;
  wire  _EVAL_113;
  wire  _EVAL_254;
  wire [72:0] _EVAL_134;
  wire [72:0] _EVAL_33;
  wire  _EVAL_130;
  wire  _EVAL_274;
  wire  _EVAL_219;
  wire  _EVAL_112;
  wire  _EVAL_199;
  wire  _EVAL_51;
  wire  _EVAL_163;
  wire  _EVAL_165;
  wire  _EVAL_214;
  wire  _EVAL_65;
  wire  _EVAL_240;
  wire  _EVAL_63;
  wire  _EVAL_42;
  wire [3:0] _EVAL_234;
  wire  _EVAL_121;
  wire [72:0] _EVAL_173;
  wire  _EVAL_252;
  wire  _EVAL_38;
  wire [3:0] _EVAL_110;
  wire  _EVAL_258;
  wire  _EVAL_176;
  wire  _EVAL_74;
  wire  _EVAL_84;
  wire  _EVAL_102;
  wire  _EVAL_78;
  wire  _EVAL_257;
  wire  _EVAL_26;
  wire  _EVAL_277;
  wire  _EVAL_127;
  wire  _EVAL_69;
  wire  _EVAL_120;
  wire  _EVAL_155;
  wire  _EVAL_167;
  wire  _EVAL_223;
  wire [3:0] _EVAL_31;
  wire [3:0] _EVAL_142;
  wire [3:0] _EVAL_228;
  wire  _EVAL_30;
  wire  _EVAL_15;
  wire  _EVAL_190;
  wire  _EVAL_97;
  wire [31:0] _EVAL_143;
  wire [3:0] _EVAL_177;
  wire  _EVAL_145;
  wire  _EVAL_210;
  wire [14:0] _EVAL_131;
  wire [15:0] _EVAL_25;
  wire [15:0] _EVAL_189;
  wire [15:0] _EVAL_259;
  wire  _EVAL_179;
  wire  _EVAL_58;
  wire  _EVAL_104;
  wire  _EVAL_186;
  wire  _EVAL_212;
  wire [12:0] _EVAL_148;
  wire [5:0] _EVAL_16;
  wire [5:0] _EVAL_182;
  wire [3:0] _EVAL_147;
  wire [3:0] _EVAL_226;
  wire  _EVAL_150;
  wire  _EVAL_32;
  wire  _EVAL_91;
  wire [3:0] _EVAL_100;
  wire  _EVAL_217;
  wire  _EVAL_136;
  wire  _EVAL_286;
  wire  _EVAL_260;
  wire  _EVAL_244;
  wire  _EVAL_133;
  wire  _EVAL_114;
  wire  _EVAL_197;
  wire  _EVAL_64;
  wire  _EVAL_59;
  wire  _EVAL_194;
  wire  _EVAL_141;
  wire  _EVAL_94;
  wire  _EVAL_227;
  wire  _EVAL_144;
  wire [2:0] _EVAL_19;
  wire  _EVAL_122;
  wire  _EVAL_192;
  wire  _EVAL_196;
  wire  _EVAL_253;
  wire  _EVAL_49;
  wire  _EVAL_128;
  wire  _EVAL_288;
  wire  _EVAL_79;
  wire  _EVAL_201;
  wire  _EVAL_23;
  wire  _EVAL_218;
  wire  _EVAL_109;
  wire  _EVAL_171;
  wire  _EVAL_52;
  wire  _EVAL_61;
  wire  _EVAL_67;
  wire  _EVAL_106;
  wire  _EVAL_168;
  wire  _EVAL_280;
  wire  _EVAL_239;
  wire  _EVAL_44;
  wire  _EVAL_246;
  wire  _EVAL_215;
  wire  _EVAL_236;
  wire  _EVAL_211;
  wire  _EVAL_151;
  wire  _EVAL_178;
  wire  _EVAL_281;
  wire  _EVAL_169;
  wire  _EVAL_156;
  wire  _EVAL_73;
  wire  _EVAL_283;
  wire  _EVAL_243;
  wire  _EVAL_205;
  wire  _EVAL_103;
  wire  _EVAL_54;
  wire  _EVAL_132;
  wire  _EVAL_99;
  wire  _EVAL_126;
  wire  _EVAL_166;
  wire  _EVAL_238;
  wire  _EVAL_18;
  wire  _EVAL_85;
  wire  _EVAL_188;
  wire  _EVAL_55;
  wire  _EVAL_60;
  wire  _EVAL_237;
  wire  _EVAL_29;
  wire  _EVAL_249;
  wire  _EVAL_123;
  wire  _EVAL_46;
  wire  _EVAL_241;
  wire  _EVAL_93;
  wire  _EVAL_213;
  wire  _EVAL_47;
  wire  _EVAL_187;
  wire  _EVAL_247;
  wire  _EVAL_174;
  wire  _EVAL_235;
  wire  _EVAL_37;
  wire  _EVAL_271;
  wire [72:0] _EVAL_224;
  wire [72:0] _EVAL_202;
  wire  _EVAL_27;
  wire  _EVAL_57;
  wire  _EVAL_198;
  wire  _EVAL_248;
  wire  _EVAL_250;
  wire  _EVAL_17;
  wire  _EVAL_101;
  wire  _EVAL_36;
  wire  _EVAL_107;
  wire  _EVAL_86;
  wire  _EVAL_232;
  wire  _EVAL_21;
  wire  _EVAL_116;
  wire  _EVAL_264;
  wire  _EVAL_88;
  wire  _EVAL_62;
  wire  _EVAL_255;
  wire  _EVAL_111;
  wire  _EVAL_82;
  wire  _EVAL_105;
  wire  _EVAL_270;
  wire  _EVAL_71;
  wire  _EVAL_159;
  wire  _EVAL_285;
  wire  _EVAL_56;
  wire  _EVAL_181;
  wire  _EVAL_207;
  wire  _EVAL_230;
  wire  _EVAL_185;
  wire  _EVAL_225;
  wire  _EVAL_28;
  wire  _EVAL_124;
  wire  _EVAL_172;
  wire  _EVAL_119;
  wire  _EVAL_108;
  wire  _EVAL_206;
  wire  _EVAL_76;
  wire  _EVAL_117;
  wire  _EVAL_96;
  wire  _EVAL_157;
  wire  _EVAL_87;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_39 = 13'h3f << _EVAL_13;
  assign _EVAL_233 = _EVAL_39[5:0];
  assign _EVAL_175 = ~ _EVAL_233;
  assign _EVAL_22 = {{9'd0}, _EVAL_175};
  assign _EVAL_276 = _EVAL_8 & _EVAL_22;
  assign _EVAL_282 = _EVAL_276 == 15'h0;
  assign _EVAL_92 = _EVAL == _EVAL_278;
  assign _EVAL_195 = _EVAL_92 | _EVAL_5;
  assign _EVAL_183 = _EVAL_195 == 1'h0;
  assign _EVAL_41 = _EVAL_4 == 3'h2;
  assign _EVAL_135 = _EVAL_7 & _EVAL_41;
  assign _EVAL_48 = _EVAL >= 3'h2;
  assign _EVAL_221 = _EVAL_0 == 7'h48;
  assign _EVAL_75 = _EVAL_0 == 7'h40;
  assign _EVAL_265 = _EVAL_221 | _EVAL_75;
  assign _EVAL_43 = _EVAL_0[6:3];
  assign _EVAL_146 = _EVAL_43 == 4'h8;
  assign _EVAL_68 = _EVAL_0[2:0];
  assign _EVAL_24 = 3'h1 <= _EVAL_68;
  assign _EVAL_180 = _EVAL_146 & _EVAL_24;
  assign _EVAL_269 = _EVAL_265 | _EVAL_180;
  assign _EVAL_263 = _EVAL_0 == 7'h20;
  assign _EVAL_193 = _EVAL_269 | _EVAL_263;
  assign _EVAL_279 = _EVAL_191 - 4'h1;
  assign _EVAL_216 = _EVAL_13 >= 3'h2;
  assign _EVAL_262 = _EVAL_13[0];
  assign _EVAL_80 = 2'h1 << _EVAL_262;
  assign _EVAL_203 = _EVAL_80 | 2'h1;
  assign _EVAL_72 = _EVAL_203[1];
  assign _EVAL_272 = _EVAL_8[1];
  assign _EVAL_242 = _EVAL_72 & _EVAL_272;
  assign _EVAL_34 = _EVAL_216 | _EVAL_242;
  assign _EVAL_81 = _EVAL_2 <= 3'h2;
  assign _EVAL_170 = _EVAL_81 | _EVAL_5;
  assign _EVAL_125 = _EVAL_10 & _EVAL_7;
  assign _EVAL_209 = _EVAL_129 == 4'h0;
  assign _EVAL_53 = _EVAL_125 & _EVAL_209;
  assign _EVAL_266 = 128'h1 << _EVAL_0;
  assign _EVAL_160 = _EVAL_53 ? _EVAL_266 : 128'h0;
  assign _EVAL_95 = _EVAL_160[72:0];
  assign _EVAL_245 = _EVAL_11 & _EVAL_6;
  assign _EVAL_229 = _EVAL_191 == 4'h0;
  assign _EVAL_204 = _EVAL_245 & _EVAL_229;
  assign _EVAL_267 = _EVAL_12 == 3'h6;
  assign _EVAL_164 = _EVAL_267 == 1'h0;
  assign _EVAL_90 = _EVAL_204 & _EVAL_164;
  assign _EVAL_220 = 128'h1 << _EVAL_14;
  assign _EVAL_287 = _EVAL_90 ? _EVAL_220 : 128'h0;
  assign _EVAL_89 = _EVAL_287[72:0];
  assign _EVAL_154 = _EVAL_95 != _EVAL_89;
  assign _EVAL_118 = _EVAL_95 != 73'h0;
  assign _EVAL_35 = _EVAL_118 == 1'h0;
  assign _EVAL_222 = _EVAL_154 | _EVAL_35;
  assign _EVAL_162 = _EVAL_222 | _EVAL_5;
  assign _EVAL_138 = _EVAL_175[5:2];
  assign _EVAL_261 = _EVAL_115 == 4'h0;
  assign _EVAL_70 = _EVAL_184 >> _EVAL_0;
  assign _EVAL_113 = _EVAL_70[0];
  assign _EVAL_254 = _EVAL_113 == 1'h0;
  assign _EVAL_134 = _EVAL_95 | _EVAL_184;
  assign _EVAL_33 = _EVAL_134 >> _EVAL_14;
  assign _EVAL_130 = _EVAL_33[0];
  assign _EVAL_274 = _EVAL_130 | _EVAL_5;
  assign _EVAL_219 = _EVAL_274 == 1'h0;
  assign _EVAL_112 = _EVAL_12 == _EVAL_140;
  assign _EVAL_199 = _EVAL_12[0];
  assign _EVAL_51 = _EVAL_8[0];
  assign _EVAL_163 = _EVAL_51 == 1'h0;
  assign _EVAL_165 = _EVAL_272 & _EVAL_163;
  assign _EVAL_214 = _EVAL_2 <= 3'h3;
  assign _EVAL_65 = _EVAL_203[0];
  assign _EVAL_240 = _EVAL_272 == 1'h0;
  assign _EVAL_63 = _EVAL_240 & _EVAL_163;
  assign _EVAL_42 = _EVAL_65 & _EVAL_63;
  assign _EVAL_234 = _EVAL_14[6:3];
  assign _EVAL_121 = _EVAL_234 == 4'h0;
  assign _EVAL_173 = _EVAL_184 | _EVAL_95;
  assign _EVAL_252 = _EVAL_4[2];
  assign _EVAL_38 = _EVAL_252 == 1'h0;
  assign _EVAL_110 = _EVAL_115 - 4'h1;
  assign _EVAL_258 = _EVAL_272 & _EVAL_51;
  assign _EVAL_176 = _EVAL_216 | _EVAL_5;
  assign _EVAL_74 = _EVAL_12 == 3'h1;
  assign _EVAL_84 = _EVAL_6 & _EVAL_74;
  assign _EVAL_102 = _EVAL_4 == 3'h3;
  assign _EVAL_78 = _EVAL_65 & _EVAL_258;
  assign _EVAL_257 = _EVAL_34 | _EVAL_78;
  assign _EVAL_26 = _EVAL_65 & _EVAL_165;
  assign _EVAL_277 = _EVAL_34 | _EVAL_26;
  assign _EVAL_127 = _EVAL_72 & _EVAL_240;
  assign _EVAL_69 = _EVAL_216 | _EVAL_127;
  assign _EVAL_120 = _EVAL_240 & _EVAL_51;
  assign _EVAL_155 = _EVAL_65 & _EVAL_120;
  assign _EVAL_167 = _EVAL_69 | _EVAL_155;
  assign _EVAL_223 = _EVAL_69 | _EVAL_42;
  assign _EVAL_31 = {_EVAL_257,_EVAL_277,_EVAL_167,_EVAL_223};
  assign _EVAL_142 = ~ _EVAL_31;
  assign _EVAL_228 = _EVAL_9 & _EVAL_142;
  assign _EVAL_30 = _EVAL_228 == 4'h0;
  assign _EVAL_15 = _EVAL_282 | _EVAL_5;
  assign _EVAL_190 = _EVAL_112 | _EVAL_5;
  assign _EVAL_97 = _EVAL_190 == 1'h0;
  assign _EVAL_143 = _EVAL_208 + 32'h1;
  assign _EVAL_177 = ~ _EVAL_9;
  assign _EVAL_145 = _EVAL_4 == 3'h5;
  assign _EVAL_210 = _EVAL_13 <= 3'h6;
  assign _EVAL_131 = _EVAL_8 ^ 15'h4000;
  assign _EVAL_25 = {1'b0,$signed(_EVAL_131)};
  assign _EVAL_189 = $signed(_EVAL_25) & $signed(-16'sh1000);
  assign _EVAL_259 = $signed(_EVAL_189);
  assign _EVAL_179 = $signed(_EVAL_259) == $signed(16'sh0);
  assign _EVAL_58 = _EVAL_210 & _EVAL_179;
  assign _EVAL_104 = _EVAL_58 | _EVAL_5;
  assign _EVAL_186 = _EVAL_104 == 1'h0;
  assign _EVAL_212 = _EVAL_200 == 4'h0;
  assign _EVAL_148 = 13'h3f << _EVAL;
  assign _EVAL_16 = _EVAL_148[5:0];
  assign _EVAL_182 = ~ _EVAL_16;
  assign _EVAL_147 = _EVAL_182[5:2];
  assign _EVAL_226 = _EVAL_200 - 4'h1;
  assign _EVAL_150 = _EVAL_245 & _EVAL_212;
  assign _EVAL_32 = _EVAL_43 == 4'h3;
  assign _EVAL_91 = _EVAL_13 == _EVAL_83;
  assign _EVAL_100 = _EVAL_129 - 4'h1;
  assign _EVAL_217 = _EVAL_212 == 1'h0;
  assign _EVAL_136 = _EVAL_12 == 3'h5;
  assign _EVAL_286 = _EVAL_8 == _EVAL_284;
  assign _EVAL_260 = _EVAL_286 | _EVAL_5;
  assign _EVAL_244 = _EVAL_260 == 1'h0;
  assign _EVAL_133 = _EVAL_0 == _EVAL_152;
  assign _EVAL_114 = _EVAL_133 | _EVAL_5;
  assign _EVAL_197 = _EVAL_91 | _EVAL_5;
  assign _EVAL_64 = _EVAL_2 <= 3'h4;
  assign _EVAL_59 = _EVAL_64 | _EVAL_5;
  assign _EVAL_194 = _EVAL_59 == 1'h0;
  assign _EVAL_141 = _EVAL_14 == 7'h48;
  assign _EVAL_94 = _EVAL_14 == 7'h40;
  assign _EVAL_227 = _EVAL_141 | _EVAL_94;
  assign _EVAL_144 = _EVAL_234 == 4'h8;
  assign _EVAL_19 = _EVAL_14[2:0];
  assign _EVAL_122 = 3'h1 <= _EVAL_19;
  assign _EVAL_192 = _EVAL_144 & _EVAL_122;
  assign _EVAL_196 = _EVAL_227 | _EVAL_192;
  assign _EVAL_253 = _EVAL_2 == 3'h0;
  assign _EVAL_49 = _EVAL_253 | _EVAL_5;
  assign _EVAL_128 = _EVAL_49 == 1'h0;
  assign _EVAL_288 = _EVAL_176 == 1'h0;
  assign _EVAL_79 = _EVAL_14 == 7'h20;
  assign _EVAL_201 = _EVAL_196 | _EVAL_79;
  assign _EVAL_23 = _EVAL_201 | _EVAL_121;
  assign _EVAL_218 = _EVAL_234 == 4'h1;
  assign _EVAL_109 = _EVAL_23 | _EVAL_218;
  assign _EVAL_171 = _EVAL_254 | _EVAL_5;
  assign _EVAL_52 = _EVAL_9 == _EVAL_31;
  assign _EVAL_61 = _EVAL_52 | _EVAL_5;
  assign _EVAL_67 = _EVAL_4 == 3'h4;
  assign _EVAL_106 = _EVAL_4 == 3'h7;
  assign _EVAL_168 = _EVAL_7 & _EVAL_106;
  assign _EVAL_280 = _EVAL_197 == 1'h0;
  assign _EVAL_239 = _EVAL_2 == _EVAL_149;
  assign _EVAL_44 = _EVAL_239 | _EVAL_5;
  assign _EVAL_246 = _EVAL_162 == 1'h0;
  assign _EVAL_215 = 3'h6 == _EVAL_13;
  assign _EVAL_236 = _EVAL_75 ? _EVAL_215 : 1'h0;
  assign _EVAL_211 = _EVAL_236 | _EVAL_5;
  assign _EVAL_151 = _EVAL_211 == 1'h0;
  assign _EVAL_178 = _EVAL_234 == 4'h2;
  assign _EVAL_281 = _EVAL_43 == 4'h0;
  assign _EVAL_169 = _EVAL_193 | _EVAL_281;
  assign _EVAL_156 = _EVAL_43 == 4'h1;
  assign _EVAL_73 = _EVAL_169 | _EVAL_156;
  assign _EVAL_283 = _EVAL_43 == 4'h2;
  assign _EVAL_243 = _EVAL_73 | _EVAL_283;
  assign _EVAL_205 = _EVAL_243 | _EVAL_32;
  assign _EVAL_103 = _EVAL_205 | _EVAL_5;
  assign _EVAL_54 = _EVAL_6 & _EVAL_136;
  assign _EVAL_132 = _EVAL_6 & _EVAL_267;
  assign _EVAL_99 = _EVAL_1 == 1'h0;
  assign _EVAL_126 = _EVAL_99 | _EVAL_5;
  assign _EVAL_166 = _EVAL_126 == 1'h0;
  assign _EVAL_238 = _EVAL_214 | _EVAL_5;
  assign _EVAL_18 = _EVAL_4 == 3'h6;
  assign _EVAL_85 = _EVAL_7 & _EVAL_18;
  assign _EVAL_188 = plusarg_reader_out == 32'h0;
  assign _EVAL_55 = _EVAL_114 == 1'h0;
  assign _EVAL_60 = _EVAL_61 == 1'h0;
  assign _EVAL_237 = _EVAL_7 & _EVAL_102;
  assign _EVAL_29 = _EVAL_170 == 1'h0;
  assign _EVAL_249 = _EVAL_238 == 1'h0;
  assign _EVAL_123 = _EVAL_14 == _EVAL_161;
  assign _EVAL_46 = _EVAL_123 | _EVAL_5;
  assign _EVAL_241 = _EVAL_109 | _EVAL_178;
  assign _EVAL_93 = _EVAL_234 == 4'h3;
  assign _EVAL_213 = _EVAL_241 | _EVAL_93;
  assign _EVAL_47 = _EVAL_213 | _EVAL_5;
  assign _EVAL_187 = _EVAL_47 == 1'h0;
  assign _EVAL_247 = _EVAL_12 == 3'h4;
  assign _EVAL_174 = _EVAL_48 | _EVAL_5;
  assign _EVAL_235 = _EVAL_12 == 3'h2;
  assign _EVAL_37 = _EVAL_6 & _EVAL_235;
  assign _EVAL_271 = _EVAL_30 | _EVAL_5;
  assign _EVAL_224 = ~ _EVAL_89;
  assign _EVAL_202 = _EVAL_173 & _EVAL_224;
  assign _EVAL_27 = _EVAL_208 < plusarg_reader_out;
  assign _EVAL_57 = _EVAL_184 != 73'h0;
  assign _EVAL_198 = _EVAL_12 <= 3'h6;
  assign _EVAL_248 = _EVAL_198 | _EVAL_5;
  assign _EVAL_250 = _EVAL_46 == 1'h0;
  assign _EVAL_17 = _EVAL_261 == 1'h0;
  assign _EVAL_101 = _EVAL_7 & _EVAL_17;
  assign _EVAL_36 = _EVAL_4 == _EVAL_153;
  assign _EVAL_107 = _EVAL_248 == 1'h0;
  assign _EVAL_86 = _EVAL_174 == 1'h0;
  assign _EVAL_232 = _EVAL_125 | _EVAL_245;
  assign _EVAL_21 = _EVAL_4 == 3'h1;
  assign _EVAL_116 = _EVAL_7 & _EVAL_21;
  assign _EVAL_264 = _EVAL_57 == 1'h0;
  assign _EVAL_88 = _EVAL_264 | _EVAL_188;
  assign _EVAL_62 = _EVAL_7 & _EVAL_67;
  assign _EVAL_255 = _EVAL_36 | _EVAL_5;
  assign _EVAL_111 = _EVAL_255 == 1'h0;
  assign _EVAL_82 = _EVAL_6 & _EVAL_247;
  assign _EVAL_105 = _EVAL_88 | _EVAL_27;
  assign _EVAL_270 = _EVAL_105 | _EVAL_5;
  assign _EVAL_71 = _EVAL_270 == 1'h0;
  assign _EVAL_159 = _EVAL_12 == 3'h0;
  assign _EVAL_285 = _EVAL_6 & _EVAL_159;
  assign _EVAL_56 = _EVAL_7 & _EVAL_145;
  assign _EVAL_181 = _EVAL_171 == 1'h0;
  assign _EVAL_207 = _EVAL_271 == 1'h0;
  assign _EVAL_230 = _EVAL_4 == 3'h0;
  assign _EVAL_185 = _EVAL_7 & _EVAL_230;
  assign _EVAL_225 = _EVAL_177 == 4'h0;
  assign _EVAL_28 = _EVAL_225 | _EVAL_5;
  assign _EVAL_124 = _EVAL_28 == 1'h0;
  assign _EVAL_172 = _EVAL_6 & _EVAL_217;
  assign _EVAL_119 = _EVAL_103 == 1'h0;
  assign _EVAL_108 = _EVAL_2 != 3'h0;
  assign _EVAL_206 = _EVAL_5 == 1'h0;
  assign _EVAL_76 = _EVAL_125 & _EVAL_261;
  assign _EVAL_117 = _EVAL_108 | _EVAL_5;
  assign _EVAL_96 = _EVAL_117 == 1'h0;
  assign _EVAL_157 = _EVAL_15 == 1'h0;
  assign _EVAL_87 = _EVAL_44 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_83 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_115 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_129 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_140 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_149 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_152 = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_153 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_161 = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {3{`RANDOM}};
  _EVAL_184 = _RAND_8[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_191 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_200 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_208 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_278 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_284 = _RAND_13[14:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_76) begin
      _EVAL_83 <= _EVAL_13;
    end
    if (_EVAL_5) begin
      _EVAL_115 <= 4'h0;
    end else begin
      if (_EVAL_125) begin
        if (_EVAL_261) begin
          if (_EVAL_38) begin
            _EVAL_115 <= _EVAL_138;
          end else begin
            _EVAL_115 <= 4'h0;
          end
        end else begin
          _EVAL_115 <= _EVAL_110;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_129 <= 4'h0;
    end else begin
      if (_EVAL_125) begin
        if (_EVAL_209) begin
          if (_EVAL_38) begin
            _EVAL_129 <= _EVAL_138;
          end else begin
            _EVAL_129 <= 4'h0;
          end
        end else begin
          _EVAL_129 <= _EVAL_100;
        end
      end
    end
    if (_EVAL_150) begin
      _EVAL_140 <= _EVAL_12;
    end
    if (_EVAL_76) begin
      _EVAL_149 <= _EVAL_2;
    end
    if (_EVAL_76) begin
      _EVAL_152 <= _EVAL_0;
    end
    if (_EVAL_76) begin
      _EVAL_153 <= _EVAL_4;
    end
    if (_EVAL_150) begin
      _EVAL_161 <= _EVAL_14;
    end
    if (_EVAL_5) begin
      _EVAL_184 <= 73'h0;
    end else begin
      _EVAL_184 <= _EVAL_202;
    end
    if (_EVAL_5) begin
      _EVAL_191 <= 4'h0;
    end else begin
      if (_EVAL_245) begin
        if (_EVAL_229) begin
          if (_EVAL_199) begin
            _EVAL_191 <= _EVAL_147;
          end else begin
            _EVAL_191 <= 4'h0;
          end
        end else begin
          _EVAL_191 <= _EVAL_279;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_200 <= 4'h0;
    end else begin
      if (_EVAL_245) begin
        if (_EVAL_212) begin
          if (_EVAL_199) begin
            _EVAL_200 <= _EVAL_147;
          end else begin
            _EVAL_200 <= 4'h0;
          end
        end else begin
          _EVAL_200 <= _EVAL_226;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_208 <= 32'h0;
    end else begin
      if (_EVAL_232) begin
        _EVAL_208 <= 32'h0;
      end else begin
        _EVAL_208 <= _EVAL_143;
      end
    end
    if (_EVAL_150) begin
      _EVAL_278 <= _EVAL;
    end
    if (_EVAL_76) begin
      _EVAL_284 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4027df3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(771c47ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f9020d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3eea788c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4679263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b130778)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afc073f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93fd1d94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b262002)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db11c694)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98c1bc6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32df592a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e526e688)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f015a34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48448815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d9abc4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a47ea0f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1adbf90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9701da2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f2bb20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d782445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3df62d0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c634cdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d96683ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbf655f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(939ea251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd157be9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3835074)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfdcf6e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb3fb31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64f83a64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfc42334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46d81049)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81159400)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c431fe0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86317108)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57659896)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a36e304d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfe5f439)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8c0ea15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36b4b7a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63518571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(859d8bbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b687fe2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6512125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb04b185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54d0f4f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ef3387)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c98f142a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99c2f937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7492210)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(688fbb0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4812e572)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae068806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acd5ef42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b0e1763)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5076db74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55099fb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7ed5525)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a07f93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f99d7797)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226296df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c458325)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4100419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ead844c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a908d7de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7659973)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2da8e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc92ae82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1af40618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6faa3a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d11ecc47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
