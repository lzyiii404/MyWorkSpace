//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_1_assert(
  input  [5:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [5:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [7:0]  _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [1:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_19;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_56;
  reg [31:0] _RAND_1;
  reg [4:0] _EVAL_65;
  reg [31:0] _RAND_2;
  reg [4:0] _EVAL_86;
  reg [31:0] _RAND_3;
  reg [5:0] _EVAL_108;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_119;
  reg [31:0] _RAND_5;
  reg  _EVAL_131;
  reg [31:0] _RAND_6;
  reg [32:0] _EVAL_136;
  reg [63:0] _RAND_7;
  reg [4:0] _EVAL_159;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_201;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_221;
  reg [31:0] _RAND_10;
  reg  _EVAL_225;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_241;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_310;
  reg [31:0] _RAND_13;
  reg [31:0] _EVAL_311;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_335;
  reg [31:0] _RAND_15;
  reg [4:0] _EVAL_370;
  reg [31:0] _RAND_16;
  wire [31:0] _EVAL_44;
  wire [32:0] _EVAL_350;
  wire  _EVAL_338;
  wire  _EVAL_328;
  wire [31:0] _EVAL_27;
  wire  _EVAL_285;
  wire  _EVAL_191;
  wire  _EVAL_317;
  wire  _EVAL_170;
  wire  _EVAL_61;
  wire  _EVAL_381;
  wire [2:0] _EVAL_222;
  wire  _EVAL_176;
  wire [1:0] _EVAL_261;
  wire [3:0] _EVAL_24;
  wire [2:0] _EVAL_239;
  wire [2:0] _EVAL_278;
  wire  _EVAL_28;
  wire  _EVAL_122;
  wire  _EVAL_72;
  wire  _EVAL_265;
  wire  _EVAL_172;
  wire  _EVAL_229;
  wire  _EVAL_187;
  wire  _EVAL_20;
  wire  _EVAL_321;
  wire  _EVAL_192;
  wire [63:0] _EVAL_341;
  wire [63:0] _EVAL_237;
  wire [32:0] _EVAL_208;
  wire [32:0] _EVAL_312;
  wire  _EVAL_35;
  wire [32:0] _EVAL_257;
  wire [32:0] _EVAL_134;
  wire  _EVAL_142;
  wire  _EVAL_264;
  wire  _EVAL_304;
  wire  _EVAL_135;
  wire  _EVAL_147;
  wire  _EVAL_333;
  wire  _EVAL_141;
  wire  _EVAL_322;
  wire  _EVAL_305;
  wire  _EVAL_160;
  wire  _EVAL_34;
  wire  _EVAL_352;
  wire  _EVAL_71;
  wire  _EVAL_23;
  wire [31:0] _EVAL_167;
  wire [32:0] _EVAL_79;
  wire [32:0] _EVAL_244;
  wire  _EVAL_291;
  wire [2:0] _EVAL_375;
  wire  _EVAL_342;
  wire  _EVAL_383;
  wire  _EVAL_26;
  wire  _EVAL_288;
  wire  _EVAL_190;
  wire  _EVAL_168;
  wire  _EVAL_110;
  wire  _EVAL_88;
  wire  _EVAL_374;
  wire  _EVAL_41;
  wire  _EVAL_174;
  wire  _EVAL_292;
  wire  _EVAL_140;
  wire  _EVAL_157;
  wire  _EVAL_224;
  wire  _EVAL_175;
  wire  _EVAL_143;
  wire  _EVAL_206;
  wire  _EVAL_145;
  wire  _EVAL_346;
  wire  _EVAL_217;
  wire  _EVAL_242;
  wire  _EVAL_76;
  wire  _EVAL_369;
  wire  _EVAL_318;
  wire  _EVAL_234;
  wire  _EVAL_207;
  wire  _EVAL_194;
  wire  _EVAL_280;
  wire  _EVAL_371;
  wire  _EVAL_180;
  wire  _EVAL_380;
  wire  _EVAL_126;
  wire  _EVAL_334;
  wire  _EVAL_254;
  wire  _EVAL_215;
  wire  _EVAL_327;
  wire  _EVAL_232;
  wire  _EVAL_247;
  wire  _EVAL_59;
  wire  _EVAL_296;
  wire  _EVAL_343;
  wire [7:0] _EVAL_273;
  wire  _EVAL_227;
  wire [32:0] _EVAL_315;
  wire [31:0] _EVAL_358;
  wire [32:0] _EVAL_51;
  wire [32:0] _EVAL_40;
  wire [32:0] _EVAL_63;
  wire  _EVAL_281;
  wire  _EVAL_91;
  wire  _EVAL_382;
  wire  _EVAL_138;
  wire  _EVAL_385;
  wire  _EVAL_129;
  wire  _EVAL_103;
  wire  _EVAL_316;
  wire [22:0] _EVAL_29;
  wire [7:0] _EVAL_284;
  wire [7:0] _EVAL_260;
  wire [4:0] _EVAL_218;
  wire  _EVAL_228;
  wire [31:0] _EVAL_363;
  wire [32:0] _EVAL_246;
  wire [32:0] _EVAL_256;
  wire [32:0] _EVAL_213;
  wire  _EVAL_367;
  wire [31:0] _EVAL_22;
  wire [32:0] _EVAL_301;
  wire [32:0] _EVAL_85;
  wire [32:0] _EVAL_57;
  wire  _EVAL_161;
  wire  _EVAL_379;
  wire  _EVAL_101;
  wire [31:0] _EVAL_70;
  wire [32:0] _EVAL_47;
  wire [32:0] _EVAL_100;
  wire [32:0] _EVAL_104;
  wire  _EVAL_289;
  wire  _EVAL_282;
  wire [32:0] _EVAL_255;
  wire [32:0] _EVAL_287;
  wire [32:0] _EVAL_33;
  wire  _EVAL_73;
  wire  _EVAL_362;
  wire [31:0] _EVAL_355;
  wire [32:0] _EVAL_214;
  wire [32:0] _EVAL_162;
  wire [32:0] _EVAL_200;
  wire  _EVAL_107;
  wire  _EVAL_36;
  wire [32:0] _EVAL_96;
  wire  _EVAL_196;
  wire  _EVAL_74;
  wire [31:0] _EVAL_53;
  wire [32:0] _EVAL_181;
  wire [32:0] _EVAL_357;
  wire [32:0] _EVAL_306;
  wire  _EVAL_275;
  wire  _EVAL_67;
  wire  _EVAL_25;
  wire  _EVAL_184;
  wire [32:0] _EVAL_339;
  wire  _EVAL_307;
  wire  _EVAL_290;
  wire  _EVAL_111;
  wire  _EVAL_249;
  wire  _EVAL_378;
  wire  _EVAL_392;
  wire  _EVAL_178;
  wire  _EVAL_156;
  wire  _EVAL_64;
  wire  _EVAL_236;
  wire  _EVAL_48;
  wire  _EVAL_263;
  wire  _EVAL_98;
  wire  _EVAL_114;
  wire  _EVAL_347;
  wire  _EVAL_389;
  wire  _EVAL_164;
  wire [63:0] _EVAL_197;
  wire [63:0] _EVAL_69;
  wire [32:0] _EVAL_186;
  wire [32:0] _EVAL_148;
  wire [32:0] _EVAL_80;
  wire  _EVAL_340;
  wire  _EVAL_146;
  wire  _EVAL_368;
  wire  _EVAL_268;
  wire  _EVAL_31;
  wire  _EVAL_144;
  wire  _EVAL_349;
  wire  _EVAL_271;
  wire  _EVAL_293;
  wire  _EVAL_299;
  wire  _EVAL_121;
  wire  _EVAL_95;
  wire  _EVAL_251;
  wire  _EVAL_120;
  wire  _EVAL_203;
  wire  _EVAL_154;
  wire [7:0] _EVAL_177;
  wire  _EVAL_253;
  wire  _EVAL_43;
  wire  _EVAL_39;
  wire  _EVAL_297;
  wire  _EVAL_105;
  wire  _EVAL_169;
  wire  _EVAL_331;
  wire [22:0] _EVAL_165;
  wire [7:0] _EVAL_279;
  wire [7:0] _EVAL_388;
  wire [4:0] _EVAL_84;
  wire  _EVAL_81;
  wire  _EVAL_118;
  wire  _EVAL_283;
  wire  _EVAL_151;
  wire [31:0] _EVAL_83;
  wire [31:0] _EVAL_276;
  wire  _EVAL_252;
  wire  _EVAL_300;
  wire [4:0] _EVAL_269;
  wire  _EVAL_376;
  wire  _EVAL_124;
  wire  _EVAL_152;
  wire [4:0] _EVAL_198;
  wire  _EVAL_308;
  wire  _EVAL_223;
  wire  _EVAL_245;
  wire  _EVAL_231;
  wire  _EVAL_37;
  wire  _EVAL_226;
  wire  _EVAL_330;
  wire  _EVAL_66;
  wire  _EVAL_361;
  wire  _EVAL_259;
  wire  _EVAL_195;
  wire  _EVAL_220;
  wire  _EVAL_391;
  wire  _EVAL_302;
  wire  _EVAL_99;
  wire  _EVAL_326;
  wire  _EVAL_212;
  wire  _EVAL_45;
  wire  _EVAL_117;
  wire  _EVAL_360;
  wire  _EVAL_32;
  wire  _EVAL_202;
  wire  _EVAL_386;
  wire  _EVAL_364;
  wire  _EVAL_272;
  wire  _EVAL_387;
  wire  _EVAL_130;
  wire  _EVAL_235;
  wire  _EVAL_113;
  wire  _EVAL_78;
  wire  _EVAL_87;
  wire  _EVAL_62;
  wire  _EVAL_97;
  wire  _EVAL_323;
  wire  _EVAL_128;
  wire  _EVAL_204;
  wire [4:0] _EVAL_356;
  wire  _EVAL_270;
  wire  _EVAL_90;
  wire  _EVAL_351;
  wire  _EVAL_294;
  wire  _EVAL_345;
  wire  _EVAL_193;
  wire  _EVAL_52;
  wire  _EVAL_153;
  wire  _EVAL_365;
  wire  _EVAL_106;
  wire  _EVAL_188;
  wire [32:0] _EVAL_377;
  wire  _EVAL_205;
  wire  _EVAL_182;
  wire  _EVAL_267;
  wire  _EVAL_274;
  wire  _EVAL_354;
  wire  _EVAL_337;
  wire  _EVAL_262;
  wire  _EVAL_199;
  wire  _EVAL_277;
  wire  _EVAL_94;
  wire  _EVAL_173;
  wire  _EVAL_238;
  wire  _EVAL_233;
  wire  _EVAL_133;
  wire  _EVAL_77;
  wire  _EVAL_139;
  wire  _EVAL_258;
  wire  _EVAL_166;
  wire  _EVAL_54;
  wire  _EVAL_38;
  wire  _EVAL_295;
  wire  _EVAL_210;
  wire  _EVAL_42;
  wire  _EVAL_309;
  wire [7:0] _EVAL_68;
  wire [7:0] _EVAL_344;
  wire  _EVAL_149;
  wire  _EVAL_93;
  wire  _EVAL_336;
  wire  _EVAL_183;
  wire  _EVAL_216;
  wire  _EVAL_313;
  wire  _EVAL_60;
  wire  _EVAL_373;
  wire  _EVAL_266;
  wire  _EVAL_189;
  wire  _EVAL_132;
  wire  _EVAL_329;
  wire  _EVAL_155;
  wire  _EVAL_58;
  wire  _EVAL_348;
  wire  _EVAL_179;
  wire [4:0] _EVAL_390;
  wire  _EVAL_303;
  wire  _EVAL_137;
  wire  _EVAL_158;
  wire  _EVAL_49;
  wire  _EVAL_102;
  wire  _EVAL_123;
  wire  _EVAL_209;
  wire  _EVAL_366;
  wire  _EVAL_286;
  wire  _EVAL_116;
  wire  _EVAL_112;
  wire  _EVAL_314;
  wire  _EVAL_75;
  wire  _EVAL_250;
  wire  _EVAL_115;
  wire  _EVAL_243;
  wire  _EVAL_219;
  wire  _EVAL_372;
  wire  _EVAL_125;
  wire  _EVAL_324;
  wire  _EVAL_163;
  wire  _EVAL_127;
  wire  _EVAL_230;
  wire  _EVAL_89;
  wire  _EVAL_46;
  wire  _EVAL_320;
  wire  _EVAL_55;
  wire  _EVAL_211;
  wire  _EVAL_21;
  wire  _EVAL_240;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_44 = _EVAL_17 ^ 32'h1900000;
  assign _EVAL_350 = {1'b0,$signed(_EVAL_44)};
  assign _EVAL_338 = _EVAL_7 >= 4'h3;
  assign _EVAL_328 = _EVAL_338 | _EVAL_4;
  assign _EVAL_27 = _EVAL_56 + 32'h1;
  assign _EVAL_285 = _EVAL_1 == _EVAL_221;
  assign _EVAL_191 = _EVAL_3 == 3'h0;
  assign _EVAL_317 = _EVAL_3 == _EVAL_335;
  assign _EVAL_170 = _EVAL_2 == _EVAL_201;
  assign _EVAL_61 = _EVAL_170 | _EVAL_4;
  assign _EVAL_381 = _EVAL_61 == 1'h0;
  assign _EVAL_222 = _EVAL_2[5:3];
  assign _EVAL_176 = _EVAL_222 == 3'h0;
  assign _EVAL_261 = _EVAL_7[1:0];
  assign _EVAL_24 = 4'h1 << _EVAL_261;
  assign _EVAL_239 = _EVAL_24[2:0];
  assign _EVAL_278 = _EVAL_239 | 3'h1;
  assign _EVAL_28 = _EVAL_278[1];
  assign _EVAL_122 = _EVAL_17[2];
  assign _EVAL_72 = _EVAL_122 == 1'h0;
  assign _EVAL_265 = _EVAL_17[1];
  assign _EVAL_172 = _EVAL_265 == 1'h0;
  assign _EVAL_229 = _EVAL_72 & _EVAL_172;
  assign _EVAL_187 = _EVAL_28 & _EVAL_229;
  assign _EVAL_20 = _EVAL_12 & _EVAL_14;
  assign _EVAL_321 = _EVAL_159 == 5'h0;
  assign _EVAL_192 = _EVAL_20 & _EVAL_321;
  assign _EVAL_341 = 64'h1 << _EVAL;
  assign _EVAL_237 = _EVAL_192 ? _EVAL_341 : 64'h0;
  assign _EVAL_208 = _EVAL_237[32:0];
  assign _EVAL_312 = _EVAL_136 | _EVAL_208;
  assign _EVAL_35 = _EVAL_0 & _EVAL_191;
  assign _EVAL_257 = _EVAL_208 | _EVAL_136;
  assign _EVAL_134 = _EVAL_257 >> _EVAL_2;
  assign _EVAL_142 = _EVAL_134[0];
  assign _EVAL_264 = _EVAL_142 | _EVAL_4;
  assign _EVAL_304 = _EVAL_264 == 1'h0;
  assign _EVAL_135 = _EVAL_278[2];
  assign _EVAL_147 = _EVAL_135 & _EVAL_72;
  assign _EVAL_333 = _EVAL_338 | _EVAL_147;
  assign _EVAL_141 = _EVAL_72 & _EVAL_265;
  assign _EVAL_322 = _EVAL_28 & _EVAL_141;
  assign _EVAL_305 = _EVAL_333 | _EVAL_322;
  assign _EVAL_160 = _EVAL_278[0];
  assign _EVAL_34 = _EVAL_17[0];
  assign _EVAL_352 = _EVAL_141 & _EVAL_34;
  assign _EVAL_71 = _EVAL_160 & _EVAL_352;
  assign _EVAL_23 = _EVAL_305 | _EVAL_71;
  assign _EVAL_167 = _EVAL_17 ^ 32'h3000;
  assign _EVAL_79 = {1'b0,$signed(_EVAL_167)};
  assign _EVAL_244 = $signed(_EVAL_79) & $signed(-33'sh1000);
  assign _EVAL_291 = _EVAL == 6'h20;
  assign _EVAL_375 = _EVAL[5:3];
  assign _EVAL_342 = _EVAL_375 == 3'h0;
  assign _EVAL_383 = _EVAL_291 | _EVAL_342;
  assign _EVAL_26 = _EVAL_375 == 3'h1;
  assign _EVAL_288 = _EVAL_383 | _EVAL_26;
  assign _EVAL_190 = _EVAL_375 == 3'h2;
  assign _EVAL_168 = _EVAL_288 | _EVAL_190;
  assign _EVAL_110 = _EVAL_375 == 3'h3;
  assign _EVAL_88 = _EVAL_168 | _EVAL_110;
  assign _EVAL_374 = _EVAL_88 | _EVAL_4;
  assign _EVAL_41 = _EVAL_374 == 1'h0;
  assign _EVAL_174 = _EVAL_136 != 33'h0;
  assign _EVAL_292 = _EVAL_135 & _EVAL_122;
  assign _EVAL_140 = _EVAL_338 | _EVAL_292;
  assign _EVAL_157 = _EVAL_122 & _EVAL_265;
  assign _EVAL_224 = _EVAL_28 & _EVAL_157;
  assign _EVAL_175 = _EVAL_140 | _EVAL_224;
  assign _EVAL_143 = _EVAL_157 & _EVAL_34;
  assign _EVAL_206 = _EVAL_160 & _EVAL_143;
  assign _EVAL_145 = _EVAL_175 | _EVAL_206;
  assign _EVAL_346 = _EVAL_34 == 1'h0;
  assign _EVAL_217 = _EVAL_157 & _EVAL_346;
  assign _EVAL_242 = _EVAL_160 & _EVAL_217;
  assign _EVAL_76 = _EVAL_175 | _EVAL_242;
  assign _EVAL_369 = _EVAL_122 & _EVAL_172;
  assign _EVAL_318 = _EVAL_28 & _EVAL_369;
  assign _EVAL_234 = _EVAL_140 | _EVAL_318;
  assign _EVAL_207 = _EVAL_369 & _EVAL_34;
  assign _EVAL_194 = _EVAL_160 & _EVAL_207;
  assign _EVAL_280 = _EVAL_234 | _EVAL_194;
  assign _EVAL_371 = _EVAL_369 & _EVAL_346;
  assign _EVAL_180 = _EVAL_160 & _EVAL_371;
  assign _EVAL_380 = _EVAL_234 | _EVAL_180;
  assign _EVAL_126 = _EVAL_141 & _EVAL_346;
  assign _EVAL_334 = _EVAL_160 & _EVAL_126;
  assign _EVAL_254 = _EVAL_305 | _EVAL_334;
  assign _EVAL_215 = _EVAL_333 | _EVAL_187;
  assign _EVAL_327 = _EVAL_229 & _EVAL_34;
  assign _EVAL_232 = _EVAL_160 & _EVAL_327;
  assign _EVAL_247 = _EVAL_215 | _EVAL_232;
  assign _EVAL_59 = _EVAL_229 & _EVAL_346;
  assign _EVAL_296 = _EVAL_160 & _EVAL_59;
  assign _EVAL_343 = _EVAL_215 | _EVAL_296;
  assign _EVAL_273 = {_EVAL_145,_EVAL_76,_EVAL_280,_EVAL_380,_EVAL_23,_EVAL_254,_EVAL_247,_EVAL_343};
  assign _EVAL_227 = _EVAL_1 == 3'h3;
  assign _EVAL_315 = $signed(_EVAL_350) & $signed(-33'sh2000);
  assign _EVAL_358 = _EVAL_17 ^ 32'hc000000;
  assign _EVAL_51 = {1'b0,$signed(_EVAL_358)};
  assign _EVAL_40 = $signed(_EVAL_51) & $signed(-33'sh4000000);
  assign _EVAL_63 = $signed(_EVAL_40);
  assign _EVAL_281 = $signed(_EVAL_63) == $signed(33'sh0);
  assign _EVAL_91 = _EVAL_15 <= 3'h3;
  assign _EVAL_382 = _EVAL_91 | _EVAL_4;
  assign _EVAL_138 = _EVAL_382 == 1'h0;
  assign _EVAL_385 = _EVAL_6 == 1'h0;
  assign _EVAL_129 = _EVAL_3 <= 3'h6;
  assign _EVAL_103 = _EVAL_129 | _EVAL_4;
  assign _EVAL_316 = _EVAL_103 == 1'h0;
  assign _EVAL_29 = 23'hff << _EVAL_18;
  assign _EVAL_284 = _EVAL_29[7:0];
  assign _EVAL_260 = ~ _EVAL_284;
  assign _EVAL_218 = _EVAL_260[7:3];
  assign _EVAL_228 = _EVAL_7 <= 4'h6;
  assign _EVAL_363 = _EVAL_17 ^ 32'h40000000;
  assign _EVAL_246 = {1'b0,$signed(_EVAL_363)};
  assign _EVAL_256 = $signed(_EVAL_246) & $signed(-33'sh2000);
  assign _EVAL_213 = $signed(_EVAL_256);
  assign _EVAL_367 = $signed(_EVAL_213) == $signed(33'sh0);
  assign _EVAL_22 = _EVAL_17 ^ 32'h80000000;
  assign _EVAL_301 = {1'b0,$signed(_EVAL_22)};
  assign _EVAL_85 = $signed(_EVAL_301) & $signed(-33'sh20000);
  assign _EVAL_57 = $signed(_EVAL_85);
  assign _EVAL_161 = $signed(_EVAL_57) == $signed(33'sh0);
  assign _EVAL_379 = _EVAL_367 | _EVAL_161;
  assign _EVAL_101 = _EVAL_379 | _EVAL_281;
  assign _EVAL_70 = _EVAL_17 ^ 32'h2000000;
  assign _EVAL_47 = {1'b0,$signed(_EVAL_70)};
  assign _EVAL_100 = $signed(_EVAL_47) & $signed(-33'sh10000);
  assign _EVAL_104 = $signed(_EVAL_100);
  assign _EVAL_289 = $signed(_EVAL_104) == $signed(33'sh0);
  assign _EVAL_282 = _EVAL_101 | _EVAL_289;
  assign _EVAL_255 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_287 = $signed(_EVAL_255) & $signed(-33'sh5000);
  assign _EVAL_33 = $signed(_EVAL_287);
  assign _EVAL_73 = $signed(_EVAL_33) == $signed(33'sh0);
  assign _EVAL_362 = _EVAL_282 | _EVAL_73;
  assign _EVAL_355 = _EVAL_17 ^ 32'h1800000;
  assign _EVAL_214 = {1'b0,$signed(_EVAL_355)};
  assign _EVAL_162 = $signed(_EVAL_214) & $signed(-33'sh8000);
  assign _EVAL_200 = $signed(_EVAL_162);
  assign _EVAL_107 = $signed(_EVAL_200) == $signed(33'sh0);
  assign _EVAL_36 = _EVAL_362 | _EVAL_107;
  assign _EVAL_96 = $signed(_EVAL_315);
  assign _EVAL_196 = $signed(_EVAL_96) == $signed(33'sh0);
  assign _EVAL_74 = _EVAL_36 | _EVAL_196;
  assign _EVAL_53 = _EVAL_17 ^ 32'h20000000;
  assign _EVAL_181 = {1'b0,$signed(_EVAL_53)};
  assign _EVAL_357 = $signed(_EVAL_181) & $signed(-33'sh2000);
  assign _EVAL_306 = $signed(_EVAL_357);
  assign _EVAL_275 = $signed(_EVAL_306) == $signed(33'sh0);
  assign _EVAL_67 = _EVAL_74 | _EVAL_275;
  assign _EVAL_25 = _EVAL_228 & _EVAL_67;
  assign _EVAL_184 = _EVAL_7 <= 4'h8;
  assign _EVAL_339 = $signed(_EVAL_244);
  assign _EVAL_307 = $signed(_EVAL_339) == $signed(33'sh0);
  assign _EVAL_290 = _EVAL_184 & _EVAL_307;
  assign _EVAL_111 = _EVAL_25 | _EVAL_290;
  assign _EVAL_249 = _EVAL_111 | _EVAL_4;
  assign _EVAL_378 = _EVAL_249 == 1'h0;
  assign _EVAL_392 = _EVAL_228 & _EVAL_161;
  assign _EVAL_178 = _EVAL_392 | _EVAL_4;
  assign _EVAL_156 = _EVAL_178 == 1'h0;
  assign _EVAL_64 = _EVAL_385 | _EVAL_11;
  assign _EVAL_236 = _EVAL_64 | _EVAL_4;
  assign _EVAL_48 = _EVAL_236 == 1'h0;
  assign _EVAL_263 = _EVAL_5 & _EVAL_0;
  assign _EVAL_98 = _EVAL_370 == 5'h0;
  assign _EVAL_114 = _EVAL_263 & _EVAL_98;
  assign _EVAL_347 = _EVAL_3 == 3'h6;
  assign _EVAL_389 = _EVAL_347 == 1'h0;
  assign _EVAL_164 = _EVAL_114 & _EVAL_389;
  assign _EVAL_197 = 64'h1 << _EVAL_2;
  assign _EVAL_69 = _EVAL_164 ? _EVAL_197 : 64'h0;
  assign _EVAL_186 = _EVAL_69[32:0];
  assign _EVAL_148 = ~ _EVAL_186;
  assign _EVAL_80 = _EVAL_312 & _EVAL_148;
  assign _EVAL_340 = _EVAL_15 != 3'h0;
  assign _EVAL_146 = _EVAL_11 == 1'h0;
  assign _EVAL_368 = _EVAL_385 | _EVAL_4;
  assign _EVAL_268 = _EVAL_18 == _EVAL_19;
  assign _EVAL_31 = _EVAL_317 | _EVAL_4;
  assign _EVAL_144 = _EVAL_31 == 1'h0;
  assign _EVAL_349 = _EVAL_17 == _EVAL_311;
  assign _EVAL_271 = _EVAL_9 == _EVAL_131;
  assign _EVAL_293 = _EVAL_271 | _EVAL_4;
  assign _EVAL_299 = _EVAL_293 == 1'h0;
  assign _EVAL_121 = _EVAL_174 == 1'h0;
  assign _EVAL_95 = plusarg_reader_out == 32'h0;
  assign _EVAL_251 = _EVAL_121 | _EVAL_95;
  assign _EVAL_120 = _EVAL_56 < plusarg_reader_out;
  assign _EVAL_203 = _EVAL_251 | _EVAL_120;
  assign _EVAL_154 = _EVAL_203 | _EVAL_4;
  assign _EVAL_177 = ~ _EVAL_13;
  assign _EVAL_253 = _EVAL_177 == 8'h0;
  assign _EVAL_43 = _EVAL_253 | _EVAL_4;
  assign _EVAL_39 = _EVAL_43 == 1'h0;
  assign _EVAL_297 = _EVAL_222 == 3'h1;
  assign _EVAL_105 = _EVAL_1 == 3'h6;
  assign _EVAL_169 = _EVAL_14 & _EVAL_105;
  assign _EVAL_331 = _EVAL_3 == 3'h4;
  assign _EVAL_165 = 23'hff << _EVAL_7;
  assign _EVAL_279 = _EVAL_165[7:0];
  assign _EVAL_388 = ~ _EVAL_279;
  assign _EVAL_84 = _EVAL_388[7:3];
  assign _EVAL_81 = _EVAL_15 == _EVAL_241;
  assign _EVAL_118 = _EVAL_81 | _EVAL_4;
  assign _EVAL_283 = _EVAL_3[0];
  assign _EVAL_151 = _EVAL_1 == 3'h7;
  assign _EVAL_83 = {{24'd0}, _EVAL_388};
  assign _EVAL_276 = _EVAL_17 & _EVAL_83;
  assign _EVAL_252 = _EVAL_276 == 32'h0;
  assign _EVAL_300 = _EVAL_86 == 5'h0;
  assign _EVAL_269 = _EVAL_86 - 5'h1;
  assign _EVAL_376 = _EVAL_6 == _EVAL_225;
  assign _EVAL_124 = _EVAL_1[2];
  assign _EVAL_152 = _EVAL_124 == 1'h0;
  assign _EVAL_198 = _EVAL_159 - 5'h1;
  assign _EVAL_308 = _EVAL_376 | _EVAL_4;
  assign _EVAL_223 = _EVAL_2 == 6'h20;
  assign _EVAL_245 = _EVAL_223 | _EVAL_176;
  assign _EVAL_231 = _EVAL_245 | _EVAL_297;
  assign _EVAL_37 = _EVAL_222 == 3'h2;
  assign _EVAL_226 = _EVAL_231 | _EVAL_37;
  assign _EVAL_330 = _EVAL_7 <= 4'h2;
  assign _EVAL_66 = _EVAL_307 | _EVAL_281;
  assign _EVAL_361 = _EVAL_66 | _EVAL_289;
  assign _EVAL_259 = _EVAL_361 | _EVAL_73;
  assign _EVAL_195 = _EVAL_259 | _EVAL_107;
  assign _EVAL_220 = _EVAL_195 | _EVAL_196;
  assign _EVAL_391 = _EVAL_220 | _EVAL_275;
  assign _EVAL_302 = _EVAL_330 & _EVAL_391;
  assign _EVAL_99 = _EVAL_302 | _EVAL_4;
  assign _EVAL_326 = _EVAL_252 | _EVAL_4;
  assign _EVAL_212 = _EVAL_349 | _EVAL_4;
  assign _EVAL_45 = _EVAL_212 == 1'h0;
  assign _EVAL_117 = _EVAL_300 == 1'h0;
  assign _EVAL_360 = _EVAL_0 & _EVAL_117;
  assign _EVAL_32 = _EVAL == _EVAL_108;
  assign _EVAL_202 = _EVAL_208 != 33'h0;
  assign _EVAL_386 = _EVAL_1 == 3'h0;
  assign _EVAL_364 = _EVAL_7 == _EVAL_119;
  assign _EVAL_272 = _EVAL_364 | _EVAL_4;
  assign _EVAL_387 = _EVAL_15 == 3'h0;
  assign _EVAL_130 = _EVAL_14 & _EVAL_227;
  assign _EVAL_235 = _EVAL_13 == _EVAL_273;
  assign _EVAL_113 = _EVAL_235 | _EVAL_4;
  assign _EVAL_78 = _EVAL_113 == 1'h0;
  assign _EVAL_87 = _EVAL_154 == 1'h0;
  assign _EVAL_62 = _EVAL_3 == 3'h5;
  assign _EVAL_97 = _EVAL_146 | _EVAL_4;
  assign _EVAL_323 = _EVAL_97 == 1'h0;
  assign _EVAL_128 = _EVAL_16 == 2'h0;
  assign _EVAL_204 = _EVAL_128 | _EVAL_4;
  assign _EVAL_356 = _EVAL_370 - 5'h1;
  assign _EVAL_270 = _EVAL_32 | _EVAL_4;
  assign _EVAL_90 = _EVAL_16 <= 2'h2;
  assign _EVAL_351 = _EVAL_340 | _EVAL_4;
  assign _EVAL_294 = _EVAL_351 == 1'h0;
  assign _EVAL_345 = _EVAL_0 & _EVAL_331;
  assign _EVAL_193 = _EVAL_15 <= 3'h4;
  assign _EVAL_52 = _EVAL_193 | _EVAL_4;
  assign _EVAL_153 = _EVAL_52 == 1'h0;
  assign _EVAL_365 = _EVAL_1 == 3'h1;
  assign _EVAL_106 = _EVAL_118 == 1'h0;
  assign _EVAL_188 = _EVAL_15 <= 3'h2;
  assign _EVAL_377 = _EVAL_136 >> _EVAL;
  assign _EVAL_205 = _EVAL_377[0];
  assign _EVAL_182 = _EVAL_205 == 1'h0;
  assign _EVAL_267 = _EVAL_182 | _EVAL_4;
  assign _EVAL_274 = _EVAL_308 == 1'h0;
  assign _EVAL_354 = _EVAL_18 >= 4'h3;
  assign _EVAL_337 = _EVAL_354 | _EVAL_4;
  assign _EVAL_262 = _EVAL_8 == 1'h0;
  assign _EVAL_199 = _EVAL_3 == 3'h1;
  assign _EVAL_277 = _EVAL_1 == 3'h4;
  assign _EVAL_94 = _EVAL_285 | _EVAL_4;
  assign _EVAL_173 = _EVAL_208 != _EVAL_186;
  assign _EVAL_238 = _EVAL_202 == 1'h0;
  assign _EVAL_233 = _EVAL_173 | _EVAL_238;
  assign _EVAL_133 = _EVAL_233 | _EVAL_4;
  assign _EVAL_77 = _EVAL_133 == 1'h0;
  assign _EVAL_139 = _EVAL_387 | _EVAL_4;
  assign _EVAL_258 = _EVAL_139 == 1'h0;
  assign _EVAL_166 = _EVAL_272 == 1'h0;
  assign _EVAL_54 = _EVAL_65 == 5'h0;
  assign _EVAL_38 = _EVAL_54 == 1'h0;
  assign _EVAL_295 = _EVAL_16 != 2'h2;
  assign _EVAL_210 = _EVAL_295 | _EVAL_4;
  assign _EVAL_42 = _EVAL_94 == 1'h0;
  assign _EVAL_309 = _EVAL_0 & _EVAL_62;
  assign _EVAL_68 = ~ _EVAL_273;
  assign _EVAL_344 = _EVAL_13 & _EVAL_68;
  assign _EVAL_149 = _EVAL_337 == 1'h0;
  assign _EVAL_93 = _EVAL_222 == 3'h3;
  assign _EVAL_336 = _EVAL_226 | _EVAL_93;
  assign _EVAL_183 = _EVAL_14 & _EVAL_38;
  assign _EVAL_216 = _EVAL_0 & _EVAL_199;
  assign _EVAL_313 = _EVAL_344 == 8'h0;
  assign _EVAL_60 = _EVAL_90 | _EVAL_4;
  assign _EVAL_373 = _EVAL_368 == 1'h0;
  assign _EVAL_266 = _EVAL_20 & _EVAL_54;
  assign _EVAL_189 = _EVAL_270 == 1'h0;
  assign _EVAL_132 = _EVAL_0 & _EVAL_347;
  assign _EVAL_329 = _EVAL_188 | _EVAL_4;
  assign _EVAL_155 = _EVAL_99 == 1'h0;
  assign _EVAL_58 = _EVAL_328 == 1'h0;
  assign _EVAL_348 = _EVAL_3 == 3'h2;
  assign _EVAL_179 = _EVAL_0 & _EVAL_348;
  assign _EVAL_390 = _EVAL_65 - 5'h1;
  assign _EVAL_303 = _EVAL_1 == 3'h2;
  assign _EVAL_137 = _EVAL_14 & _EVAL_303;
  assign _EVAL_158 = _EVAL_4 == 1'h0;
  assign _EVAL_49 = _EVAL_313 | _EVAL_4;
  assign _EVAL_102 = _EVAL_204 == 1'h0;
  assign _EVAL_123 = _EVAL_268 | _EVAL_4;
  assign _EVAL_209 = _EVAL_123 == 1'h0;
  assign _EVAL_366 = _EVAL_336 | _EVAL_4;
  assign _EVAL_286 = _EVAL_366 == 1'h0;
  assign _EVAL_116 = _EVAL_14 & _EVAL_365;
  assign _EVAL_112 = _EVAL_20 | _EVAL_263;
  assign _EVAL_314 = _EVAL_290 | _EVAL_4;
  assign _EVAL_75 = _EVAL_326 == 1'h0;
  assign _EVAL_250 = _EVAL_267 == 1'h0;
  assign _EVAL_115 = _EVAL_329 == 1'h0;
  assign _EVAL_243 = _EVAL_16 == _EVAL_310;
  assign _EVAL_219 = _EVAL_243 | _EVAL_4;
  assign _EVAL_372 = _EVAL_262 | _EVAL_4;
  assign _EVAL_125 = _EVAL_1 == 3'h5;
  assign _EVAL_324 = _EVAL_14 & _EVAL_125;
  assign _EVAL_163 = _EVAL_14 & _EVAL_151;
  assign _EVAL_127 = _EVAL_263 & _EVAL_300;
  assign _EVAL_230 = _EVAL_14 & _EVAL_386;
  assign _EVAL_89 = _EVAL_314 == 1'h0;
  assign _EVAL_46 = _EVAL_60 == 1'h0;
  assign _EVAL_320 = _EVAL_14 & _EVAL_277;
  assign _EVAL_55 = _EVAL_219 == 1'h0;
  assign _EVAL_211 = _EVAL_210 == 1'h0;
  assign _EVAL_21 = _EVAL_49 == 1'h0;
  assign _EVAL_240 = _EVAL_372 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_19 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_56 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_65 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_86 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_108 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_119 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_131 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _EVAL_136 = _RAND_7[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_159 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_201 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_221 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_225 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_241 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_310 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_311 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_335 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_370 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_10) begin
    if (_EVAL_127) begin
      _EVAL_19 <= _EVAL_18;
    end
    if (_EVAL_4) begin
      _EVAL_56 <= 32'h0;
    end else begin
      if (_EVAL_112) begin
        _EVAL_56 <= 32'h0;
      end else begin
        _EVAL_56 <= _EVAL_27;
      end
    end
    if (_EVAL_4) begin
      _EVAL_65 <= 5'h0;
    end else begin
      if (_EVAL_20) begin
        if (_EVAL_54) begin
          if (_EVAL_152) begin
            _EVAL_65 <= _EVAL_84;
          end else begin
            _EVAL_65 <= 5'h0;
          end
        end else begin
          _EVAL_65 <= _EVAL_390;
        end
      end
    end
    if (_EVAL_4) begin
      _EVAL_86 <= 5'h0;
    end else begin
      if (_EVAL_263) begin
        if (_EVAL_300) begin
          if (_EVAL_283) begin
            _EVAL_86 <= _EVAL_218;
          end else begin
            _EVAL_86 <= 5'h0;
          end
        end else begin
          _EVAL_86 <= _EVAL_269;
        end
      end
    end
    if (_EVAL_266) begin
      _EVAL_108 <= _EVAL;
    end
    if (_EVAL_266) begin
      _EVAL_119 <= _EVAL_7;
    end
    if (_EVAL_127) begin
      _EVAL_131 <= _EVAL_9;
    end
    if (_EVAL_4) begin
      _EVAL_136 <= 33'h0;
    end else begin
      _EVAL_136 <= _EVAL_80;
    end
    if (_EVAL_4) begin
      _EVAL_159 <= 5'h0;
    end else begin
      if (_EVAL_20) begin
        if (_EVAL_321) begin
          if (_EVAL_152) begin
            _EVAL_159 <= _EVAL_84;
          end else begin
            _EVAL_159 <= 5'h0;
          end
        end else begin
          _EVAL_159 <= _EVAL_198;
        end
      end
    end
    if (_EVAL_127) begin
      _EVAL_201 <= _EVAL_2;
    end
    if (_EVAL_266) begin
      _EVAL_221 <= _EVAL_1;
    end
    if (_EVAL_127) begin
      _EVAL_225 <= _EVAL_6;
    end
    if (_EVAL_266) begin
      _EVAL_241 <= _EVAL_15;
    end
    if (_EVAL_127) begin
      _EVAL_310 <= _EVAL_16;
    end
    if (_EVAL_266) begin
      _EVAL_311 <= _EVAL_17;
    end
    if (_EVAL_127) begin
      _EVAL_335 <= _EVAL_3;
    end
    if (_EVAL_4) begin
      _EVAL_370 <= 5'h0;
    end else begin
      if (_EVAL_263) begin
        if (_EVAL_98) begin
          if (_EVAL_283) begin
            _EVAL_370 <= _EVAL_218;
          end else begin
            _EVAL_370 <= 5'h0;
          end
        end else begin
          _EVAL_370 <= _EVAL_356;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68b25e53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e7ddd17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73a91688)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85cd7a97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5c18702)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(688dc0eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c69b076)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c310c99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(419b2a65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0b44ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(622cd2f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dacddda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed0d6bc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4108c1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ec0a32a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e8ea312)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad07c15b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(577c73ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c64f57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33d501a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e34af18f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fe5b7a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0582d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f5926fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b49de310)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb769034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b994c250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a32aa384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db0bfc20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7ec3103)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fdc622a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(562bace3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ab990b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_373) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(790ee0e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d01872d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49d9e4ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43bd5bb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8086acbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf57e81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b58db2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0ffc1aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(444cb54a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d138bcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53142e10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9da2117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7da8618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cffd54c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(121f3237)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4ba40ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9a5c0b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_381) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee62f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f9a4b6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78583369)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_373) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0a1c6c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a424b0c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf98f33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1148063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db93af4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa746c2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca49e7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea388ff1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ae1777)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60b6bf51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd1dac85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b84859e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e3a0bb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66c2b345)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4657efe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20fca5e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67373b09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(766e5c97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1b1d3d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dac28db3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce3bf98a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e596e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7526b6b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1011f292)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e17152f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80be1468)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0152d3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dd3ec89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39ca995e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1625bcf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d863aada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6094b18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(242e8249)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e90deac9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a88e044a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_381) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
