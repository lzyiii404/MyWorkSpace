//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_232(
  output  _EVAL,
  output  _EVAL_0,
  output  _EVAL_1,
  output  _EVAL_2,
  output  _EVAL_3,
  output  _EVAL_4,
  output  _EVAL_5,
  output  _EVAL_6,
  output  _EVAL_7,
  output  _EVAL_8,
  input   _EVAL_9,
  output  _EVAL_10,
  output  _EVAL_11,
  output  _EVAL_12,
  input   _EVAL_13,
  output  _EVAL_14,
  input   _EVAL_15,
  output  _EVAL_16,
  output  _EVAL_17
);
  reg  _EVAL_18;
  reg [31:0] _RAND_0;
  reg  _EVAL_19;
  reg [31:0] _RAND_1;
  reg  _EVAL_20;
  reg [31:0] _RAND_2;
  reg  _EVAL_21;
  reg [31:0] _RAND_3;
  reg  _EVAL_22;
  reg [31:0] _RAND_4;
  reg  _EVAL_23;
  reg [31:0] _RAND_5;
  reg  _EVAL_26;
  reg [31:0] _RAND_6;
  reg  _EVAL_31;
  reg [31:0] _RAND_7;
  reg  _EVAL_33;
  reg [31:0] _RAND_8;
  reg  _EVAL_36;
  reg [31:0] _RAND_9;
  reg  _EVAL_39;
  reg [31:0] _RAND_10;
  reg  _EVAL_40;
  reg [31:0] _RAND_11;
  reg  _EVAL_42;
  reg [31:0] _RAND_12;
  reg  _EVAL_48;
  reg [31:0] _RAND_13;
  reg  _EVAL_50;
  reg [31:0] _RAND_14;
  reg  _EVAL_51;
  reg [31:0] _RAND_15;
  wire  _EVAL_52;
  wire  _EVAL_41;
  wire  _EVAL_34;
  assign _EVAL_52 = _EVAL_50 ^ _EVAL_19;
  assign _EVAL_41 = _EVAL_52 ^ _EVAL_39;
  assign _EVAL_34 = _EVAL_41 ^ _EVAL_23;
  assign _EVAL = _EVAL_39;
  assign _EVAL_2 = _EVAL_31;
  assign _EVAL_17 = _EVAL_36;
  assign _EVAL_8 = _EVAL_40;
  assign _EVAL_6 = _EVAL_51;
  assign _EVAL_12 = _EVAL_42;
  assign _EVAL_10 = _EVAL_26;
  assign _EVAL_14 = _EVAL_48;
  assign _EVAL_1 = _EVAL_19;
  assign _EVAL_5 = _EVAL_20;
  assign _EVAL_16 = _EVAL_21;
  assign _EVAL_4 = _EVAL_23;
  assign _EVAL_11 = _EVAL_18;
  assign _EVAL_3 = _EVAL_22;
  assign _EVAL_0 = _EVAL_50;
  assign _EVAL_7 = _EVAL_33;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_18 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_19 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_20 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_21 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_22 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_23 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_26 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_31 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_33 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_36 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_39 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_40 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_42 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_48 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_50 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_51 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_15) begin
    if (_EVAL_13) begin
      _EVAL_18 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_18 <= _EVAL_22;
      end
    end
    if (_EVAL_13) begin
      _EVAL_19 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_19 <= _EVAL_39;
      end
    end
    if (_EVAL_13) begin
      _EVAL_20 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_20 <= _EVAL_23;
      end
    end
    if (_EVAL_13) begin
      _EVAL_21 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_21 <= _EVAL_40;
      end
    end
    if (_EVAL_13) begin
      _EVAL_22 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_22 <= _EVAL_21;
      end
    end
    if (_EVAL_13) begin
      _EVAL_23 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_23 <= _EVAL_51;
      end
    end
    if (_EVAL_13) begin
      _EVAL_26 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_26 <= _EVAL_48;
      end
    end
    if (_EVAL_13) begin
      _EVAL_31 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_31 <= _EVAL_42;
      end
    end
    if (_EVAL_13) begin
      _EVAL_33 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_33 <= _EVAL_34;
      end
    end
    if (_EVAL_13) begin
      _EVAL_36 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_36 <= _EVAL_19;
      end
    end
    if (_EVAL_13) begin
      _EVAL_39 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_39 <= _EVAL_20;
      end
    end
    if (_EVAL_13) begin
      _EVAL_40 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_40 <= _EVAL_26;
      end
    end
    if (_EVAL_13) begin
      _EVAL_42 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_42 <= _EVAL_18;
      end
    end
    if (_EVAL_13) begin
      _EVAL_48 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_48 <= _EVAL_33;
      end
    end
    if (_EVAL_13) begin
      _EVAL_50 <= 1'h1;
    end else begin
      if (_EVAL_9) begin
        _EVAL_50 <= _EVAL_36;
      end
    end
    if (_EVAL_13) begin
      _EVAL_51 <= 1'h0;
    end else begin
      if (_EVAL_9) begin
        _EVAL_51 <= _EVAL_31;
      end
    end
  end
endmodule
