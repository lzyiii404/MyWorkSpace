//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL(
  input   _EVAL,
  output  _EVAL_0,
  input   _EVAL_1,
  input   _EVAL_2,
  input   _EVAL_3,
  input   _EVAL_4,
  input   _EVAL_5,
  output  _EVAL_6,
  input   _EVAL_7,
  input   _EVAL_8,
  input   _EVAL_9,
  output  _EVAL_10,
  input   _EVAL_11,
  output  _EVAL_12,
  input   _EVAL_13,
  input   _EVAL_14,
  output  _EVAL_15,
  output  _EVAL_16,
  input   _EVAL_17,
  input   _EVAL_18,
  input   _EVAL_19,
  input   _EVAL_20,
  input   _EVAL_21,
  output  _EVAL_22,
  input   _EVAL_23,
  input   _EVAL_24,
  input   _EVAL_25,
  output  _EVAL_26,
  input   _EVAL_27,
  input   _EVAL_28,
  input   _EVAL_29,
  input   _EVAL_30,
  output  _EVAL_31,
  output  _EVAL_32,
  input   _EVAL_33,
  output  _EVAL_34,
  output  _EVAL_35,
  input   _EVAL_36,
  input   _EVAL_37,
  output  _EVAL_38,
  output  _EVAL_39,
  input   _EVAL_40,
  input   _EVAL_41,
  input   _EVAL_42,
  input   _EVAL_43,
  output  _EVAL_44,
  output  _EVAL_45,
  output  _EVAL_46,
  output  _EVAL_47,
  input   _EVAL_48,
  input   _EVAL_49,
  input   _EVAL_50,
  output  _EVAL_51,
  input   _EVAL_52,
  input   _EVAL_53,
  input   _EVAL_54,
  input   _EVAL_55,
  input   _EVAL_56,
  output  _EVAL_57,
  output  _EVAL_58,
  output  _EVAL_59,
  input   _EVAL_60,
  input   _EVAL_61,
  input   _EVAL_62,
  output  _EVAL_63,
  input   _EVAL_64,
  input   _EVAL_65,
  output  _EVAL_66,
  input   _EVAL_67,
  input   _EVAL_68,
  input   _EVAL_69,
  input   _EVAL_70,
  output  _EVAL_71,
  input   _EVAL_72,
  input   _EVAL_73,
  output  _EVAL_74,
  output  _EVAL_75,
  output  _EVAL_76,
  input   _EVAL_77,
  output  _EVAL_78,
  input   _EVAL_79,
  output  _EVAL_80,
  input   _EVAL_81,
  input   _EVAL_82,
  input   _EVAL_83,
  output  _EVAL_84,
  output  _EVAL_85,
  output  _EVAL_86,
  output  _EVAL_87,
  output  _EVAL_88,
  input   _EVAL_89,
  output  _EVAL_90,
  output  _EVAL_91,
  input   _EVAL_92,
  output  _EVAL_93,
  output  _EVAL_94,
  input   _EVAL_95,
  input   _EVAL_96,
  output  _EVAL_97,
  input   _EVAL_98,
  output  _EVAL_99,
  input   _EVAL_100,
  input   _EVAL_101,
  output  _EVAL_102,
  input   _EVAL_103,
  output  _EVAL_104,
  input   _EVAL_105,
  output  _EVAL_106,
  output  _EVAL_107,
  output  _EVAL_108,
  output  _EVAL_109,
  input   _EVAL_110,
  output  _EVAL_111,
  output  _EVAL_112,
  output  _EVAL_113,
  input   _EVAL_114,
  output  _EVAL_115,
  input   _EVAL_116,
  input   _EVAL_117,
  output  _EVAL_118,
  output  _EVAL_119,
  input   _EVAL_120,
  input   _EVAL_121,
  input   _EVAL_122,
  input   _EVAL_123,
  input   _EVAL_124,
  output  _EVAL_125,
  output  _EVAL_126,
  output  _EVAL_127,
  output  _EVAL_128,
  output  _EVAL_129,
  input   _EVAL_130,
  input   _EVAL_131,
  input   _EVAL_132,
  output  _EVAL_133,
  input   _EVAL_134,
  output  _EVAL_135,
  input   _EVAL_136,
  output  _EVAL_137,
  output  _EVAL_138,
  input   _EVAL_139,
  output  _EVAL_140,
  output  _EVAL_141,
  input   _EVAL_142,
  output  _EVAL_143,
  output  _EVAL_144,
  output  _EVAL_145,
  input   _EVAL_146,
  output  _EVAL_147,
  output  _EVAL_148,
  input   _EVAL_149,
  output  _EVAL_150,
  output  _EVAL_151,
  output  _EVAL_152,
  input   _EVAL_153,
  output  _EVAL_154,
  output  _EVAL_155,
  output  _EVAL_156,
  output  _EVAL_157,
  input   _EVAL_158,
  output  _EVAL_159,
  output  _EVAL_160,
  input   _EVAL_161,
  input   _EVAL_162,
  input   _EVAL_163,
  output  _EVAL_164,
  output  _EVAL_165,
  input   _EVAL_166,
  output  _EVAL_167,
  input   _EVAL_168,
  output  _EVAL_169,
  output  _EVAL_170,
  input   _EVAL_171,
  output  _EVAL_172,
  input   _EVAL_173,
  output  _EVAL_174,
  input   _EVAL_175,
  output  _EVAL_176,
  output  _EVAL_177,
  input   _EVAL_178,
  output  _EVAL_179,
  output  _EVAL_180,
  output  _EVAL_181,
  input   _EVAL_182,
  output  _EVAL_183,
  input   _EVAL_184,
  output  _EVAL_185,
  output  _EVAL_186,
  output  _EVAL_187,
  output  _EVAL_188,
  input   _EVAL_189,
  output  _EVAL_190,
  output  _EVAL_191,
  output  _EVAL_192,
  input   _EVAL_193,
  input   _EVAL_194,
  output  _EVAL_195,
  output  _EVAL_196,
  input   _EVAL_197,
  output  _EVAL_198,
  input   _EVAL_199,
  output  _EVAL_200,
  output  _EVAL_201,
  output  _EVAL_202,
  output  _EVAL_203,
  input   _EVAL_204,
  input   _EVAL_205,
  output  _EVAL_206,
  input   _EVAL_207,
  output  _EVAL_208,
  input   _EVAL_209,
  input   _EVAL_210,
  input   _EVAL_211,
  input   _EVAL_212,
  output  _EVAL_213,
  input   _EVAL_214,
  input   _EVAL_215,
  input   _EVAL_216,
  input   _EVAL_217,
  output  _EVAL_218,
  output  _EVAL_219,
  output  _EVAL_220,
  input   _EVAL_221,
  input   _EVAL_222,
  output  _EVAL_223,
  output  _EVAL_224,
  input   _EVAL_225,
  input   _EVAL_226,
  input   _EVAL_227,
  input   _EVAL_228,
  input   _EVAL_229,
  output  _EVAL_230,
  output  _EVAL_231,
  output  _EVAL_232,
  input   _EVAL_233,
  output  _EVAL_234,
  input   _EVAL_235,
  output  _EVAL_236,
  output  _EVAL_237,
  input   _EVAL_238,
  output  _EVAL_239,
  output  _EVAL_240,
  output  _EVAL_241,
  output  _EVAL_242,
  output  _EVAL_243,
  input   _EVAL_244,
  input   _EVAL_245,
  input   _EVAL_246,
  output  _EVAL_247,
  input   _EVAL_248,
  output  _EVAL_249,
  input   _EVAL_250,
  input   _EVAL_251,
  output  _EVAL_252
);
  assign _EVAL_141 = _EVAL_62;
  assign _EVAL_58 = _EVAL_5;
  assign _EVAL_22 = _EVAL_101;
  assign _EVAL_12 = _EVAL_211;
  assign _EVAL_113 = _EVAL_229;
  assign _EVAL_118 = _EVAL_123;
  assign _EVAL_180 = _EVAL_4;
  assign _EVAL_94 = _EVAL_42;
  assign _EVAL_247 = _EVAL_146;
  assign _EVAL_39 = _EVAL_64;
  assign _EVAL_181 = _EVAL_184;
  assign _EVAL_150 = _EVAL_134;
  assign _EVAL_172 = _EVAL_228;
  assign _EVAL_97 = _EVAL_121;
  assign _EVAL_170 = _EVAL_20;
  assign _EVAL_16 = _EVAL_162;
  assign _EVAL_35 = _EVAL_238;
  assign _EVAL_156 = _EVAL_227;
  assign _EVAL_243 = _EVAL_2;
  assign _EVAL_34 = _EVAL_182;
  assign _EVAL_191 = _EVAL_13;
  assign _EVAL_85 = _EVAL_48;
  assign _EVAL_157 = _EVAL_161;
  assign _EVAL_183 = _EVAL_60;
  assign _EVAL_231 = _EVAL_193;
  assign _EVAL_32 = _EVAL_149;
  assign _EVAL_230 = _EVAL_122;
  assign _EVAL_176 = _EVAL_50;
  assign _EVAL_203 = _EVAL_37;
  assign _EVAL_84 = _EVAL_70;
  assign _EVAL_240 = _EVAL_226;
  assign _EVAL_144 = _EVAL_173;
  assign _EVAL_138 = _EVAL_212;
  assign _EVAL_249 = _EVAL_53;
  assign _EVAL_127 = _EVAL_69;
  assign _EVAL_87 = _EVAL_49;
  assign _EVAL_202 = _EVAL_21;
  assign _EVAL_223 = _EVAL_110;
  assign _EVAL_167 = _EVAL_61;
  assign _EVAL_76 = _EVAL_205;
  assign _EVAL_195 = _EVAL_81;
  assign _EVAL_78 = _EVAL_3;
  assign _EVAL_86 = _EVAL_72;
  assign _EVAL_125 = _EVAL_24;
  assign _EVAL_140 = _EVAL_210;
  assign _EVAL_188 = _EVAL_158;
  assign _EVAL_126 = _EVAL_83;
  assign _EVAL_174 = _EVAL_139;
  assign _EVAL_99 = _EVAL_95;
  assign _EVAL_187 = _EVAL_142;
  assign _EVAL_135 = _EVAL_251;
  assign _EVAL_239 = _EVAL_194;
  assign _EVAL_145 = _EVAL_25;
  assign _EVAL_38 = _EVAL_92;
  assign _EVAL_63 = _EVAL_73;
  assign _EVAL_152 = _EVAL_215;
  assign _EVAL_224 = _EVAL_67;
  assign _EVAL_6 = _EVAL_163;
  assign _EVAL_104 = _EVAL_79;
  assign _EVAL_15 = _EVAL_136;
  assign _EVAL_74 = _EVAL_120;
  assign _EVAL_219 = _EVAL_222;
  assign _EVAL_213 = _EVAL_153;
  assign _EVAL_208 = _EVAL_105;
  assign _EVAL_165 = _EVAL;
  assign _EVAL_169 = _EVAL_199;
  assign _EVAL_71 = _EVAL_68;
  assign _EVAL_236 = _EVAL_8;
  assign _EVAL_232 = _EVAL_221;
  assign _EVAL_107 = _EVAL_1;
  assign _EVAL_0 = _EVAL_29;
  assign _EVAL_133 = _EVAL_225;
  assign _EVAL_129 = _EVAL_248;
  assign _EVAL_128 = _EVAL_214;
  assign _EVAL_234 = _EVAL_168;
  assign _EVAL_159 = _EVAL_116;
  assign _EVAL_160 = _EVAL_178;
  assign _EVAL_93 = _EVAL_244;
  assign _EVAL_31 = _EVAL_124;
  assign _EVAL_119 = _EVAL_18;
  assign _EVAL_179 = _EVAL_98;
  assign _EVAL_198 = _EVAL_77;
  assign _EVAL_109 = _EVAL_100;
  assign _EVAL_137 = _EVAL_52;
  assign _EVAL_90 = _EVAL_41;
  assign _EVAL_154 = _EVAL_197;
  assign _EVAL_51 = _EVAL_65;
  assign _EVAL_59 = _EVAL_28;
  assign _EVAL_112 = _EVAL_11;
  assign _EVAL_186 = _EVAL_56;
  assign _EVAL_111 = _EVAL_245;
  assign _EVAL_177 = _EVAL_89;
  assign _EVAL_190 = _EVAL_117;
  assign _EVAL_200 = _EVAL_36;
  assign _EVAL_164 = _EVAL_114;
  assign _EVAL_108 = _EVAL_246;
  assign _EVAL_75 = _EVAL_17;
  assign _EVAL_220 = _EVAL_54;
  assign _EVAL_148 = _EVAL_33;
  assign _EVAL_218 = _EVAL_96;
  assign _EVAL_206 = _EVAL_189;
  assign _EVAL_10 = _EVAL_14;
  assign _EVAL_44 = _EVAL_40;
  assign _EVAL_45 = _EVAL_9;
  assign _EVAL_102 = _EVAL_43;
  assign _EVAL_185 = _EVAL_132;
  assign _EVAL_115 = _EVAL_131;
  assign _EVAL_88 = _EVAL_19;
  assign _EVAL_242 = _EVAL_130;
  assign _EVAL_143 = _EVAL_103;
  assign _EVAL_151 = _EVAL_82;
  assign _EVAL_196 = _EVAL_233;
  assign _EVAL_241 = _EVAL_171;
  assign _EVAL_201 = _EVAL_216;
  assign _EVAL_57 = _EVAL_209;
  assign _EVAL_46 = _EVAL_7;
  assign _EVAL_91 = _EVAL_27;
  assign _EVAL_66 = _EVAL_30;
  assign _EVAL_147 = _EVAL_250;
  assign _EVAL_106 = _EVAL_204;
  assign _EVAL_26 = _EVAL_55;
  assign _EVAL_192 = _EVAL_175;
  assign _EVAL_47 = _EVAL_166;
  assign _EVAL_237 = _EVAL_235;
  assign _EVAL_80 = _EVAL_23;
  assign _EVAL_252 = _EVAL_207;
  assign _EVAL_155 = _EVAL_217;
endmodule
