//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_322(
  input  [8:0]  _EVAL,
  output [8:0]  _EVAL_0,
  input  [8:0]  _EVAL_1,
  input  [7:0]  _EVAL_2,
  output [8:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  output [2:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  output [63:0] _EVAL_10,
  output        _EVAL_11,
  input  [2:0]  _EVAL_12,
  output        _EVAL_13,
  input  [63:0] _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input  [2:0]  _EVAL_17,
  output [2:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  input  [63:0] _EVAL_23,
  output [2:0]  _EVAL_24,
  output [7:0]  _EVAL_25,
  input  [2:0]  _EVAL_26,
  output [2:0]  _EVAL_27,
  output        _EVAL_28,
  output [63:0] _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  output [2:0]  _EVAL_34,
  output [31:0] _EVAL_35,
  input         _EVAL_36
);
  assign _EVAL_10 = _EVAL_14;
  assign _EVAL_18 = _EVAL_26;
  assign _EVAL_11 = _EVAL_6;
  assign _EVAL_24 = _EVAL_5;
  assign _EVAL_28 = _EVAL_36;
  assign _EVAL_7 = _EVAL_12;
  assign _EVAL_22 = _EVAL_33;
  assign _EVAL_0 = _EVAL;
  assign _EVAL_27 = _EVAL_17;
  assign _EVAL_16 = _EVAL_4;
  assign _EVAL_34 = _EVAL_19;
  assign _EVAL_25 = _EVAL_2;
  assign _EVAL_13 = _EVAL_32;
  assign _EVAL_29 = _EVAL_23;
  assign _EVAL_3 = _EVAL_1;
  assign _EVAL_35 = _EVAL_8;
  assign _EVAL_31 = _EVAL_21;
  assign _EVAL_20 = _EVAL_30;
endmodule
