//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_165(
  output        _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output [7:0]  _EVAL_4,
  input         _EVAL_5,
  output [1:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  output [1:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [3:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  input  [1:0]  _EVAL_17,
  input  [31:0] _EVAL_18,
  output [3:0]  _EVAL_19,
  output [2:0]  _EVAL_20,
  input         _EVAL_21,
  input  [1:0]  _EVAL_22,
  output [3:0]  _EVAL_23,
  output [3:0]  _EVAL_24,
  input  [3:0]  _EVAL_25,
  output [29:0] _EVAL_26,
  output [31:0] _EVAL_27,
  input         _EVAL_28,
  input  [2:0]  _EVAL_29,
  input         _EVAL_30,
  output [29:0] _EVAL_31,
  input  [1:0]  _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  output [2:0]  _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  output        _EVAL_40,
  output        _EVAL_41,
  input  [2:0]  _EVAL_42,
  input         _EVAL_43,
  output [2:0]  _EVAL_44,
  output        _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  output [2:0]  _EVAL_49,
  input  [29:0] _EVAL_50,
  output [3:0]  _EVAL_51,
  output [3:0]  _EVAL_52,
  input         _EVAL_53,
  output [1:0]  _EVAL_54,
  output        _EVAL_55,
  input  [7:0]  _EVAL_56,
  input         _EVAL_57,
  input  [7:0]  _EVAL_58,
  input  [2:0]  _EVAL_59,
  output        _EVAL_60,
  output        _EVAL_61,
  output [1:0]  _EVAL_62,
  input  [3:0]  _EVAL_63,
  output        _EVAL_64,
  input  [3:0]  _EVAL_65,
  input  [1:0]  _EVAL_66,
  output [7:0]  _EVAL_67,
  output        _EVAL_68,
  output        _EVAL_69,
  input  [29:0] _EVAL_70
);
  wire [31:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire [31:0] Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire [3:0] Queue_1__EVAL_8;
  wire  Queue_1__EVAL_9;
  wire [3:0] Queue_1__EVAL_10;
  wire [31:0] Queue_4__EVAL;
  wire [1:0] Queue_4__EVAL_0;
  wire  Queue_4__EVAL_1;
  wire [1:0] Queue_4__EVAL_2;
  wire  Queue_4__EVAL_3;
  wire  Queue_4__EVAL_4;
  wire  Queue_4__EVAL_5;
  wire  Queue_4__EVAL_6;
  wire  Queue_4__EVAL_7;
  wire  Queue_4__EVAL_8;
  wire  Queue_4__EVAL_9;
  wire [31:0] Queue_4__EVAL_10;
  wire [1:0] Queue_2__EVAL;
  wire  Queue_2__EVAL_0;
  wire [1:0] Queue_2__EVAL_1;
  wire  Queue_2__EVAL_2;
  wire  Queue_2__EVAL_3;
  wire  Queue_2__EVAL_4;
  wire  Queue_2__EVAL_5;
  wire  Queue_2__EVAL_6;
  wire [7:0] Queue_3__EVAL;
  wire [3:0] Queue_3__EVAL_0;
  wire  Queue_3__EVAL_1;
  wire  Queue_3__EVAL_2;
  wire [2:0] Queue_3__EVAL_3;
  wire  Queue_3__EVAL_4;
  wire [29:0] Queue_3__EVAL_5;
  wire  Queue_3__EVAL_6;
  wire  Queue_3__EVAL_7;
  wire [2:0] Queue_3__EVAL_8;
  wire [7:0] Queue_3__EVAL_9;
  wire  Queue_3__EVAL_10;
  wire [2:0] Queue_3__EVAL_11;
  wire [29:0] Queue_3__EVAL_12;
  wire  Queue_3__EVAL_13;
  wire  Queue_3__EVAL_14;
  wire [3:0] Queue_3__EVAL_15;
  wire [3:0] Queue_3__EVAL_16;
  wire [1:0] Queue_3__EVAL_17;
  wire [2:0] Queue_3__EVAL_18;
  wire [3:0] Queue_3__EVAL_19;
  wire  Queue_3__EVAL_20;
  wire [1:0] Queue_3__EVAL_21;
  wire  Queue_3__EVAL_22;
  wire [7:0] Queue__EVAL;
  wire [3:0] Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire [2:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire [29:0] Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire [2:0] Queue__EVAL_8;
  wire [7:0] Queue__EVAL_9;
  wire  Queue__EVAL_10;
  wire [2:0] Queue__EVAL_11;
  wire [29:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire [3:0] Queue__EVAL_15;
  wire [3:0] Queue__EVAL_16;
  wire [1:0] Queue__EVAL_17;
  wire [2:0] Queue__EVAL_18;
  wire [3:0] Queue__EVAL_19;
  wire  Queue__EVAL_20;
  wire [1:0] Queue__EVAL_21;
  wire  Queue__EVAL_22;
  SiFive__EVAL_22 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10)
  );
  SiFive__EVAL_164 Queue_4 (
    ._EVAL(Queue_4__EVAL),
    ._EVAL_0(Queue_4__EVAL_0),
    ._EVAL_1(Queue_4__EVAL_1),
    ._EVAL_2(Queue_4__EVAL_2),
    ._EVAL_3(Queue_4__EVAL_3),
    ._EVAL_4(Queue_4__EVAL_4),
    ._EVAL_5(Queue_4__EVAL_5),
    ._EVAL_6(Queue_4__EVAL_6),
    ._EVAL_7(Queue_4__EVAL_7),
    ._EVAL_8(Queue_4__EVAL_8),
    ._EVAL_9(Queue_4__EVAL_9),
    ._EVAL_10(Queue_4__EVAL_10)
  );
  SiFive__EVAL_163 Queue_2 (
    ._EVAL(Queue_2__EVAL),
    ._EVAL_0(Queue_2__EVAL_0),
    ._EVAL_1(Queue_2__EVAL_1),
    ._EVAL_2(Queue_2__EVAL_2),
    ._EVAL_3(Queue_2__EVAL_3),
    ._EVAL_4(Queue_2__EVAL_4),
    ._EVAL_5(Queue_2__EVAL_5),
    ._EVAL_6(Queue_2__EVAL_6)
  );
  SiFive__EVAL_162 Queue_3 (
    ._EVAL(Queue_3__EVAL),
    ._EVAL_0(Queue_3__EVAL_0),
    ._EVAL_1(Queue_3__EVAL_1),
    ._EVAL_2(Queue_3__EVAL_2),
    ._EVAL_3(Queue_3__EVAL_3),
    ._EVAL_4(Queue_3__EVAL_4),
    ._EVAL_5(Queue_3__EVAL_5),
    ._EVAL_6(Queue_3__EVAL_6),
    ._EVAL_7(Queue_3__EVAL_7),
    ._EVAL_8(Queue_3__EVAL_8),
    ._EVAL_9(Queue_3__EVAL_9),
    ._EVAL_10(Queue_3__EVAL_10),
    ._EVAL_11(Queue_3__EVAL_11),
    ._EVAL_12(Queue_3__EVAL_12),
    ._EVAL_13(Queue_3__EVAL_13),
    ._EVAL_14(Queue_3__EVAL_14),
    ._EVAL_15(Queue_3__EVAL_15),
    ._EVAL_16(Queue_3__EVAL_16),
    ._EVAL_17(Queue_3__EVAL_17),
    ._EVAL_18(Queue_3__EVAL_18),
    ._EVAL_19(Queue_3__EVAL_19),
    ._EVAL_20(Queue_3__EVAL_20),
    ._EVAL_21(Queue_3__EVAL_21),
    ._EVAL_22(Queue_3__EVAL_22)
  );
  SiFive__EVAL_162 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18),
    ._EVAL_19(Queue__EVAL_19),
    ._EVAL_20(Queue__EVAL_20),
    ._EVAL_21(Queue__EVAL_21),
    ._EVAL_22(Queue__EVAL_22)
  );
  assign Queue_3__EVAL_5 = _EVAL_50;
  assign Queue_3__EVAL_11 = _EVAL_29;
  assign _EVAL_51 = Queue_3__EVAL_16;
  assign Queue__EVAL = _EVAL_58;
  assign Queue_4__EVAL_10 = _EVAL_18;
  assign _EVAL = Queue__EVAL_4;
  assign Queue__EVAL_11 = _EVAL_42;
  assign _EVAL_60 = Queue_2__EVAL_4;
  assign _EVAL_55 = Queue_1__EVAL_7;
  assign Queue_1__EVAL_8 = _EVAL_65;
  assign _EVAL_33 = Queue__EVAL_13;
  assign Queue__EVAL_17 = _EVAL_66;
  assign _EVAL_24 = Queue__EVAL_16;
  assign _EVAL_41 = Queue_4__EVAL_3;
  assign _EVAL_47 = Queue__EVAL_20;
  assign Queue_3__EVAL_6 = _EVAL_28;
  assign Queue_3__EVAL_14 = _EVAL_43;
  assign _EVAL_19 = Queue_1__EVAL_10;
  assign _EVAL_16 = Queue_4__EVAL;
  assign Queue_3__EVAL_22 = _EVAL_36;
  assign Queue_4__EVAL_4 = _EVAL_0;
  assign _EVAL_11 = Queue_3__EVAL_21;
  assign _EVAL_20 = Queue_3__EVAL_8;
  assign Queue_4__EVAL_1 = _EVAL_35;
  assign Queue__EVAL_14 = _EVAL_39;
  assign _EVAL_64 = Queue_3__EVAL_4;
  assign Queue_3__EVAL_2 = _EVAL_35;
  assign _EVAL_26 = Queue__EVAL_12;
  assign Queue_1__EVAL_2 = _EVAL_35;
  assign Queue_2__EVAL_1 = _EVAL_22;
  assign _EVAL_23 = Queue_3__EVAL_0;
  assign Queue_4__EVAL_9 = _EVAL_2;
  assign _EVAL_61 = Queue_3__EVAL_13;
  assign Queue_2__EVAL_6 = _EVAL_36;
  assign _EVAL_7 = Queue_2__EVAL_0;
  assign Queue_1__EVAL = _EVAL_14;
  assign _EVAL_40 = Queue_3__EVAL_20;
  assign Queue__EVAL_2 = _EVAL_35;
  assign Queue_3__EVAL_19 = _EVAL_12;
  assign _EVAL_67 = Queue__EVAL_9;
  assign _EVAL_68 = Queue_4__EVAL_7;
  assign Queue_1__EVAL_0 = _EVAL_3;
  assign _EVAL_69 = Queue_1__EVAL_6;
  assign Queue__EVAL_22 = _EVAL_36;
  assign Queue__EVAL_5 = _EVAL_70;
  assign _EVAL_62 = Queue_4__EVAL_2;
  assign _EVAL_9 = Queue__EVAL_10;
  assign Queue_3__EVAL = _EVAL_56;
  assign Queue_2__EVAL_2 = _EVAL_35;
  assign Queue__EVAL_1 = _EVAL_13;
  assign _EVAL_6 = Queue_2__EVAL;
  assign Queue_3__EVAL_1 = _EVAL_38;
  assign Queue_2__EVAL_5 = _EVAL_8;
  assign _EVAL_48 = Queue_1__EVAL_5;
  assign Queue__EVAL_6 = _EVAL_10;
  assign Queue_4__EVAL_8 = _EVAL_57;
  assign Queue_2__EVAL_3 = _EVAL_5;
  assign Queue__EVAL_19 = _EVAL_15;
  assign _EVAL_34 = Queue_4__EVAL_5;
  assign Queue_3__EVAL_3 = _EVAL_1;
  assign Queue_1__EVAL_9 = _EVAL_46;
  assign Queue_3__EVAL_17 = _EVAL_32;
  assign _EVAL_44 = Queue__EVAL_8;
  assign _EVAL_31 = Queue_3__EVAL_12;
  assign _EVAL_27 = Queue_1__EVAL_3;
  assign Queue__EVAL_15 = _EVAL_63;
  assign Queue_4__EVAL_6 = _EVAL_36;
  assign Queue__EVAL_7 = _EVAL_21;
  assign _EVAL_45 = Queue_3__EVAL_10;
  assign Queue__EVAL_3 = _EVAL_59;
  assign _EVAL_49 = Queue__EVAL_18;
  assign Queue_1__EVAL_4 = _EVAL_36;
  assign _EVAL_4 = Queue_3__EVAL_9;
  assign Queue_4__EVAL_0 = _EVAL_17;
  assign _EVAL_37 = Queue_3__EVAL_18;
  assign _EVAL_54 = Queue__EVAL_21;
  assign Queue_3__EVAL_15 = _EVAL_25;
  assign _EVAL_52 = Queue__EVAL_0;
  assign Queue_3__EVAL_7 = _EVAL_30;
  assign Queue_1__EVAL_1 = _EVAL_53;
endmodule
