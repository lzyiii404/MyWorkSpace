//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_328(
  output        _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  output [6:0]  _EVAL_2,
  output        _EVAL_3,
  input  [6:0]  _EVAL_4,
  input  [31:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [1:0]  _EVAL_11,
  output [1:0]  _EVAL_12,
  output [31:0] _EVAL_13
);
  reg  _EVAL_14;
  reg [31:0] _RAND_0;
  reg  _EVAL_23;
  reg [31:0] _RAND_1;
  reg  _EVAL_28;
  reg [31:0] _RAND_2;
  reg  _EVAL_38;
  reg [31:0] _RAND_3;
  reg  _EVAL_39;
  reg [31:0] _RAND_4;
  reg  _EVAL_40;
  reg [31:0] _RAND_5;
  reg  _EVAL_41;
  reg [31:0] _RAND_6;
  reg  _EVAL_49;
  reg [31:0] _RAND_7;
  reg  _EVAL_51;
  reg [31:0] _RAND_8;
  reg  _EVAL_52;
  reg [31:0] _RAND_9;
  reg  _EVAL_61;
  reg [31:0] _RAND_10;
  reg  _EVAL_64;
  reg [31:0] _RAND_11;
  reg  _EVAL_68;
  reg [31:0] _RAND_12;
  reg  _EVAL_73;
  reg [31:0] _RAND_13;
  reg  _EVAL_78;
  reg [31:0] _RAND_14;
  reg  _EVAL_82;
  reg [31:0] _RAND_15;
  reg  _EVAL_84;
  reg [31:0] _RAND_16;
  reg  _EVAL_86;
  reg [31:0] _RAND_17;
  reg  _EVAL_87;
  reg [31:0] _RAND_18;
  reg  _EVAL_89;
  reg [31:0] _RAND_19;
  reg  _EVAL_93;
  reg [31:0] _RAND_20;
  reg  _EVAL_94;
  reg [31:0] _RAND_21;
  reg  _EVAL_95;
  reg [31:0] _RAND_22;
  reg  _EVAL_100;
  reg [31:0] _RAND_23;
  reg  _EVAL_101;
  reg [31:0] _RAND_24;
  reg  _EVAL_111;
  reg [31:0] _RAND_25;
  reg  _EVAL_115;
  reg [31:0] _RAND_26;
  reg  _EVAL_118;
  reg [31:0] _RAND_27;
  reg  _EVAL_126;
  reg [31:0] _RAND_28;
  reg  _EVAL_127;
  reg [31:0] _RAND_29;
  reg  _EVAL_128;
  reg [31:0] _RAND_30;
  reg  _EVAL_131;
  reg [31:0] _RAND_31;
  reg  _EVAL_135;
  reg [31:0] _RAND_32;
  reg  _EVAL_140;
  reg [31:0] _RAND_33;
  reg  _EVAL_148;
  reg [31:0] _RAND_34;
  reg  _EVAL_149;
  reg [31:0] _RAND_35;
  reg  _EVAL_167;
  reg [31:0] _RAND_36;
  reg  _EVAL_168;
  reg [31:0] _RAND_37;
  reg  _EVAL_181;
  reg [31:0] _RAND_38;
  reg  _EVAL_187;
  reg [31:0] _RAND_39;
  reg  _EVAL_188;
  reg [31:0] _RAND_40;
  wire [9:0] _EVAL_66;
  wire [40:0] _EVAL_193;
  wire  _EVAL_129;
  wire  _EVAL_88;
  wire  _EVAL_170;
  wire  _EVAL_99;
  wire  _EVAL_136;
  wire  _EVAL_50;
  wire  _EVAL_34;
  wire [4:0] _EVAL_183;
  wire [9:0] _EVAL_43;
  wire [9:0] _EVAL_130;
  wire [40:0] _EVAL_116;
  wire  _EVAL_108;
  wire  _EVAL_145;
  wire  _EVAL_60;
  wire  _EVAL_133;
  wire  _EVAL_46;
  wire  _EVAL_21;
  wire  _EVAL_81;
  wire  _EVAL_109;
  wire  _EVAL_143;
  wire  _EVAL_158;
  wire  _EVAL_150;
  wire  _EVAL_110;
  wire  _EVAL_83;
  wire  _EVAL_25;
  wire  _EVAL_124;
  wire  _EVAL_65;
  wire  _EVAL_74;
  wire  _EVAL_32;
  wire  _EVAL_62;
  wire  _EVAL_142;
  wire  _EVAL_26;
  wire  _EVAL_185;
  wire  _EVAL_161;
  wire  _EVAL_72;
  wire  _EVAL_117;
  wire  _EVAL_75;
  wire  _EVAL_113;
  wire  _EVAL_105;
  wire  _EVAL_119;
  wire  _EVAL_91;
  wire  _EVAL_165;
  wire  _EVAL_70;
  wire  _EVAL_125;
  wire  _EVAL_59;
  assign _EVAL_66 = {_EVAL_168,_EVAL_111,_EVAL_40,_EVAL_135,_EVAL_94,_EVAL_73,_EVAL_23,_EVAL_131,_EVAL_41,_EVAL_149};
  assign _EVAL_193 = {_EVAL_4,_EVAL_5,_EVAL_11};
  assign _EVAL_129 = _EVAL_193[3];
  assign _EVAL_88 = _EVAL_193[27];
  assign _EVAL_170 = _EVAL_193[18];
  assign _EVAL_99 = _EVAL_193[28];
  assign _EVAL_136 = _EVAL_193[13];
  assign _EVAL_50 = _EVAL_193[12];
  assign _EVAL_34 = _EVAL_193[17];
  assign _EVAL_183 = {_EVAL_64,_EVAL_127,_EVAL_39,_EVAL_38,_EVAL_93};
  assign _EVAL_43 = {_EVAL_87,_EVAL_101,_EVAL_148,_EVAL_188,_EVAL_28,_EVAL_68,_EVAL_49,_EVAL_128,_EVAL_82,_EVAL_14};
  assign _EVAL_130 = {_EVAL_52,_EVAL_187,_EVAL_61,_EVAL_89,_EVAL_167,_EVAL_78,_EVAL_115,_EVAL_181,_EVAL_118,_EVAL_126};
  assign _EVAL_116 = {_EVAL_100,_EVAL_86,_EVAL_95,_EVAL_84,_EVAL_140,_EVAL_51,_EVAL_183,_EVAL_43,_EVAL_130,_EVAL_66};
  assign _EVAL_108 = _EVAL_193[2];
  assign _EVAL_145 = _EVAL_193[16];
  assign _EVAL_60 = _EVAL_193[24];
  assign _EVAL_133 = _EVAL_193[40];
  assign _EVAL_46 = _EVAL_193[0];
  assign _EVAL_21 = _EVAL_193[1];
  assign _EVAL_81 = _EVAL_193[36];
  assign _EVAL_109 = _EVAL_193[8];
  assign _EVAL_143 = _EVAL_193[25];
  assign _EVAL_158 = _EVAL_193[23];
  assign _EVAL_150 = _EVAL_193[38];
  assign _EVAL_110 = _EVAL_193[11];
  assign _EVAL_83 = _EVAL_193[14];
  assign _EVAL_25 = _EVAL_193[19];
  assign _EVAL_124 = _EVAL_193[31];
  assign _EVAL_65 = _EVAL_193[29];
  assign _EVAL_74 = _EVAL_193[15];
  assign _EVAL_32 = _EVAL_193[7];
  assign _EVAL_62 = _EVAL_193[34];
  assign _EVAL_142 = _EVAL_193[39];
  assign _EVAL_26 = _EVAL_193[9];
  assign _EVAL_185 = _EVAL_193[26];
  assign _EVAL_161 = _EVAL_193[37];
  assign _EVAL_72 = _EVAL_193[6];
  assign _EVAL_117 = _EVAL_193[32];
  assign _EVAL_75 = _EVAL_193[10];
  assign _EVAL_113 = _EVAL_193[20];
  assign _EVAL_105 = _EVAL_193[33];
  assign _EVAL_119 = _EVAL_193[21];
  assign _EVAL_91 = _EVAL_193[30];
  assign _EVAL_165 = _EVAL_193[35];
  assign _EVAL_70 = _EVAL_193[22];
  assign _EVAL_125 = _EVAL_193[5];
  assign _EVAL_59 = _EVAL_193[4];
  assign _EVAL = _EVAL_0;
  assign _EVAL_12 = _EVAL_116[1:0];
  assign _EVAL_13 = _EVAL_116[33:2];
  assign _EVAL_3 = _EVAL_149;
  assign _EVAL_1 = _EVAL_0 ? 1'h0 : _EVAL_9;
  assign _EVAL_2 = _EVAL_116[40:34];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_14 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_23 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_28 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_38 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_39 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_40 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_41 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_49 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_51 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_52 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_61 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_64 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_68 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_73 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_78 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_82 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_84 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_86 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_87 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_89 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_93 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_94 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_95 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_100 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_101 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_111 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_115 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_118 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_126 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_127 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_128 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_131 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_135 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_140 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_148 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_149 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_167 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_168 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_181 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_187 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_188 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_8) begin
    if (_EVAL_0) begin
      _EVAL_14 <= _EVAL_113;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_14 <= _EVAL_82;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_23 <= _EVAL_129;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_23 <= _EVAL_73;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_28 <= _EVAL_143;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_28 <= _EVAL_188;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_38 <= _EVAL_124;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_38 <= _EVAL_39;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_39 <= _EVAL_117;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_39 <= _EVAL_127;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_40 <= _EVAL_32;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_40 <= _EVAL_111;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_41 <= _EVAL_21;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_41 <= _EVAL_131;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_49 <= _EVAL_158;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_49 <= _EVAL_68;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_51 <= _EVAL_165;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_51 <= _EVAL_140;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_52 <= _EVAL_25;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_52 <= _EVAL_14;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_61 <= _EVAL_34;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_61 <= _EVAL_187;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_64 <= _EVAL_62;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_64 <= _EVAL_51;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_68 <= _EVAL_60;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_68 <= _EVAL_28;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_73 <= _EVAL_59;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_73 <= _EVAL_94;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_78 <= _EVAL_83;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_78 <= _EVAL_167;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_82 <= _EVAL_119;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_82 <= _EVAL_128;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_84 <= _EVAL_161;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_84 <= _EVAL_95;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_86 <= _EVAL_142;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_86 <= _EVAL_100;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_87 <= _EVAL_65;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_87 <= _EVAL_93;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_89 <= _EVAL_145;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_89 <= _EVAL_61;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_93 <= _EVAL_91;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_93 <= _EVAL_38;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_94 <= _EVAL_125;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_94 <= _EVAL_135;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_95 <= _EVAL_150;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_95 <= _EVAL_86;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_100 <= _EVAL_133;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_100 <= _EVAL_7;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_101 <= _EVAL_99;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_101 <= _EVAL_87;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_111 <= _EVAL_109;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_111 <= _EVAL_168;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_115 <= _EVAL_136;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_115 <= _EVAL_78;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_118 <= _EVAL_110;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_118 <= _EVAL_181;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_126 <= _EVAL_75;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_126 <= _EVAL_118;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_127 <= _EVAL_105;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_127 <= _EVAL_64;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_128 <= _EVAL_70;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_128 <= _EVAL_49;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_131 <= _EVAL_108;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_131 <= _EVAL_23;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_135 <= _EVAL_72;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_135 <= _EVAL_40;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_140 <= _EVAL_81;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_140 <= _EVAL_84;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_148 <= _EVAL_88;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_148 <= _EVAL_101;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_149 <= _EVAL_46;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_149 <= _EVAL_41;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_167 <= _EVAL_74;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_167 <= _EVAL_89;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_168 <= _EVAL_26;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_168 <= _EVAL_126;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_181 <= _EVAL_50;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_181 <= _EVAL_115;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_187 <= _EVAL_170;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_187 <= _EVAL_52;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_188 <= _EVAL_185;
    end else begin
      if (!(_EVAL_9)) begin
        if (_EVAL_10) begin
          _EVAL_188 <= _EVAL_148;
        end
      end
    end
  end
endmodule
