//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_65_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [4:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [4:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [5:0] _EVAL_25;
  reg [31:0] _RAND_0;
  reg [5:0] _EVAL_33;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_50;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_74;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_79;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_86;
  reg [31:0] _RAND_5;
  reg [5:0] _EVAL_133;
  reg [31:0] _RAND_6;
  reg [4:0] _EVAL_134;
  reg [31:0] _RAND_7;
  reg [31:0] _EVAL_150;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_156;
  reg [31:0] _RAND_9;
  reg  _EVAL_175;
  reg [31:0] _RAND_10;
  reg  _EVAL_192;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_268;
  reg [31:0] _RAND_12;
  reg [5:0] _EVAL_287;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_288;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_326;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_355;
  reg [31:0] _RAND_16;
  wire  _EVAL_146;
  wire  _EVAL_84;
  wire  _EVAL_154;
  wire [31:0] _EVAL_53;
  wire [31:0] _EVAL_271;
  wire  _EVAL_77;
  wire  _EVAL_210;
  wire  _EVAL_75;
  wire  _EVAL_168;
  wire  _EVAL_119;
  wire  _EVAL_318;
  wire [31:0] _EVAL_334;
  wire [31:0] _EVAL_121;
  wire  _EVAL_98;
  wire  _EVAL_26;
  wire  _EVAL_108;
  wire  _EVAL_65;
  wire  _EVAL_219;
  wire  _EVAL_96;
  wire  _EVAL_137;
  wire  _EVAL_63;
  wire  _EVAL_322;
  wire  _EVAL_293;
  wire  _EVAL_236;
  wire [22:0] _EVAL_350;
  wire [7:0] _EVAL_78;
  wire [7:0] _EVAL_60;
  wire [31:0] _EVAL_329;
  wire [31:0] _EVAL_282;
  wire  _EVAL_55;
  wire  _EVAL_214;
  wire  _EVAL_52;
  wire [32:0] _EVAL_352;
  wire [32:0] _EVAL_218;
  wire [1:0] _EVAL_278;
  wire  _EVAL_159;
  wire  _EVAL_142;
  wire  _EVAL_317;
  wire  _EVAL_224;
  wire  _EVAL_70;
  wire  _EVAL_131;
  wire  _EVAL_196;
  wire  _EVAL_321;
  wire  _EVAL_62;
  wire  _EVAL_124;
  wire  _EVAL_103;
  wire  _EVAL_111;
  wire  _EVAL_182;
  wire  _EVAL_128;
  wire  _EVAL_266;
  wire  _EVAL_127;
  wire  _EVAL_190;
  wire  _EVAL_209;
  wire  _EVAL_306;
  wire  _EVAL_347;
  wire  _EVAL_183;
  wire  _EVAL_311;
  wire [22:0] _EVAL_163;
  wire [7:0] _EVAL_240;
  wire [7:0] _EVAL_221;
  wire [5:0] _EVAL_171;
  wire [31:0] _EVAL_216;
  wire [32:0] _EVAL_202;
  wire [32:0] _EVAL_76;
  wire [32:0] _EVAL_247;
  wire  _EVAL_47;
  wire  _EVAL_90;
  wire  _EVAL_297;
  wire [1:0] _EVAL_177;
  wire [1:0] _EVAL_195;
  wire  _EVAL_258;
  wire  _EVAL_116;
  wire  _EVAL_298;
  wire  _EVAL_349;
  wire  _EVAL_260;
  wire  _EVAL_290;
  wire  _EVAL_237;
  wire  _EVAL_275;
  wire  _EVAL_158;
  wire  _EVAL_264;
  wire  _EVAL_105;
  wire  _EVAL_301;
  wire  _EVAL_178;
  wire  _EVAL_173;
  wire  _EVAL_130;
  wire  _EVAL_102;
  wire  _EVAL_341;
  wire [3:0] _EVAL_144;
  wire  _EVAL_45;
  wire [3:0] _EVAL_339;
  wire [3:0] _EVAL_204;
  wire  _EVAL_68;
  wire  _EVAL_136;
  wire  _EVAL_57;
  wire  _EVAL_256;
  wire  _EVAL_205;
  wire  _EVAL_338;
  wire  _EVAL_106;
  wire  _EVAL_348;
  wire  _EVAL_38;
  wire [31:0] _EVAL_233;
  wire [32:0] _EVAL_155;
  wire [32:0] _EVAL_346;
  wire [32:0] _EVAL_340;
  wire  _EVAL_49;
  wire  _EVAL_143;
  wire [31:0] _EVAL_324;
  wire [32:0] _EVAL_176;
  wire [32:0] _EVAL_91;
  wire [32:0] _EVAL_284;
  wire  _EVAL_153;
  wire  _EVAL_165;
  wire [31:0] _EVAL_118;
  wire [32:0] _EVAL_342;
  wire [32:0] _EVAL_43;
  wire [32:0] _EVAL_245;
  wire  _EVAL_331;
  wire  _EVAL_35;
  wire  _EVAL_302;
  wire [31:0] _EVAL_295;
  wire [32:0] _EVAL_343;
  wire [32:0] _EVAL_29;
  wire [32:0] _EVAL_208;
  wire  _EVAL_48;
  wire  _EVAL_114;
  wire  _EVAL_328;
  wire [32:0] _EVAL_252;
  wire  _EVAL_251;
  wire  _EVAL_194;
  wire [31:0] _EVAL_200;
  wire [32:0] _EVAL_32;
  wire [32:0] _EVAL_310;
  wire [32:0] _EVAL_235;
  wire  _EVAL_313;
  wire  _EVAL_241;
  wire [31:0] _EVAL_64;
  wire [32:0] _EVAL_39;
  wire [32:0] _EVAL_296;
  wire [32:0] _EVAL_54;
  wire  _EVAL_274;
  wire  _EVAL_291;
  wire [31:0] _EVAL_198;
  wire [32:0] _EVAL_117;
  wire [32:0] _EVAL_327;
  wire [32:0] _EVAL_259;
  wire  _EVAL_253;
  wire  _EVAL_123;
  wire  _EVAL_132;
  wire  _EVAL_44;
  wire [31:0] _EVAL_263;
  wire [31:0] _EVAL_344;
  wire  _EVAL_185;
  wire  _EVAL_174;
  wire  _EVAL_169;
  wire  _EVAL_307;
  wire [5:0] _EVAL_167;
  wire [3:0] _EVAL_184;
  wire  _EVAL_170;
  wire  _EVAL_335;
  wire  _EVAL_248;
  wire  _EVAL_161;
  wire  _EVAL_58;
  wire  _EVAL_110;
  wire  _EVAL_61;
  wire  _EVAL_228;
  wire  _EVAL_267;
  wire  _EVAL_262;
  wire  _EVAL_89;
  wire [5:0] _EVAL_332;
  wire  _EVAL_23;
  wire  _EVAL_303;
  wire  _EVAL_356;
  wire  _EVAL_211;
  wire [31:0] _EVAL_187;
  wire  _EVAL_101;
  wire  _EVAL_160;
  wire  _EVAL_239;
  wire  _EVAL_299;
  wire  _EVAL_42;
  wire  _EVAL_265;
  wire  _EVAL_238;
  wire  _EVAL_292;
  wire  _EVAL_227;
  wire  _EVAL_166;
  wire  _EVAL_191;
  wire  _EVAL_312;
  wire  _EVAL_85;
  wire  _EVAL_149;
  wire  _EVAL_270;
  wire  _EVAL_222;
  wire  _EVAL_243;
  wire  _EVAL_115;
  wire  _EVAL_325;
  wire [5:0] _EVAL_80;
  wire  _EVAL_99;
  wire  _EVAL_280;
  wire  _EVAL_285;
  wire  _EVAL_107;
  wire  _EVAL_277;
  wire  _EVAL_289;
  wire  _EVAL_37;
  wire  _EVAL_152;
  wire  _EVAL_92;
  wire  _EVAL_206;
  wire  _EVAL_314;
  wire  _EVAL_24;
  wire  _EVAL_88;
  wire  _EVAL_294;
  wire  _EVAL_300;
  wire  _EVAL_125;
  wire  _EVAL_31;
  wire  _EVAL_223;
  wire  _EVAL_351;
  wire  _EVAL_113;
  wire  _EVAL_97;
  wire  _EVAL_286;
  wire  _EVAL_213;
  wire  _EVAL_82;
  wire  _EVAL_66;
  wire [1:0] _EVAL_353;
  wire  _EVAL_272;
  wire  _EVAL_129;
  wire  _EVAL_40;
  wire  _EVAL_120;
  wire  _EVAL_104;
  wire  _EVAL_93;
  wire  _EVAL_157;
  wire  _EVAL_30;
  wire  _EVAL_181;
  wire  _EVAL_100;
  wire  _EVAL_20;
  wire  _EVAL_323;
  wire  _EVAL_95;
  wire [5:0] _EVAL_232;
  wire [31:0] _EVAL_46;
  wire  _EVAL_330;
  wire  _EVAL_122;
  wire  _EVAL_109;
  wire  _EVAL_242;
  wire  _EVAL_207;
  wire  _EVAL_316;
  wire  _EVAL_234;
  wire  _EVAL_226;
  wire  _EVAL_27;
  wire  _EVAL_345;
  wire  _EVAL_255;
  wire [31:0] _EVAL_56;
  wire [31:0] _EVAL_230;
  wire [31:0] _EVAL_145;
  wire  _EVAL_112;
  wire  _EVAL_315;
  wire  _EVAL_336;
  wire  _EVAL_279;
  wire  _EVAL_197;
  wire  _EVAL_308;
  wire  _EVAL_305;
  wire  _EVAL_81;
  wire  _EVAL_34;
  wire  _EVAL_354;
  wire  _EVAL_164;
  wire  _EVAL_180;
  wire  _EVAL_147;
  wire  _EVAL_201;
  wire  _EVAL_41;
  wire  _EVAL_220;
  wire  _EVAL_269;
  wire  _EVAL_21;
  wire  _EVAL_141;
  wire  _EVAL_215;
  wire  _EVAL_179;
  wire  _EVAL_333;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_71;
  wire  _EVAL_283;
  wire  _EVAL_229;
  wire  _EVAL_19;
  wire  _EVAL_28;
  wire  _EVAL_273;
  wire  _EVAL_73;
  wire  _EVAL_51;
  wire [5:0] _EVAL_203;
  wire  _EVAL_151;
  wire  _EVAL_140;
  wire  _EVAL_138;
  wire  _EVAL_126;
  wire  _EVAL_337;
  wire  _EVAL_320;
  wire  _EVAL_22;
  wire  _EVAL_231;
  wire  _EVAL_72;
  wire  _EVAL_199;
  wire  _EVAL_217;
  wire  _EVAL_304;
  wire  _EVAL_139;
  wire  _EVAL_193;
  wire  _EVAL_276;
  wire  _EVAL_87;
  wire  _EVAL_94;
  wire  _EVAL_69;
  wire  _EVAL_319;
  wire  _EVAL_67;
  wire  _EVAL_257;
  wire  _EVAL_281;
  wire  _EVAL_189;
  wire  _EVAL_244;
  wire  _EVAL_186;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_146 = _EVAL_16 & _EVAL_14;
  assign _EVAL_84 = _EVAL_133 == 6'h0;
  assign _EVAL_154 = _EVAL_146 & _EVAL_84;
  assign _EVAL_53 = 32'h1 << _EVAL_6;
  assign _EVAL_271 = _EVAL_154 ? _EVAL_53 : 32'h0;
  assign _EVAL_77 = _EVAL_12 & _EVAL_18;
  assign _EVAL_210 = _EVAL_25 == 6'h0;
  assign _EVAL_75 = _EVAL_77 & _EVAL_210;
  assign _EVAL_168 = _EVAL == 3'h6;
  assign _EVAL_119 = _EVAL_168 == 1'h0;
  assign _EVAL_318 = _EVAL_75 & _EVAL_119;
  assign _EVAL_334 = 32'h1 << _EVAL_10;
  assign _EVAL_121 = _EVAL_318 ? _EVAL_334 : 32'h0;
  assign _EVAL_98 = _EVAL_271 != _EVAL_121;
  assign _EVAL_26 = _EVAL_271 != 32'h0;
  assign _EVAL_108 = _EVAL_26 == 1'h0;
  assign _EVAL_65 = _EVAL_98 | _EVAL_108;
  assign _EVAL_219 = _EVAL_65 | _EVAL_5;
  assign _EVAL_96 = _EVAL_9 <= 3'h3;
  assign _EVAL_137 = _EVAL_96 | _EVAL_5;
  assign _EVAL_63 = _EVAL_137 == 1'h0;
  assign _EVAL_322 = _EVAL_287 == 6'h0;
  assign _EVAL_293 = _EVAL_322 == 1'h0;
  assign _EVAL_236 = _EVAL_14 & _EVAL_293;
  assign _EVAL_350 = 23'hff << _EVAL_4;
  assign _EVAL_78 = _EVAL_350[7:0];
  assign _EVAL_60 = ~ _EVAL_78;
  assign _EVAL_329 = {{24'd0}, _EVAL_60};
  assign _EVAL_282 = _EVAL_2 & _EVAL_329;
  assign _EVAL_55 = _EVAL_282 == 32'h0;
  assign _EVAL_214 = _EVAL_55 | _EVAL_5;
  assign _EVAL_52 = _EVAL_214 == 1'h0;
  assign _EVAL_352 = {1'b0,$signed(_EVAL_2)};
  assign _EVAL_218 = $signed(_EVAL_352) & $signed(-33'sh5000);
  assign _EVAL_278 = _EVAL_6[4:3];
  assign _EVAL_159 = _EVAL_278 == 2'h0;
  assign _EVAL_142 = _EVAL_278 == 2'h1;
  assign _EVAL_317 = _EVAL_159 | _EVAL_142;
  assign _EVAL_224 = _EVAL_278 == 2'h2;
  assign _EVAL_70 = _EVAL_317 | _EVAL_224;
  assign _EVAL_131 = _EVAL_1 == 2'h0;
  assign _EVAL_196 = _EVAL_131 | _EVAL_5;
  assign _EVAL_321 = _EVAL_196 == 1'h0;
  assign _EVAL_62 = _EVAL_268 != 32'h0;
  assign _EVAL_124 = _EVAL_62 == 1'h0;
  assign _EVAL_103 = _EVAL_3 == _EVAL_355;
  assign _EVAL_111 = _EVAL_103 | _EVAL_5;
  assign _EVAL_182 = _EVAL_111 == 1'h0;
  assign _EVAL_128 = _EVAL_2[1];
  assign _EVAL_266 = _EVAL_128 == 1'h0;
  assign _EVAL_127 = _EVAL_2[0];
  assign _EVAL_190 = _EVAL_127 == 1'h0;
  assign _EVAL_209 = _EVAL_266 & _EVAL_190;
  assign _EVAL_306 = _EVAL_15 == 3'h2;
  assign _EVAL_347 = _EVAL_1 != 2'h2;
  assign _EVAL_183 = _EVAL_347 | _EVAL_5;
  assign _EVAL_311 = _EVAL[0];
  assign _EVAL_163 = 23'hff << _EVAL_3;
  assign _EVAL_240 = _EVAL_163[7:0];
  assign _EVAL_221 = ~ _EVAL_240;
  assign _EVAL_171 = _EVAL_221[7:2];
  assign _EVAL_216 = _EVAL_2 ^ 32'h80000000;
  assign _EVAL_202 = {1'b0,$signed(_EVAL_216)};
  assign _EVAL_76 = $signed(_EVAL_202) & $signed(-33'sh20000);
  assign _EVAL_247 = $signed(_EVAL_76);
  assign _EVAL_47 = _EVAL_4 == _EVAL_50;
  assign _EVAL_90 = _EVAL_4 >= 4'h2;
  assign _EVAL_297 = _EVAL_4[0];
  assign _EVAL_177 = 2'h1 << _EVAL_297;
  assign _EVAL_195 = _EVAL_177 | 2'h1;
  assign _EVAL_258 = _EVAL_195[1];
  assign _EVAL_116 = _EVAL_258 & _EVAL_128;
  assign _EVAL_298 = _EVAL_90 | _EVAL_116;
  assign _EVAL_349 = _EVAL_195[0];
  assign _EVAL_260 = _EVAL_128 & _EVAL_127;
  assign _EVAL_290 = _EVAL_349 & _EVAL_260;
  assign _EVAL_237 = _EVAL_298 | _EVAL_290;
  assign _EVAL_275 = _EVAL_128 & _EVAL_190;
  assign _EVAL_158 = _EVAL_349 & _EVAL_275;
  assign _EVAL_264 = _EVAL_298 | _EVAL_158;
  assign _EVAL_105 = _EVAL_258 & _EVAL_266;
  assign _EVAL_301 = _EVAL_90 | _EVAL_105;
  assign _EVAL_178 = _EVAL_266 & _EVAL_127;
  assign _EVAL_173 = _EVAL_349 & _EVAL_178;
  assign _EVAL_130 = _EVAL_301 | _EVAL_173;
  assign _EVAL_102 = _EVAL_349 & _EVAL_209;
  assign _EVAL_341 = _EVAL_301 | _EVAL_102;
  assign _EVAL_144 = {_EVAL_237,_EVAL_264,_EVAL_130,_EVAL_341};
  assign _EVAL_45 = _EVAL_17 == _EVAL_144;
  assign _EVAL_339 = ~ _EVAL_144;
  assign _EVAL_204 = _EVAL_17 & _EVAL_339;
  assign _EVAL_68 = _EVAL_204 == 4'h0;
  assign _EVAL_136 = _EVAL_68 | _EVAL_5;
  assign _EVAL_57 = _EVAL_2 == _EVAL_79;
  assign _EVAL_256 = _EVAL_57 | _EVAL_5;
  assign _EVAL_205 = _EVAL_256 == 1'h0;
  assign _EVAL_338 = _EVAL_4 <= 4'h6;
  assign _EVAL_106 = $signed(_EVAL_247) == $signed(33'sh0);
  assign _EVAL_348 = _EVAL_338 & _EVAL_106;
  assign _EVAL_38 = _EVAL_348 | _EVAL_5;
  assign _EVAL_233 = _EVAL_2 ^ 32'h40000000;
  assign _EVAL_155 = {1'b0,$signed(_EVAL_233)};
  assign _EVAL_346 = $signed(_EVAL_155) & $signed(-33'sh2000);
  assign _EVAL_340 = $signed(_EVAL_346);
  assign _EVAL_49 = $signed(_EVAL_340) == $signed(33'sh0);
  assign _EVAL_143 = _EVAL_49 | _EVAL_106;
  assign _EVAL_324 = _EVAL_2 ^ 32'hc000000;
  assign _EVAL_176 = {1'b0,$signed(_EVAL_324)};
  assign _EVAL_91 = $signed(_EVAL_176) & $signed(-33'sh4000000);
  assign _EVAL_284 = $signed(_EVAL_91);
  assign _EVAL_153 = $signed(_EVAL_284) == $signed(33'sh0);
  assign _EVAL_165 = _EVAL_143 | _EVAL_153;
  assign _EVAL_118 = _EVAL_2 ^ 32'h2000000;
  assign _EVAL_342 = {1'b0,$signed(_EVAL_118)};
  assign _EVAL_43 = $signed(_EVAL_342) & $signed(-33'sh10000);
  assign _EVAL_245 = $signed(_EVAL_43);
  assign _EVAL_331 = $signed(_EVAL_245) == $signed(33'sh0);
  assign _EVAL_35 = _EVAL_165 | _EVAL_331;
  assign _EVAL_302 = _EVAL_90 | _EVAL_5;
  assign _EVAL_295 = _EVAL_2 ^ 32'h3000;
  assign _EVAL_343 = {1'b0,$signed(_EVAL_295)};
  assign _EVAL_29 = $signed(_EVAL_343) & $signed(-33'sh1000);
  assign _EVAL_208 = $signed(_EVAL_29);
  assign _EVAL_48 = $signed(_EVAL_208) == $signed(33'sh0);
  assign _EVAL_114 = _EVAL_48 | _EVAL_153;
  assign _EVAL_328 = _EVAL_114 | _EVAL_331;
  assign _EVAL_252 = $signed(_EVAL_218);
  assign _EVAL_251 = $signed(_EVAL_252) == $signed(33'sh0);
  assign _EVAL_194 = _EVAL_328 | _EVAL_251;
  assign _EVAL_200 = _EVAL_2 ^ 32'h1800000;
  assign _EVAL_32 = {1'b0,$signed(_EVAL_200)};
  assign _EVAL_310 = $signed(_EVAL_32) & $signed(-33'sh8000);
  assign _EVAL_235 = $signed(_EVAL_310);
  assign _EVAL_313 = $signed(_EVAL_235) == $signed(33'sh0);
  assign _EVAL_241 = _EVAL_194 | _EVAL_313;
  assign _EVAL_64 = _EVAL_2 ^ 32'h1900000;
  assign _EVAL_39 = {1'b0,$signed(_EVAL_64)};
  assign _EVAL_296 = $signed(_EVAL_39) & $signed(-33'sh2000);
  assign _EVAL_54 = $signed(_EVAL_296);
  assign _EVAL_274 = $signed(_EVAL_54) == $signed(33'sh0);
  assign _EVAL_291 = _EVAL_241 | _EVAL_274;
  assign _EVAL_198 = _EVAL_2 ^ 32'h20000000;
  assign _EVAL_117 = {1'b0,$signed(_EVAL_198)};
  assign _EVAL_327 = $signed(_EVAL_117) & $signed(-33'sh2000);
  assign _EVAL_259 = $signed(_EVAL_327);
  assign _EVAL_253 = $signed(_EVAL_259) == $signed(33'sh0);
  assign _EVAL_123 = _EVAL_291 | _EVAL_253;
  assign _EVAL_132 = _EVAL_13 == _EVAL_192;
  assign _EVAL_44 = _EVAL_132 | _EVAL_5;
  assign _EVAL_263 = _EVAL_271 | _EVAL_268;
  assign _EVAL_344 = _EVAL_263 >> _EVAL_10;
  assign _EVAL_185 = plusarg_reader_out == 32'h0;
  assign _EVAL_174 = _EVAL_124 | _EVAL_185;
  assign _EVAL_169 = _EVAL_150 < plusarg_reader_out;
  assign _EVAL_307 = _EVAL_174 | _EVAL_169;
  assign _EVAL_167 = _EVAL_60[7:2];
  assign _EVAL_184 = ~ _EVAL_17;
  assign _EVAL_170 = _EVAL_184 == 4'h0;
  assign _EVAL_335 = _EVAL_4 <= 4'h8;
  assign _EVAL_248 = _EVAL_335 & _EVAL_48;
  assign _EVAL_161 = _EVAL_248 | _EVAL_5;
  assign _EVAL_58 = _EVAL_161 == 1'h0;
  assign _EVAL_110 = _EVAL_146 & _EVAL_322;
  assign _EVAL_61 = _EVAL_9 <= 3'h4;
  assign _EVAL_228 = _EVAL_61 | _EVAL_5;
  assign _EVAL_267 = _EVAL_228 == 1'h0;
  assign _EVAL_262 = _EVAL_15[2];
  assign _EVAL_89 = _EVAL_262 == 1'h0;
  assign _EVAL_332 = _EVAL_133 - 6'h1;
  assign _EVAL_23 = _EVAL_5 == 1'h0;
  assign _EVAL_303 = _EVAL == 3'h1;
  assign _EVAL_356 = _EVAL_18 & _EVAL_303;
  assign _EVAL_211 = _EVAL_146 | _EVAL_77;
  assign _EVAL_187 = _EVAL_150 + 32'h1;
  assign _EVAL_101 = _EVAL_35 | _EVAL_251;
  assign _EVAL_160 = _EVAL_101 | _EVAL_313;
  assign _EVAL_239 = _EVAL_160 | _EVAL_274;
  assign _EVAL_299 = _EVAL_239 | _EVAL_253;
  assign _EVAL_42 = _EVAL_338 & _EVAL_299;
  assign _EVAL_265 = _EVAL_42 | _EVAL_248;
  assign _EVAL_238 = _EVAL_265 | _EVAL_5;
  assign _EVAL_292 = _EVAL_238 == 1'h0;
  assign _EVAL_227 = _EVAL == 3'h2;
  assign _EVAL_166 = _EVAL_278 == 2'h3;
  assign _EVAL_191 = _EVAL_70 | _EVAL_166;
  assign _EVAL_312 = _EVAL_191 | _EVAL_5;
  assign _EVAL_85 = _EVAL_344[0];
  assign _EVAL_149 = _EVAL_85 | _EVAL_5;
  assign _EVAL_270 = _EVAL_149 == 1'h0;
  assign _EVAL_222 = _EVAL_33 == 6'h0;
  assign _EVAL_243 = _EVAL_312 == 1'h0;
  assign _EVAL_115 = _EVAL_18 & _EVAL_168;
  assign _EVAL_325 = _EVAL_15 == 3'h4;
  assign _EVAL_80 = _EVAL_287 - 6'h1;
  assign _EVAL_99 = _EVAL_15 == _EVAL_156;
  assign _EVAL_280 = _EVAL_99 | _EVAL_5;
  assign _EVAL_285 = _EVAL_280 == 1'h0;
  assign _EVAL_107 = _EVAL_15 == 3'h1;
  assign _EVAL_277 = _EVAL_11 == 1'h0;
  assign _EVAL_289 = _EVAL_277 | _EVAL_5;
  assign _EVAL_37 = _EVAL_289 == 1'h0;
  assign _EVAL_152 = _EVAL_47 | _EVAL_5;
  assign _EVAL_92 = _EVAL_152 == 1'h0;
  assign _EVAL_206 = _EVAL_183 == 1'h0;
  assign _EVAL_314 = _EVAL_7 == 1'h0;
  assign _EVAL_24 = _EVAL_170 | _EVAL_5;
  assign _EVAL_88 = _EVAL_24 == 1'h0;
  assign _EVAL_294 = _EVAL_1 == _EVAL_74;
  assign _EVAL_300 = _EVAL_9 == _EVAL_326;
  assign _EVAL_125 = _EVAL_8 == 1'h0;
  assign _EVAL_31 = _EVAL_125 | _EVAL_7;
  assign _EVAL_223 = _EVAL_31 | _EVAL_5;
  assign _EVAL_351 = _EVAL_9 == 3'h0;
  assign _EVAL_113 = _EVAL_351 | _EVAL_5;
  assign _EVAL_97 = _EVAL_3 >= 4'h2;
  assign _EVAL_286 = _EVAL_9 <= 3'h2;
  assign _EVAL_213 = _EVAL_286 | _EVAL_5;
  assign _EVAL_82 = _EVAL_6 == _EVAL_134;
  assign _EVAL_66 = _EVAL_125 | _EVAL_5;
  assign _EVAL_353 = _EVAL_10[4:3];
  assign _EVAL_272 = _EVAL_353 == 2'h0;
  assign _EVAL_129 = _EVAL_353 == 2'h1;
  assign _EVAL_40 = _EVAL_272 | _EVAL_129;
  assign _EVAL_120 = _EVAL_353 == 2'h2;
  assign _EVAL_104 = _EVAL_40 | _EVAL_120;
  assign _EVAL_93 = _EVAL_113 == 1'h0;
  assign _EVAL_157 = _EVAL_9 != 3'h0;
  assign _EVAL_30 = _EVAL_157 | _EVAL_5;
  assign _EVAL_181 = _EVAL_30 == 1'h0;
  assign _EVAL_100 = _EVAL_45 | _EVAL_5;
  assign _EVAL_20 = _EVAL_15 == 3'h3;
  assign _EVAL_323 = _EVAL_14 & _EVAL_20;
  assign _EVAL_95 = _EVAL_14 & _EVAL_325;
  assign _EVAL_232 = _EVAL_25 - 6'h1;
  assign _EVAL_46 = _EVAL_268 >> _EVAL_6;
  assign _EVAL_330 = _EVAL_46[0];
  assign _EVAL_122 = _EVAL_330 == 1'h0;
  assign _EVAL_109 = _EVAL_122 | _EVAL_5;
  assign _EVAL_242 = _EVAL_109 == 1'h0;
  assign _EVAL_207 = _EVAL_18 & _EVAL_227;
  assign _EVAL_316 = _EVAL_353 == 2'h3;
  assign _EVAL_234 = _EVAL_104 | _EVAL_316;
  assign _EVAL_226 = _EVAL_38 == 1'h0;
  assign _EVAL_27 = _EVAL_294 | _EVAL_5;
  assign _EVAL_345 = _EVAL_66 == 1'h0;
  assign _EVAL_255 = _EVAL_300 | _EVAL_5;
  assign _EVAL_56 = _EVAL_268 | _EVAL_271;
  assign _EVAL_230 = ~ _EVAL_121;
  assign _EVAL_145 = _EVAL_56 & _EVAL_230;
  assign _EVAL_112 = _EVAL <= 3'h6;
  assign _EVAL_315 = _EVAL_112 | _EVAL_5;
  assign _EVAL_336 = _EVAL_234 | _EVAL_5;
  assign _EVAL_279 = _EVAL_136 == 1'h0;
  assign _EVAL_197 = _EVAL_8 == _EVAL_175;
  assign _EVAL_308 = _EVAL_100 == 1'h0;
  assign _EVAL_305 = _EVAL_302 == 1'h0;
  assign _EVAL_81 = _EVAL_82 | _EVAL_5;
  assign _EVAL_34 = _EVAL_81 == 1'h0;
  assign _EVAL_354 = _EVAL_15 == 3'h6;
  assign _EVAL_164 = _EVAL_4 <= 4'h2;
  assign _EVAL_180 = _EVAL_164 & _EVAL_123;
  assign _EVAL_147 = _EVAL_180 | _EVAL_5;
  assign _EVAL_201 = _EVAL_15 == 3'h7;
  assign _EVAL_41 = _EVAL_14 & _EVAL_201;
  assign _EVAL_220 = _EVAL == 3'h4;
  assign _EVAL_269 = _EVAL_18 & _EVAL_220;
  assign _EVAL_21 = _EVAL == 3'h5;
  assign _EVAL_141 = _EVAL_18 & _EVAL_21;
  assign _EVAL_215 = _EVAL_223 == 1'h0;
  assign _EVAL_179 = _EVAL == 3'h0;
  assign _EVAL_333 = _EVAL_1 <= 2'h2;
  assign _EVAL_249 = _EVAL_333 | _EVAL_5;
  assign _EVAL_250 = _EVAL_15 == 3'h5;
  assign _EVAL_71 = _EVAL_314 | _EVAL_5;
  assign _EVAL_283 = _EVAL_71 == 1'h0;
  assign _EVAL_229 = _EVAL == _EVAL_288;
  assign _EVAL_19 = _EVAL_229 | _EVAL_5;
  assign _EVAL_28 = _EVAL_19 == 1'h0;
  assign _EVAL_273 = _EVAL_15 == 3'h0;
  assign _EVAL_73 = _EVAL_307 | _EVAL_5;
  assign _EVAL_51 = _EVAL_14 & _EVAL_306;
  assign _EVAL_203 = _EVAL_33 - 6'h1;
  assign _EVAL_151 = _EVAL_27 == 1'h0;
  assign _EVAL_140 = _EVAL_77 & _EVAL_222;
  assign _EVAL_138 = _EVAL_14 & _EVAL_354;
  assign _EVAL_126 = _EVAL_18 & _EVAL_179;
  assign _EVAL_337 = _EVAL_97 | _EVAL_5;
  assign _EVAL_320 = _EVAL_337 == 1'h0;
  assign _EVAL_22 = _EVAL_14 & _EVAL_107;
  assign _EVAL_231 = _EVAL_197 | _EVAL_5;
  assign _EVAL_72 = _EVAL_231 == 1'h0;
  assign _EVAL_199 = _EVAL_10 == _EVAL_86;
  assign _EVAL_217 = _EVAL_199 | _EVAL_5;
  assign _EVAL_304 = _EVAL_249 == 1'h0;
  assign _EVAL_139 = _EVAL_147 == 1'h0;
  assign _EVAL_193 = _EVAL_213 == 1'h0;
  assign _EVAL_276 = _EVAL_219 == 1'h0;
  assign _EVAL_87 = _EVAL_222 == 1'h0;
  assign _EVAL_94 = _EVAL_18 & _EVAL_87;
  assign _EVAL_69 = _EVAL_14 & _EVAL_273;
  assign _EVAL_319 = _EVAL_217 == 1'h0;
  assign _EVAL_67 = _EVAL_14 & _EVAL_250;
  assign _EVAL_257 = _EVAL_336 == 1'h0;
  assign _EVAL_281 = _EVAL_73 == 1'h0;
  assign _EVAL_189 = _EVAL_44 == 1'h0;
  assign _EVAL_244 = _EVAL_255 == 1'h0;
  assign _EVAL_186 = _EVAL_315 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_25 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_33 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_50 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_74 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_79 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_86 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_133 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_134 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_150 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_156 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_175 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_192 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_268 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_287 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_288 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_326 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_355 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_5) begin
      _EVAL_25 <= 6'h0;
    end else begin
      if (_EVAL_77) begin
        if (_EVAL_210) begin
          if (_EVAL_311) begin
            _EVAL_25 <= _EVAL_171;
          end else begin
            _EVAL_25 <= 6'h0;
          end
        end else begin
          _EVAL_25 <= _EVAL_232;
        end
      end
    end
    if (_EVAL_5) begin
      _EVAL_33 <= 6'h0;
    end else begin
      if (_EVAL_77) begin
        if (_EVAL_222) begin
          if (_EVAL_311) begin
            _EVAL_33 <= _EVAL_171;
          end else begin
            _EVAL_33 <= 6'h0;
          end
        end else begin
          _EVAL_33 <= _EVAL_203;
        end
      end
    end
    if (_EVAL_110) begin
      _EVAL_50 <= _EVAL_4;
    end
    if (_EVAL_140) begin
      _EVAL_74 <= _EVAL_1;
    end
    if (_EVAL_110) begin
      _EVAL_79 <= _EVAL_2;
    end
    if (_EVAL_140) begin
      _EVAL_86 <= _EVAL_10;
    end
    if (_EVAL_5) begin
      _EVAL_133 <= 6'h0;
    end else begin
      if (_EVAL_146) begin
        if (_EVAL_84) begin
          if (_EVAL_89) begin
            _EVAL_133 <= _EVAL_167;
          end else begin
            _EVAL_133 <= 6'h0;
          end
        end else begin
          _EVAL_133 <= _EVAL_332;
        end
      end
    end
    if (_EVAL_110) begin
      _EVAL_134 <= _EVAL_6;
    end
    if (_EVAL_5) begin
      _EVAL_150 <= 32'h0;
    end else begin
      if (_EVAL_211) begin
        _EVAL_150 <= 32'h0;
      end else begin
        _EVAL_150 <= _EVAL_187;
      end
    end
    if (_EVAL_110) begin
      _EVAL_156 <= _EVAL_15;
    end
    if (_EVAL_140) begin
      _EVAL_175 <= _EVAL_8;
    end
    if (_EVAL_140) begin
      _EVAL_192 <= _EVAL_13;
    end
    if (_EVAL_5) begin
      _EVAL_268 <= 32'h0;
    end else begin
      _EVAL_268 <= _EVAL_145;
    end
    if (_EVAL_5) begin
      _EVAL_287 <= 6'h0;
    end else begin
      if (_EVAL_146) begin
        if (_EVAL_322) begin
          if (_EVAL_89) begin
            _EVAL_287 <= _EVAL_167;
          end else begin
            _EVAL_287 <= 6'h0;
          end
        end else begin
          _EVAL_287 <= _EVAL_80;
        end
      end
    end
    if (_EVAL_140) begin
      _EVAL_288 <= _EVAL;
    end
    if (_EVAL_110) begin
      _EVAL_326 <= _EVAL_9;
    end
    if (_EVAL_140) begin
      _EVAL_355 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56dcff8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b7e33e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5b4ab6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98484894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f539813)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee3aef3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d8a1d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(855c639a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a67caa09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52237df5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0e7825f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d2f19af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_320) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b03da70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a662767f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9335e51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_320) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba9bc68d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb9b2bcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9fc8ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(573cf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90c32e52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13b115e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fecb599f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29a1ec80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8cdb8cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(230da648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48bbeddc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39f356a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74c39d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf89f73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f99edd92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62f79ad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a85d862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98a6174d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8f3a520)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(498ad28d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8cec8b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ce1de84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f41c62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff201b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7dbb1bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26c72129)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcb691cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1639e21b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33beb8d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41628c06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(535b1614)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(159627f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a7061a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1301b013)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_320) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f2d13aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e401d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc228f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cb244e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4681931)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c7bd1fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fcc244)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5c7ec30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_345) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b27a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44dc0834)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d809ffd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f410713a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19b271c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9348c238)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_320) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5380a151)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_320) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(646da68f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ca62692)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_345) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c536856)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(808b2f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae3248e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8035fc3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5afaa238)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4d5e8b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a4d20fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e4901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce2c841d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(509795b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2799494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c181062)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_320) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7232c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbbed7db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ba3e40b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1790b822)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(922baba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fe9491c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e992f94e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc95fd3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96e94300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b383cbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
