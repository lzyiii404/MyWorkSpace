//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_83(
  input  [1:0]  _EVAL,
  output [31:0] _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input  [3:0]  _EVAL_10,
  output [3:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  output [2:0]  _EVAL_14,
  output [5:0]  _EVAL_15,
  input         _EVAL_16,
  output [1:0]  _EVAL_17,
  input  [5:0]  _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20
);
  reg [3:0] _EVAL_26 [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] _EVAL_26__EVAL_27_data;
  wire  _EVAL_26__EVAL_27_addr;
  wire [3:0] _EVAL_26__EVAL_28_data;
  wire  _EVAL_26__EVAL_28_addr;
  wire  _EVAL_26__EVAL_28_mask;
  wire  _EVAL_26__EVAL_28_en;
  reg  _EVAL_29 [0:1];
  reg [31:0] _RAND_1;
  wire  _EVAL_29__EVAL_30_data;
  wire  _EVAL_29__EVAL_30_addr;
  wire  _EVAL_29__EVAL_31_data;
  wire  _EVAL_29__EVAL_31_addr;
  wire  _EVAL_29__EVAL_31_mask;
  wire  _EVAL_29__EVAL_31_en;
  reg  _EVAL_34 [0:1];
  reg [31:0] _RAND_2;
  wire  _EVAL_34__EVAL_35_data;
  wire  _EVAL_34__EVAL_35_addr;
  wire  _EVAL_34__EVAL_36_data;
  wire  _EVAL_34__EVAL_36_addr;
  wire  _EVAL_34__EVAL_36_mask;
  wire  _EVAL_34__EVAL_36_en;
  reg [1:0] _EVAL_37 [0:1];
  reg [31:0] _RAND_3;
  wire [1:0] _EVAL_37__EVAL_38_data;
  wire  _EVAL_37__EVAL_38_addr;
  wire [1:0] _EVAL_37__EVAL_39_data;
  wire  _EVAL_37__EVAL_39_addr;
  wire  _EVAL_37__EVAL_39_mask;
  wire  _EVAL_37__EVAL_39_en;
  reg  _EVAL_41 [0:1];
  reg [31:0] _RAND_4;
  wire  _EVAL_41__EVAL_42_data;
  wire  _EVAL_41__EVAL_42_addr;
  wire  _EVAL_41__EVAL_43_data;
  wire  _EVAL_41__EVAL_43_addr;
  wire  _EVAL_41__EVAL_43_mask;
  wire  _EVAL_41__EVAL_43_en;
  reg [31:0] _EVAL_44 [0:1];
  reg [31:0] _RAND_5;
  wire [31:0] _EVAL_44__EVAL_45_data;
  wire  _EVAL_44__EVAL_45_addr;
  wire [31:0] _EVAL_44__EVAL_46_data;
  wire  _EVAL_44__EVAL_46_addr;
  wire  _EVAL_44__EVAL_46_mask;
  wire  _EVAL_44__EVAL_46_en;
  reg [2:0] _EVAL_50 [0:1];
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_50__EVAL_51_data;
  wire  _EVAL_50__EVAL_51_addr;
  wire [2:0] _EVAL_50__EVAL_52_data;
  wire  _EVAL_50__EVAL_52_addr;
  wire  _EVAL_50__EVAL_52_mask;
  wire  _EVAL_50__EVAL_52_en;
  reg [5:0] _EVAL_53 [0:1];
  reg [31:0] _RAND_7;
  wire [5:0] _EVAL_53__EVAL_54_data;
  wire  _EVAL_53__EVAL_54_addr;
  wire [5:0] _EVAL_53__EVAL_55_data;
  wire  _EVAL_53__EVAL_55_addr;
  wire  _EVAL_53__EVAL_55_mask;
  wire  _EVAL_53__EVAL_55_en;
  reg  _EVAL_24;
  reg [31:0] _RAND_8;
  reg  _EVAL_48;
  reg [31:0] _RAND_9;
  reg  _EVAL_59;
  reg [31:0] _RAND_10;
  wire  _EVAL_21;
  wire  _EVAL_57;
  wire  _EVAL_33;
  wire  _EVAL_49;
  wire  _EVAL_32;
  wire  _EVAL_58;
  wire  _EVAL_25;
  wire  _EVAL_61;
  wire  _EVAL_40;
  assign _EVAL_26__EVAL_27_addr = _EVAL_24;
  assign _EVAL_26__EVAL_27_data = _EVAL_26[_EVAL_26__EVAL_27_addr];
  assign _EVAL_26__EVAL_28_data = _EVAL_10;
  assign _EVAL_26__EVAL_28_addr = _EVAL_59;
  assign _EVAL_26__EVAL_28_mask = 1'h1;
  assign _EVAL_26__EVAL_28_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_29__EVAL_30_addr = _EVAL_24;
  assign _EVAL_29__EVAL_30_data = _EVAL_29[_EVAL_29__EVAL_30_addr];
  assign _EVAL_29__EVAL_31_data = _EVAL_20;
  assign _EVAL_29__EVAL_31_addr = _EVAL_59;
  assign _EVAL_29__EVAL_31_mask = 1'h1;
  assign _EVAL_29__EVAL_31_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_34__EVAL_35_addr = _EVAL_24;
  assign _EVAL_34__EVAL_35_data = _EVAL_34[_EVAL_34__EVAL_35_addr];
  assign _EVAL_34__EVAL_36_data = _EVAL_12;
  assign _EVAL_34__EVAL_36_addr = _EVAL_59;
  assign _EVAL_34__EVAL_36_mask = 1'h1;
  assign _EVAL_34__EVAL_36_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_37__EVAL_38_addr = _EVAL_24;
  assign _EVAL_37__EVAL_38_data = _EVAL_37[_EVAL_37__EVAL_38_addr];
  assign _EVAL_37__EVAL_39_data = _EVAL;
  assign _EVAL_37__EVAL_39_addr = _EVAL_59;
  assign _EVAL_37__EVAL_39_mask = 1'h1;
  assign _EVAL_37__EVAL_39_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_41__EVAL_42_addr = _EVAL_24;
  assign _EVAL_41__EVAL_42_data = _EVAL_41[_EVAL_41__EVAL_42_addr];
  assign _EVAL_41__EVAL_43_data = _EVAL_1;
  assign _EVAL_41__EVAL_43_addr = _EVAL_59;
  assign _EVAL_41__EVAL_43_mask = 1'h1;
  assign _EVAL_41__EVAL_43_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_44__EVAL_45_addr = _EVAL_24;
  assign _EVAL_44__EVAL_45_data = _EVAL_44[_EVAL_44__EVAL_45_addr];
  assign _EVAL_44__EVAL_46_data = _EVAL_2;
  assign _EVAL_44__EVAL_46_addr = _EVAL_59;
  assign _EVAL_44__EVAL_46_mask = 1'h1;
  assign _EVAL_44__EVAL_46_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_50__EVAL_51_addr = _EVAL_24;
  assign _EVAL_50__EVAL_51_data = _EVAL_50[_EVAL_50__EVAL_51_addr];
  assign _EVAL_50__EVAL_52_data = _EVAL_7;
  assign _EVAL_50__EVAL_52_addr = _EVAL_59;
  assign _EVAL_50__EVAL_52_mask = 1'h1;
  assign _EVAL_50__EVAL_52_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_53__EVAL_54_addr = _EVAL_24;
  assign _EVAL_53__EVAL_54_data = _EVAL_53[_EVAL_53__EVAL_54_addr];
  assign _EVAL_53__EVAL_55_data = _EVAL_18;
  assign _EVAL_53__EVAL_55_addr = _EVAL_59;
  assign _EVAL_53__EVAL_55_mask = 1'h1;
  assign _EVAL_53__EVAL_55_en = _EVAL_8 & _EVAL_13;
  assign _EVAL_21 = _EVAL_24 + 1'h1;
  assign _EVAL_57 = _EVAL_59 == _EVAL_24;
  assign _EVAL_33 = _EVAL_48 == 1'h0;
  assign _EVAL_49 = _EVAL_57 & _EVAL_33;
  assign _EVAL_32 = _EVAL_57 & _EVAL_48;
  assign _EVAL_58 = _EVAL_8 & _EVAL_13;
  assign _EVAL_25 = _EVAL_6 & _EVAL_4;
  assign _EVAL_61 = _EVAL_58 != _EVAL_25;
  assign _EVAL_40 = _EVAL_59 + 1'h1;
  assign _EVAL_8 = _EVAL_32 == 1'h0;
  assign _EVAL_17 = _EVAL_37__EVAL_38_data;
  assign _EVAL_0 = _EVAL_44__EVAL_45_data;
  assign _EVAL_5 = _EVAL_41__EVAL_42_data;
  assign _EVAL_3 = _EVAL_34__EVAL_35_data;
  assign _EVAL_14 = _EVAL_50__EVAL_51_data;
  assign _EVAL_4 = _EVAL_49 == 1'h0;
  assign _EVAL_15 = _EVAL_53__EVAL_54_data;
  assign _EVAL_9 = _EVAL_29__EVAL_30_data;
  assign _EVAL_11 = _EVAL_26__EVAL_27_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_26[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_29[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_34[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_37[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_41[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_44[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_50[initvar] = _RAND_6[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_53[initvar] = _RAND_7[5:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_24 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_48 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_59 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_16) begin
    if(_EVAL_26__EVAL_28_en & _EVAL_26__EVAL_28_mask) begin
      _EVAL_26[_EVAL_26__EVAL_28_addr] <= _EVAL_26__EVAL_28_data;
    end
    if(_EVAL_29__EVAL_31_en & _EVAL_29__EVAL_31_mask) begin
      _EVAL_29[_EVAL_29__EVAL_31_addr] <= _EVAL_29__EVAL_31_data;
    end
    if(_EVAL_34__EVAL_36_en & _EVAL_34__EVAL_36_mask) begin
      _EVAL_34[_EVAL_34__EVAL_36_addr] <= _EVAL_34__EVAL_36_data;
    end
    if(_EVAL_37__EVAL_39_en & _EVAL_37__EVAL_39_mask) begin
      _EVAL_37[_EVAL_37__EVAL_39_addr] <= _EVAL_37__EVAL_39_data;
    end
    if(_EVAL_41__EVAL_43_en & _EVAL_41__EVAL_43_mask) begin
      _EVAL_41[_EVAL_41__EVAL_43_addr] <= _EVAL_41__EVAL_43_data;
    end
    if(_EVAL_44__EVAL_46_en & _EVAL_44__EVAL_46_mask) begin
      _EVAL_44[_EVAL_44__EVAL_46_addr] <= _EVAL_44__EVAL_46_data;
    end
    if(_EVAL_50__EVAL_52_en & _EVAL_50__EVAL_52_mask) begin
      _EVAL_50[_EVAL_50__EVAL_52_addr] <= _EVAL_50__EVAL_52_data;
    end
    if(_EVAL_53__EVAL_55_en & _EVAL_53__EVAL_55_mask) begin
      _EVAL_53[_EVAL_53__EVAL_55_addr] <= _EVAL_53__EVAL_55_data;
    end
    if (_EVAL_19) begin
      _EVAL_24 <= 1'h0;
    end else begin
      if (_EVAL_25) begin
        _EVAL_24 <= _EVAL_21;
      end
    end
    if (_EVAL_19) begin
      _EVAL_48 <= 1'h0;
    end else begin
      if (_EVAL_61) begin
        _EVAL_48 <= _EVAL_58;
      end
    end
    if (_EVAL_19) begin
      _EVAL_59 <= 1'h0;
    end else begin
      if (_EVAL_58) begin
        _EVAL_59 <= _EVAL_40;
      end
    end
  end
endmodule
