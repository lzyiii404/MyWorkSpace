//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_56(
  output [31:0] _EVAL,
  input  [3:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [2:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  output [31:0] _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  output [31:0] _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  input  [1:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  input  [31:0] _EVAL_22,
  output [3:0]  _EVAL_23,
  output        _EVAL_24,
  output [3:0]  _EVAL_25,
  input  [3:0]  _EVAL_26,
  output [1:0]  _EVAL_27,
  output        _EVAL_28,
  input  [31:0] _EVAL_29,
  input  [2:0]  _EVAL_30,
  output [3:0]  _EVAL_31,
  output        _EVAL_32
);
  assign _EVAL_13 = _EVAL_2;
  assign _EVAL = _EVAL_22;
  assign _EVAL_21 = _EVAL_30;
  assign _EVAL_25 = _EVAL_1;
  assign _EVAL_32 = _EVAL_18;
  assign _EVAL_31 = _EVAL_0;
  assign _EVAL_17 = _EVAL_12;
  assign _EVAL_4 = _EVAL_3;
  assign _EVAL_28 = _EVAL_8;
  assign _EVAL_14 = _EVAL_5;
  assign _EVAL_19 = _EVAL_7;
  assign _EVAL_10 = _EVAL_29;
  assign _EVAL_24 = _EVAL_15;
  assign _EVAL_27 = _EVAL_20;
  assign _EVAL_9 = _EVAL_16;
  assign _EVAL_23 = _EVAL_26;
endmodule
