//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_266(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  output [2:0]  _EVAL_5,
  output        _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [7:0]  _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [63:0] _EVAL_11,
  output        _EVAL_12,
  output [2:0]  _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  output [63:0] _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  output [31:0] _EVAL_22,
  output [7:0]  _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [3:0]  _EVAL_26,
  output        _EVAL_27,
  output [1:0]  _EVAL_28,
  output [3:0]  _EVAL_29,
  input         _EVAL_30,
  output [2:0]  _EVAL_31,
  input  [1:0]  _EVAL_32,
  output        _EVAL_33,
  output [2:0]  _EVAL_34,
  input  [3:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  input  [31:0] _EVAL_40,
  output [3:0]  _EVAL_41,
  input  [63:0] _EVAL_42,
  output [63:0] _EVAL_43,
  input         _EVAL_44,
  output [31:0] _EVAL_45,
  output        _EVAL_46,
  output        _EVAL_47,
  input         _EVAL_48,
  output [1:0]  _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  output        _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  output [3:0]  _EVAL_57,
  input  [3:0]  _EVAL_58,
  output [31:0] _EVAL_59,
  input  [3:0]  _EVAL_60,
  input  [2:0]  _EVAL_61,
  output [3:0]  _EVAL_62,
  output        _EVAL_63,
  output [63:0] _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  input  [2:0]  _EVAL_67,
  input  [63:0] _EVAL_68,
  output [3:0]  _EVAL_69,
  output        _EVAL_70,
  input  [2:0]  _EVAL_71,
  input         _EVAL_72
);
  assign _EVAL_27 = _EVAL_53;
  assign _EVAL_70 = _EVAL_30;
  assign _EVAL_29 = _EVAL_15;
  assign _EVAL_34 = _EVAL_71;
  assign _EVAL_66 = _EVAL_21;
  assign _EVAL = _EVAL_19;
  assign _EVAL_5 = _EVAL_7;
  assign _EVAL_6 = _EVAL_56;
  assign _EVAL_63 = _EVAL_55;
  assign _EVAL_52 = _EVAL_54;
  assign _EVAL_23 = _EVAL_9;
  assign _EVAL_57 = _EVAL_58;
  assign _EVAL_26 = _EVAL_35;
  assign _EVAL_17 = _EVAL_68;
  assign _EVAL_64 = _EVAL_42;
  assign _EVAL_22 = _EVAL_2;
  assign _EVAL_45 = _EVAL_0;
  assign _EVAL_36 = _EVAL_67;
  assign _EVAL_13 = _EVAL_61;
  assign _EVAL_65 = _EVAL_48;
  assign _EVAL_33 = _EVAL_51;
  assign _EVAL_31 = _EVAL_25;
  assign _EVAL_46 = _EVAL_38;
  assign _EVAL_20 = _EVAL_1;
  assign _EVAL_12 = _EVAL_44;
  assign _EVAL_43 = _EVAL_11;
  assign _EVAL_4 = _EVAL_14;
  assign _EVAL_49 = _EVAL_10;
  assign _EVAL_62 = _EVAL_8;
  assign _EVAL_69 = _EVAL_60;
  assign _EVAL_41 = _EVAL_16;
  assign _EVAL_24 = _EVAL_3;
  assign _EVAL_59 = _EVAL_40;
  assign _EVAL_39 = _EVAL_50;
  assign _EVAL_47 = _EVAL_18;
  assign _EVAL_28 = _EVAL_32;
endmodule
