//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_43(
  input         _EVAL,
  output [3:0]  _EVAL_0,
  output [6:0]  _EVAL_1,
  output [3:0]  _EVAL_2,
  input  [6:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  output [1:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  output [6:0]  _EVAL_9,
  input  [63:0] _EVAL_10,
  output [63:0] _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  output [2:0]  _EVAL_14,
  input  [7:0]  _EVAL_15,
  input         _EVAL_16,
  output [2:0]  _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  output [29:0] _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  output        _EVAL_23,
  input  [31:0] _EVAL_24,
  input  [1:0]  _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [29:0] _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  output [31:0] _EVAL_32,
  input  [3:0]  _EVAL_33,
  input  [6:0]  _EVAL_34,
  output        _EVAL_35,
  output [3:0]  _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  output        _EVAL_39,
  input  [2:0]  _EVAL_40
);
  wire  Repeater__EVAL;
  wire  Repeater__EVAL_0;
  wire [2:0] Repeater__EVAL_1;
  wire  Repeater__EVAL_2;
  wire  Repeater__EVAL_3;
  wire [6:0] Repeater__EVAL_4;
  wire  Repeater__EVAL_5;
  wire [2:0] Repeater__EVAL_6;
  wire [29:0] Repeater__EVAL_7;
  wire [3:0] Repeater__EVAL_8;
  wire [63:0] Repeater__EVAL_9;
  wire [63:0] Repeater__EVAL_10;
  wire [2:0] Repeater__EVAL_11;
  wire [7:0] Repeater__EVAL_12;
  wire [3:0] Repeater__EVAL_13;
  wire [29:0] Repeater__EVAL_14;
  wire  Repeater__EVAL_15;
  wire  Repeater__EVAL_16;
  wire  Repeater__EVAL_17;
  wire [6:0] Repeater__EVAL_18;
  wire [2:0] Repeater__EVAL_19;
  wire  Repeater__EVAL_20;
  wire [7:0] Repeater__EVAL_21;
  reg [31:0] _EVAL_65;
  reg [31:0] _RAND_0;
  reg  _EVAL_70;
  reg [31:0] _RAND_1;
  reg  _EVAL_72;
  reg [31:0] _RAND_2;
  reg  _EVAL_91;
  reg [31:0] _RAND_3;
  wire [29:0] _EVAL_60;
  wire  _EVAL_83;
  wire  _EVAL_79;
  wire [3:0] _EVAL_76;
  wire [31:0] _EVAL_90;
  wire [31:0] _EVAL_78;
  wire [63:0] _EVAL_86;
  wire [31:0] _EVAL_54;
  wire  _EVAL_77;
  wire [17:0] _EVAL_74;
  wire [2:0] _EVAL_41;
  wire [2:0] _EVAL_88;
  wire  _EVAL_75;
  wire  _EVAL_89;
  wire  _EVAL_64;
  wire  _EVAL_61;
  wire  _EVAL_68;
  wire  _EVAL_57;
  wire  _EVAL_47;
  wire [2:0] _EVAL_87;
  wire  _EVAL_51;
  wire  _EVAL_82;
  wire  _EVAL_84;
  wire [17:0] _EVAL_66;
  wire [2:0] _EVAL_94;
  wire [2:0] _EVAL_71;
  wire  _EVAL_49;
  wire  _EVAL_52;
  wire  _EVAL_93;
  wire  _EVAL_85;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_48;
  wire [31:0] _EVAL_50;
  wire [31:0] _EVAL_59;
  wire  _EVAL_81;
  wire  _EVAL_62;
  wire  _EVAL_73;
  wire [7:0] _EVAL_58;
  wire [3:0] _EVAL_63;
  wire [3:0] _EVAL_69;
  SiFive__EVAL_42 Repeater (
    ._EVAL(Repeater__EVAL),
    ._EVAL_0(Repeater__EVAL_0),
    ._EVAL_1(Repeater__EVAL_1),
    ._EVAL_2(Repeater__EVAL_2),
    ._EVAL_3(Repeater__EVAL_3),
    ._EVAL_4(Repeater__EVAL_4),
    ._EVAL_5(Repeater__EVAL_5),
    ._EVAL_6(Repeater__EVAL_6),
    ._EVAL_7(Repeater__EVAL_7),
    ._EVAL_8(Repeater__EVAL_8),
    ._EVAL_9(Repeater__EVAL_9),
    ._EVAL_10(Repeater__EVAL_10),
    ._EVAL_11(Repeater__EVAL_11),
    ._EVAL_12(Repeater__EVAL_12),
    ._EVAL_13(Repeater__EVAL_13),
    ._EVAL_14(Repeater__EVAL_14),
    ._EVAL_15(Repeater__EVAL_15),
    ._EVAL_16(Repeater__EVAL_16),
    ._EVAL_17(Repeater__EVAL_17),
    ._EVAL_18(Repeater__EVAL_18),
    ._EVAL_19(Repeater__EVAL_19),
    ._EVAL_20(Repeater__EVAL_20),
    ._EVAL_21(Repeater__EVAL_21)
  );
  assign _EVAL_60 = Repeater__EVAL_14;
  assign _EVAL_83 = _EVAL_60[2];
  assign _EVAL_79 = _EVAL_83 | _EVAL_91;
  assign _EVAL_76 = Repeater__EVAL_13;
  assign _EVAL_90 = Repeater__EVAL_10[63:32];
  assign _EVAL_78 = _EVAL_10[31:0];
  assign _EVAL_86 = {_EVAL_90,_EVAL_78};
  assign _EVAL_54 = _EVAL_86[31:0];
  assign _EVAL_77 = Repeater__EVAL_2;
  assign _EVAL_74 = 18'h7 << _EVAL_33;
  assign _EVAL_41 = _EVAL_74[2:0];
  assign _EVAL_88 = ~ _EVAL_41;
  assign _EVAL_75 = _EVAL_88[2:2];
  assign _EVAL_89 = _EVAL_72 == _EVAL_75;
  assign _EVAL_64 = _EVAL_40[0];
  assign _EVAL_61 = _EVAL_64 == 1'h0;
  assign _EVAL_68 = _EVAL_89 | _EVAL_61;
  assign _EVAL_57 = _EVAL_68 == 1'h0;
  assign _EVAL_47 = _EVAL | _EVAL_57;
  assign _EVAL_87 = Repeater__EVAL_11;
  assign _EVAL_51 = _EVAL_87[2];
  assign _EVAL_82 = _EVAL_12 | _EVAL_70;
  assign _EVAL_84 = _EVAL_6 & _EVAL_77;
  assign _EVAL_66 = 18'h7 << _EVAL_76;
  assign _EVAL_94 = _EVAL_66[2:0];
  assign _EVAL_71 = ~ _EVAL_94;
  assign _EVAL_49 = _EVAL_71[2:2];
  assign _EVAL_52 = _EVAL_91 == _EVAL_49;
  assign _EVAL_93 = _EVAL_51 == 1'h0;
  assign _EVAL_85 = _EVAL_93 == 1'h0;
  assign _EVAL_43 = _EVAL_52 | _EVAL_85;
  assign _EVAL_44 = _EVAL_91 + 1'h1;
  assign _EVAL_46 = _EVAL_72 & _EVAL_75;
  assign _EVAL_48 = _EVAL_46 == 1'h0;
  assign _EVAL_50 = _EVAL_48 ? _EVAL_24 : _EVAL_65;
  assign _EVAL_59 = _EVAL_86[63:32];
  assign _EVAL_81 = _EVAL_47 & _EVAL_26;
  assign _EVAL_62 = _EVAL_72 + 1'h1;
  assign _EVAL_73 = _EVAL_81 & _EVAL_57;
  assign _EVAL_58 = Repeater__EVAL_12;
  assign _EVAL_63 = _EVAL_58[3:0];
  assign _EVAL_69 = _EVAL_58[7:4];
  assign _EVAL_32 = _EVAL_79 ? _EVAL_59 : _EVAL_54;
  assign _EVAL_9 = _EVAL_34;
  assign Repeater__EVAL_16 = _EVAL_16;
  assign _EVAL_5 = _EVAL_25;
  assign _EVAL_23 = Repeater__EVAL_15;
  assign _EVAL_39 = _EVAL_29;
  assign _EVAL_17 = Repeater__EVAL_11;
  assign Repeater__EVAL_5 = _EVAL_43 == 1'h0;
  assign Repeater__EVAL_4 = _EVAL_3;
  assign _EVAL_14 = Repeater__EVAL_6;
  assign Repeater__EVAL_8 = _EVAL_4;
  assign _EVAL_0 = _EVAL_33;
  assign Repeater__EVAL = _EVAL_7;
  assign _EVAL_37 = _EVAL_12 | _EVAL_70;
  assign Repeater__EVAL_20 = _EVAL_8;
  assign Repeater__EVAL_3 = _EVAL_31;
  assign _EVAL_11 = {_EVAL_24,_EVAL_50};
  assign _EVAL_30 = _EVAL_27;
  assign Repeater__EVAL_7 = _EVAL_28;
  assign Repeater__EVAL_1 = _EVAL_13;
  assign _EVAL_20 = Repeater__EVAL_14;
  assign _EVAL_36 = Repeater__EVAL_13;
  assign _EVAL_1 = Repeater__EVAL_18;
  assign _EVAL_38 = Repeater__EVAL_17;
  assign Repeater__EVAL_21 = _EVAL_15;
  assign _EVAL_2 = _EVAL_79 ? _EVAL_69 : _EVAL_63;
  assign _EVAL_18 = _EVAL | _EVAL_57;
  assign Repeater__EVAL_9 = _EVAL_10;
  assign Repeater__EVAL_19 = _EVAL_21;
  assign _EVAL_19 = Repeater__EVAL_2;
  assign _EVAL_22 = _EVAL_40;
  assign _EVAL_35 = _EVAL_26 & _EVAL_68;
  assign Repeater__EVAL_0 = _EVAL_6;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_65 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_70 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_72 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_91 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_7) begin
    if (_EVAL_73) begin
      if (_EVAL_48) begin
        _EVAL_65 <= _EVAL_24;
      end
    end
    if (_EVAL_31) begin
      _EVAL_70 <= 1'h0;
    end else begin
      if (_EVAL_81) begin
        if (_EVAL_68) begin
          _EVAL_70 <= 1'h0;
        end else begin
          _EVAL_70 <= _EVAL_82;
        end
      end
    end
    if (_EVAL_31) begin
      _EVAL_72 <= 1'h0;
    end else begin
      if (_EVAL_81) begin
        if (_EVAL_68) begin
          _EVAL_72 <= 1'h0;
        end else begin
          _EVAL_72 <= _EVAL_62;
        end
      end
    end
    if (_EVAL_31) begin
      _EVAL_91 <= 1'h0;
    end else begin
      if (_EVAL_84) begin
        if (_EVAL_43) begin
          _EVAL_91 <= 1'h0;
        end else begin
          _EVAL_91 <= _EVAL_44;
        end
      end
    end
  end
endmodule
