//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_259(
  output        _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [29:0] _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output [5:0]  _EVAL_17,
  input         _EVAL_18,
  input  [29:0] _EVAL_19,
  input  [31:0] _EVAL_20,
  input         _EVAL_21,
  input  [31:0] _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input         _EVAL_25,
  input  [29:0] _EVAL_26,
  input         _EVAL_27,
  input  [29:0] _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  output [1:0]  _EVAL_34,
  output        _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input  [63:0] _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  output [2:0]  _EVAL_41,
  output        _EVAL_42,
  output        _EVAL_43,
  output        _EVAL_44,
  input         _EVAL_45,
  output [7:0]  _EVAL_46,
  output [5:0]  _EVAL_47,
  output        _EVAL_48,
  input  [1:0]  _EVAL_49,
  output [31:0] _EVAL_50,
  input  [1:0]  _EVAL_51,
  input  [31:0] _EVAL_52,
  input  [1:0]  _EVAL_53,
  input         _EVAL_54,
  input  [31:0] _EVAL_55,
  input  [1:0]  _EVAL_56,
  output [2:0]  _EVAL_57,
  input         _EVAL_58,
  output [63:0] _EVAL_59,
  input  [31:0] _EVAL_60,
  output        _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  output        _EVAL_64,
  output [3:0]  _EVAL_65,
  input  [2:0]  _EVAL_66,
  input  [29:0] _EVAL_67,
  output [31:0] _EVAL_68,
  input  [31:0] _EVAL_69,
  output        _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  output [31:0] _EVAL_73,
  input         _EVAL_74,
  output        _EVAL_75,
  output        _EVAL_76,
  input  [3:0]  _EVAL_77,
  input         _EVAL_78,
  input  [31:0] _EVAL_79,
  output [3:0]  _EVAL_80,
  input         _EVAL_81,
  output        _EVAL_82,
  input         _EVAL_83,
  output        _EVAL_84,
  input  [1:0]  _EVAL_85,
  input         _EVAL_86,
  input         _EVAL_87,
  input         _EVAL_88,
  input  [1:0]  _EVAL_89,
  input         _EVAL_90,
  output        _EVAL_91,
  output [63:0] _EVAL_92,
  input  [1:0]  _EVAL_93,
  output [31:0] _EVAL_94,
  input  [29:0] _EVAL_95,
  input         _EVAL_96,
  input         _EVAL_97,
  input         _EVAL_98,
  input  [3:0]  _EVAL_99,
  output        _EVAL_100,
  input         _EVAL_101,
  input  [29:0] _EVAL_102,
  output        _EVAL_103,
  input         _EVAL_104,
  output        _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  output        _EVAL_108,
  input  [31:0] _EVAL_109,
  output        _EVAL_110,
  output        _EVAL_111,
  input  [1:0]  _EVAL_112,
  input         _EVAL_113,
  input  [1:0]  _EVAL_114,
  input         _EVAL_115,
  input  [31:0] _EVAL_116,
  input         _EVAL_117,
  input         _EVAL_118,
  output [4:0]  _EVAL_119,
  input         _EVAL_120,
  output [31:0] _EVAL_121,
  input  [31:0] _EVAL_122,
  output [2:0]  _EVAL_123,
  input         _EVAL_124,
  input  [31:0] _EVAL_125,
  output [2:0]  _EVAL_126,
  output [31:0] _EVAL_127,
  output        _EVAL_128,
  output        _EVAL_129,
  output [31:0] _EVAL_130,
  input         _EVAL_131,
  input  [1:0]  _EVAL_132,
  input  [5:0]  _EVAL_133,
  output [2:0]  _EVAL_134,
  input  [4:0]  _EVAL_135,
  output [31:0] _EVAL_136,
  input         _EVAL_137,
  output        _EVAL_138,
  input  [31:0] _EVAL_139,
  input  [1:0]  _EVAL_140,
  input  [1:0]  _EVAL_141,
  input         _EVAL_142,
  output        _EVAL_143,
  input         _EVAL_144,
  input         _EVAL_145,
  output        _EVAL_146,
  output        _EVAL_147,
  input         _EVAL_148,
  output        _EVAL_149,
  input  [29:0] _EVAL_150
);
  wire [63:0] data__EVAL;
  wire  data__EVAL_0;
  wire [63:0] data__EVAL_1;
  wire [3:0] data__EVAL_2;
  wire  data__EVAL_3;
  wire [11:0] data__EVAL_4;
  wire [63:0] data__EVAL_5;
  wire [3:0] data__EVAL_6;
  wire [63:0] data__EVAL_7;
  wire [63:0] data__EVAL_8;
  wire [1:0] data__EVAL_9;
  wire  data__EVAL_10;
  wire  dcache_clock_gate_in;
  wire  dcache_clock_gate_en;
  wire  dcache_clock_gate_out;
  wire  tlb__EVAL;
  wire  tlb__EVAL_0;
  wire  tlb__EVAL_1;
  wire [1:0] tlb__EVAL_2;
  wire [31:0] tlb__EVAL_3;
  wire [29:0] tlb__EVAL_4;
  wire  tlb__EVAL_5;
  wire  tlb__EVAL_6;
  wire  tlb__EVAL_7;
  wire  tlb__EVAL_8;
  wire  tlb__EVAL_9;
  wire  tlb__EVAL_10;
  wire  tlb__EVAL_11;
  wire [1:0] tlb__EVAL_12;
  wire [31:0] tlb__EVAL_13;
  wire  tlb__EVAL_14;
  wire [29:0] tlb__EVAL_15;
  wire  tlb__EVAL_16;
  wire [29:0] tlb__EVAL_17;
  wire  tlb__EVAL_18;
  wire [29:0] tlb__EVAL_19;
  wire [1:0] tlb__EVAL_20;
  wire [31:0] tlb__EVAL_21;
  wire  tlb__EVAL_22;
  wire  tlb__EVAL_23;
  wire [31:0] tlb__EVAL_24;
  wire [1:0] tlb__EVAL_25;
  wire  tlb__EVAL_26;
  wire [31:0] tlb__EVAL_27;
  wire [29:0] tlb__EVAL_28;
  wire [31:0] tlb__EVAL_29;
  wire  tlb__EVAL_30;
  wire  tlb__EVAL_31;
  wire [1:0] tlb__EVAL_32;
  wire [31:0] tlb__EVAL_33;
  wire  tlb__EVAL_34;
  wire [29:0] tlb__EVAL_35;
  wire  tlb__EVAL_36;
  wire  tlb__EVAL_37;
  wire [31:0] tlb__EVAL_38;
  wire  tlb__EVAL_39;
  wire [1:0] tlb__EVAL_40;
  wire  tlb__EVAL_41;
  wire  tlb__EVAL_42;
  wire  tlb__EVAL_43;
  wire  tlb__EVAL_44;
  wire  tlb__EVAL_45;
  wire  tlb__EVAL_46;
  wire  tlb__EVAL_47;
  wire  tlb__EVAL_48;
  wire [4:0] tlb__EVAL_49;
  wire [29:0] tlb__EVAL_50;
  wire  tlb__EVAL_51;
  wire  tlb__EVAL_52;
  wire [1:0] tlb__EVAL_53;
  wire  tlb__EVAL_54;
  wire  tlb__EVAL_55;
  wire [1:0] tlb__EVAL_56;
  wire  tlb__EVAL_57;
  wire  tlb__EVAL_58;
  wire [31:0] tlb__EVAL_59;
  wire  tlb__EVAL_60;
  wire  tlb__EVAL_61;
  wire  tlb__EVAL_62;
  wire [1:0] tlb__EVAL_63;
  wire  tlb__EVAL_64;
  wire [29:0] tlb__EVAL_65;
  wire [31:0] tlb__EVAL_66;
  wire  tlb__EVAL_67;
  wire  tlb__EVAL_68;
  wire  tlb__EVAL_69;
  wire  tlb__EVAL_70;
  wire [1:0] tlb__EVAL_71;
  wire  q__EVAL;
  wire  q__EVAL_0;
  wire [63:0] q__EVAL_1;
  wire [2:0] q__EVAL_2;
  wire [3:0] q__EVAL_3;
  wire  q__EVAL_4;
  wire [2:0] q__EVAL_5;
  wire  q__EVAL_6;
  wire [7:0] q__EVAL_7;
  wire  q__EVAL_8;
  wire [2:0] q__EVAL_9;
  wire [7:0] q__EVAL_10;
  wire [2:0] q__EVAL_11;
  wire  q__EVAL_12;
  wire [2:0] q__EVAL_13;
  wire [31:0] q__EVAL_14;
  wire [3:0] q__EVAL_15;
  wire  q__EVAL_16;
  wire [2:0] q__EVAL_17;
  wire [31:0] q__EVAL_18;
  wire [63:0] q__EVAL_19;
  wire  MaxPeriodFibonacciLFSR__EVAL;
  wire  MaxPeriodFibonacciLFSR__EVAL_0;
  wire  MaxPeriodFibonacciLFSR__EVAL_1;
  wire  MaxPeriodFibonacciLFSR__EVAL_2;
  wire  MaxPeriodFibonacciLFSR__EVAL_3;
  wire  MaxPeriodFibonacciLFSR__EVAL_4;
  wire  MaxPeriodFibonacciLFSR__EVAL_5;
  wire  MaxPeriodFibonacciLFSR__EVAL_6;
  wire  MaxPeriodFibonacciLFSR__EVAL_7;
  wire  MaxPeriodFibonacciLFSR__EVAL_8;
  wire  MaxPeriodFibonacciLFSR__EVAL_9;
  wire  MaxPeriodFibonacciLFSR__EVAL_10;
  wire  MaxPeriodFibonacciLFSR__EVAL_11;
  wire  MaxPeriodFibonacciLFSR__EVAL_12;
  wire  MaxPeriodFibonacciLFSR__EVAL_13;
  wire  MaxPeriodFibonacciLFSR__EVAL_14;
  wire  MaxPeriodFibonacciLFSR__EVAL_15;
  wire  MaxPeriodFibonacciLFSR__EVAL_16;
  wire  MaxPeriodFibonacciLFSR__EVAL_17;
  wire [3:0] amoalu__EVAL;
  wire [31:0] amoalu__EVAL_0;
  wire [4:0] amoalu__EVAL_1;
  wire [31:0] amoalu__EVAL_2;
  wire [31:0] amoalu__EVAL_3;
  wire [21:0] tag_array__EVAL;
  wire  tag_array__EVAL_0;
  wire [21:0] tag_array__EVAL_1;
  wire  tag_array__EVAL_2;
  wire [21:0] tag_array__EVAL_3;
  wire [21:0] tag_array__EVAL_4;
  wire [21:0] tag_array__EVAL_5;
  wire [21:0] tag_array__EVAL_6;
  wire [5:0] tag_array__EVAL_7;
  wire [21:0] tag_array__EVAL_8;
  wire  tag_array__EVAL_9;
  wire  tag_array__EVAL_10;
  wire [21:0] tag_array__EVAL_11;
  wire  tag_array__EVAL_12;
  wire  tag_array__EVAL_13;
  wire  tag_array__EVAL_14;
  reg [31:0] _EVAL_155;
  reg [31:0] _RAND_0;
  reg [1:0] _EVAL_162;
  reg [31:0] _RAND_1;
  reg  _EVAL_165;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_190;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_204;
  reg [31:0] _RAND_4;
  reg [1:0] _EVAL_211;
  reg [31:0] _RAND_5;
  reg [4:0] _EVAL_239;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_254;
  reg [31:0] _RAND_7;
  reg  _EVAL_263;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_277;
  reg [31:0] _RAND_9;
  reg [31:0] _EVAL_280;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_291;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_293;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_300;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_320;
  reg [31:0] _RAND_14;
  reg  _EVAL_322;
  reg [31:0] _RAND_15;
  reg  _EVAL_332;
  reg [31:0] _RAND_16;
  reg  _EVAL_341;
  reg [31:0] _RAND_17;
  reg  _EVAL_356;
  reg [31:0] _RAND_18;
  reg  _EVAL_357;
  reg [31:0] _RAND_19;
  reg [31:0] _EVAL_359;
  reg [31:0] _RAND_20;
  reg [31:0] _EVAL_367;
  reg [31:0] _RAND_21;
  reg  _EVAL_375;
  reg [31:0] _RAND_22;
  reg  _EVAL_376;
  reg [31:0] _RAND_23;
  reg  _EVAL_377;
  reg [31:0] _RAND_24;
  reg [31:0] _EVAL_387;
  reg [31:0] _RAND_25;
  reg [31:0] _EVAL_389;
  reg [31:0] _RAND_26;
  reg [3:0] _EVAL_393;
  reg [31:0] _RAND_27;
  reg [2:0] _EVAL_396;
  reg [31:0] _RAND_28;
  reg  _EVAL_401;
  reg [31:0] _RAND_29;
  reg [31:0] _EVAL_433;
  reg [31:0] _RAND_30;
  reg [4:0] _EVAL_451;
  reg [31:0] _RAND_31;
  reg [3:0] _EVAL_461;
  reg [31:0] _RAND_32;
  reg  _EVAL_477;
  reg [31:0] _RAND_33;
  reg  _EVAL_487;
  reg [31:0] _RAND_34;
  reg [4:0] _EVAL_502;
  reg [31:0] _RAND_35;
  reg [7:0] _EVAL_506;
  reg [31:0] _RAND_36;
  reg  _EVAL_526;
  reg [31:0] _RAND_37;
  reg  _EVAL_541;
  reg [31:0] _RAND_38;
  reg [19:0] _EVAL_549;
  reg [31:0] _RAND_39;
  reg  _EVAL_559;
  reg [31:0] _RAND_40;
  reg  _EVAL_588;
  reg [31:0] _RAND_41;
  reg [1:0] _EVAL_598;
  reg [31:0] _RAND_42;
  reg  _EVAL_611;
  reg [31:0] _RAND_43;
  reg  _EVAL_612;
  reg [31:0] _RAND_44;
  reg  _EVAL_613;
  reg [31:0] _RAND_45;
  reg  _EVAL_614;
  reg [31:0] _RAND_46;
  reg [31:0] _EVAL_629;
  reg [31:0] _RAND_47;
  reg  _EVAL_631;
  reg [31:0] _RAND_48;
  reg [25:0] _EVAL_632;
  reg [31:0] _RAND_49;
  reg  _EVAL_655;
  reg [31:0] _RAND_50;
  reg [4:0] _EVAL_659;
  reg [31:0] _RAND_51;
  reg  _EVAL_700;
  reg [31:0] _RAND_52;
  reg [7:0] _EVAL_730;
  reg [31:0] _RAND_53;
  reg  _EVAL_732;
  reg [31:0] _RAND_54;
  reg [1:0] _EVAL_746;
  reg [31:0] _RAND_55;
  reg [31:0] _EVAL_753;
  reg [31:0] _RAND_56;
  reg  _EVAL_759;
  reg [31:0] _RAND_57;
  reg [7:0] _EVAL_763;
  reg [31:0] _RAND_58;
  reg [4:0] _EVAL_769;
  reg [31:0] _RAND_59;
  reg  _EVAL_800;
  reg [31:0] _RAND_60;
  reg [31:0] _EVAL_801;
  reg [31:0] _RAND_61;
  reg [3:0] _EVAL_831;
  reg [31:0] _RAND_62;
  reg [31:0] _EVAL_846;
  reg [31:0] _RAND_63;
  reg  _EVAL_872;
  reg [31:0] _RAND_64;
  reg [4:0] _EVAL_874;
  reg [31:0] _RAND_65;
  reg [6:0] _EVAL_893;
  reg [31:0] _RAND_66;
  reg  _EVAL_907;
  reg [31:0] _RAND_67;
  reg  _EVAL_918;
  reg [31:0] _RAND_68;
  reg  _EVAL_924;
  reg [31:0] _RAND_69;
  reg  _EVAL_926;
  reg [31:0] _RAND_70;
  reg  _EVAL_937;
  reg [31:0] _RAND_71;
  reg [1:0] _EVAL_951;
  reg [31:0] _RAND_72;
  reg [1:0] _EVAL_981;
  reg [31:0] _RAND_73;
  reg [31:0] _EVAL_982;
  reg [31:0] _RAND_74;
  reg  _EVAL_1001;
  reg [31:0] _RAND_75;
  reg [2:0] _EVAL_1032;
  reg [31:0] _RAND_76;
  reg  _EVAL_1049;
  reg [31:0] _RAND_77;
  reg [1:0] _EVAL_1058;
  reg [31:0] _RAND_78;
  reg [7:0] _EVAL_1060;
  reg [31:0] _RAND_79;
  reg [31:0] _EVAL_1096;
  reg [31:0] _RAND_80;
  reg  _EVAL_1100;
  reg [31:0] _RAND_81;
  reg  _EVAL_1104;
  reg [31:0] _RAND_82;
  reg [31:0] _EVAL_1107;
  reg [31:0] _RAND_83;
  reg  _EVAL_1109;
  reg [31:0] _RAND_84;
  reg [3:0] _EVAL_1121;
  reg [31:0] _RAND_85;
  reg  _EVAL_1122;
  reg [31:0] _RAND_86;
  reg [4:0] _EVAL_1134;
  reg [31:0] _RAND_87;
  reg [1:0] _EVAL_1135;
  reg [31:0] _RAND_88;
  reg  _EVAL_1140;
  reg [31:0] _RAND_89;
  reg [31:0] _EVAL_1172;
  reg [31:0] _RAND_90;
  reg [7:0] _EVAL_1195;
  reg [31:0] _RAND_91;
  reg [1:0] _EVAL_1200;
  reg [31:0] _RAND_92;
  reg [5:0] _EVAL_1213;
  reg [31:0] _RAND_93;
  reg [4:0] _EVAL_1225;
  reg [31:0] _RAND_94;
  reg [5:0] _EVAL_1240;
  reg [31:0] _RAND_95;
  reg  _EVAL_1252;
  reg [31:0] _RAND_96;
  reg  _EVAL_1269;
  reg [31:0] _RAND_97;
  reg  _EVAL_1271;
  reg [31:0] _RAND_98;
  reg  _EVAL_1278;
  reg [31:0] _RAND_99;
  reg [5:0] _EVAL_1300;
  reg [31:0] _RAND_100;
  reg [1:0] _EVAL_1316;
  reg [31:0] _RAND_101;
  reg  _EVAL_1319;
  reg [31:0] _RAND_102;
  reg [4:0] _EVAL_1325;
  reg [31:0] _RAND_103;
  reg  _EVAL_1350;
  reg [31:0] _RAND_104;
  reg [3:0] _EVAL_1366;
  reg [31:0] _RAND_105;
  reg [31:0] _EVAL_1370;
  reg [31:0] _RAND_106;
  reg [1:0] _EVAL_1373;
  reg [31:0] _RAND_107;
  reg  _EVAL_1374;
  reg [31:0] _RAND_108;
  reg [5:0] _EVAL_1387;
  reg [31:0] _RAND_109;
  reg [5:0] _EVAL_1390;
  reg [31:0] _RAND_110;
  reg [31:0] _EVAL_1417;
  reg [31:0] _RAND_111;
  reg  _EVAL_1422;
  reg [31:0] _RAND_112;
  reg [31:0] _EVAL_1431;
  reg [31:0] _RAND_113;
  reg [3:0] _EVAL_1439;
  reg [31:0] _RAND_114;
  reg [31:0] _EVAL_1441;
  reg [31:0] _RAND_115;
  reg  _EVAL_1442;
  reg [31:0] _RAND_116;
  reg [31:0] _EVAL_1444;
  reg [31:0] _RAND_117;
  reg  _EVAL_1450;
  reg [31:0] _RAND_118;
  reg  _EVAL_1486;
  reg [31:0] _RAND_119;
  reg  _EVAL_1489;
  reg [31:0] _RAND_120;
  reg [1:0] _EVAL_1500;
  reg [31:0] _RAND_121;
  reg [2:0] _EVAL_1502;
  reg [31:0] _RAND_122;
  reg  _EVAL_1506;
  reg [31:0] _RAND_123;
  reg [31:0] _EVAL_1527;
  reg [31:0] _RAND_124;
  reg [5:0] _EVAL_1541;
  reg [31:0] _RAND_125;
  reg  _EVAL_1555;
  reg [31:0] _RAND_126;
  reg [1:0] _EVAL_1569;
  reg [31:0] _RAND_127;
  reg  _EVAL_1594;
  reg [31:0] _RAND_128;
  reg  _EVAL_1595;
  reg [31:0] _RAND_129;
  reg [31:0] _EVAL_1619;
  reg [31:0] _RAND_130;
  reg  _EVAL_1620;
  reg [31:0] _RAND_131;
  reg [4:0] _EVAL_1625;
  reg [31:0] _RAND_132;
  reg [31:0] _EVAL_1626;
  reg [31:0] _RAND_133;
  reg  _EVAL_1650;
  reg [31:0] _RAND_134;
  reg [1:0] _EVAL_1661;
  reg [31:0] _RAND_135;
  reg [31:0] _EVAL_1688;
  reg [31:0] _RAND_136;
  reg  _EVAL_1697;
  reg [31:0] _RAND_137;
  reg [31:0] _EVAL_1709;
  reg [31:0] _RAND_138;
  reg  _EVAL_1716;
  reg [31:0] _RAND_139;
  reg [31:0] _EVAL_1724;
  reg [31:0] _RAND_140;
  reg  _EVAL_1733;
  reg [31:0] _RAND_141;
  reg  _EVAL_1739;
  reg [31:0] _RAND_142;
  reg [4:0] _EVAL_1740;
  reg [31:0] _RAND_143;
  reg [4:0] _EVAL_1756;
  reg [31:0] _RAND_144;
  reg [31:0] _EVAL_1774;
  reg [31:0] _RAND_145;
  reg [31:0] _EVAL_1784;
  reg [31:0] _RAND_146;
  reg  _EVAL_1800;
  reg [31:0] _RAND_147;
  reg  _EVAL_1805;
  reg [31:0] _RAND_148;
  reg [5:0] _EVAL_1810;
  reg [31:0] _RAND_149;
  reg [4:0] _EVAL_1814;
  reg [31:0] _RAND_150;
  reg [3:0] _EVAL_1827;
  reg [31:0] _RAND_151;
  reg [5:0] _EVAL_1831;
  reg [31:0] _RAND_152;
  reg  _EVAL_1832;
  reg [31:0] _RAND_153;
  reg  _EVAL_1835;
  reg [31:0] _RAND_154;
  reg [5:0] _EVAL_1844;
  reg [31:0] _RAND_155;
  reg  _EVAL_1847;
  reg [31:0] _RAND_156;
  reg [31:0] _EVAL_1851;
  reg [31:0] _RAND_157;
  wire  _EVAL_742;
  wire  _EVAL_1415;
  wire  _EVAL_1328;
  wire  _EVAL_1088;
  wire [6:0] _EVAL_762;
  wire [6:0] _EVAL_409;
  wire [7:0] _EVAL_1311;
  wire  _EVAL_770;
  wire  _EVAL_971;
  wire  _EVAL_307;
  wire  _EVAL_1715;
  wire  _EVAL_1326;
  wire  _EVAL_1303;
  wire  _EVAL_1263;
  wire [2:0] _EVAL_460;
  wire [2:0] _EVAL_885;
  wire [2:0] _EVAL_1535;
  wire [2:0] _EVAL_481;
  wire [2:0] _EVAL_1777;
  wire [2:0] _EVAL_855;
  wire [2:0] _EVAL_1117;
  wire [7:0] _EVAL_535;
  wire [6:0] _EVAL_187;
  wire  _EVAL_661;
  wire  _EVAL_1627;
  wire  _EVAL_476;
  wire  _EVAL_1609;
  wire  _EVAL_731;
  wire [2:0] _EVAL_1346;
  wire [2:0] _EVAL_1484;
  wire [2:0] _EVAL_696;
  wire  _EVAL_605;
  wire [3:0] _EVAL_647;
  wire [3:0] _EVAL_1686;
  wire [22:0] _EVAL_1022;
  wire [7:0] _EVAL_1194;
  wire [7:0] _EVAL_871;
  wire [4:0] _EVAL_908;
  wire [4:0] _EVAL_1523;
  wire [4:0] _EVAL_1526;
  wire [4:0] _EVAL_1306;
  wire [4:0] _EVAL_185;
  wire [5:0] _EVAL_551;
  wire  _EVAL_1865;
  wire  _EVAL_720;
  wire [3:0] _EVAL_1610;
  wire  _EVAL_1679;
  wire  _EVAL_1132;
  wire  _EVAL_1217;
  wire  _EVAL_1253;
  wire  _EVAL_994;
  wire  _EVAL_733;
  wire  _EVAL_418;
  wire  _EVAL_1823;
  wire  _EVAL_1007;
  wire  _EVAL_1685;
  wire  _EVAL_1861;
  wire  _EVAL_231;
  wire  _EVAL_287;
  wire  _EVAL_758;
  wire  _EVAL_1228;
  wire  _EVAL_1048;
  wire  _EVAL_1098;
  wire  _EVAL_1722;
  wire  _EVAL_398;
  wire  _EVAL_1536;
  wire  _EVAL_1458;
  wire  _EVAL_804;
  wire  _EVAL_1036;
  wire  _EVAL_1674;
  wire  _EVAL_1322;
  wire [1:0] _EVAL_1752;
  wire [1:0] _EVAL_1699;
  wire [1:0] _EVAL_787;
  wire [1:0] _EVAL_498;
  wire [5:0] _EVAL_1703;
  wire [5:0] _EVAL_1102;
  wire [2:0] _EVAL_1164;
  wire [5:0] _EVAL_660;
  wire  _EVAL_1358;
  wire  _EVAL_463;
  wire  _EVAL_439;
  wire  _EVAL_1511;
  wire  _EVAL_196;
  wire [1:0] _EVAL_977;
  wire [1:0] _EVAL_349;
  wire  _EVAL_812;
  wire [1:0] _EVAL_976;
  wire [1:0] _EVAL_1068;
  wire [1:0] _EVAL_1283;
  wire [3:0] _EVAL_1653;
  wire [3:0] _EVAL_1765;
  wire  _EVAL_314;
  wire  _EVAL_671;
  wire  _EVAL_450;
  wire [2:0] _EVAL_1186;
  wire [2:0] _EVAL_1124;
  wire [2:0] _EVAL_346;
  wire [2:0] _EVAL_449;
  wire [2:0] _EVAL_1023;
  wire [2:0] _EVAL_593;
  wire [2:0] _EVAL_1337;
  wire [2:0] _EVAL_442;
  wire  _EVAL_1110;
  wire  _EVAL_1191;
  wire  _EVAL_368;
  wire  _EVAL_548;
  wire [31:0] _EVAL_1333;
  wire [31:0] _EVAL_688;
  wire [31:0] _EVAL_806;
  wire  _EVAL_1762;
  wire  _EVAL_760;
  wire  _EVAL_530;
  wire  _EVAL_220;
  wire [31:0] _EVAL_1562;
  wire  _EVAL_552;
  wire [31:0] _EVAL_1876;
  wire  _EVAL_809;
  wire [31:0] _EVAL_567;
  wire [31:0] _EVAL_1084;
  wire  _EVAL_1214;
  wire [31:0] _EVAL_1581;
  wire [31:0] _EVAL_1792;
  wire  _EVAL_1126;
  wire [31:0] _EVAL_457;
  wire [31:0] _EVAL_1177;
  wire  _EVAL_562;
  wire [31:0] _EVAL_832;
  wire  _EVAL_1349;
  wire [31:0] _EVAL_159;
  wire [31:0] _EVAL_459;
  wire  _EVAL_735;
  wire [31:0] _EVAL_436;
  wire [31:0] _EVAL_1872;
  wire  _EVAL_1576;
  wire [31:0] _EVAL_830;
  wire [31:0] _EVAL_1423;
  wire [63:0] _EVAL_483;
  wire [7:0] _EVAL_507;
  wire [7:0] _EVAL_1143;
  wire [7:0] _EVAL_675;
  wire [7:0] _EVAL_1411;
  wire [7:0] _EVAL_525;
  wire [7:0] _EVAL_1862;
  wire [7:0] _EVAL_1236;
  wire [7:0] _EVAL_1080;
  wire [63:0] _EVAL_250;
  wire [31:0] _EVAL_680;
  wire [31:0] _EVAL_738;
  wire [31:0] _EVAL_353;
  wire [31:0] _EVAL_419;
  wire [15:0] _EVAL_1612;
  wire [15:0] _EVAL_1281;
  wire [15:0] _EVAL_623;
  wire  _EVAL_1597;
  wire  _EVAL_903;
  wire [15:0] _EVAL_601;
  wire [15:0] _EVAL_1434;
  wire [31:0] _EVAL_689;
  wire [7:0] _EVAL_1105;
  wire [7:0] _EVAL_1290;
  wire [7:0] _EVAL_912;
  wire [7:0] _EVAL_724;
  wire [5:0] _EVAL_1723;
  wire  _EVAL_878;
  wire  _EVAL_170;
  wire  _EVAL_794;
  wire  _EVAL_780;
  wire  _EVAL_404;
  wire  _EVAL_1552;
  wire  _EVAL_1871;
  wire  _EVAL_692;
  wire  _EVAL_486;
  wire  _EVAL_882;
  wire  _EVAL_805;
  wire  _EVAL_1244;
  wire  _EVAL_1384;
  wire  _EVAL_986;
  wire  _EVAL_299;
  wire  _EVAL_1368;
  wire  _EVAL_1158;
  wire  _EVAL_710;
  wire  _EVAL_440;
  wire  _EVAL_1717;
  wire  _EVAL_756;
  wire  _EVAL_1720;
  wire  _EVAL_873;
  wire  _EVAL_223;
  wire  _EVAL_925;
  wire  _EVAL_587;
  wire  _EVAL_1448;
  wire  _EVAL_1003;
  wire  _EVAL_511;
  wire  _EVAL_815;
  wire [3:0] _EVAL_840;
  wire  _EVAL_944;
  wire  _EVAL_1692;
  wire  _EVAL_1371;
  wire  _EVAL_216;
  wire  _EVAL_1667;
  wire  _EVAL_252;
  wire  _EVAL_201;
  wire  _EVAL_1247;
  wire  _EVAL_490;
  wire  _EVAL_238;
  wire  _EVAL_1364;
  wire  _EVAL_814;
  wire  _EVAL_1376;
  wire  _EVAL_1663;
  wire  _EVAL_259;
  wire  _EVAL_1826;
  wire  _EVAL_1226;
  wire  _EVAL_1018;
  wire  _EVAL_1628;
  wire  _EVAL_1850;
  wire  _EVAL_1781;
  wire  _EVAL_210;
  wire  _EVAL_394;
  wire  _EVAL_209;
  wire  _EVAL_1184;
  wire [25:0] _EVAL_714;
  wire  _EVAL_1857;
  wire  _EVAL_571;
  wire  _EVAL_1698;
  wire  _EVAL_1395;
  wire  _EVAL_1025;
  wire  _EVAL_860;
  wire  _EVAL_1753;
  wire  _EVAL_153;
  wire [21:0] _EVAL_456;
  wire [1:0] _EVAL_1561;
  wire  _EVAL_469;
  wire [19:0] _EVAL_1418;
  wire [19:0] _EVAL_1483;
  wire  _EVAL_1825;
  wire  _EVAL_424;
  wire [21:0] _EVAL_1010;
  wire [1:0] _EVAL_313;
  wire  _EVAL_1279;
  wire [19:0] _EVAL_799;
  wire  _EVAL_446;
  wire  _EVAL_1807;
  wire [21:0] _EVAL_1277;
  wire [1:0] _EVAL_1264;
  wire  _EVAL_1449;
  wire [19:0] _EVAL_1218;
  wire  _EVAL_1622;
  wire  _EVAL_1445;
  wire [21:0] _EVAL_407;
  wire [1:0] _EVAL_693;
  wire  _EVAL_437;
  wire [19:0] _EVAL_545;
  wire  _EVAL_317;
  wire  _EVAL_1242;
  wire [3:0] _EVAL_258;
  wire  _EVAL_722;
  wire [1:0] _EVAL_1858;
  wire  _EVAL_236;
  wire  _EVAL_1642;
  wire  _EVAL_564;
  wire [19:0] _EVAL_1534;
  wire [21:0] _EVAL_1258;
  wire  _EVAL_1780;
  wire  _EVAL_932;
  wire  _EVAL_1363;
  wire  _EVAL_1758;
  wire  _EVAL_1352;
  wire [1:0] _EVAL_1646;
  wire [1:0] _EVAL_334;
  wire [1:0] _EVAL_702;
  wire [1:0] _EVAL_1009;
  wire [1:0] _EVAL_1833;
  wire [1:0] _EVAL_1251;
  wire [1:0] _EVAL_1604;
  wire [1:0] _EVAL_1704;
  wire [1:0] _EVAL_662;
  wire [1:0] _EVAL_1867;
  wire [1:0] _EVAL_1701;
  wire [1:0] _EVAL_1014;
  wire  _EVAL_1478;
  wire  _EVAL_309;
  wire  _EVAL_792;
  wire [21:0] _EVAL_154;
  wire [2:0] _EVAL_1399;
  wire  _EVAL_679;
  wire  _EVAL_373;
  wire  _EVAL_1564;
  wire  _EVAL_1618;
  wire  _EVAL_1738;
  wire [3:0] _EVAL_431;
  wire [22:0] _EVAL_1745;
  wire [7:0] _EVAL_1072;
  wire [7:0] _EVAL_1557;
  wire [4:0] _EVAL_462;
  wire [4:0] _EVAL_345;
  wire  _EVAL_681;
  wire  _EVAL_553;
  wire  _EVAL_993;
  wire  _EVAL_1841;
  wire  _EVAL_990;
  wire  _EVAL_620;
  wire  _EVAL_946;
  wire  _EVAL_292;
  wire  _EVAL_1413;
  wire  _EVAL_1542;
  wire  _EVAL_400;
  wire  _EVAL_470;
  wire  _EVAL_602;
  wire  _EVAL_910;
  wire  _EVAL_1265;
  wire  _EVAL_405;
  wire  _EVAL_608;
  wire  _EVAL_697;
  wire  _EVAL_1398;
  wire  _EVAL_218;
  wire  _EVAL_1406;
  wire  _EVAL_364;
  wire  _EVAL_594;
  wire  _EVAL_1155;
  wire  _EVAL_271;
  wire  _EVAL_1845;
  wire  _EVAL_718;
  wire  _EVAL_466;
  wire  _EVAL_1660;
  wire  _EVAL_978;
  wire  _EVAL_1211;
  wire  _EVAL_172;
  wire  _EVAL_1127;
  wire  _EVAL_838;
  wire  _EVAL_1726;
  wire  _EVAL_778;
  wire  _EVAL_754;
  wire  _EVAL_590;
  wire  _EVAL_1207;
  wire  _EVAL_913;
  wire  _EVAL_261;
  wire  _EVAL_699;
  wire  _EVAL_1160;
  wire  _EVAL_194;
  wire  _EVAL_199;
  wire  _EVAL_849;
  wire  _EVAL_1118;
  wire  _EVAL_583;
  wire  _EVAL_435;
  wire  _EVAL_555;
  wire  _EVAL_822;
  wire  _EVAL_1302;
  wire  _EVAL_709;
  wire  _EVAL_1725;
  wire  _EVAL_1438;
  wire  _EVAL_1270;
  wire  _EVAL_1757;
  wire  _EVAL_816;
  wire  _EVAL_927;
  wire  _EVAL_1782;
  wire  _EVAL_1669;
  wire  _EVAL_193;
  wire  _EVAL_306;
  wire  _EVAL_1016;
  wire  _EVAL_1221;
  wire  _EVAL_1718;
  wire  _EVAL_1020;
  wire  _EVAL_1166;
  wire  _EVAL_1129;
  wire  _EVAL_1343;
  wire  _EVAL_1788;
  wire [1:0] _EVAL_448;
  wire [3:0] _EVAL_455;
  wire  _EVAL_818;
  wire  _EVAL_1241;
  wire  _EVAL_518;
  wire  _EVAL_1809;
  wire [1:0] _EVAL_572;
  wire [1:0] _EVAL_184;
  wire [1:0] _EVAL_565;
  wire [1:0] _EVAL_782;
  wire [21:0] _EVAL_1459;
  wire  _EVAL_311;
  wire  _EVAL_1273;
  wire [3:0] _EVAL_163;
  wire  _EVAL_1785;
  wire  _EVAL_687;
  wire  _EVAL_1493;
  wire  _EVAL_789;
  wire  _EVAL_179;
  wire  _EVAL_381;
  wire  _EVAL_1391;
  wire [1:0] _EVAL_727;
  wire [1:0] _EVAL_468;
  wire [1:0] _EVAL_1386;
  wire [1:0] _EVAL_1440;
  wire [1:0] _EVAL_443;
  wire [1:0] _EVAL_1039;
  wire [1:0] _EVAL_510;
  wire [1:0] _EVAL_491;
  wire [1:0] _EVAL_983;
  wire [1:0] _EVAL_1336;
  wire [1:0] _EVAL_1066;
  wire [1:0] _EVAL_1112;
  wire [1:0] _EVAL_494;
  wire [1:0] _EVAL_324;
  wire [1:0] _EVAL_1401;
  wire [31:0] _EVAL_1293;
  wire [19:0] _EVAL_707;
  wire [21:0] _EVAL_930;
  wire  _EVAL_1237;
  wire [21:0] _EVAL_788;
  wire  _EVAL_403;
  wire  _EVAL_1524;
  wire  _EVAL_694;
  wire  _EVAL_1027;
  wire  _EVAL_824;
  wire  _EVAL_509;
  wire  _EVAL_242;
  wire  _EVAL_1206;
  wire  _EVAL_1605;
  wire  _EVAL_1481;
  wire  _EVAL_1131;
  wire [21:0] _EVAL_854;
  wire [21:0] _EVAL_1354;
  wire [21:0] _EVAL_1770;
  wire [21:0] _EVAL_825;
  wire [21:0] _EVAL_1378;
  wire [21:0] _EVAL_1215;
  wire [21:0] _EVAL_972;
  wire [21:0] _EVAL_1607;
  wire  _EVAL_1430;
  wire  _EVAL_705;
  wire  _EVAL_219;
  wire  _EVAL_1086;
  wire  _EVAL_531;
  wire  _EVAL_560;
  wire  _EVAL_1601;
  wire  _EVAL_428;
  wire  _EVAL_1455;
  wire [11:0] _EVAL_561;
  wire  _EVAL_284;
  wire  _EVAL_1462;
  wire  _EVAL_791;
  wire  _EVAL_1611;
  wire  _EVAL_1687;
  wire [3:0] _EVAL_465;
  wire  _EVAL_736;
  wire [2:0] _EVAL_547;
  wire [2:0] _EVAL_169;
  wire  _EVAL_240;
  wire  _EVAL_344;
  wire  _EVAL_191;
  wire  _EVAL_1820;
  wire  _EVAL_276;
  wire [31:0] _EVAL_1151;
  wire [31:0] _EVAL_899;
  wire [63:0] _EVAL_752;
  wire [7:0] _EVAL_865;
  wire  _EVAL_331;
  wire  _EVAL_180;
  wire  _EVAL_1457;
  wire  _EVAL_796;
  wire  _EVAL_264;
  wire [2:0] _EVAL_513;
  wire [7:0] _EVAL_960;
  wire [6:0] _EVAL_1769;
  wire  _EVAL_1348;
  wire  _EVAL_176;
  wire  _EVAL_1632;
  wire  _EVAL_1736;
  wire  _EVAL_672;
  wire  _EVAL_467;
  wire  _EVAL_1475;
  wire  _EVAL_453;
  wire  _EVAL_1205;
  wire  _EVAL_1170;
  wire  _EVAL_970;
  wire  _EVAL_1464;
  wire  _EVAL_901;
  wire  _EVAL_267;
  wire  _EVAL_884;
  wire  _EVAL_870;
  wire  _EVAL_862;
  wire  _EVAL_406;
  wire  _EVAL_497;
  wire  _EVAL_568;
  wire  _EVAL_416;
  wire  _EVAL_249;
  wire  _EVAL_1672;
  wire  _EVAL_174;
  wire  _EVAL_445;
  wire  _EVAL_1005;
  wire  _EVAL_1658;
  wire [63:0] _EVAL_382;
  wire  _EVAL_935;
  wire  _EVAL_496;
  wire  _EVAL_1061;
  wire  _EVAL_813;
  wire  _EVAL_779;
  wire  _EVAL_1567;
  wire  _EVAL_1369;
  wire  _EVAL_546;
  wire  _EVAL_1520;
  wire  _EVAL_1295;
  wire  _EVAL_817;
  wire  _EVAL_784;
  wire [2:0] _EVAL_454;
  wire [2:0] _EVAL_1623;
  wire [2:0] _EVAL_622;
  wire [2:0] _EVAL_1577;
  wire [2:0] _EVAL_1299;
  wire [2:0] _EVAL_711;
  wire [2:0] _EVAL_691;
  wire [2:0] _EVAL_734;
  wire [1:0] _EVAL_615;
  wire [7:0] _EVAL_207;
  wire [15:0] _EVAL_1710;
  wire  _EVAL_606;
  wire  _EVAL_524;
  wire  _EVAL_1819;
  wire  _EVAL_1312;
  wire  _EVAL_634;
  wire  _EVAL_1267;
  wire  _EVAL_1298;
  wire  _EVAL_1517;
  wire  _EVAL_1187;
  wire  _EVAL_1389;
  wire  _EVAL_479;
  wire  _EVAL_1313;
  wire  _EVAL_1474;
  wire  _EVAL_412;
  wire  _EVAL_1063;
  wire  _EVAL_580;
  wire [7:0] _EVAL_698;
  wire [15:0] _EVAL_947;
  wire [1:0] _EVAL_1556;
  wire [1:0] _EVAL_426;
  wire  _EVAL_563;
  wire  _EVAL_1046;
  wire [3:0] _EVAL_1062;
  wire [3:0] _EVAL_1838;
  wire [5:0] _EVAL_1181;
  wire [11:0] _EVAL_658;
  wire  _EVAL_945;
  wire  _EVAL_1315;
  wire [31:0] _EVAL_1476;
  wire [31:0] _EVAL_1409;
  wire [5:0] _EVAL_851;
  wire  _EVAL_1097;
  wire  _EVAL_923;
  wire  _EVAL_217;
  wire  _EVAL_1775;
  wire  _EVAL_521;
  wire [4:0] _EVAL_900;
  wire [4:0] _EVAL_168;
  wire [4:0] _EVAL_294;
  wire [7:0] _EVAL_569;
  wire [31:0] _EVAL_785;
  wire  _EVAL_879;
  wire  _EVAL_1188;
  wire  _EVAL_641;
  wire  _EVAL_1284;
  wire  _EVAL_1821;
  wire  _EVAL_253;
  wire  _EVAL_1153;
  wire  _EVAL_1587;
  wire  _EVAL_617;
  wire [2:0] _EVAL_664;
  wire [2:0] _EVAL_954;
  wire [2:0] _EVAL_303;
  wire [2:0] _EVAL_576;
  wire [2:0] _EVAL_391;
  wire [2:0] _EVAL_523;
  wire [2:0] _EVAL_1505;
  wire [2:0] _EVAL_1367;
  wire [2:0] _EVAL_1201;
  wire [2:0] _EVAL_934;
  wire  _EVAL_1327;
  wire  _EVAL_716;
  wire [3:0] _EVAL_597;
  wire [3:0] _EVAL_619;
  wire [3:0] _EVAL_166;
  wire [3:0] _EVAL_1676;
  wire [3:0] _EVAL_996;
  wire [3:0] _EVAL_1522;
  wire [3:0] _EVAL_330;
  wire [3:0] _EVAL_1707;
  wire [3:0] _EVAL_1152;
  wire [3:0] _EVAL_297;
  wire [3:0] _EVAL_747;
  wire [3:0] _EVAL_638;
  wire [3:0] _EVAL_421;
  wire [22:0] _EVAL_1648;
  wire [7:0] _EVAL_1297;
  wire [7:0] _EVAL_420;
  wire [4:0] _EVAL_1681;
  wire [4:0] _EVAL_447;
  wire [4:0] _EVAL_1055;
  wire [9:0] _EVAL_1380;
  wire [9:0] _EVAL_1248;
  wire  _EVAL_310;
  wire  _EVAL_298;
  wire  _EVAL_1168;
  wire  _EVAL_1538;
  wire  _EVAL_1763;
  wire [3:0] _EVAL_1521;
  wire  _EVAL_1161;
  wire  _EVAL_1165;
  wire  _EVAL_1737;
  wire  _EVAL_869;
  wire [3:0] _EVAL_1631;
  wire  _EVAL_1256;
  wire  _EVAL_670;
  wire  _EVAL_1693;
  wire  _EVAL_1528;
  wire [3:0] _EVAL_1503;
  wire  _EVAL_997;
  wire  _EVAL_768;
  wire  _EVAL_1671;
  wire  _EVAL_1288;
  wire [3:0] _EVAL_1495;
  wire [3:0] _EVAL_1053;
  wire  _EVAL_1641;
  wire [3:0] _EVAL_182;
  wire  _EVAL_755;
  wire  _EVAL_399;
  wire  _EVAL_1860;
  wire  _EVAL_1394;
  wire  _EVAL_1673;
  wire  _EVAL_251;
  wire  _EVAL_1624;
  wire  _EVAL_427;
  wire  _EVAL_343;
  wire  _EVAL_1846;
  wire  _EVAL_1508;
  wire  _EVAL_296;
  wire  _EVAL_807;
  wire [7:0] _EVAL_1119;
  wire [63:0] _EVAL_512;
  wire [31:0] _EVAL_534;
  wire [3:0] _EVAL_811;
  wire [3:0] _EVAL_1185;
  wire [3:0] _EVAL_829;
  wire  _EVAL_1433;
  wire  _EVAL_175;
  wire  _EVAL_248;
  wire  _EVAL_1011;
  wire  _EVAL_1359;
  wire  _EVAL_1192;
  wire  _EVAL_1254;
  wire  _EVAL_351;
  wire [2:0] _EVAL_950;
  wire [2:0] _EVAL_422;
  wire [2:0] _EVAL_1566;
  wire [2:0] _EVAL_366;
  wire  _EVAL_1830;
  wire  _EVAL_891;
  wire  _EVAL_1519;
  wire  _EVAL_772;
  wire  _EVAL_1680;
  wire  _EVAL_1729;
  wire  _EVAL_1764;
  wire  _EVAL_1420;
  wire  _EVAL_1139;
  wire  _EVAL_957;
  wire  _EVAL_1608;
  wire  _EVAL_1323;
  wire  _EVAL_889;
  wire  _EVAL_704;
  wire  _EVAL_1818;
  wire  _EVAL_668;
  wire [2:0] _EVAL_1815;
  wire [2:0] _EVAL_347;
  wire [2:0] _EVAL_1640;
  wire [2:0] _EVAL_295;
  wire [2:0] _EVAL_1150;
  wire [2:0] _EVAL_948;
  wire [2:0] _EVAL_1559;
  wire [2:0] _EVAL_1094;
  wire [1:0] _EVAL_350;
  wire [3:0] _EVAL_1379;
  wire [2:0] _EVAL_1537;
  wire [2:0] _EVAL_235;
  wire  _EVAL_1572;
  wire  _EVAL_1246;
  wire  _EVAL_1314;
  wire  _EVAL_1092;
  wire  _EVAL_444;
  wire [63:0] _EVAL_1488;
  wire [63:0] _EVAL_765;
  wire [63:0] _EVAL_1585;
  wire [63:0] _EVAL_1848;
  wire [63:0] _EVAL_1727;
  wire [63:0] _EVAL_633;
  wire [3:0] _EVAL_434;
  wire [3:0] _EVAL_713;
  wire  _EVAL_1778;
  wire  _EVAL_939;
  wire  _EVAL_452;
  wire [1:0] _EVAL_1250;
  wire  _EVAL_195;
  wire [19:0] _EVAL_1342;
  wire [31:0] _EVAL_1694;
  wire [19:0] _EVAL_464;
  wire [11:0] _EVAL_663;
  wire [31:0] _EVAL_529;
  wire [31:0] _EVAL_1741;
  wire [11:0] _EVAL_1108;
  wire [31:0] _EVAL_1579;
  wire [5:0] _EVAL_625;
  wire [11:0] _EVAL_968;
  wire [31:0] _EVAL_1360;
  wire [32:0] _EVAL_1178;
  wire [32:0] _EVAL_304;
  wire [32:0] _EVAL_1593;
  wire [31:0] _EVAL_234;
  wire [31:0] _EVAL_1197;
  wire [31:0] _EVAL_473;
  wire [31:0] _EVAL_260;
  wire [31:0] _EVAL_522;
  wire [31:0] _EVAL_266;
  wire [31:0] _EVAL_1615;
  wire  _EVAL_1078;
  wire  _EVAL_379;
  wire  _EVAL_837;
  wire  _EVAL_676;
  wire  _EVAL_233;
  wire  _EVAL_892;
  wire  _EVAL_886;
  wire  _EVAL_1338;
  wire  _EVAL_828;
  wire  _EVAL_160;
  wire  _EVAL_1760;
  wire [31:0] _EVAL_867;
  wire [31:0] _EVAL_339;
  wire [3:0] _EVAL_283;
  wire [3:0] _EVAL_1209;
  wire [3:0] _EVAL_589;
  wire [3:0] _EVAL_1437;
  wire [9:0] _EVAL_1793;
  wire  _EVAL_1125;
  wire  _EVAL_348;
  wire  _EVAL_1750;
  wire  _EVAL_748;
  wire  _EVAL_906;
  wire [3:0] _EVAL_1432;
  wire  _EVAL_319;
  wire  _EVAL_586;
  wire  _EVAL_823;
  wire  _EVAL_197;
  wire [3:0] _EVAL_508;
  wire [3:0] _EVAL_868;
  wire  _EVAL_952;
  wire  _EVAL_1639;
  wire  _EVAL_863;
  wire  _EVAL_441;
  wire  _EVAL_1705;
  wire  _EVAL_1223;
  wire  _EVAL_1813;
  wire  _EVAL_919;
  wire  _EVAL_363;
  wire  _EVAL_1294;
  wire  _EVAL_956;
  wire  _EVAL_648;
  wire  _EVAL_876;
  wire  _EVAL_1220;
  wire  _EVAL_1568;
  wire  _EVAL_1008;
  wire  _EVAL_1662;
  wire  _EVAL_301;
  wire  _EVAL_1786;
  wire  _EVAL_1309;
  wire  _EVAL_1637;
  wire  _EVAL_1849;
  wire  _EVAL_1515;
  wire [79:0] _EVAL_810;
  wire [79:0] _EVAL_1087;
  wire [79:0] _EVAL_640;
  wire [79:0] _EVAL_1268;
  wire [79:0] _EVAL_808;
  wire [79:0] _EVAL_1000;
  wire [79:0] _EVAL_1280;
  wire [79:0] _EVAL_327;
  wire  _EVAL_1393;
  wire [79:0] _EVAL_636;
  wire [79:0] _EVAL_227;
  wire [79:0] _EVAL_1351;
  wire  _EVAL_362;
  wire [79:0] _EVAL_1245;
  wire [79:0] _EVAL_1070;
  wire [79:0] _EVAL_1447;
  wire [79:0] _EVAL_880;
  wire [79:0] _EVAL_517;
  wire [79:0] _EVAL_1093;
  wire  _EVAL_585;
  wire  _EVAL_1766;
  wire  _EVAL_1675;
  wire  _EVAL_338;
  wire  _EVAL_1123;
  wire  _EVAL_1635;
  wire  _EVAL_1017;
  wire [2:0] _EVAL_991;
  wire [2:0] _EVAL_603;
  wire [2:0] _EVAL_1308;
  wire [2:0] _EVAL_1772;
  wire [2:0] _EVAL_1282;
  wire [2:0] _EVAL_192;
  wire [2:0] _EVAL_1429;
  wire [2:0] _EVAL_500;
  wire [2:0] _EVAL_326;
  wire [2:0] _EVAL_1331;
  wire [2:0] _EVAL_539;
  wire  _EVAL_1219;
  wire [31:0] _EVAL_536;
  wire  _EVAL_843;
  wire  _EVAL_537;
  wire  _EVAL_245;
  wire  _EVAL_1580;
  wire  _EVAL_499;
  wire  _EVAL_1510;
  wire  _EVAL_669;
  wire  _EVAL_1106;
  wire  _EVAL_652;
  wire  _EVAL_1743;
  wire  _EVAL_244;
  wire  _EVAL_574;
  wire  _EVAL_1543;
  wire  _EVAL_866;
  wire  _EVAL_1836;
  wire  _EVAL_1103;
  wire  _EVAL_988;
  wire  _EVAL_1602;
  wire  _EVAL_1408;
  wire  _EVAL_262;
  wire  _EVAL_1469;
  wire  _EVAL_281;
  wire  _EVAL_1799;
  wire  _EVAL_1712;
  wire  _EVAL_1403;
  wire  _EVAL_974;
  wire [2:0] _EVAL_1529;
  wire [1:0] _EVAL_985;
  wire  _EVAL_1163;
  wire [1:0] _EVAL_857;
  wire [3:0] _EVAL_917;
  wire  _EVAL_1064;
  wire [79:0] _EVAL_1613;
  wire [79:0] _EVAL_1042;
  wire [79:0] _EVAL_1853;
  wire  _EVAL_653;
  wire [31:0] _EVAL_516;
  wire  _EVAL_358;
  wire  _EVAL_1400;
  wire [63:0] _EVAL_1362;
  wire [31:0] _EVAL_208;
  wire [31:0] _EVAL_203;
  wire [31:0] _EVAL_764;
  wire [15:0] _EVAL_856;
  wire [15:0] _EVAL_1547;
  wire [15:0] _EVAL_1045;
  wire  _EVAL_1452;
  wire  _EVAL_1210;
  wire [31:0] _EVAL_1073;
  wire [2:0] _EVAL_1514;
  wire [2:0] _EVAL_1335;
  wire [2:0] _EVAL_864;
  wire [2:0] _EVAL_965;
  wire  _EVAL_214;
  wire [7:0] _EVAL_1030;
  wire  _EVAL_392;
  wire  _EVAL_321;
  wire [63:0] _EVAL_1388;
  wire [63:0] _EVAL_964;
  wire  _EVAL_255;
  wire  _EVAL_1071;
  wire  _EVAL_1180;
  wire  _EVAL_1133;
  wire  _EVAL_673;
  wire  _EVAL_1138;
  wire  _EVAL_504;
  wire  _EVAL_1713;
  wire [19:0] _EVAL_888;
  wire  _EVAL_156;
  wire  _EVAL_1614;
  wire  _EVAL_360;
  wire  _EVAL_161;
  wire  _EVAL_833;
  wire  _EVAL_1353;
  wire  _EVAL_333;
  wire  _EVAL_929;
  wire [2:0] _EVAL_554;
  wire [2:0] _EVAL_852;
  wire [2:0] _EVAL_1130;
  wire [2:0] _EVAL_695;
  wire  _EVAL_1038;
  wire [19:0] _EVAL_1643;
  wire  _EVAL_1477;
  wire  _EVAL_1768;
  wire  _EVAL_1344;
  wire  _EVAL_1645;
  wire  _EVAL_975;
  wire  _EVAL_1728;
  wire  _EVAL_383;
  wire  _EVAL_1357;
  wire  _EVAL_757;
  wire  _EVAL_1291;
  wire [31:0] _EVAL_600;
  wire [7:0] _EVAL_432;
  wire [7:0] _EVAL_270;
  wire [7:0] _EVAL_1307;
  wire [7:0] _EVAL_1578;
  wire [31:0] _EVAL_1182;
  wire  _EVAL_581;
  wire  _EVAL_1530;
  wire [6:0] _EVAL_1652;
  wire  _EVAL_337;
  wire  _EVAL_848;
  wire  _EVAL_1321;
  wire  _EVAL_575;
  wire [25:0] _EVAL_489;
  wire [31:0] _EVAL_1732;
  wire [31:0] _EVAL_684;
  wire [11:0] _EVAL_1487;
  wire [11:0] _EVAL_1059;
  wire [11:0] _EVAL_1824;
  wire [11:0] _EVAL_1414;
  wire [11:0] _EVAL_802;
  wire [11:0] _EVAL_1385;
  wire [5:0] _EVAL_1204;
  wire [25:0] _EVAL_1301;
  wire  _EVAL_336;
  wire  _EVAL_751;
  wire  _EVAL_1747;
  wire  _EVAL_1491;
  wire  _EVAL_685;
  wire  _EVAL_1822;
  wire  _EVAL_1443;
  wire [7:0] _EVAL_781;
  wire  _EVAL_783;
  wire  _EVAL_478;
  wire  _EVAL_607;
  wire  _EVAL_1111;
  wire  _EVAL_657;
  wire  _EVAL_1549;
  wire [1:0] _EVAL_1795;
  wire [1:0] _EVAL_1397;
  wire [2:0] _EVAL_626;
  wire  _EVAL_1116;
  wire  _EVAL_936;
  wire  _EVAL_682;
  wire  _EVAL_1085;
  wire  _EVAL_323;
  wire  _EVAL_285;
  wire  _EVAL_726;
  wire  _EVAL_1216;
  wire  _EVAL_1621;
  wire  _EVAL_206;
  wire  _EVAL_570;
  wire  _EVAL_378;
  wire  _EVAL_649;
  wire  _EVAL_1149;
  wire  _EVAL_318;
  wire  _EVAL_1142;
  wire  _EVAL_1199;
  wire  _EVAL_1573;
  wire  _EVAL_578;
  wire  _EVAL_173;
  wire  _EVAL_1790;
  wire  _EVAL_237;
  wire  _EVAL_1260;
  wire  _EVAL_803;
  wire  _EVAL_1162;
  wire  _EVAL_1383;
  wire  _EVAL_1099;
  wire  _EVAL_1659;
  wire  _EVAL_385;
  wire [7:0] _EVAL_501;
  wire [7:0] _EVAL_1599;
  wire [7:0] _EVAL_599;
  wire [7:0] _EVAL_834;
  wire  _EVAL_1345;
  wire  _EVAL_1050;
  wire [2:0] _EVAL_1451;
  wire [1:0] _EVAL_1719;
  wire [3:0] _EVAL_630;
  wire [8:0] _EVAL_1539;
  wire [2:0] _EVAL_157;
  wire  _EVAL_881;
  wire [25:0] _EVAL_1339;
  wire [5:0] _EVAL_1859;
  wire [31:0] _EVAL_1606;
  wire [2:0] _EVAL_797;
  wire [2:0] _EVAL_1787;
  wire [2:0] _EVAL_256;
  wire [2:0] _EVAL_1532;
  wire [2:0] _EVAL_243;
  wire [2:0] _EVAL_1683;
  wire [2:0] _EVAL_1305;
  wire [2:0] _EVAL_1571;
  wire  _EVAL_335;
  wire [1:0] _EVAL_520;
  wire  _EVAL_743;
  wire [15:0] _EVAL_1012;
  wire [15:0] _EVAL_1179;
  wire [31:0] _EVAL_550;
  wire [7:0] _EVAL_1468;
  wire [7:0] _EVAL_1276;
  wire [7:0] _EVAL_505;
  wire  _EVAL_1224;
  wire  _EVAL_1289;
  wire [23:0] _EVAL_1504;
  wire [7:0] _EVAL_844;
  wire [7:0] _EVAL_1654;
  wire [7:0] _EVAL_1144;
  wire [7:0] _EVAL_1320;
  wire [7:0] _EVAL_1173;
  wire [7:0] _EVAL_920;
  wire [2:0] _EVAL_1075;
  wire  _EVAL_229;
  wire [1:0] _EVAL_200;
  wire [1:0] _EVAL_423;
  wire  _EVAL_315;
  wire  _EVAL_1136;
  wire  _EVAL_1866;
  wire  _EVAL_1591;
  wire  _EVAL_706;
  wire  _EVAL_1081;
  wire  _EVAL_528;
  wire  _EVAL_1249;
  wire  _EVAL_1629;
  wire  _EVAL_246;
  wire  _EVAL_610;
  wire  _EVAL_1137;
  wire  _EVAL_1424;
  wire  _EVAL_415;
  wire  _EVAL_1551;
  wire  _EVAL_1834;
  wire  _EVAL_1347;
  wire  _EVAL_958;
  wire  _EVAL_515;
  wire  _EVAL_729;
  wire  _EVAL_1175;
  wire  _EVAL_941;
  wire  _EVAL_1159;
  wire [3:0] _EVAL_1052;
  wire [3:0] _EVAL_495;
  wire [3:0] _EVAL_1148;
  wire [3:0] _EVAL_850;
  wire [3:0] _EVAL_1575;
  wire [3:0] _EVAL_1381;
  wire [31:0] _EVAL_1708;
  wire [31:0] _EVAL_1545;
  wire [31:0] _EVAL_1146;
  wire [31:0] _EVAL_1574;
  wire  _EVAL_411;
  wire  _EVAL_798;
  wire [23:0] _EVAL_1095;
  wire  _EVAL_1657;
  wire  _EVAL_1113;
  wire [31:0] _EVAL_628;
  wire [7:0] _EVAL_1533;
  wire [4:0] _EVAL_371;
  wire [3:0] _EVAL_527;
  wire [3:0] _EVAL_340;
  wire [3:0] _EVAL_1029;
  wire [3:0] _EVAL_222;
  wire [5:0] _EVAL_916;
  wire [5:0] _EVAL_1304;
  wire [5:0] _EVAL_842;
  wire [5:0] _EVAL_1425;
  wire [5:0] _EVAL_914;
  wire [5:0] _EVAL_1021;
  wire [31:0] _EVAL_1655;
  wire [7:0] _EVAL_305;
  wire  _EVAL_1019;
  wire  _EVAL_1497;
  wire  _EVAL_1617;
  wire  _EVAL_1771;
  wire  _EVAL_744;
  wire [2:0] _EVAL_845;
  wire  _EVAL_1463;
  wire [2:0] _EVAL_183;
  wire [2:0] _EVAL_1446;
  wire [2:0] _EVAL_894;
  wire [2:0] _EVAL_1157;
  wire  _EVAL_767;
  wire [7:0] _EVAL_213;
  wire [7:0] _EVAL_717;
  wire [7:0] _EVAL_540;
  wire [31:0] _EVAL_940;
  wire [7:0] _EVAL_998;
  wire [7:0] _EVAL_188;
  wire [7:0] _EVAL_616;
  wire [31:0] _EVAL_579;
  wire [63:0] _EVAL_1702;
  wire  _EVAL_963;
  wire [1:0] _EVAL_1695;
  wire [1:0] _EVAL_1435;
  wire [1:0] _EVAL_1461;
  wire  _EVAL_1616;
  wire [3:0] _EVAL_312;
  wire [3:0] _EVAL_1811;
  wire  _EVAL_635;
  wire  _EVAL_643;
  wire [2:0] _EVAL_1412;
  wire [2:0] _EVAL_1589;
  wire  _EVAL_1261;
  wire  _EVAL_1649;
  wire [23:0] _EVAL_995;
  wire [5:0] _EVAL_1665;
  wire [5:0] _EVAL_835;
  wire [5:0] _EVAL_275;
  wire [5:0] _EVAL_1794;
  wire [5:0] _EVAL_609;
  wire [63:0] _EVAL_905;
  wire [63:0] _EVAL_1115;
  wire [8:0] _EVAL_1518;
  wire [8:0] _EVAL_883;
  wire [8:0] _EVAL_890;
  wire [3:0] _EVAL_279;
  wire [63:0] _EVAL_1330;
  wire [2:0] _EVAL_771;
  wire [2:0] _EVAL_151;
  wire [2:0] _EVAL_1198;
  wire  _EVAL_1466;
  wire [1:0] _EVAL_966;
  wire [1:0] _EVAL_177;
  wire  _EVAL_1202;
  wire [1:0] _EVAL_268;
  wire [1:0] _EVAL_793;
  wire  _EVAL_1332;
  wire  _EVAL_683;
  wire  _EVAL_646;
  wire [7:0] _EVAL_1499;
  wire [7:0] _EVAL_774;
  wire [7:0] _EVAL_1754;
  wire [31:0] _EVAL_566;
  wire [63:0] _EVAL_761;
  wire  _EVAL_665;
  wire  _EVAL_1749;
  wire  _EVAL_1426;
  wire  _EVAL_979;
  wire [31:0] _EVAL_984;
  wire [31:0] _EVAL_750;
  wire [31:0] _EVAL_1791;
  wire [31:0] _EVAL_1798;
  wire [7:0] _EVAL_1091;
  wire [63:0] _EVAL_482;
  wire [63:0] _EVAL_1040;
  wire [63:0] _EVAL_402;
  wire [63:0] _EVAL_1208;
  wire [63:0] _EVAL_604;
  wire  _EVAL_1467;
  wire  _EVAL_164;
  wire  _EVAL_1803;
  wire  _EVAL_1812;
  wire [2:0] _EVAL_1318;
  wire  _EVAL_961;
  wire [7:0] _EVAL_425;
  wire [7:0] _EVAL_1840;
  wire  _EVAL_577;
  wire  _EVAL_484;
  wire  _EVAL_1230;
  wire  _EVAL_708;
  wire  _EVAL_325;
  wire  _EVAL_241;
  wire [3:0] _EVAL_931;
  wire  _EVAL_969;
  wire [1:0] _EVAL_1582;
  wire [1:0] _EVAL_654;
  wire [1:0] _EVAL_773;
  wire [5:0] _EVAL_288;
  wire [5:0] _EVAL_384;
  wire [5:0] _EVAL_395;
  wire  _EVAL_1839;
  wire  _EVAL_667;
  wire [63:0] _EVAL_1069;
  wire [31:0] _EVAL_1077;
  wire  _EVAL_1243;
  wire  _EVAL_1516;
  wire  _EVAL_1404;
  wire  _EVAL_1668;
  wire [63:0] _EVAL_1141;
  wire [31:0] _EVAL_962;
  wire  _EVAL_1666;
  wire  _EVAL_224;
  wire  _EVAL_1465;
  wire  _EVAL_1748;
  wire [23:0] _EVAL_225;
  wire [23:0] _EVAL_1806;
  wire  _EVAL_973;
  wire [31:0] _EVAL_1183;
  wire  _EVAL_1233;
  wire  _EVAL_1512;
  wire  _EVAL_1751;
  wire [31:0] _EVAL_493;
  wire [11:0] _EVAL_1636;
  wire [63:0] _EVAL_1340;
  wire  _EVAL_618;
  wire [63:0] _EVAL_1473;
  wire [31:0] _EVAL_1761;
  wire [31:0] _EVAL_532;
  wire [2:0] _EVAL_328;
  wire  _EVAL_1711;
  wire [2:0] _EVAL_1065;
  wire  _EVAL_1863;
  wire [23:0] _EVAL_226;
  wire [63:0] _EVAL_1402;
  wire  _EVAL_959;
  wire  _EVAL_627;
  wire [31:0] _EVAL_1507;
  wire [1:0] _EVAL_949;
  wire  _EVAL_1190;
  wire  _EVAL_1082;
  wire  _EVAL_1588;
  wire [2:0] _EVAL_1600;
  wire  _EVAL_167;
  wire  _EVAL_591;
  wire  _EVAL_1498;
  wire  _EVAL_1272;
  wire  _EVAL_380;
  wire [7:0] _EVAL_820;
  wire [2:0] _EVAL_1596;
  wire  _EVAL_584;
  wire  _EVAL_430;
  wire  _EVAL_1193;
  wire [3:0] _EVAL_721;
  wire  _EVAL_492;
  wire  _EVAL_186;
  wire  _EVAL_841;
  wire [31:0] _EVAL_417;
  wire [63:0] _EVAL_1076;
  wire  _EVAL_374;
  wire [3:0] _EVAL_1691;
  wire  _EVAL_1334;
  wire [31:0] _EVAL_458;
  wire  _EVAL_278;
  wire  _EVAL_1361;
  wire  _EVAL_686;
  wire  _EVAL_1456;
  wire  _EVAL_967;
  wire  _EVAL_1570;
  wire [7:0] _EVAL_839;
  wire  _EVAL_895;
  wire [11:0] _EVAL_666;
  wire  _EVAL_1407;
  wire  _EVAL_471;
  wire [31:0] _EVAL_1682;
  wire  _EVAL_1416;
  wire  _EVAL_1329;
  wire  _EVAL_677;
  SiFive__EVAL_254 data (
    ._EVAL(data__EVAL),
    ._EVAL_0(data__EVAL_0),
    ._EVAL_1(data__EVAL_1),
    ._EVAL_2(data__EVAL_2),
    ._EVAL_3(data__EVAL_3),
    ._EVAL_4(data__EVAL_4),
    ._EVAL_5(data__EVAL_5),
    ._EVAL_6(data__EVAL_6),
    ._EVAL_7(data__EVAL_7),
    ._EVAL_8(data__EVAL_8),
    ._EVAL_9(data__EVAL_9),
    ._EVAL_10(data__EVAL_10)
  );
  EICG_wrapper dcache_clock_gate (
    .in(dcache_clock_gate_in),
    .en(dcache_clock_gate_en),
    .out(dcache_clock_gate_out)
  );
  SiFive__EVAL_257 tlb (
    ._EVAL(tlb__EVAL),
    ._EVAL_0(tlb__EVAL_0),
    ._EVAL_1(tlb__EVAL_1),
    ._EVAL_2(tlb__EVAL_2),
    ._EVAL_3(tlb__EVAL_3),
    ._EVAL_4(tlb__EVAL_4),
    ._EVAL_5(tlb__EVAL_5),
    ._EVAL_6(tlb__EVAL_6),
    ._EVAL_7(tlb__EVAL_7),
    ._EVAL_8(tlb__EVAL_8),
    ._EVAL_9(tlb__EVAL_9),
    ._EVAL_10(tlb__EVAL_10),
    ._EVAL_11(tlb__EVAL_11),
    ._EVAL_12(tlb__EVAL_12),
    ._EVAL_13(tlb__EVAL_13),
    ._EVAL_14(tlb__EVAL_14),
    ._EVAL_15(tlb__EVAL_15),
    ._EVAL_16(tlb__EVAL_16),
    ._EVAL_17(tlb__EVAL_17),
    ._EVAL_18(tlb__EVAL_18),
    ._EVAL_19(tlb__EVAL_19),
    ._EVAL_20(tlb__EVAL_20),
    ._EVAL_21(tlb__EVAL_21),
    ._EVAL_22(tlb__EVAL_22),
    ._EVAL_23(tlb__EVAL_23),
    ._EVAL_24(tlb__EVAL_24),
    ._EVAL_25(tlb__EVAL_25),
    ._EVAL_26(tlb__EVAL_26),
    ._EVAL_27(tlb__EVAL_27),
    ._EVAL_28(tlb__EVAL_28),
    ._EVAL_29(tlb__EVAL_29),
    ._EVAL_30(tlb__EVAL_30),
    ._EVAL_31(tlb__EVAL_31),
    ._EVAL_32(tlb__EVAL_32),
    ._EVAL_33(tlb__EVAL_33),
    ._EVAL_34(tlb__EVAL_34),
    ._EVAL_35(tlb__EVAL_35),
    ._EVAL_36(tlb__EVAL_36),
    ._EVAL_37(tlb__EVAL_37),
    ._EVAL_38(tlb__EVAL_38),
    ._EVAL_39(tlb__EVAL_39),
    ._EVAL_40(tlb__EVAL_40),
    ._EVAL_41(tlb__EVAL_41),
    ._EVAL_42(tlb__EVAL_42),
    ._EVAL_43(tlb__EVAL_43),
    ._EVAL_44(tlb__EVAL_44),
    ._EVAL_45(tlb__EVAL_45),
    ._EVAL_46(tlb__EVAL_46),
    ._EVAL_47(tlb__EVAL_47),
    ._EVAL_48(tlb__EVAL_48),
    ._EVAL_49(tlb__EVAL_49),
    ._EVAL_50(tlb__EVAL_50),
    ._EVAL_51(tlb__EVAL_51),
    ._EVAL_52(tlb__EVAL_52),
    ._EVAL_53(tlb__EVAL_53),
    ._EVAL_54(tlb__EVAL_54),
    ._EVAL_55(tlb__EVAL_55),
    ._EVAL_56(tlb__EVAL_56),
    ._EVAL_57(tlb__EVAL_57),
    ._EVAL_58(tlb__EVAL_58),
    ._EVAL_59(tlb__EVAL_59),
    ._EVAL_60(tlb__EVAL_60),
    ._EVAL_61(tlb__EVAL_61),
    ._EVAL_62(tlb__EVAL_62),
    ._EVAL_63(tlb__EVAL_63),
    ._EVAL_64(tlb__EVAL_64),
    ._EVAL_65(tlb__EVAL_65),
    ._EVAL_66(tlb__EVAL_66),
    ._EVAL_67(tlb__EVAL_67),
    ._EVAL_68(tlb__EVAL_68),
    ._EVAL_69(tlb__EVAL_69),
    ._EVAL_70(tlb__EVAL_70),
    ._EVAL_71(tlb__EVAL_71)
  );
  SiFive__EVAL_255 q (
    ._EVAL(q__EVAL),
    ._EVAL_0(q__EVAL_0),
    ._EVAL_1(q__EVAL_1),
    ._EVAL_2(q__EVAL_2),
    ._EVAL_3(q__EVAL_3),
    ._EVAL_4(q__EVAL_4),
    ._EVAL_5(q__EVAL_5),
    ._EVAL_6(q__EVAL_6),
    ._EVAL_7(q__EVAL_7),
    ._EVAL_8(q__EVAL_8),
    ._EVAL_9(q__EVAL_9),
    ._EVAL_10(q__EVAL_10),
    ._EVAL_11(q__EVAL_11),
    ._EVAL_12(q__EVAL_12),
    ._EVAL_13(q__EVAL_13),
    ._EVAL_14(q__EVAL_14),
    ._EVAL_15(q__EVAL_15),
    ._EVAL_16(q__EVAL_16),
    ._EVAL_17(q__EVAL_17),
    ._EVAL_18(q__EVAL_18),
    ._EVAL_19(q__EVAL_19)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR (
    ._EVAL(MaxPeriodFibonacciLFSR__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR__EVAL_17)
  );
  SiFive__EVAL_258 amoalu (
    ._EVAL(amoalu__EVAL),
    ._EVAL_0(amoalu__EVAL_0),
    ._EVAL_1(amoalu__EVAL_1),
    ._EVAL_2(amoalu__EVAL_2),
    ._EVAL_3(amoalu__EVAL_3)
  );
  SiFive__EVAL_344 tag_array (
    ._EVAL(tag_array__EVAL),
    ._EVAL_0(tag_array__EVAL_0),
    ._EVAL_1(tag_array__EVAL_1),
    ._EVAL_2(tag_array__EVAL_2),
    ._EVAL_3(tag_array__EVAL_3),
    ._EVAL_4(tag_array__EVAL_4),
    ._EVAL_5(tag_array__EVAL_5),
    ._EVAL_6(tag_array__EVAL_6),
    ._EVAL_7(tag_array__EVAL_7),
    ._EVAL_8(tag_array__EVAL_8),
    ._EVAL_9(tag_array__EVAL_9),
    ._EVAL_10(tag_array__EVAL_10),
    ._EVAL_11(tag_array__EVAL_11),
    ._EVAL_12(tag_array__EVAL_12),
    ._EVAL_13(tag_array__EVAL_13),
    ._EVAL_14(tag_array__EVAL_14)
  );
  assign _EVAL_742 = _EVAL_872 == 1'h0;
  assign _EVAL_1415 = _EVAL_526 == 1'h0;
  assign _EVAL_1328 = _EVAL_1832 & _EVAL_1415;
  assign _EVAL_1088 = _EVAL_742 | _EVAL_1328;
  assign _EVAL_762 = {_EVAL_1122,_EVAL_655,_EVAL_357,_EVAL_1271,_EVAL_1350,_EVAL_613,_EVAL_332};
  assign _EVAL_409 = ~ _EVAL_762;
  assign _EVAL_1311 = {_EVAL_409, 1'h0};
  assign _EVAL_770 = _EVAL_1311[0];
  assign _EVAL_971 = _EVAL_1311[1];
  assign _EVAL_307 = _EVAL_1311[2];
  assign _EVAL_1715 = _EVAL_1311[3];
  assign _EVAL_1326 = _EVAL_1311[4];
  assign _EVAL_1303 = _EVAL_1311[5];
  assign _EVAL_1263 = _EVAL_1311[6];
  assign _EVAL_460 = _EVAL_1263 ? 3'h6 : 3'h7;
  assign _EVAL_885 = _EVAL_1303 ? 3'h5 : _EVAL_460;
  assign _EVAL_1535 = _EVAL_1326 ? 3'h4 : _EVAL_885;
  assign _EVAL_481 = _EVAL_1715 ? 3'h3 : _EVAL_1535;
  assign _EVAL_1777 = _EVAL_307 ? 3'h2 : _EVAL_481;
  assign _EVAL_855 = _EVAL_971 ? 3'h1 : _EVAL_1777;
  assign _EVAL_1117 = _EVAL_770 ? 3'h0 : _EVAL_855;
  assign _EVAL_535 = 8'h1 << _EVAL_1117;
  assign _EVAL_187 = _EVAL_535[7:1];
  assign _EVAL_661 = _EVAL_187[5];
  assign _EVAL_1627 = _EVAL_396 == 3'h1;
  assign _EVAL_476 = _EVAL_396 == 3'h6;
  assign _EVAL_1609 = _EVAL_1627 | _EVAL_476;
  assign _EVAL_731 = _EVAL_396 == 3'h2;
  assign _EVAL_1346 = _EVAL_731 ? 3'h5 : 3'h4;
  assign _EVAL_1484 = _EVAL_1609 ? 3'h7 : _EVAL_1346;
  assign _EVAL_696 = _EVAL_1484;
  assign _EVAL_605 = _EVAL_696[0];
  assign _EVAL_647 = _EVAL_1609 ? 4'h6 : _EVAL_1366;
  assign _EVAL_1686 = _EVAL_647;
  assign _EVAL_1022 = 23'hff << _EVAL_1686;
  assign _EVAL_1194 = _EVAL_1022[7:0];
  assign _EVAL_871 = ~ _EVAL_1194;
  assign _EVAL_908 = _EVAL_871[7:3];
  assign _EVAL_1523 = _EVAL_605 ? _EVAL_908 : 5'h0;
  assign _EVAL_1526 = _EVAL_502 - 5'h1;
  assign _EVAL_1306 = ~ _EVAL_1526;
  assign _EVAL_185 = _EVAL_1523 & _EVAL_1306;
  assign _EVAL_551 = {1'h0,_EVAL_185};
  assign _EVAL_1865 = _EVAL_396 == 3'h3;
  assign _EVAL_720 = _EVAL_396 == 3'h5;
  assign _EVAL_1610 = {_EVAL_598,_EVAL_1373};
  assign _EVAL_1679 = 4'h3 == _EVAL_1610;
  assign _EVAL_1132 = 4'h2 == _EVAL_1610;
  assign _EVAL_1217 = 4'h1 == _EVAL_1610;
  assign _EVAL_1253 = 4'h0 == _EVAL_1610;
  assign _EVAL_994 = 4'h7 == _EVAL_1610;
  assign _EVAL_733 = 4'h6 == _EVAL_1610;
  assign _EVAL_418 = 4'h5 == _EVAL_1610;
  assign _EVAL_1823 = 4'h4 == _EVAL_1610;
  assign _EVAL_1007 = 4'hb == _EVAL_1610;
  assign _EVAL_1685 = _EVAL_1823 ? 1'h0 : _EVAL_1007;
  assign _EVAL_1861 = _EVAL_418 ? 1'h0 : _EVAL_1685;
  assign _EVAL_231 = _EVAL_733 ? 1'h0 : _EVAL_1861;
  assign _EVAL_287 = _EVAL_994 ? 1'h1 : _EVAL_231;
  assign _EVAL_758 = _EVAL_1253 ? 1'h0 : _EVAL_287;
  assign _EVAL_1228 = _EVAL_1217 ? 1'h0 : _EVAL_758;
  assign _EVAL_1048 = _EVAL_1132 ? 1'h0 : _EVAL_1228;
  assign _EVAL_1098 = _EVAL_1679 ? 1'h1 : _EVAL_1048;
  assign _EVAL_1722 = _EVAL_1098 ? _EVAL_1104 : 1'h1;
  assign _EVAL_398 = _EVAL_1450 ? _EVAL_1722 : _EVAL_1104;
  assign _EVAL_1536 = _EVAL_720 ? 1'h1 : _EVAL_398;
  assign _EVAL_1458 = _EVAL_1865 ? 1'h1 : _EVAL_1536;
  assign _EVAL_804 = _EVAL_1458;
  assign _EVAL_1036 = _EVAL_86;
  assign _EVAL_1674 = _EVAL_1036 == 1'h0;
  assign _EVAL_1322 = _EVAL_804 & _EVAL_1674;
  assign _EVAL_1752 = {{1'd0}, _EVAL_356};
  assign _EVAL_1699 = {1'h0,_EVAL_1104};
  assign _EVAL_787 = _EVAL_1752 + _EVAL_1699;
  assign _EVAL_498 = _EVAL_1322 ? 2'h0 : _EVAL_787;
  assign _EVAL_1703 = {{4'd0}, _EVAL_498};
  assign _EVAL_1102 = _EVAL_551 + _EVAL_1703;
  assign _EVAL_1164 = _EVAL_1102[2:0];
  assign _EVAL_660 = {_EVAL_1164, 3'h0};
  assign _EVAL_1358 = _EVAL_155[1];
  assign _EVAL_463 = _EVAL_155[0];
  assign _EVAL_439 = _EVAL_1661 >= 2'h1;
  assign _EVAL_1511 = _EVAL_463 | _EVAL_439;
  assign _EVAL_196 = _EVAL_463 ? 1'h0 : 1'h1;
  assign _EVAL_977 = {_EVAL_1511,_EVAL_196};
  assign _EVAL_349 = _EVAL_1358 ? _EVAL_977 : 2'h0;
  assign _EVAL_812 = _EVAL_1661 >= 2'h2;
  assign _EVAL_976 = _EVAL_812 ? 2'h3 : 2'h0;
  assign _EVAL_1068 = _EVAL_349 | _EVAL_976;
  assign _EVAL_1283 = _EVAL_1358 ? 2'h0 : _EVAL_977;
  assign _EVAL_1653 = {_EVAL_1068,_EVAL_1283};
  assign _EVAL_1765 = _EVAL_1121 & _EVAL_1653;
  assign _EVAL_314 = 4'ha == _EVAL_1610;
  assign _EVAL_671 = 4'h9 == _EVAL_1610;
  assign _EVAL_450 = 4'h8 == _EVAL_1610;
  assign _EVAL_1186 = _EVAL_450 ? 3'h5 : 3'h0;
  assign _EVAL_1124 = _EVAL_671 ? 3'h2 : _EVAL_1186;
  assign _EVAL_346 = _EVAL_314 ? 3'h1 : _EVAL_1124;
  assign _EVAL_449 = _EVAL_1007 ? 3'h1 : _EVAL_346;
  assign _EVAL_1023 = _EVAL_1823 ? 3'h2 : _EVAL_449;
  assign _EVAL_593 = _EVAL_418 ? 3'h4 : _EVAL_1023;
  assign _EVAL_1337 = _EVAL_733 ? 3'h0 : _EVAL_593;
  assign _EVAL_442 = _EVAL_994 ? 3'h0 : _EVAL_1337;
  assign _EVAL_1110 = _EVAL_187[6];
  assign _EVAL_1191 = 5'hd == _EVAL_1325;
  assign _EVAL_368 = 5'he == _EVAL_1325;
  assign _EVAL_548 = 5'hf == _EVAL_1325;
  assign _EVAL_1333 = _EVAL_548 ? _EVAL_389 : 32'h0;
  assign _EVAL_688 = _EVAL_368 ? _EVAL_389 : _EVAL_1333;
  assign _EVAL_806 = _EVAL_1191 ? _EVAL_389 : _EVAL_688;
  assign _EVAL_1762 = _EVAL_1325 == 5'h7;
  assign _EVAL_760 = _EVAL_389[0];
  assign _EVAL_530 = _EVAL_981 == 2'h1;
  assign _EVAL_220 = _EVAL_389[1];
  assign _EVAL_1562 = _EVAL_1442 ? _EVAL_254 : 32'h0;
  assign _EVAL_552 = _EVAL_320[0];
  assign _EVAL_1876 = _EVAL_552 ? _EVAL_1709 : 32'h0;
  assign _EVAL_809 = _EVAL_320[1];
  assign _EVAL_567 = _EVAL_809 ? _EVAL_1527 : 32'h0;
  assign _EVAL_1084 = _EVAL_1876 | _EVAL_567;
  assign _EVAL_1214 = _EVAL_320[2];
  assign _EVAL_1581 = _EVAL_1214 ? _EVAL_1619 : 32'h0;
  assign _EVAL_1792 = _EVAL_1084 | _EVAL_1581;
  assign _EVAL_1126 = _EVAL_320[3];
  assign _EVAL_457 = _EVAL_1126 ? _EVAL_1431 : 32'h0;
  assign _EVAL_1177 = _EVAL_1792 | _EVAL_457;
  assign _EVAL_562 = _EVAL_1827[0];
  assign _EVAL_832 = _EVAL_562 ? _EVAL_367 : 32'h0;
  assign _EVAL_1349 = _EVAL_1827[1];
  assign _EVAL_159 = _EVAL_1349 ? _EVAL_359 : 32'h0;
  assign _EVAL_459 = _EVAL_832 | _EVAL_159;
  assign _EVAL_735 = _EVAL_1827[2];
  assign _EVAL_436 = _EVAL_735 ? _EVAL_293 : 32'h0;
  assign _EVAL_1872 = _EVAL_459 | _EVAL_436;
  assign _EVAL_1576 = _EVAL_1827[3];
  assign _EVAL_830 = _EVAL_1576 ? _EVAL_433 : 32'h0;
  assign _EVAL_1423 = _EVAL_1872 | _EVAL_830;
  assign _EVAL_483 = {_EVAL_1177,_EVAL_1423};
  assign _EVAL_507 = _EVAL_483[63:56];
  assign _EVAL_1143 = _EVAL_483[55:48];
  assign _EVAL_675 = _EVAL_483[47:40];
  assign _EVAL_1411 = _EVAL_483[39:32];
  assign _EVAL_525 = _EVAL_483[31:24];
  assign _EVAL_1862 = _EVAL_483[23:16];
  assign _EVAL_1236 = _EVAL_483[15:8];
  assign _EVAL_1080 = _EVAL_483[7:0];
  assign _EVAL_250 = {_EVAL_507,_EVAL_1143,_EVAL_675,_EVAL_1411,_EVAL_525,_EVAL_1862,_EVAL_1236,_EVAL_1080};
  assign _EVAL_680 = _EVAL_250[31:0];
  assign _EVAL_738 = _EVAL_250[63:32];
  assign _EVAL_353 = _EVAL_680 | _EVAL_738;
  assign _EVAL_419 = _EVAL_1562 | _EVAL_353;
  assign _EVAL_1612 = _EVAL_419[31:16];
  assign _EVAL_1281 = _EVAL_419[15:0];
  assign _EVAL_623 = _EVAL_220 ? _EVAL_1612 : _EVAL_1281;
  assign _EVAL_1597 = _EVAL_623[15];
  assign _EVAL_903 = _EVAL_165 & _EVAL_1597;
  assign _EVAL_601 = _EVAL_903 ? 16'hffff : 16'h0;
  assign _EVAL_1434 = _EVAL_530 ? _EVAL_601 : _EVAL_1612;
  assign _EVAL_689 = {_EVAL_1434,_EVAL_623};
  assign _EVAL_1105 = _EVAL_689[15:8];
  assign _EVAL_1290 = _EVAL_689[7:0];
  assign _EVAL_912 = _EVAL_760 ? _EVAL_1105 : _EVAL_1290;
  assign _EVAL_724 = _EVAL_1762 ? 8'h0 : _EVAL_912;
  assign _EVAL_1723 = {_EVAL_64,_EVAL_143,_EVAL_110,_EVAL_111,_EVAL_31,_EVAL_33};
  assign _EVAL_878 = _EVAL_1723 != 6'h0;
  assign _EVAL_170 = _EVAL_878 == 1'h0;
  assign _EVAL_794 = _EVAL_1109 & _EVAL_170;
  assign _EVAL_780 = _EVAL_794 & _EVAL_263;
  assign _EVAL_404 = _EVAL_1325 == 5'h1;
  assign _EVAL_1552 = _EVAL_1325 == 5'h11;
  assign _EVAL_1871 = _EVAL_404 | _EVAL_1552;
  assign _EVAL_692 = _EVAL_1871 | _EVAL_1762;
  assign _EVAL_486 = _EVAL_1325 == 5'h4;
  assign _EVAL_882 = _EVAL_1325 == 5'h9;
  assign _EVAL_805 = _EVAL_486 | _EVAL_882;
  assign _EVAL_1244 = _EVAL_1325 == 5'ha;
  assign _EVAL_1384 = _EVAL_805 | _EVAL_1244;
  assign _EVAL_986 = _EVAL_1325 == 5'hb;
  assign _EVAL_299 = _EVAL_1384 | _EVAL_986;
  assign _EVAL_1368 = _EVAL_1325 == 5'h8;
  assign _EVAL_1158 = _EVAL_1325 == 5'hc;
  assign _EVAL_710 = _EVAL_1368 | _EVAL_1158;
  assign _EVAL_440 = _EVAL_1325 == 5'hd;
  assign _EVAL_1717 = _EVAL_710 | _EVAL_440;
  assign _EVAL_756 = _EVAL_1325 == 5'he;
  assign _EVAL_1720 = _EVAL_1717 | _EVAL_756;
  assign _EVAL_873 = _EVAL_1325 == 5'hf;
  assign _EVAL_223 = _EVAL_1720 | _EVAL_873;
  assign _EVAL_925 = _EVAL_299 | _EVAL_223;
  assign _EVAL_587 = _EVAL_692 | _EVAL_925;
  assign _EVAL_1448 = _EVAL_1325 == 5'h3;
  assign _EVAL_1003 = _EVAL_587 | _EVAL_1448;
  assign _EVAL_511 = _EVAL_1325 == 5'h6;
  assign _EVAL_815 = _EVAL_1003 | _EVAL_511;
  assign _EVAL_840 = {_EVAL_587,_EVAL_815,_EVAL_951};
  assign _EVAL_944 = 4'h3 == _EVAL_840;
  assign _EVAL_1692 = 4'h2 == _EVAL_840;
  assign _EVAL_1371 = 4'h1 == _EVAL_840;
  assign _EVAL_216 = 4'h7 == _EVAL_840;
  assign _EVAL_1667 = 4'h6 == _EVAL_840;
  assign _EVAL_252 = 4'hf == _EVAL_840;
  assign _EVAL_201 = 4'he == _EVAL_840;
  assign _EVAL_1247 = _EVAL_252 ? 1'h1 : _EVAL_201;
  assign _EVAL_490 = _EVAL_1667 ? 1'h1 : _EVAL_1247;
  assign _EVAL_238 = _EVAL_216 ? 1'h1 : _EVAL_490;
  assign _EVAL_1364 = _EVAL_1371 ? 1'h1 : _EVAL_238;
  assign _EVAL_814 = _EVAL_1692 ? 1'h1 : _EVAL_1364;
  assign _EVAL_1376 = _EVAL_944 ? 1'h1 : _EVAL_814;
  assign _EVAL_1663 = _EVAL_780 & _EVAL_1376;
  assign _EVAL_259 = _EVAL_1325 == 5'h0;
  assign _EVAL_1826 = _EVAL_259 | _EVAL_511;
  assign _EVAL_1226 = _EVAL_1826 | _EVAL_1762;
  assign _EVAL_1018 = _EVAL_1226 | _EVAL_925;
  assign _EVAL_1628 = _EVAL_1018 | _EVAL_587;
  assign _EVAL_1850 = _EVAL_1663 & _EVAL_1628;
  assign _EVAL_1781 = _EVAL_1850 & _EVAL_587;
  assign _EVAL_210 = _EVAL_54 == 1'h0;
  assign _EVAL_394 = _EVAL_1781 & _EVAL_210;
  assign _EVAL_209 = _EVAL_394 | _EVAL_1252;
  assign _EVAL_1184 = _EVAL_893 > 7'h3;
  assign _EVAL_714 = _EVAL_389[31:6];
  assign _EVAL_1857 = _EVAL_632 == _EVAL_714;
  assign _EVAL_571 = _EVAL_1184 & _EVAL_1857;
  assign _EVAL_1698 = _EVAL_571 == 1'h0;
  assign _EVAL_1395 = _EVAL_1762 & _EVAL_1698;
  assign _EVAL_1025 = _EVAL_1395 == 1'h0;
  assign _EVAL_860 = _EVAL_1781 & _EVAL_1025;
  assign _EVAL_1753 = _EVAL_860 & _EVAL_210;
  assign _EVAL_153 = _EVAL_1753 | _EVAL_1252;
  assign _EVAL_456 = tag_array__EVAL;
  assign _EVAL_1561 = _EVAL_456[21:20];
  assign _EVAL_469 = _EVAL_1561 > 2'h0;
  assign _EVAL_1418 = _EVAL_456[19:0];
  assign _EVAL_1483 = tlb__EVAL_38[31:12];
  assign _EVAL_1825 = _EVAL_1418 == _EVAL_1483;
  assign _EVAL_424 = _EVAL_469 & _EVAL_1825;
  assign _EVAL_1010 = tag_array__EVAL_5;
  assign _EVAL_313 = _EVAL_1010[21:20];
  assign _EVAL_1279 = _EVAL_313 > 2'h0;
  assign _EVAL_799 = _EVAL_1010[19:0];
  assign _EVAL_446 = _EVAL_799 == _EVAL_1483;
  assign _EVAL_1807 = _EVAL_1279 & _EVAL_446;
  assign _EVAL_1277 = tag_array__EVAL_3;
  assign _EVAL_1264 = _EVAL_1277[21:20];
  assign _EVAL_1449 = _EVAL_1264 > 2'h0;
  assign _EVAL_1218 = _EVAL_1277[19:0];
  assign _EVAL_1622 = _EVAL_1218 == _EVAL_1483;
  assign _EVAL_1445 = _EVAL_1449 & _EVAL_1622;
  assign _EVAL_407 = tag_array__EVAL_11;
  assign _EVAL_693 = _EVAL_407[21:20];
  assign _EVAL_437 = _EVAL_693 > 2'h0;
  assign _EVAL_545 = _EVAL_407[19:0];
  assign _EVAL_317 = _EVAL_545 == _EVAL_1483;
  assign _EVAL_1242 = _EVAL_437 & _EVAL_317;
  assign _EVAL_258 = {_EVAL_424,_EVAL_1807,_EVAL_1445,_EVAL_1242};
  assign _EVAL_722 = _EVAL_951 > 2'h0;
  assign _EVAL_1858 = _EVAL_722 ? _EVAL_951 : _EVAL_1200;
  assign _EVAL_236 = _EVAL_1100 == 1'h0;
  assign _EVAL_1642 = _EVAL_236 & _EVAL_210;
  assign _EVAL_564 = _EVAL_800;
  assign _EVAL_1534 = _EVAL_389[31:12];
  assign _EVAL_1258 = {2'h0,_EVAL_1534};
  assign _EVAL_1780 = 4'h0 == _EVAL_840;
  assign _EVAL_932 = 4'h5 == _EVAL_840;
  assign _EVAL_1363 = 4'h4 == _EVAL_840;
  assign _EVAL_1758 = 4'hd == _EVAL_840;
  assign _EVAL_1352 = 4'hc == _EVAL_840;
  assign _EVAL_1646 = _EVAL_1352 ? 2'h1 : 2'h0;
  assign _EVAL_334 = _EVAL_1758 ? 2'h2 : _EVAL_1646;
  assign _EVAL_702 = _EVAL_1363 ? 2'h1 : _EVAL_334;
  assign _EVAL_1009 = _EVAL_932 ? 2'h2 : _EVAL_702;
  assign _EVAL_1833 = _EVAL_1780 ? 2'h0 : _EVAL_1009;
  assign _EVAL_1251 = _EVAL_201 ? 2'h3 : _EVAL_1833;
  assign _EVAL_1604 = _EVAL_252 ? 2'h3 : _EVAL_1251;
  assign _EVAL_1704 = _EVAL_1667 ? 2'h2 : _EVAL_1604;
  assign _EVAL_662 = _EVAL_216 ? 2'h3 : _EVAL_1704;
  assign _EVAL_1867 = _EVAL_1371 ? 2'h1 : _EVAL_662;
  assign _EVAL_1701 = _EVAL_1692 ? 2'h2 : _EVAL_1867;
  assign _EVAL_1014 = _EVAL_944 ? 2'h3 : _EVAL_1701;
  assign _EVAL_1478 = _EVAL_951 == _EVAL_1014;
  assign _EVAL_309 = _EVAL_1478 == 1'h0;
  assign _EVAL_792 = _EVAL_1850 & _EVAL_309;
  assign _EVAL_154 = {_EVAL_1014,_EVAL_1534};
  assign _EVAL_1399 = _EVAL_5;
  assign _EVAL_679 = _EVAL_1399 == 3'h4;
  assign _EVAL_373 = _EVAL_1399 == 3'h5;
  assign _EVAL_1564 = _EVAL_679 | _EVAL_373;
  assign _EVAL_1618 = _EVAL_659 == 5'h1;
  assign _EVAL_1738 = _EVAL_1399[0];
  assign _EVAL_431 = _EVAL_99;
  assign _EVAL_1745 = 23'hff << _EVAL_431;
  assign _EVAL_1072 = _EVAL_1745[7:0];
  assign _EVAL_1557 = ~ _EVAL_1072;
  assign _EVAL_462 = _EVAL_1557[7:3];
  assign _EVAL_345 = _EVAL_1738 ? _EVAL_462 : 5'h0;
  assign _EVAL_681 = _EVAL_345 == 5'h0;
  assign _EVAL_553 = _EVAL_1618 | _EVAL_681;
  assign _EVAL_993 = _EVAL_1399 == 3'h1;
  assign _EVAL_1841 = _EVAL_124 == 1'h0;
  assign _EVAL_990 = _EVAL_993 & _EVAL_1841;
  assign _EVAL_620 = _EVAL_1109 & _EVAL_587;
  assign _EVAL_946 = _EVAL_620 | _EVAL_1252;
  assign _EVAL_292 = _EVAL_946 & _EVAL_322;
  assign _EVAL_1413 = _EVAL_204 == 5'h1;
  assign _EVAL_1542 = _EVAL_204 == 5'h11;
  assign _EVAL_400 = _EVAL_1413 | _EVAL_1542;
  assign _EVAL_470 = _EVAL_204 == 5'h7;
  assign _EVAL_602 = _EVAL_400 | _EVAL_470;
  assign _EVAL_910 = _EVAL_204 == 5'h4;
  assign _EVAL_1265 = _EVAL_204 == 5'h9;
  assign _EVAL_405 = _EVAL_910 | _EVAL_1265;
  assign _EVAL_608 = _EVAL_204 == 5'ha;
  assign _EVAL_697 = _EVAL_405 | _EVAL_608;
  assign _EVAL_1398 = _EVAL_204 == 5'hb;
  assign _EVAL_218 = _EVAL_697 | _EVAL_1398;
  assign _EVAL_1406 = _EVAL_204 == 5'h8;
  assign _EVAL_364 = _EVAL_204 == 5'hc;
  assign _EVAL_594 = _EVAL_1406 | _EVAL_364;
  assign _EVAL_1155 = _EVAL_204 == 5'hd;
  assign _EVAL_271 = _EVAL_594 | _EVAL_1155;
  assign _EVAL_1845 = _EVAL_204 == 5'he;
  assign _EVAL_718 = _EVAL_271 | _EVAL_1845;
  assign _EVAL_466 = _EVAL_204 == 5'hf;
  assign _EVAL_1660 = _EVAL_718 | _EVAL_466;
  assign _EVAL_978 = _EVAL_218 | _EVAL_1660;
  assign _EVAL_1211 = _EVAL_602 | _EVAL_978;
  assign _EVAL_172 = _EVAL_1697 & _EVAL_1211;
  assign _EVAL_1127 = _EVAL_172 | _EVAL_1486;
  assign _EVAL_838 = _EVAL_292 & _EVAL_1127;
  assign _EVAL_1726 = _EVAL_1781 | _EVAL_1252;
  assign _EVAL_778 = _EVAL_1486 == 1'h0;
  assign _EVAL_754 = _EVAL_1726 & _EVAL_778;
  assign _EVAL_590 = _EVAL_754 | _EVAL_322;
  assign _EVAL_1207 = _EVAL_135 == 5'h1;
  assign _EVAL_913 = _EVAL_135 == 5'h3;
  assign _EVAL_261 = _EVAL_1207 | _EVAL_913;
  assign _EVAL_699 = _EVAL_261 == 1'h0;
  assign _EVAL_1160 = _EVAL_37 & _EVAL_699;
  assign _EVAL_194 = _EVAL_1160 == 1'h0;
  assign _EVAL_199 = _EVAL_926 | _EVAL_1450;
  assign _EVAL_849 = _EVAL_396 != 3'h0;
  assign _EVAL_1118 = _EVAL_199 | _EVAL_849;
  assign _EVAL_583 = _EVAL_1118 | _EVAL_907;
  assign _EVAL_435 = _EVAL_194 | _EVAL_583;
  assign _EVAL_555 = _EVAL_590 & _EVAL_435;
  assign _EVAL_822 = _EVAL_838 | _EVAL_555;
  assign _EVAL_1302 = _EVAL_822 == 1'h0;
  assign _EVAL_709 = _EVAL_1302 == 1'h0;
  assign _EVAL_1725 = _EVAL_373 & _EVAL_709;
  assign _EVAL_1438 = _EVAL_659 == 5'h0;
  assign _EVAL_1270 = _EVAL_1438 == 1'h0;
  assign _EVAL_1757 = _EVAL_10;
  assign _EVAL_816 = _EVAL_1270 | _EVAL_1757;
  assign _EVAL_927 = _EVAL_1609 == 1'h0;
  assign _EVAL_1782 = _EVAL_816 & _EVAL_927;
  assign _EVAL_1669 = _EVAL_1564 ? _EVAL_1782 : 1'h1;
  assign _EVAL_193 = _EVAL_1725 ? 1'h0 : _EVAL_1669;
  assign _EVAL_306 = _EVAL_990 ? 1'h0 : _EVAL_193;
  assign _EVAL_1016 = _EVAL_306;
  assign _EVAL_1221 = _EVAL_107;
  assign _EVAL_1718 = _EVAL_1016 & _EVAL_1221;
  assign _EVAL_1020 = _EVAL_553 & _EVAL_1718;
  assign _EVAL_1166 = _EVAL_1564 & _EVAL_1020;
  assign _EVAL_1129 = _EVAL_36;
  assign _EVAL_1343 = _EVAL_1129 == 1'h0;
  assign _EVAL_1788 = _EVAL_1166 & _EVAL_1343;
  assign _EVAL_448 = _EVAL_112;
  assign _EVAL_455 = {_EVAL_587,_EVAL_815,_EVAL_448};
  assign _EVAL_818 = 4'h1 == _EVAL_455;
  assign _EVAL_1241 = 4'h0 == _EVAL_455;
  assign _EVAL_518 = 4'h4 == _EVAL_455;
  assign _EVAL_1809 = 4'hc == _EVAL_455;
  assign _EVAL_572 = _EVAL_1809 ? 2'h3 : 2'h0;
  assign _EVAL_184 = _EVAL_518 ? 2'h2 : _EVAL_572;
  assign _EVAL_565 = _EVAL_1241 ? 2'h2 : _EVAL_184;
  assign _EVAL_782 = _EVAL_818 ? 2'h1 : _EVAL_565;
  assign _EVAL_1459 = {_EVAL_782,_EVAL_1534};
  assign _EVAL_311 = _EVAL_396 == 3'h7;
  assign _EVAL_1273 = _EVAL_476 | _EVAL_311;
  assign _EVAL_163 = {2'h2,_EVAL_1858};
  assign _EVAL_1785 = 4'h3 == _EVAL_163;
  assign _EVAL_687 = 4'h2 == _EVAL_163;
  assign _EVAL_1493 = 4'h1 == _EVAL_163;
  assign _EVAL_789 = 4'h0 == _EVAL_163;
  assign _EVAL_179 = 4'h7 == _EVAL_163;
  assign _EVAL_381 = 4'h6 == _EVAL_163;
  assign _EVAL_1391 = 4'h5 == _EVAL_163;
  assign _EVAL_727 = _EVAL_1391 ? 2'h1 : 2'h0;
  assign _EVAL_468 = _EVAL_381 ? 2'h1 : _EVAL_727;
  assign _EVAL_1386 = _EVAL_179 ? 2'h1 : _EVAL_468;
  assign _EVAL_1440 = _EVAL_789 ? 2'h0 : _EVAL_1386;
  assign _EVAL_443 = _EVAL_1493 ? 2'h1 : _EVAL_1440;
  assign _EVAL_1039 = _EVAL_687 ? 2'h2 : _EVAL_443;
  assign _EVAL_510 = _EVAL_1785 ? 2'h2 : _EVAL_1039;
  assign _EVAL_491 = _EVAL_418 ? 2'h1 : 2'h0;
  assign _EVAL_983 = _EVAL_733 ? 2'h1 : _EVAL_491;
  assign _EVAL_1336 = _EVAL_994 ? 2'h1 : _EVAL_983;
  assign _EVAL_1066 = _EVAL_1253 ? 2'h0 : _EVAL_1336;
  assign _EVAL_1112 = _EVAL_1217 ? 2'h1 : _EVAL_1066;
  assign _EVAL_494 = _EVAL_1132 ? 2'h2 : _EVAL_1112;
  assign _EVAL_324 = _EVAL_1679 ? 2'h2 : _EVAL_494;
  assign _EVAL_1401 = _EVAL_1609 ? _EVAL_510 : _EVAL_324;
  assign _EVAL_1293 = _EVAL_1107;
  assign _EVAL_707 = _EVAL_1293[31:12];
  assign _EVAL_930 = {_EVAL_1401,_EVAL_707};
  assign _EVAL_1237 = _EVAL_1422 & _EVAL_236;
  assign _EVAL_788 = _EVAL_930;
  assign _EVAL_403 = _EVAL_396 == 3'h4;
  assign _EVAL_1524 = _EVAL_14;
  assign _EVAL_694 = _EVAL_1032 > 3'h0;
  assign _EVAL_1027 = _EVAL_694 | _EVAL_1184;
  assign _EVAL_824 = _EVAL_1027 == 1'h0;
  assign _EVAL_509 = _EVAL_893 > 7'h0;
  assign _EVAL_242 = _EVAL_1184 == 1'h0;
  assign _EVAL_1206 = _EVAL_509 & _EVAL_242;
  assign _EVAL_1605 = _EVAL_824 | _EVAL_1206;
  assign _EVAL_1481 = _EVAL_1524 & _EVAL_1605;
  assign _EVAL_1131 = _EVAL_403 ? 1'h1 : _EVAL_1481;
  assign _EVAL_854 = _EVAL_930;
  assign _EVAL_1354 = _EVAL_930;
  assign _EVAL_1770 = _EVAL_1131 ? _EVAL_854 : _EVAL_1354;
  assign _EVAL_825 = _EVAL_1237 ? _EVAL_788 : _EVAL_1770;
  assign _EVAL_1378 = _EVAL_1273 ? _EVAL_930 : _EVAL_825;
  assign _EVAL_1215 = _EVAL_1788 ? _EVAL_1459 : _EVAL_1378;
  assign _EVAL_972 = _EVAL_792 ? _EVAL_154 : _EVAL_1215;
  assign _EVAL_1607 = _EVAL_564 ? _EVAL_1258 : _EVAL_972;
  assign _EVAL_1430 = _EVAL_1373 > 2'h0;
  assign _EVAL_705 = _EVAL_502 == 5'h1;
  assign _EVAL_219 = _EVAL_1523 == 5'h0;
  assign _EVAL_1086 = _EVAL_705 | _EVAL_219;
  assign _EVAL_531 = _EVAL_1036 & _EVAL_804;
  assign _EVAL_560 = _EVAL_1086 & _EVAL_531;
  assign _EVAL_1601 = _EVAL_560 == 1'h0;
  assign _EVAL_428 = _EVAL_1430 ? 1'h1 : _EVAL_1601;
  assign _EVAL_1455 = _EVAL_187[4];
  assign _EVAL_561 = _EVAL_389[11:0];
  assign _EVAL_284 = _EVAL_780 & _EVAL_1628;
  assign _EVAL_1462 = _EVAL_1376 == 1'h0;
  assign _EVAL_791 = _EVAL_284 & _EVAL_1462;
  assign _EVAL_1611 = _EVAL_559 == 1'h0;
  assign _EVAL_1687 = _EVAL_791 & _EVAL_1611;
  assign _EVAL_465 = _EVAL_322 ? _EVAL_1121 : _EVAL_393;
  assign _EVAL_736 = _EVAL_465[2];
  assign _EVAL_547 = _EVAL_548 ? 3'h2 : 3'h0;
  assign _EVAL_169 = _EVAL_368 ? 3'h2 : _EVAL_547;
  assign _EVAL_240 = _EVAL_1221 & _EVAL_1438;
  assign _EVAL_344 = _EVAL_240 & _EVAL_1564;
  assign _EVAL_191 = _EVAL_344 & _EVAL_927;
  assign _EVAL_1820 = _EVAL_1725 ? 1'h0 : _EVAL_191;
  assign _EVAL_276 = _EVAL_1820;
  assign _EVAL_1151 = {_EVAL_506,_EVAL_730,_EVAL_1195,_EVAL_763};
  assign _EVAL_899 = _EVAL_322 ? _EVAL_1151 : _EVAL_1096;
  assign _EVAL_752 = {_EVAL_899,_EVAL_899};
  assign _EVAL_865 = _EVAL_752[7:0];
  assign _EVAL_331 = _EVAL_187[1];
  assign _EVAL_180 = _EVAL_1399 == 3'h0;
  assign _EVAL_1457 = _EVAL_993 | _EVAL_180;
  assign _EVAL_796 = _EVAL_1399 == 3'h2;
  assign _EVAL_264 = _EVAL_1457 | _EVAL_796;
  assign _EVAL_513 = _EVAL_66;
  assign _EVAL_960 = 8'h1 << _EVAL_513;
  assign _EVAL_1769 = _EVAL_960[7:1];
  assign _EVAL_1348 = _EVAL_1769[1];
  assign _EVAL_176 = _EVAL_1348 & _EVAL_553;
  assign _EVAL_1632 = q__EVAL_8;
  assign _EVAL_1736 = _EVAL_1088 == 1'h0;
  assign _EVAL_672 = _EVAL_1687 & _EVAL_1736;
  assign _EVAL_467 = _EVAL_762 != 7'h0;
  assign _EVAL_1475 = _EVAL_467 == 1'h0;
  assign _EVAL_453 = _EVAL_672 & _EVAL_1475;
  assign _EVAL_1205 = 4'h4 == _EVAL_163;
  assign _EVAL_1170 = 4'hb == _EVAL_163;
  assign _EVAL_970 = _EVAL_1205 ? 1'h0 : _EVAL_1170;
  assign _EVAL_1464 = _EVAL_1391 ? 1'h0 : _EVAL_970;
  assign _EVAL_901 = _EVAL_381 ? 1'h0 : _EVAL_1464;
  assign _EVAL_267 = _EVAL_179 ? 1'h1 : _EVAL_901;
  assign _EVAL_884 = _EVAL_789 ? 1'h0 : _EVAL_267;
  assign _EVAL_870 = _EVAL_1493 ? 1'h0 : _EVAL_884;
  assign _EVAL_862 = _EVAL_687 ? 1'h0 : _EVAL_870;
  assign _EVAL_406 = _EVAL_1785 ? 1'h1 : _EVAL_862;
  assign _EVAL_497 = _EVAL_406 == 1'h0;
  assign _EVAL_568 = _EVAL_453 & _EVAL_497;
  assign _EVAL_416 = _EVAL_1687 & _EVAL_1088;
  assign _EVAL_249 = _EVAL_762 == 7'h7f;
  assign _EVAL_1672 = _EVAL_249 == 1'h0;
  assign _EVAL_174 = _EVAL_416 & _EVAL_1672;
  assign _EVAL_445 = _EVAL_568 | _EVAL_174;
  assign _EVAL_1005 = _EVAL_210 & _EVAL_445;
  assign _EVAL_1658 = _EVAL_1632 & _EVAL_1005;
  assign _EVAL_382 = _EVAL_250;
  assign _EVAL_935 = _EVAL_1221 & _EVAL_373;
  assign _EVAL_496 = _EVAL_935 & _EVAL_927;
  assign _EVAL_1061 = _EVAL_822 | _EVAL_496;
  assign _EVAL_813 = _EVAL_1627 | _EVAL_731;
  assign _EVAL_779 = _EVAL_1102 < 6'h8;
  assign _EVAL_1567 = _EVAL_813 & _EVAL_779;
  assign _EVAL_1369 = _EVAL_1061 | _EVAL_1567;
  assign _EVAL_546 = _EVAL_1369 == 1'h0;
  assign _EVAL_1520 = _EVAL_546 == 1'h0;
  assign _EVAL_1295 = 4'ha == _EVAL_163;
  assign _EVAL_817 = 4'h9 == _EVAL_163;
  assign _EVAL_784 = 4'h8 == _EVAL_163;
  assign _EVAL_454 = _EVAL_784 ? 3'h5 : 3'h0;
  assign _EVAL_1623 = _EVAL_817 ? 3'h2 : _EVAL_454;
  assign _EVAL_622 = _EVAL_1295 ? 3'h1 : _EVAL_1623;
  assign _EVAL_1577 = _EVAL_1170 ? 3'h1 : _EVAL_622;
  assign _EVAL_1299 = _EVAL_1205 ? 3'h2 : _EVAL_1577;
  assign _EVAL_711 = _EVAL_1391 ? 3'h4 : _EVAL_1299;
  assign _EVAL_691 = _EVAL_381 ? 3'h0 : _EVAL_711;
  assign _EVAL_734 = _EVAL_179 ? 3'h0 : _EVAL_691;
  assign _EVAL_615 = _EVAL_1060[7:6];
  assign _EVAL_207 = {MaxPeriodFibonacciLFSR__EVAL_12,MaxPeriodFibonacciLFSR__EVAL_11,MaxPeriodFibonacciLFSR__EVAL_3,MaxPeriodFibonacciLFSR__EVAL_16,MaxPeriodFibonacciLFSR__EVAL_8,MaxPeriodFibonacciLFSR__EVAL_10,MaxPeriodFibonacciLFSR__EVAL_14,MaxPeriodFibonacciLFSR__EVAL_7};
  assign _EVAL_1710 = {MaxPeriodFibonacciLFSR__EVAL_0,MaxPeriodFibonacciLFSR__EVAL_17,MaxPeriodFibonacciLFSR__EVAL_1,MaxPeriodFibonacciLFSR__EVAL,MaxPeriodFibonacciLFSR__EVAL_5,MaxPeriodFibonacciLFSR__EVAL_4,MaxPeriodFibonacciLFSR__EVAL_6,MaxPeriodFibonacciLFSR__EVAL_2,_EVAL_207};
  assign _EVAL_606 = _EVAL_1710[0];
  assign _EVAL_524 = _EVAL_1710[1];
  assign _EVAL_1819 = _EVAL_1710[2];
  assign _EVAL_1312 = _EVAL_1710[3];
  assign _EVAL_634 = _EVAL_1710[4];
  assign _EVAL_1267 = _EVAL_1710[5];
  assign _EVAL_1298 = _EVAL_1710[6];
  assign _EVAL_1517 = _EVAL_1710[7];
  assign _EVAL_1187 = _EVAL_1710[8];
  assign _EVAL_1389 = _EVAL_1710[9];
  assign _EVAL_479 = _EVAL_1710[10];
  assign _EVAL_1313 = _EVAL_1710[11];
  assign _EVAL_1474 = _EVAL_1710[12];
  assign _EVAL_412 = _EVAL_1710[13];
  assign _EVAL_1063 = _EVAL_1710[14];
  assign _EVAL_580 = _EVAL_1710[15];
  assign _EVAL_698 = {_EVAL_1187,_EVAL_1389,_EVAL_479,_EVAL_1313,_EVAL_1474,_EVAL_412,_EVAL_1063,_EVAL_580};
  assign _EVAL_947 = {_EVAL_606,_EVAL_524,_EVAL_1819,_EVAL_1312,_EVAL_634,_EVAL_1267,_EVAL_1298,_EVAL_1517,_EVAL_698};
  assign _EVAL_1556 = _EVAL_947[1:0];
  assign _EVAL_426 = _EVAL_1422 ? _EVAL_615 : _EVAL_1556;
  assign _EVAL_563 = _EVAL_426 == 2'h1;
  assign _EVAL_1046 = _EVAL_187[3];
  assign _EVAL_1062 = 4'h1 << _EVAL_746;
  assign _EVAL_1838 = _EVAL_722 ? _EVAL_277 : _EVAL_1062;
  assign _EVAL_1181 = _EVAL_1107[11:6];
  assign _EVAL_658 = {_EVAL_1181, 6'h0};
  assign _EVAL_945 = _EVAL_71 == 1'h0;
  assign _EVAL_1315 = _EVAL_1697 & _EVAL_945;
  assign _EVAL_1476 = _EVAL_20;
  assign _EVAL_1409 = _EVAL_1476 ^ _EVAL_982;
  assign _EVAL_851 = _EVAL_1409[11:6];
  assign _EVAL_1097 = _EVAL_851 == 6'h0;
  assign _EVAL_923 = _EVAL_559 & _EVAL_1097;
  assign _EVAL_217 = _EVAL_1118 | _EVAL_923;
  assign _EVAL_1775 = _EVAL_217 | _EVAL_1319;
  assign _EVAL_521 = _EVAL_1027 | _EVAL_1775;
  assign _EVAL_900 = _EVAL_659 - 5'h1;
  assign _EVAL_168 = ~ _EVAL_900;
  assign _EVAL_294 = _EVAL_345 & _EVAL_168;
  assign _EVAL_569 = {_EVAL_294, 3'h0};
  assign _EVAL_785 = {{24'd0}, _EVAL_569};
  assign _EVAL_879 = _EVAL_1814 == 5'h0;
  assign _EVAL_1188 = _EVAL_587 == 1'h0;
  assign _EVAL_641 = _EVAL_1018 == 1'h0;
  assign _EVAL_1284 = 5'h4 == _EVAL_1325;
  assign _EVAL_1821 = 5'h9 == _EVAL_1325;
  assign _EVAL_253 = 5'ha == _EVAL_1325;
  assign _EVAL_1153 = 5'hb == _EVAL_1325;
  assign _EVAL_1587 = 5'h8 == _EVAL_1325;
  assign _EVAL_617 = 5'hc == _EVAL_1325;
  assign _EVAL_664 = _EVAL_1191 ? 3'h2 : _EVAL_169;
  assign _EVAL_954 = _EVAL_617 ? 3'h2 : _EVAL_664;
  assign _EVAL_303 = _EVAL_1587 ? 3'h2 : _EVAL_954;
  assign _EVAL_576 = _EVAL_1153 ? 3'h3 : _EVAL_303;
  assign _EVAL_391 = _EVAL_253 ? 3'h3 : _EVAL_576;
  assign _EVAL_523 = _EVAL_1821 ? 3'h3 : _EVAL_391;
  assign _EVAL_1505 = _EVAL_1284 ? 3'h3 : _EVAL_523;
  assign _EVAL_1367 = _EVAL_641 ? 3'h0 : _EVAL_1505;
  assign _EVAL_1201 = _EVAL_1188 ? 3'h4 : _EVAL_1367;
  assign _EVAL_934 = _EVAL_1736 ? 3'h6 : _EVAL_1201;
  assign _EVAL_1327 = _EVAL_934[2];
  assign _EVAL_716 = _EVAL_1327 == 1'h0;
  assign _EVAL_597 = {{2'd0}, _EVAL_981};
  assign _EVAL_619 = _EVAL_548 ? _EVAL_597 : 4'h0;
  assign _EVAL_166 = _EVAL_368 ? _EVAL_597 : _EVAL_619;
  assign _EVAL_1676 = _EVAL_1191 ? _EVAL_597 : _EVAL_166;
  assign _EVAL_996 = _EVAL_617 ? _EVAL_597 : _EVAL_1676;
  assign _EVAL_1522 = _EVAL_1587 ? _EVAL_597 : _EVAL_996;
  assign _EVAL_330 = _EVAL_1153 ? _EVAL_597 : _EVAL_1522;
  assign _EVAL_1707 = _EVAL_253 ? _EVAL_597 : _EVAL_330;
  assign _EVAL_1152 = _EVAL_1821 ? _EVAL_597 : _EVAL_1707;
  assign _EVAL_297 = _EVAL_1284 ? _EVAL_597 : _EVAL_1152;
  assign _EVAL_747 = _EVAL_641 ? _EVAL_597 : _EVAL_297;
  assign _EVAL_638 = _EVAL_1188 ? _EVAL_597 : _EVAL_747;
  assign _EVAL_421 = _EVAL_1736 ? 4'h6 : _EVAL_638;
  assign _EVAL_1648 = 23'hff << _EVAL_421;
  assign _EVAL_1297 = _EVAL_1648[7:0];
  assign _EVAL_420 = ~ _EVAL_1297;
  assign _EVAL_1681 = _EVAL_420[7:3];
  assign _EVAL_447 = _EVAL_716 ? _EVAL_1681 : 5'h0;
  assign _EVAL_1055 = _EVAL_1814 - 5'h1;
  assign _EVAL_1380 = _EVAL_1774[11:2];
  assign _EVAL_1248 = _EVAL_155[11:2];
  assign _EVAL_310 = _EVAL_1380 == _EVAL_1248;
  assign _EVAL_298 = _EVAL_393[3];
  assign _EVAL_1168 = _EVAL_393[2];
  assign _EVAL_1538 = _EVAL_393[1];
  assign _EVAL_1763 = _EVAL_393[0];
  assign _EVAL_1521 = {_EVAL_298,_EVAL_1168,_EVAL_1538,_EVAL_1763};
  assign _EVAL_1161 = _EVAL_1521[3];
  assign _EVAL_1165 = _EVAL_1521[2];
  assign _EVAL_1737 = _EVAL_1521[1];
  assign _EVAL_869 = _EVAL_1521[0];
  assign _EVAL_1631 = {_EVAL_1161,_EVAL_1165,_EVAL_1737,_EVAL_869};
  assign _EVAL_1256 = _EVAL_1653[3];
  assign _EVAL_670 = _EVAL_1653[2];
  assign _EVAL_1693 = _EVAL_1653[1];
  assign _EVAL_1528 = _EVAL_1653[0];
  assign _EVAL_1503 = {_EVAL_1256,_EVAL_670,_EVAL_1693,_EVAL_1528};
  assign _EVAL_997 = _EVAL_1503[3];
  assign _EVAL_768 = _EVAL_1503[2];
  assign _EVAL_1671 = _EVAL_1503[1];
  assign _EVAL_1288 = _EVAL_1503[0];
  assign _EVAL_1495 = {_EVAL_997,_EVAL_768,_EVAL_1671,_EVAL_1288};
  assign _EVAL_1053 = _EVAL_1631 & _EVAL_1495;
  assign _EVAL_1641 = _EVAL_1053 != 4'h0;
  assign _EVAL_182 = _EVAL_393 & _EVAL_1653;
  assign _EVAL_755 = _EVAL_182 != 4'h0;
  assign _EVAL_399 = _EVAL_1211 ? _EVAL_1641 : _EVAL_755;
  assign _EVAL_1860 = _EVAL_310 & _EVAL_399;
  assign _EVAL_1394 = _EVAL_465[3];
  assign _EVAL_1673 = _EVAL_187[2];
  assign _EVAL_251 = _EVAL_1769[2];
  assign _EVAL_1624 = _EVAL_251 & _EVAL_553;
  assign _EVAL_427 = _EVAL_1325 == 5'h5;
  assign _EVAL_343 = _EVAL_981[0];
  assign _EVAL_1846 = _EVAL_343 == 1'h0;
  assign _EVAL_1508 = _EVAL_427 & _EVAL_1846;
  assign _EVAL_296 = _EVAL_1769[5];
  assign _EVAL_807 = _EVAL_296 & _EVAL_553;
  assign _EVAL_1119 = q__EVAL_10;
  assign _EVAL_512 = data__EVAL_1;
  assign _EVAL_534 = _EVAL_512[31:0];
  assign _EVAL_811 = _EVAL_722 ? _EVAL_277 : _EVAL_1062;
  assign _EVAL_1185 = _EVAL_1609 ? _EVAL_811 : _EVAL_1439;
  assign _EVAL_829 = _EVAL_1185;
  assign _EVAL_1433 = _EVAL_465[0];
  assign _EVAL_175 = _EVAL_564 | _EVAL_792;
  assign _EVAL_248 = _EVAL_175 | _EVAL_1788;
  assign _EVAL_1011 = _EVAL_248 | _EVAL_1273;
  assign _EVAL_1359 = _EVAL_1011 | _EVAL_1237;
  assign _EVAL_1192 = _EVAL_1359 == 1'h0;
  assign _EVAL_1254 = _EVAL_759;
  assign _EVAL_351 = _EVAL_1192 & _EVAL_1254;
  assign _EVAL_950 = _EVAL_560 ? 3'h7 : 3'h3;
  assign _EVAL_422 = _EVAL_560 ? 3'h0 : 3'h5;
  assign _EVAL_1566 = _EVAL_1430 ? _EVAL_950 : _EVAL_422;
  assign _EVAL_366 = _EVAL_1098 ? 3'h2 : _EVAL_1566;
  assign _EVAL_1830 = _EVAL_427 & _EVAL_343;
  assign _EVAL_891 = _EVAL_1663 & _EVAL_1830;
  assign _EVAL_1519 = _EVAL_891 & _EVAL_1611;
  assign _EVAL_772 = _EVAL_453 | _EVAL_1519;
  assign _EVAL_1680 = _EVAL_772 | _EVAL_1278;
  assign _EVAL_1729 = _EVAL_1278 == 1'h0;
  assign _EVAL_1764 = _EVAL_1729 & _EVAL_54;
  assign _EVAL_1420 = _EVAL_1764 == 1'h0;
  assign _EVAL_1139 = _EVAL_1680 & _EVAL_1420;
  assign _EVAL_957 = _EVAL_981[1];
  assign _EVAL_1608 = _EVAL_1519 & _EVAL_957;
  assign _EVAL_1323 = _EVAL_1058[1];
  assign _EVAL_889 = _EVAL_1278 & _EVAL_1323;
  assign _EVAL_704 = _EVAL_1608 | _EVAL_889;
  assign _EVAL_1818 = _EVAL_704 == 1'h0;
  assign _EVAL_668 = _EVAL_406 & _EVAL_1818;
  assign _EVAL_1815 = _EVAL_668 ? 3'h1 : 3'h6;
  assign _EVAL_347 = _EVAL_1139 ? _EVAL_1815 : _EVAL_396;
  assign _EVAL_1640 = _EVAL_1450 ? _EVAL_366 : _EVAL_347;
  assign _EVAL_295 = _EVAL_351 ? 3'h0 : _EVAL_1640;
  assign _EVAL_1150 = _EVAL_403 ? _EVAL_295 : _EVAL_1640;
  assign _EVAL_948 = _EVAL_560 ? 3'h0 : _EVAL_1150;
  assign _EVAL_1559 = _EVAL_720 ? _EVAL_948 : _EVAL_1150;
  assign _EVAL_1094 = {{1'd0}, _EVAL_981};
  assign _EVAL_350 = _EVAL_1094[1:0];
  assign _EVAL_1379 = 4'h1 << _EVAL_350;
  assign _EVAL_1537 = _EVAL_1379[2:0];
  assign _EVAL_235 = _EVAL_1537 | 3'h1;
  assign _EVAL_1572 = _EVAL_235[1];
  assign _EVAL_1246 = _EVAL_389[2];
  assign _EVAL_1314 = _EVAL_1246 == 1'h0;
  assign _EVAL_1092 = _EVAL_1314 & _EVAL_220;
  assign _EVAL_444 = _EVAL_1572 & _EVAL_1092;
  assign _EVAL_1488 = {_EVAL_1096,_EVAL_1096};
  assign _EVAL_765 = _EVAL_548 ? _EVAL_1488 : 64'h0;
  assign _EVAL_1585 = _EVAL_368 ? _EVAL_1488 : _EVAL_765;
  assign _EVAL_1848 = _EVAL_1191 ? _EVAL_1488 : _EVAL_1585;
  assign _EVAL_1727 = _EVAL_617 ? _EVAL_1488 : _EVAL_1848;
  assign _EVAL_633 = _EVAL_1587 ? _EVAL_1488 : _EVAL_1727;
  assign _EVAL_434 = _EVAL_1185;
  assign _EVAL_713 = _EVAL_1131 ? _EVAL_434 : _EVAL_829;
  assign _EVAL_1778 = _EVAL_187[0];
  assign _EVAL_939 = _EVAL_1733 == 1'h0;
  assign _EVAL_452 = _EVAL_1622 & _EVAL_939;
  assign _EVAL_1250 = _EVAL_452 ? _EVAL_1264 : 2'h0;
  assign _EVAL_195 = _EVAL_760 == 1'h0;
  assign _EVAL_1342 = _EVAL_1417[31:12];
  assign _EVAL_1694 = {_EVAL_1342,_EVAL_561};
  assign _EVAL_464 = _EVAL_52[31:12];
  assign _EVAL_663 = _EVAL_1694[11:0];
  assign _EVAL_529 = {_EVAL_464,_EVAL_663};
  assign _EVAL_1741 = {_EVAL_464,_EVAL_663};
  assign _EVAL_1108 = _EVAL_1107[11:0];
  assign _EVAL_1579 = {_EVAL_464,_EVAL_1108};
  assign _EVAL_625 = _EVAL_1060[5:0];
  assign _EVAL_968 = {_EVAL_625, 6'h0};
  assign _EVAL_1360 = {_EVAL_464,_EVAL_968};
  assign _EVAL_1178 = {1'h0,_EVAL_1107};
  assign _EVAL_304 = {1'h0,_EVAL_1476};
  assign _EVAL_1593 = _EVAL_403 ? _EVAL_1178 : _EVAL_304;
  assign _EVAL_234 = _EVAL_1593[31:0];
  assign _EVAL_1197 = _EVAL_52;
  assign _EVAL_473 = _EVAL_1131 ? _EVAL_234 : _EVAL_1197;
  assign _EVAL_260 = _EVAL_1237 ? _EVAL_1360 : _EVAL_473;
  assign _EVAL_522 = _EVAL_1273 ? _EVAL_1579 : _EVAL_260;
  assign _EVAL_266 = _EVAL_1788 ? _EVAL_1741 : _EVAL_522;
  assign _EVAL_1615 = _EVAL_792 ? _EVAL_529 : _EVAL_266;
  assign _EVAL_1078 = _EVAL_1769[0];
  assign _EVAL_379 = _EVAL_1359 | _EVAL_1131;
  assign _EVAL_837 = _EVAL_379 == 1'h0;
  assign _EVAL_676 = _EVAL_837 == 1'h0;
  assign _EVAL_233 = _EVAL_37;
  assign _EVAL_892 = _EVAL_676 | _EVAL_233;
  assign _EVAL_886 = _EVAL_54 == 1'h0;
  assign _EVAL_1338 = _EVAL_1788 ? 1'h1 : _EVAL_1273;
  assign _EVAL_828 = _EVAL_792 ? _EVAL_886 : _EVAL_1338;
  assign _EVAL_160 = _EVAL_564 ? 1'h1 : _EVAL_828;
  assign _EVAL_1760 = _EVAL_892 & _EVAL_160;
  assign _EVAL_867 = _EVAL_1360;
  assign _EVAL_339 = _EVAL_564 ? _EVAL_867 : _EVAL_1615;
  assign _EVAL_283 = 4'hf;
  assign _EVAL_1209 = _EVAL_283;
  assign _EVAL_589 = _EVAL_283;
  assign _EVAL_1437 = _EVAL_1567 ? _EVAL_1209 : _EVAL_589;
  assign _EVAL_1793 = _EVAL_291[11:2];
  assign _EVAL_1125 = _EVAL_1793 == _EVAL_1248;
  assign _EVAL_348 = _EVAL_1121[3];
  assign _EVAL_1750 = _EVAL_1121[2];
  assign _EVAL_748 = _EVAL_1121[1];
  assign _EVAL_906 = _EVAL_1121[0];
  assign _EVAL_1432 = {_EVAL_348,_EVAL_1750,_EVAL_748,_EVAL_906};
  assign _EVAL_319 = _EVAL_1432[3];
  assign _EVAL_586 = _EVAL_1432[2];
  assign _EVAL_823 = _EVAL_1432[1];
  assign _EVAL_197 = _EVAL_1432[0];
  assign _EVAL_508 = {_EVAL_319,_EVAL_586,_EVAL_823,_EVAL_197};
  assign _EVAL_868 = _EVAL_508 & _EVAL_1495;
  assign _EVAL_952 = _EVAL_868 != 4'h0;
  assign _EVAL_1639 = _EVAL_1765 != 4'h0;
  assign _EVAL_863 = _EVAL_1211 ? _EVAL_952 : _EVAL_1639;
  assign _EVAL_441 = _EVAL_1125 & _EVAL_863;
  assign _EVAL_1705 = _EVAL_322 & _EVAL_441;
  assign _EVAL_1223 = _EVAL_248 == 1'h0;
  assign _EVAL_1813 = _EVAL_1011 == 1'h0;
  assign _EVAL_919 = _EVAL_1813 & _EVAL_1254;
  assign _EVAL_363 = _EVAL_204 == 5'h0;
  assign _EVAL_1294 = _EVAL_204 == 5'h6;
  assign _EVAL_956 = _EVAL_363 | _EVAL_1294;
  assign _EVAL_648 = _EVAL_956 | _EVAL_470;
  assign _EVAL_876 = _EVAL_648 | _EVAL_978;
  assign _EVAL_1220 = _EVAL_1211 & _EVAL_1542;
  assign _EVAL_1568 = _EVAL_876 | _EVAL_1220;
  assign _EVAL_1008 = _EVAL_172 & _EVAL_1568;
  assign _EVAL_1662 = q__EVAL_16;
  assign _EVAL_301 = _EVAL_1508 & _EVAL_1100;
  assign _EVAL_1786 = _EVAL_1422 == 1'h0;
  assign _EVAL_1309 = _EVAL_301 & _EVAL_1786;
  assign _EVAL_1637 = _EVAL_1830 & _EVAL_1462;
  assign _EVAL_1849 = _EVAL_1309 | _EVAL_1637;
  assign _EVAL_1515 = _EVAL_780 & _EVAL_1849;
  assign _EVAL_810 = {_EVAL_1626,_EVAL_1300,_EVAL_1134,_EVAL_211,_EVAL_401,_EVAL_487,_EVAL_1049,_EVAL_1851};
  assign _EVAL_1087 = _EVAL_1078 ? _EVAL_810 : 80'h0;
  assign _EVAL_640 = {_EVAL_801,_EVAL_1387,_EVAL_451,_EVAL_1569,_EVAL_937,_EVAL_1269,_EVAL_732,_EVAL_753};
  assign _EVAL_1268 = _EVAL_1348 ? _EVAL_640 : 80'h0;
  assign _EVAL_808 = _EVAL_1087 | _EVAL_1268;
  assign _EVAL_1000 = {_EVAL_1441,_EVAL_1810,_EVAL_874,_EVAL_1316,_EVAL_918,_EVAL_377,_EVAL_1001,_EVAL_280};
  assign _EVAL_1280 = _EVAL_251 ? _EVAL_1000 : 80'h0;
  assign _EVAL_327 = _EVAL_808 | _EVAL_1280;
  assign _EVAL_1393 = _EVAL_1769[3];
  assign _EVAL_636 = {_EVAL_1172,_EVAL_1240,_EVAL_1740,_EVAL_1500,_EVAL_376,_EVAL_1739,_EVAL_1800,_EVAL_1688};
  assign _EVAL_227 = _EVAL_1393 ? _EVAL_636 : 80'h0;
  assign _EVAL_1351 = _EVAL_327 | _EVAL_227;
  assign _EVAL_362 = _EVAL_1769[4];
  assign _EVAL_1245 = {_EVAL_1724,_EVAL_1831,_EVAL_1625,_EVAL_300,_EVAL_1140,_EVAL_614,_EVAL_477,_EVAL_1444};
  assign _EVAL_1070 = _EVAL_362 ? _EVAL_1245 : 80'h0;
  assign _EVAL_1447 = _EVAL_1351 | _EVAL_1070;
  assign _EVAL_880 = {_EVAL_1784,_EVAL_1213,_EVAL_1756,_EVAL_162,_EVAL_1847,_EVAL_1489,_EVAL_541,_EVAL_387};
  assign _EVAL_517 = _EVAL_296 ? _EVAL_880 : 80'h0;
  assign _EVAL_1093 = _EVAL_1447 | _EVAL_517;
  assign _EVAL_585 = _EVAL_946 & _EVAL_1860;
  assign _EVAL_1766 = _EVAL_585 | _EVAL_1705;
  assign _EVAL_1675 = _EVAL_876 & _EVAL_1766;
  assign _EVAL_338 = _EVAL_1697 & _EVAL_1675;
  assign _EVAL_1123 = _EVAL_1850 & _EVAL_309;
  assign _EVAL_1635 = _EVAL_42 | _EVAL_1123;
  assign _EVAL_1017 = _EVAL_338 ? 1'h1 : _EVAL_1635;
  assign _EVAL_991 = _EVAL_548 ? 3'h3 : 3'h0;
  assign _EVAL_603 = _EVAL_368 ? 3'h2 : _EVAL_991;
  assign _EVAL_1308 = _EVAL_1191 ? 3'h1 : _EVAL_603;
  assign _EVAL_1772 = _EVAL_617 ? 3'h0 : _EVAL_1308;
  assign _EVAL_1282 = _EVAL_1587 ? 3'h4 : _EVAL_1772;
  assign _EVAL_192 = _EVAL_1153 ? 3'h2 : _EVAL_1282;
  assign _EVAL_1429 = _EVAL_253 ? 3'h1 : _EVAL_192;
  assign _EVAL_500 = _EVAL_1821 ? 3'h0 : _EVAL_1429;
  assign _EVAL_326 = _EVAL_1284 ? 3'h3 : _EVAL_500;
  assign _EVAL_1331 = _EVAL_641 ? 3'h0 : _EVAL_326;
  assign _EVAL_539 = _EVAL_1188 ? 3'h0 : _EVAL_1331;
  assign _EVAL_1219 = _EVAL_919 & _EVAL_1237;
  assign _EVAL_536 = _EVAL_322 ? _EVAL_291 : _EVAL_1774;
  assign _EVAL_843 = _EVAL_981 >= 2'h3;
  assign _EVAL_537 = _EVAL_235[2];
  assign _EVAL_245 = _EVAL_537 & _EVAL_1246;
  assign _EVAL_1580 = _EVAL_843 | _EVAL_245;
  assign _EVAL_499 = _EVAL_220 == 1'h0;
  assign _EVAL_1510 = _EVAL_1246 & _EVAL_499;
  assign _EVAL_669 = _EVAL_1572 & _EVAL_1510;
  assign _EVAL_1106 = _EVAL_1580 | _EVAL_669;
  assign _EVAL_652 = _EVAL_235[0];
  assign _EVAL_1743 = _EVAL_1510 & _EVAL_760;
  assign _EVAL_244 = _EVAL_652 & _EVAL_1743;
  assign _EVAL_574 = _EVAL_1106 | _EVAL_244;
  assign _EVAL_1543 = _EVAL_396 == 3'h0;
  assign _EVAL_866 = _EVAL_1835 == 1'h0;
  assign _EVAL_1836 = _EVAL_1543 & _EVAL_866;
  assign _EVAL_1103 = _EVAL_1098 ? 1'h1 : _EVAL_428;
  assign _EVAL_988 = _EVAL_1103 ? 1'h1 : _EVAL_1017;
  assign _EVAL_1602 = _EVAL_1450 ? _EVAL_988 : _EVAL_1017;
  assign _EVAL_1408 = _EVAL_1602 == 1'h0;
  assign _EVAL_262 = _EVAL_1836 & _EVAL_1408;
  assign _EVAL_1469 = _EVAL_521 | _EVAL_1697;
  assign _EVAL_281 = _EVAL_1469 | _EVAL_1109;
  assign _EVAL_1799 = _EVAL_281 == 1'h0;
  assign _EVAL_1712 = _EVAL_351 & _EVAL_1799;
  assign _EVAL_1403 = _EVAL_1712;
  assign _EVAL_974 = _EVAL_1403 & _EVAL_1524;
  assign _EVAL_1529 = 3'h0;
  assign _EVAL_985 = {_EVAL_1394,_EVAL_736};
  assign _EVAL_1163 = _EVAL_465[1];
  assign _EVAL_857 = {_EVAL_1163,_EVAL_1433};
  assign _EVAL_917 = {_EVAL_985,_EVAL_857};
  assign _EVAL_1064 = _EVAL_1769[6];
  assign _EVAL_1613 = {_EVAL_846,_EVAL_1541,_EVAL_239,_EVAL_1135,_EVAL_700,_EVAL_375,_EVAL_1595,_EVAL_629};
  assign _EVAL_1042 = _EVAL_1064 ? _EVAL_1613 : 80'h0;
  assign _EVAL_1853 = _EVAL_1093 | _EVAL_1042;
  assign _EVAL_653 = _EVAL_1853[34];
  assign _EVAL_516 = _EVAL_1853[79:48];
  assign _EVAL_358 = _EVAL_516[1];
  assign _EVAL_1400 = _EVAL_516[2];
  assign _EVAL_1362 = _EVAL_38;
  assign _EVAL_208 = _EVAL_1362[63:32];
  assign _EVAL_203 = _EVAL_1362[31:0];
  assign _EVAL_764 = _EVAL_1400 ? _EVAL_208 : _EVAL_203;
  assign _EVAL_856 = _EVAL_764[31:16];
  assign _EVAL_1547 = _EVAL_764[15:0];
  assign _EVAL_1045 = _EVAL_358 ? _EVAL_856 : _EVAL_1547;
  assign _EVAL_1452 = _EVAL_1045[15];
  assign _EVAL_1210 = _EVAL_653 & _EVAL_1452;
  assign _EVAL_1073 = amoalu__EVAL_0;
  assign _EVAL_1514 = _EVAL_548 ? _EVAL_1117 : 3'h0;
  assign _EVAL_1335 = _EVAL_368 ? _EVAL_1117 : _EVAL_1514;
  assign _EVAL_864 = _EVAL_1191 ? _EVAL_1117 : _EVAL_1335;
  assign _EVAL_965 = _EVAL_617 ? _EVAL_1117 : _EVAL_864;
  assign _EVAL_214 = _EVAL_160 == 1'h0;
  assign _EVAL_1030 = _EVAL_1073[7:0];
  assign _EVAL_392 = _EVAL_946 | _EVAL_322;
  assign _EVAL_321 = _EVAL_1008 & _EVAL_392;
  assign _EVAL_1388 = _EVAL_1153 ? _EVAL_1488 : _EVAL_633;
  assign _EVAL_964 = _EVAL_253 ? _EVAL_1488 : _EVAL_1388;
  assign _EVAL_255 = _EVAL_125[0];
  assign _EVAL_1071 = _EVAL_255 | _EVAL_96;
  assign _EVAL_1180 = _EVAL_1071 | _EVAL_892;
  assign _EVAL_1133 = _EVAL_1180 | _EVAL_926;
  assign _EVAL_673 = _EVAL_1133 | _EVAL_1450;
  assign _EVAL_1138 = _EVAL_673 | _EVAL_1697;
  assign _EVAL_504 = _EVAL_1138 | _EVAL_1109;
  assign _EVAL_1713 = _EVAL_504 | _EVAL_1252;
  assign _EVAL_888 = _EVAL_389[31:12];
  assign _EVAL_156 = _EVAL_537 & _EVAL_1314;
  assign _EVAL_1614 = _EVAL_843 | _EVAL_156;
  assign _EVAL_360 = _EVAL_1314 & _EVAL_499;
  assign _EVAL_161 = _EVAL_1572 & _EVAL_360;
  assign _EVAL_833 = _EVAL_1614 | _EVAL_161;
  assign _EVAL_1353 = _EVAL_360 & _EVAL_760;
  assign _EVAL_333 = _EVAL_652 & _EVAL_1353;
  assign _EVAL_929 = _EVAL_833 | _EVAL_333;
  assign _EVAL_554 = _EVAL_1587 ? _EVAL_1117 : _EVAL_965;
  assign _EVAL_852 = _EVAL_1153 ? _EVAL_1117 : _EVAL_554;
  assign _EVAL_1130 = _EVAL_253 ? _EVAL_1117 : _EVAL_852;
  assign _EVAL_695 = _EVAL_1821 ? _EVAL_1117 : _EVAL_1130;
  assign _EVAL_1038 = _EVAL_536[2];
  assign _EVAL_1643 = _EVAL_1519 ? _EVAL_888 : _EVAL_549;
  assign _EVAL_1477 = _EVAL_1399 == 3'h6;
  assign _EVAL_1768 = _EVAL_1246 & _EVAL_220;
  assign _EVAL_1344 = _EVAL_1768 & _EVAL_195;
  assign _EVAL_1645 = _EVAL_652 & _EVAL_1344;
  assign _EVAL_975 = _EVAL_362 & _EVAL_553;
  assign _EVAL_1728 = _EVAL_135 == 5'h0;
  assign _EVAL_383 = _EVAL_135 == 5'h6;
  assign _EVAL_1357 = _EVAL_1728 | _EVAL_383;
  assign _EVAL_757 = _EVAL_135 == 5'h7;
  assign _EVAL_1291 = _EVAL_1357 | _EVAL_757;
  assign _EVAL_600 = _EVAL_512[63:32];
  assign _EVAL_432 = _EVAL_1362[55:48];
  assign _EVAL_270 = _EVAL_1362[63:56];
  assign _EVAL_1307 = _EVAL_1362[47:40];
  assign _EVAL_1578 = _EVAL_1362[39:32];
  assign _EVAL_1182 = {_EVAL_270,_EVAL_432,_EVAL_1307,_EVAL_1578};
  assign _EVAL_581 = _EVAL_780 & _EVAL_210;
  assign _EVAL_1530 = _EVAL_581 & _EVAL_1184;
  assign _EVAL_1652 = _EVAL_893 - 7'h1;
  assign _EVAL_337 = _EVAL_1850 & _EVAL_511;
  assign _EVAL_848 = _EVAL_337 & _EVAL_866;
  assign _EVAL_1321 = _EVAL_848 | _EVAL_453;
  assign _EVAL_575 = _EVAL_1321 & _EVAL_210;
  assign _EVAL_489 = _EVAL_1694[31:6];
  assign _EVAL_1732 = {_EVAL_489, 6'h0};
  assign _EVAL_684 = _EVAL_1732 | _EVAL_785;
  assign _EVAL_1487 = _EVAL_684[11:0];
  assign _EVAL_1059 = {{6'd0}, _EVAL_660};
  assign _EVAL_1824 = _EVAL_658 | _EVAL_1059;
  assign _EVAL_1414 = _EVAL_52[11:0];
  assign _EVAL_802 = _EVAL_1567 ? _EVAL_1824 : _EVAL_1414;
  assign _EVAL_1385 = _EVAL_496 ? _EVAL_1487 : _EVAL_802;
  assign _EVAL_1204 = _EVAL_389[11:6];
  assign _EVAL_1301 = {_EVAL_1643,_EVAL_1204};
  assign _EVAL_336 = _EVAL_892 & _EVAL_214;
  assign _EVAL_751 = _EVAL_135 == 5'h11;
  assign _EVAL_1747 = _EVAL_1100 & _EVAL_1543;
  assign _EVAL_1491 = _EVAL_1747 & _EVAL_1611;
  assign _EVAL_685 = _EVAL_780 & _EVAL_1508;
  assign _EVAL_1822 = _EVAL_1642 & _EVAL_1611;
  assign _EVAL_1443 = _EVAL_1822 & _EVAL_1475;
  assign _EVAL_781 = _EVAL_1073[31:24];
  assign _EVAL_783 = _EVAL_620 & _EVAL_1486;
  assign _EVAL_478 = _EVAL_783 & _EVAL_172;
  assign _EVAL_607 = _EVAL_1697 | _EVAL_1109;
  assign _EVAL_1111 = _EVAL_607 | _EVAL_1835;
  assign _EVAL_657 = _EVAL_135 == 5'hf;
  assign _EVAL_1549 = _EVAL_317 & _EVAL_939;
  assign _EVAL_1795 = _EVAL_1549 ? _EVAL_693 : 2'h0;
  assign _EVAL_1397 = _EVAL_1795 | _EVAL_1250;
  assign _EVAL_626 = _EVAL_1502;
  assign _EVAL_1116 = _EVAL_172 | _EVAL_946;
  assign _EVAL_936 = _EVAL_1116 | _EVAL_322;
  assign _EVAL_682 = _EVAL_502 == 5'h0;
  assign _EVAL_1085 = _EVAL_531 & _EVAL_682;
  assign _EVAL_323 = _EVAL_209 & _EVAL_778;
  assign _EVAL_285 = _EVAL_323 | _EVAL_322;
  assign _EVAL_726 = _EVAL_285 & _EVAL_435;
  assign _EVAL_1216 = _EVAL_838 | _EVAL_726;
  assign _EVAL_1621 = _EVAL_1216 == 1'h0;
  assign _EVAL_206 = _EVAL_322 & _EVAL_1621;
  assign _EVAL_570 = _EVAL_1572 & _EVAL_1768;
  assign _EVAL_378 = _EVAL_1580 | _EVAL_570;
  assign _EVAL_649 = _EVAL_1768 & _EVAL_760;
  assign _EVAL_1149 = _EVAL_652 & _EVAL_649;
  assign _EVAL_318 = _EVAL_378 | _EVAL_1149;
  assign _EVAL_1142 = _EVAL_378 | _EVAL_1645;
  assign _EVAL_1199 = _EVAL_1510 & _EVAL_195;
  assign _EVAL_1573 = _EVAL_652 & _EVAL_1199;
  assign _EVAL_578 = _EVAL_1106 | _EVAL_1573;
  assign _EVAL_173 = _EVAL_1614 | _EVAL_444;
  assign _EVAL_1790 = _EVAL_1092 & _EVAL_760;
  assign _EVAL_237 = _EVAL_652 & _EVAL_1790;
  assign _EVAL_1260 = _EVAL_173 | _EVAL_237;
  assign _EVAL_803 = _EVAL_1092 & _EVAL_195;
  assign _EVAL_1162 = _EVAL_652 & _EVAL_803;
  assign _EVAL_1383 = _EVAL_173 | _EVAL_1162;
  assign _EVAL_1099 = _EVAL_360 & _EVAL_195;
  assign _EVAL_1659 = _EVAL_652 & _EVAL_1099;
  assign _EVAL_385 = _EVAL_833 | _EVAL_1659;
  assign _EVAL_501 = {_EVAL_318,_EVAL_1142,_EVAL_574,_EVAL_578,_EVAL_1260,_EVAL_1383,_EVAL_929,_EVAL_385};
  assign _EVAL_1599 = _EVAL_548 ? _EVAL_501 : 8'h0;
  assign _EVAL_599 = _EVAL_368 ? _EVAL_501 : _EVAL_1599;
  assign _EVAL_834 = _EVAL_1191 ? _EVAL_501 : _EVAL_599;
  assign _EVAL_1345 = _EVAL_145;
  assign _EVAL_1050 = _EVAL_1345;
  assign _EVAL_1451 = _EVAL_1032 - 3'h1;
  assign _EVAL_1719 = 2'h1 << _EVAL_1038;
  assign _EVAL_630 = _EVAL_722 ? _EVAL_277 : _EVAL_1062;
  assign _EVAL_1539 = _EVAL_1060 + 8'h1;
  assign _EVAL_157 = _EVAL_1539[8:6];
  assign _EVAL_881 = _EVAL_157 == 3'h4;
  assign _EVAL_1339 = _EVAL_339[31:6];
  assign _EVAL_1859 = _EVAL_52[5:0];
  assign _EVAL_1606 = {_EVAL_1339,_EVAL_1859};
  assign _EVAL_797 = _EVAL_1253 ? 3'h5 : _EVAL_442;
  assign _EVAL_1787 = _EVAL_1217 ? 3'h4 : _EVAL_797;
  assign _EVAL_256 = _EVAL_1132 ? 3'h3 : _EVAL_1787;
  assign _EVAL_1532 = _EVAL_1679 ? 3'h3 : _EVAL_256;
  assign _EVAL_243 = _EVAL_1430 ? _EVAL_1532 : 3'h5;
  assign _EVAL_1683 = _EVAL_1098 ? 3'h5 : _EVAL_243;
  assign _EVAL_1305 = _EVAL_1450 ? _EVAL_1683 : 3'h5;
  assign _EVAL_1571 = _EVAL_1865 ? _EVAL_1532 : _EVAL_1305;
  assign _EVAL_335 = _EVAL_516[0];
  assign _EVAL_520 = _EVAL_1853[36:35];
  assign _EVAL_743 = _EVAL_520 == 2'h1;
  assign _EVAL_1012 = _EVAL_1210 ? 16'hffff : 16'h0;
  assign _EVAL_1179 = _EVAL_743 ? _EVAL_1012 : _EVAL_856;
  assign _EVAL_550 = {_EVAL_1179,_EVAL_1045};
  assign _EVAL_1468 = _EVAL_550[15:8];
  assign _EVAL_1276 = _EVAL_550[7:0];
  assign _EVAL_505 = _EVAL_335 ? _EVAL_1468 : _EVAL_1276;
  assign _EVAL_1224 = _EVAL_505[7];
  assign _EVAL_1289 = _EVAL_653 & _EVAL_1224;
  assign _EVAL_1504 = _EVAL_1289 ? 24'hffffff : 24'h0;
  assign _EVAL_844 = _EVAL_617 ? _EVAL_501 : _EVAL_834;
  assign _EVAL_1654 = _EVAL_1587 ? _EVAL_501 : _EVAL_844;
  assign _EVAL_1144 = _EVAL_1153 ? _EVAL_501 : _EVAL_1654;
  assign _EVAL_1320 = _EVAL_253 ? _EVAL_501 : _EVAL_1144;
  assign _EVAL_1173 = _EVAL_1821 ? _EVAL_501 : _EVAL_1320;
  assign _EVAL_920 = _EVAL_1284 ? _EVAL_501 : _EVAL_1173;
  assign _EVAL_1075 = _EVAL_731 ? _EVAL_1532 : _EVAL_1571;
  assign _EVAL_229 = _EVAL_52[2];
  assign _EVAL_200 = 2'h1 << _EVAL_229;
  assign _EVAL_423 = _EVAL_1567 ? 2'h3 : _EVAL_200;
  assign _EVAL_315 = _EVAL_135 == 5'h4;
  assign _EVAL_1136 = _EVAL_135 == 5'h9;
  assign _EVAL_1866 = _EVAL_315 | _EVAL_1136;
  assign _EVAL_1591 = _EVAL_135 == 5'ha;
  assign _EVAL_706 = _EVAL_1866 | _EVAL_1591;
  assign _EVAL_1081 = _EVAL_135 == 5'hb;
  assign _EVAL_528 = _EVAL_706 | _EVAL_1081;
  assign _EVAL_1249 = _EVAL_135 == 5'h8;
  assign _EVAL_1629 = _EVAL_135 == 5'hc;
  assign _EVAL_246 = _EVAL_1249 | _EVAL_1629;
  assign _EVAL_610 = _EVAL_135 == 5'hd;
  assign _EVAL_1137 = _EVAL_246 | _EVAL_610;
  assign _EVAL_1424 = _EVAL_135 == 5'he;
  assign _EVAL_415 = _EVAL_1137 | _EVAL_1424;
  assign _EVAL_1551 = _EVAL_415 | _EVAL_657;
  assign _EVAL_1834 = _EVAL_528 | _EVAL_1551;
  assign _EVAL_1347 = _EVAL_1291 | _EVAL_1834;
  assign _EVAL_958 = _EVAL_1520 & _EVAL_1347;
  assign _EVAL_515 = _EVAL_958 ? 1'h0 : _EVAL_262;
  assign _EVAL_729 = _EVAL_1393 & _EVAL_553;
  assign _EVAL_1175 = _EVAL_1713 | _EVAL_322;
  assign _EVAL_941 = _EVAL_1175 | _EVAL_849;
  assign _EVAL_1159 = _EVAL_941 | _EVAL_559;
  assign _EVAL_1052 = _EVAL_722 ? _EVAL_277 : _EVAL_1062;
  assign _EVAL_495 = _EVAL_1185;
  assign _EVAL_1148 = _EVAL_1237 ? _EVAL_495 : _EVAL_713;
  assign _EVAL_850 = _EVAL_1273 ? _EVAL_1185 : _EVAL_1148;
  assign _EVAL_1575 = _EVAL_1788 ? _EVAL_630 : _EVAL_850;
  assign _EVAL_1381 = _EVAL_792 ? _EVAL_1052 : _EVAL_1575;
  assign _EVAL_1708 = _EVAL_617 ? _EVAL_389 : _EVAL_806;
  assign _EVAL_1545 = _EVAL_1587 ? _EVAL_389 : _EVAL_1708;
  assign _EVAL_1146 = _EVAL_1153 ? _EVAL_389 : _EVAL_1545;
  assign _EVAL_1574 = _EVAL_253 ? _EVAL_389 : _EVAL_1146;
  assign _EVAL_411 = _EVAL_724[7];
  assign _EVAL_798 = _EVAL_165 & _EVAL_411;
  assign _EVAL_1095 = _EVAL_798 ? 24'hffffff : 24'h0;
  assign _EVAL_1657 = _EVAL_981 == 2'h0;
  assign _EVAL_1113 = _EVAL_1657 | _EVAL_1762;
  assign _EVAL_628 = {_EVAL_1301, 6'h0};
  assign _EVAL_1533 = _EVAL_752[39:32];
  assign _EVAL_371 = _EVAL_1225 - 5'h1;
  assign _EVAL_527 = _EVAL_322 ? _EVAL_461 : _EVAL_831;
  assign _EVAL_340 = _EVAL_496 ? _EVAL_1838 : 4'hf;
  assign _EVAL_1029 = _EVAL_822 ? _EVAL_527 : _EVAL_340;
  assign _EVAL_222 = ~ _EVAL_393;
  assign _EVAL_916 = _EVAL_1694[11:6];
  assign _EVAL_1304 = _EVAL_1476[11:6];
  assign _EVAL_842 = _EVAL_403 ? _EVAL_1181 : _EVAL_1304;
  assign _EVAL_1425 = _EVAL_52[11:6];
  assign _EVAL_914 = _EVAL_1131 ? _EVAL_842 : _EVAL_1425;
  assign _EVAL_1021 = _EVAL_1237 ? _EVAL_625 : _EVAL_914;
  assign _EVAL_1655 = {{31'd0}, _EVAL_1395};
  assign _EVAL_305 = _EVAL_1362[7:0];
  assign _EVAL_1019 = _EVAL_322 & _EVAL_946;
  assign _EVAL_1497 = _EVAL_1019 & _EVAL_172;
  assign _EVAL_1617 = _EVAL_1159 | _EVAL_1835;
  assign _EVAL_1771 = _EVAL_1617 | _EVAL_467;
  assign _EVAL_744 = _EVAL_1771 | _EVAL_509;
  assign _EVAL_845 = _EVAL_1502;
  assign _EVAL_1463 = _EVAL_155[2];
  assign _EVAL_183 = _EVAL_789 ? 3'h5 : _EVAL_734;
  assign _EVAL_1446 = _EVAL_1493 ? 3'h4 : _EVAL_183;
  assign _EVAL_894 = _EVAL_687 ? 3'h3 : _EVAL_1446;
  assign _EVAL_1157 = _EVAL_1785 ? 3'h3 : _EVAL_894;
  assign _EVAL_767 = _EVAL_1369 == 1'h0;
  assign _EVAL_213 = _EVAL_752[63:56];
  assign _EVAL_717 = _EVAL_752[55:48];
  assign _EVAL_540 = _EVAL_752[47:40];
  assign _EVAL_940 = {_EVAL_213,_EVAL_717,_EVAL_540,_EVAL_1533};
  assign _EVAL_998 = _EVAL_752[31:24];
  assign _EVAL_188 = _EVAL_752[23:16];
  assign _EVAL_616 = _EVAL_752[15:8];
  assign _EVAL_579 = {_EVAL_998,_EVAL_188,_EVAL_616,_EVAL_865};
  assign _EVAL_1702 = {_EVAL_940,_EVAL_579};
  assign _EVAL_963 = _EVAL_341 == 1'h0;
  assign _EVAL_1695 = 2'h1 << _EVAL_1463;
  assign _EVAL_1435 = _EVAL_963 ? 2'h0 : _EVAL_1695;
  assign _EVAL_1461 = _EVAL_813 ? 2'h3 : _EVAL_1435;
  assign _EVAL_1616 = _EVAL_1697 & _EVAL_1408;
  assign _EVAL_312 = _EVAL_496 ? 4'hf : _EVAL_1437;
  assign _EVAL_1811 = _EVAL_822 ? _EVAL_917 : _EVAL_312;
  assign _EVAL_635 = _EVAL_1078 & _EVAL_553;
  assign _EVAL_643 = _EVAL_1061 == 1'h0;
  assign _EVAL_1412 = _EVAL_1609 ? _EVAL_1157 : _EVAL_1075;
  assign _EVAL_1589 = _EVAL_1412;
  assign _EVAL_1261 = _EVAL_172 | _EVAL_783;
  assign _EVAL_1649 = _EVAL_1261 | _EVAL_292;
  assign _EVAL_995 = _EVAL_550[31:8];
  assign _EVAL_1665 = _EVAL_1694[11:6];
  assign _EVAL_835 = _EVAL_1107[11:6];
  assign _EVAL_275 = _EVAL_1273 ? _EVAL_835 : _EVAL_1021;
  assign _EVAL_1794 = _EVAL_1788 ? _EVAL_916 : _EVAL_275;
  assign _EVAL_609 = _EVAL_792 ? _EVAL_1665 : _EVAL_1794;
  assign _EVAL_905 = _EVAL_1821 ? _EVAL_1488 : _EVAL_964;
  assign _EVAL_1115 = _EVAL_1284 ? _EVAL_1488 : _EVAL_905;
  assign _EVAL_1518 = _EVAL_1278 ? _EVAL_1539 : {{1'd0}, _EVAL_1060};
  assign _EVAL_883 = _EVAL_1422 ? _EVAL_1518 : {{1'd0}, _EVAL_1060};
  assign _EVAL_890 = _EVAL_800 ? _EVAL_1539 : _EVAL_883;
  assign _EVAL_279 = q__EVAL_15;
  assign _EVAL_1330 = q__EVAL_19;
  assign _EVAL_771 = _EVAL_1284 ? _EVAL_1117 : _EVAL_695;
  assign _EVAL_151 = _EVAL_641 ? _EVAL_1117 : _EVAL_771;
  assign _EVAL_1198 = _EVAL_1188 ? _EVAL_1117 : _EVAL_151;
  assign _EVAL_1466 = _EVAL_446 & _EVAL_939;
  assign _EVAL_966 = _EVAL_1466 ? _EVAL_313 : 2'h0;
  assign _EVAL_177 = _EVAL_1397 | _EVAL_966;
  assign _EVAL_1202 = _EVAL_1825 & _EVAL_939;
  assign _EVAL_268 = _EVAL_1202 ? _EVAL_1561 : 2'h0;
  assign _EVAL_793 = _EVAL_177 | _EVAL_268;
  assign _EVAL_1332 = _EVAL_1616 | _EVAL_1733;
  assign _EVAL_683 = _EVAL_204 == 5'h14;
  assign _EVAL_646 = _EVAL_683 == 1'h0;
  assign _EVAL_1499 = _EVAL_1362[31:24];
  assign _EVAL_774 = _EVAL_1362[23:16];
  assign _EVAL_1754 = _EVAL_1362[15:8];
  assign _EVAL_566 = {_EVAL_1499,_EVAL_774,_EVAL_1754,_EVAL_305};
  assign _EVAL_761 = {_EVAL_1182,_EVAL_566};
  assign _EVAL_665 = _EVAL_1850 == 1'h0;
  assign _EVAL_1749 = _EVAL_876 | _EVAL_1211;
  assign _EVAL_1426 = _EVAL_1225 == 5'h0;
  assign _EVAL_979 = _EVAL_204 == 5'h5;
  assign _EVAL_984 = _EVAL_1821 ? _EVAL_389 : _EVAL_1574;
  assign _EVAL_750 = _EVAL_1284 ? _EVAL_389 : _EVAL_984;
  assign _EVAL_1791 = _EVAL_641 ? _EVAL_389 : _EVAL_750;
  assign _EVAL_1798 = _EVAL_1188 ? _EVAL_389 : _EVAL_1791;
  assign _EVAL_1091 = 8'hff;
  assign _EVAL_482 = _EVAL_761;
  assign _EVAL_1040 = _EVAL_761;
  assign _EVAL_402 = _EVAL_1567 ? _EVAL_482 : _EVAL_1040;
  assign _EVAL_1208 = _EVAL_496 ? _EVAL_761 : _EVAL_402;
  assign _EVAL_604 = _EVAL_822 ? _EVAL_1702 : _EVAL_1208;
  assign _EVAL_1467 = _EVAL_1345;
  assign _EVAL_164 = _EVAL_1814 == 5'h1;
  assign _EVAL_1803 = _EVAL_447 == 5'h0;
  assign _EVAL_1812 = _EVAL_164 | _EVAL_1803;
  assign _EVAL_1318 = {{1'd0}, _EVAL_1014};
  assign _EVAL_961 = _EVAL_1658 & _EVAL_1736;
  assign _EVAL_425 = _EVAL_641 ? _EVAL_501 : _EVAL_920;
  assign _EVAL_1840 = _EVAL_1188 ? _EVAL_501 : _EVAL_425;
  assign _EVAL_577 = _EVAL_1207 | _EVAL_751;
  assign _EVAL_484 = _EVAL_577 | _EVAL_757;
  assign _EVAL_1230 = _EVAL_484 | _EVAL_1834;
  assign _EVAL_708 = _EVAL_1230 & _EVAL_751;
  assign _EVAL_325 = _EVAL_1347 | _EVAL_708;
  assign _EVAL_241 = _EVAL_37 & _EVAL_325;
  assign _EVAL_931 = 4'h6;
  assign _EVAL_969 = _EVAL_1661[0];
  assign _EVAL_1582 = _EVAL_496 ? 2'h3 : _EVAL_423;
  assign _EVAL_654 = _EVAL_822 ? _EVAL_1719 : _EVAL_1582;
  assign _EVAL_773 = _EVAL_49;
  assign _EVAL_288 = _EVAL_625;
  assign _EVAL_384 = _EVAL_564 ? _EVAL_288 : _EVAL_609;
  assign _EVAL_395 = _EVAL_384;
  assign _EVAL_1839 = _EVAL_90;
  assign _EVAL_667 = _EVAL_1129 | _EVAL_1839;
  assign _EVAL_1069 = data__EVAL_5;
  assign _EVAL_1077 = _EVAL_1069[31:0];
  assign _EVAL_1243 = _EVAL_837 & _EVAL_1254;
  assign _EVAL_1516 = _EVAL_1243 == 1'h0;
  assign _EVAL_1404 = _EVAL_1315 & _EVAL_646;
  assign _EVAL_1668 = _EVAL_1064 & _EVAL_553;
  assign _EVAL_1141 = data__EVAL;
  assign _EVAL_962 = _EVAL_1141[31:0];
  assign _EVAL_1666 = _EVAL_426 == 2'h2;
  assign _EVAL_224 = _EVAL_153 & _EVAL_322;
  assign _EVAL_1465 = _EVAL_1564 ? _EVAL_553 : 1'h0;
  assign _EVAL_1748 = q__EVAL_12;
  assign _EVAL_225 = _EVAL_689[31:8];
  assign _EVAL_1806 = _EVAL_1113 ? _EVAL_1095 : _EVAL_225;
  assign _EVAL_973 = _EVAL_426 == 2'h3;
  assign _EVAL_1183 = {_EVAL_1806,_EVAL_724};
  assign _EVAL_1233 = _EVAL_1219 & _EVAL_939;
  assign _EVAL_1512 = _EVAL_1233 & _EVAL_1729;
  assign _EVAL_1751 = _EVAL_174 & _EVAL_1632;
  assign _EVAL_493 = _EVAL_1069[63:32];
  assign _EVAL_1636 = _EVAL_536[11:0];
  assign _EVAL_1340 = _EVAL_641 ? _EVAL_1488 : _EVAL_1115;
  assign _EVAL_618 = _EVAL_979 & _EVAL_969;
  assign _EVAL_1473 = data__EVAL_7;
  assign _EVAL_1761 = _EVAL_1473[63:32];
  assign _EVAL_532 = q__EVAL_18;
  assign _EVAL_328 = q__EVAL_13;
  assign _EVAL_1711 = _EVAL_1515 == 1'h0;
  assign _EVAL_1065 = q__EVAL_9;
  assign _EVAL_1863 = _EVAL_520 == 2'h0;
  assign _EVAL_226 = _EVAL_1863 ? _EVAL_1504 : _EVAL_995;
  assign _EVAL_1402 = 64'h0;
  assign _EVAL_959 = _EVAL_1322 == 1'h0;
  assign _EVAL_627 = _EVAL_1512 & _EVAL_1543;
  assign _EVAL_1507 = _EVAL_1141[63:32];
  assign _EVAL_949 = _EVAL_16 ? 2'h0 : _EVAL_1461;
  assign _EVAL_1190 = _EVAL_949[0];
  assign _EVAL_1082 = 1'h0;
  assign _EVAL_1588 = _EVAL_569 < 8'h38;
  assign _EVAL_1600 = q__EVAL_2;
  assign _EVAL_167 = _EVAL_322 == _EVAL_1216;
  assign _EVAL_591 = _EVAL_153 & _EVAL_167;
  assign _EVAL_1498 = _EVAL_546 & _EVAL_241;
  assign _EVAL_1272 = _EVAL_1697 | _EVAL_813;
  assign _EVAL_380 = _EVAL_767 == 1'h0;
  assign _EVAL_820 = _EVAL_1073[23:16];
  assign _EVAL_1596 = 3'h6;
  assign _EVAL_584 = _EVAL_1225 == 5'h1;
  assign _EVAL_430 = _EVAL_1616 & _EVAL_1211;
  assign _EVAL_1193 = _EVAL_838 | _EVAL_726;
  assign _EVAL_721 = ~ _EVAL_222;
  assign _EVAL_492 = _EVAL_1751 == 1'h0;
  assign _EVAL_186 = _EVAL_1111 | _EVAL_467;
  assign _EVAL_841 = _EVAL_584 | _EVAL_219;
  assign _EVAL_417 = _EVAL_1107;
  assign _EVAL_1076 = _EVAL_1188 ? 64'h0 : _EVAL_1340;
  assign _EVAL_374 = _EVAL_1272 | _EVAL_16;
  assign _EVAL_1691 = _EVAL_564 ? 4'hf : _EVAL_1381;
  assign _EVAL_1334 = _EVAL_1223 & _EVAL_1254;
  assign _EVAL_458 = _EVAL_1473[31:0];
  assign _EVAL_278 = _EVAL_37 & _EVAL_699;
  assign _EVAL_1361 = _EVAL_949[1];
  assign _EVAL_686 = _EVAL_822 ? _EVAL_1193 : _EVAL_496;
  assign _EVAL_1456 = _EVAL & _EVAL_37;
  assign _EVAL_967 = _EVAL_137;
  assign _EVAL_1570 = _EVAL_478 | _EVAL_1497;
  assign _EVAL_839 = _EVAL_1073[15:8];
  assign _EVAL_895 = _EVAL_380 | _EVAL_278;
  assign _EVAL_666 = _EVAL_822 ? _EVAL_1636 : _EVAL_1385;
  assign _EVAL_1407 = _EVAL_794 & _EVAL_492;
  assign _EVAL_471 = _EVAL_1407 & _EVAL_1711;
  assign _EVAL_1682 = {_EVAL_714, 6'h0};
  assign _EVAL_1416 = _EVAL_1334 & _EVAL_1273;
  assign _EVAL_1329 = 1'h0;
  assign _EVAL_677 = _EVAL_1749 | _EVAL_618;
  assign tlb__EVAL_7 = _EVAL_142;
  assign q__EVAL_6 = _EVAL_18;
  assign tlb__EVAL_54 = _EVAL_97;
  assign _EVAL_34 = _EVAL_981;
  assign _EVAL_130 = _EVAL_1562 | _EVAL_353;
  assign tag_array__EVAL_2 = _EVAL_336 | _EVAL_1760;
  assign MaxPeriodFibonacciLFSR__EVAL_9 = _EVAL_1718 ? _EVAL_1465 : 1'h0;
  assign tag_array__EVAL_1 = _EVAL_1607;
  assign amoalu__EVAL_1 = _EVAL_769;
  assign data__EVAL_0 = dcache_clock_gate_out;
  assign q__EVAL_5 = _EVAL_1736 ? _EVAL_1318 : _EVAL_539;
  assign _EVAL_32 = _EVAL_1088 & _EVAL_1462;
  assign q__EVAL_4 = _EVAL_967;
  assign _EVAL_68 = _EVAL_1183 | _EVAL_1655;
  assign data__EVAL_3 = _EVAL_895;
  assign tlb__EVAL_12 = _EVAL_51;
  assign _EVAL_91 = _EVAL_553 & _EVAL_1718;
  assign tlb__EVAL_71 = _EVAL_141;
  assign tlb__EVAL_46 = _EVAL_62;
  assign data__EVAL_8 = _EVAL_604;
  assign _EVAL_30 = _EVAL_1065;
  assign dcache_clock_gate_en = _EVAL_759;
  assign _EVAL_105 = _EVAL_1570 == 1'h0;
  assign _EVAL_59 = _EVAL_1330;
  assign tlb__EVAL_56 = _EVAL_114;
  assign _EVAL_76 = _EVAL_1403;
  assign tlb__EVAL_48 = _EVAL_11;
  assign tlb__EVAL_20 = _EVAL_89;
  assign tlb__EVAL_25 = _EVAL_140;
  assign tlb__EVAL_2 = _EVAL_1661;
  assign _EVAL_46 = _EVAL_1119;
  assign tlb__EVAL_14 = _EVAL_63;
  assign _EVAL_92 = _EVAL_382;
  assign tlb__EVAL_35 = _EVAL_28;
  assign data__EVAL_4 = _EVAL_666;
  assign tag_array__EVAL_12 = _EVAL_1691[2];
  assign _EVAL_16 = 1'h0;
  assign _EVAL_146 = _EVAL_759;
  assign _EVAL_80 = _EVAL_279;
  assign tlb__EVAL_63 = _EVAL_53;
  assign _EVAL_47 = _EVAL_1390;
  assign tlb__EVAL_29 = _EVAL_155;
  assign _EVAL_70 = _EVAL_1662;
  assign _EVAL_136 = _EVAL_1442 ? 32'h0 : _EVAL_389;
  assign tlb__EVAL_13 = _EVAL_116;
  assign tlb__EVAL_70 = _EVAL_101;
  assign tag_array__EVAL_14 = _EVAL_1691[1];
  assign _EVAL_108 = _EVAL_1649 == 1'h0;
  assign tag_array__EVAL_6 = _EVAL_1607;
  assign tlb__EVAL_28 = _EVAL_2;
  assign tag_array__EVAL_0 = _EVAL_160;
  assign tlb__EVAL_10 = _EVAL_21;
  assign _EVAL_31 = _EVAL_588 ? _EVAL_612 : 1'h0;
  assign amoalu__EVAL_3 = _EVAL_1096;
  assign tlb__EVAL_67 = _EVAL_83;
  assign _EVAL_149 = _EVAL_841 & _EVAL_531;
  assign tlb__EVAL_60 = _EVAL_18;
  assign _EVAL_110 = _EVAL_588 ? _EVAL_1506 : 1'h0;
  assign _EVAL_121 = _EVAL_532;
  assign tlb__EVAL_65 = _EVAL_19;
  assign _EVAL_33 = _EVAL_588 ? _EVAL_1716 : 1'h0;
  assign tlb__EVAL_59 = _EVAL_22;
  assign tlb__EVAL_15 = _EVAL_95;
  assign _EVAL_13 = _EVAL_1748;
  assign _EVAL_24 = _EVAL_1226 | _EVAL_925;
  assign tlb__EVAL_61 = _EVAL_40;
  assign tlb__EVAL_21 = _EVAL_122;
  assign _EVAL_15 = _EVAL_1082;
  assign tlb__EVAL_66 = _EVAL_55;
  assign _EVAL_17 = _EVAL_1853[47:42];
  assign _EVAL_138 = 1'h0;
  assign _EVAL_1 = _EVAL_1718 & _EVAL_667;
  assign tlb__EVAL_49 = _EVAL_204;
  assign tlb__EVAL = _EVAL_118;
  assign tlb__EVAL_37 = _EVAL_144;
  assign tlb__EVAL_26 = _EVAL_58;
  assign tlb__EVAL_45 = _EVAL_23;
  assign tlb__EVAL_36 = _EVAL_9;
  assign tlb__EVAL_30 = _EVAL_45;
  assign tlb__EVAL_27 = _EVAL_69;
  assign tlb__EVAL_1 = _EVAL_25;
  assign tlb__EVAL_11 = dcache_clock_gate_out;
  assign tlb__EVAL_24 = _EVAL_60;
  assign _EVAL_143 = _EVAL_588 ? _EVAL_1805 : 1'h0;
  assign q__EVAL_7 = _EVAL_1736 ? 8'hff : _EVAL_1840;
  assign tlb__EVAL_31 = _EVAL_39;
  assign q__EVAL_0 = dcache_clock_gate_out;
  assign data__EVAL_9 = _EVAL_654;
  assign q__EVAL_3 = _EVAL_1736 ? 4'h6 : _EVAL_638;
  assign _EVAL_48 = _EVAL_321 == 1'h0;
  assign _EVAL_127 = {_EVAL_226,_EVAL_505};
  assign _EVAL_111 = _EVAL_588 ? _EVAL_611 : 1'h0;
  assign tag_array__EVAL_7 = _EVAL_1760 ? _EVAL_395 : _EVAL_395;
  assign q__EVAL_17 = _EVAL_1736 ? 3'h6 : _EVAL_1201;
  assign tlb__EVAL_5 = _EVAL_88;
  assign tlb__EVAL_41 = _EVAL_1315 & _EVAL_677;
  assign _EVAL_100 = _EVAL_276;
  assign _EVAL_73 = _EVAL_680 | _EVAL_738;
  assign _EVAL_134 = _EVAL_626;
  assign tlb__EVAL_39 = _EVAL_115;
  assign data__EVAL_10 = _EVAL_686;
  assign q__EVAL_11 = _EVAL_1736 ? 3'h0 : _EVAL_1198;
  assign _EVAL_103 = _EVAL_804;
  assign _EVAL_61 = _EVAL_1221 & _EVAL_993;
  assign tlb__EVAL_0 = _EVAL_106;
  assign _EVAL_50 = _EVAL_1293;
  assign tlb__EVAL_53 = _EVAL_93;
  assign tlb__EVAL_34 = _EVAL_4;
  assign tlb__EVAL_22 = _EVAL_29;
  assign data__EVAL_2 = _EVAL_1811;
  assign tlb__EVAL_50 = _EVAL_150;
  assign tag_array__EVAL_9 = dcache_clock_gate_out;
  assign dcache_clock_gate_in = _EVAL_72;
  assign _EVAL_41 = _EVAL_328;
  assign tag_array__EVAL_8 = _EVAL_1607;
  assign tag_array__EVAL_10 = _EVAL_1691[0];
  assign data__EVAL_6 = _EVAL_1029;
  assign _EVAL_126 = _EVAL_1589;
  assign tlb__EVAL_47 = _EVAL_74;
  assign tag_array__EVAL_13 = _EVAL_1691[3];
  assign _EVAL = _EVAL_1516 ? 1'h0 : _EVAL_515;
  assign _EVAL_123 = _EVAL_696;
  assign MaxPeriodFibonacciLFSR__EVAL_15 = dcache_clock_gate_out;
  assign _EVAL_82 = _EVAL_186 == 1'h0;
  assign _EVAL_84 = _EVAL_1812 & _EVAL_1658;
  assign _EVAL_6 = _EVAL_1467;
  assign _EVAL_129 = _EVAL_1835 & _EVAL_1588;
  assign tlb__EVAL_62 = _EVAL_81;
  assign tlb__EVAL_3 = _EVAL_79;
  assign amoalu__EVAL_2 = _EVAL_680 | _EVAL_738;
  assign tlb__EVAL_57 = _EVAL_87;
  assign tlb__EVAL_16 = _EVAL_78;
  assign _EVAL_43 = _EVAL_1850 | _EVAL_1442;
  assign q__EVAL_1 = _EVAL_1736 ? 64'h0 : _EVAL_1076;
  assign tlb__EVAL_44 = _EVAL_27;
  assign tlb__EVAL_19 = _EVAL_26;
  assign _EVAL_65 = _EVAL_1686;
  assign tlb__EVAL_42 = _EVAL_131;
  assign tlb__EVAL_40 = _EVAL_132;
  assign _EVAL_64 = _EVAL_588 ? _EVAL_631 : 1'h0;
  assign amoalu__EVAL = _EVAL_393;
  assign _EVAL_44 = _EVAL_165;
  assign _EVAL_147 = _EVAL_1016;
  assign MaxPeriodFibonacciLFSR__EVAL_13 = _EVAL_18;
  assign tag_array__EVAL_4 = _EVAL_1607;
  assign tlb__EVAL_8 = _EVAL_98;
  assign tlb__EVAL_33 = _EVAL_109;
  assign _EVAL_57 = _EVAL_1600;
  assign tlb__EVAL_6 = _EVAL_113;
  assign tlb__EVAL_51 = _EVAL_12;
  assign tlb__EVAL_55 = _EVAL_120;
  assign q__EVAL_14 = _EVAL_1736 ? _EVAL_1682 : _EVAL_1798;
  assign _EVAL_128 = _EVAL_7 & _EVAL_138;
  assign tlb__EVAL_32 = _EVAL_85;
  assign tlb__EVAL_43 = _EVAL_0;
  assign q__EVAL = _EVAL_210 & _EVAL_445;
  assign _EVAL_94 = _EVAL_1096;
  assign _EVAL_75 = _EVAL_936 == 1'h0;
  assign _EVAL_35 = _EVAL_924;
  assign _EVAL_42 = _EVAL_471 & _EVAL_665;
  assign tlb__EVAL_17 = _EVAL_67;
  assign tlb__EVAL_4 = _EVAL_102;
  assign _EVAL_119 = _EVAL_1325;
  assign _EVAL_3 = _EVAL_1442;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_155 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_162 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_165 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_190 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_204 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_211 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_239 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_254 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_263 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_277 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_280 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_291 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_293 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_300 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_320 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_322 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_332 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_341 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_356 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_357 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_359 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_367 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_375 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_376 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_377 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_387 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_389 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_393 = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_396 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_401 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_433 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_451 = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_461 = _RAND_32[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_477 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_487 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_502 = _RAND_35[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_506 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_526 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_541 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_549 = _RAND_39[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_559 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_588 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_598 = _RAND_42[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_611 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_612 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_613 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_614 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_629 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_631 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_632 = _RAND_49[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_655 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_659 = _RAND_51[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_700 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_730 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_732 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_746 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_753 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_759 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_763 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_769 = _RAND_59[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_800 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_801 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_831 = _RAND_62[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_846 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_872 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_874 = _RAND_65[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_893 = _RAND_66[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_907 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_918 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_924 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_926 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_937 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_951 = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_981 = _RAND_73[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_982 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1001 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1032 = _RAND_76[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1049 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1058 = _RAND_78[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1060 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1096 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1100 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1104 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1107 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1109 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1121 = _RAND_85[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1122 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1134 = _RAND_87[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1135 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1140 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1172 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1195 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1200 = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1213 = _RAND_93[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1225 = _RAND_94[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1240 = _RAND_95[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1252 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1269 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1271 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1278 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1300 = _RAND_100[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1316 = _RAND_101[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1319 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1325 = _RAND_103[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1350 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1366 = _RAND_105[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1370 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_1373 = _RAND_107[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1374 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_1387 = _RAND_109[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1390 = _RAND_110[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1417 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1422 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1431 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _EVAL_1439 = _RAND_114[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_1441 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1442 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1444 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1450 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_1486 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1489 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1500 = _RAND_121[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1502 = _RAND_122[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1506 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_1527 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_1541 = _RAND_125[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_1555 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_1569 = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_1594 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_1595 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_1619 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_1620 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_1625 = _RAND_132[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_1626 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_1650 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_1661 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_1688 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_1697 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_1709 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_1716 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_1724 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_1733 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _EVAL_1739 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_1740 = _RAND_143[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _EVAL_1756 = _RAND_144[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _EVAL_1774 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_1784 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _EVAL_1800 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _EVAL_1805 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _EVAL_1810 = _RAND_149[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _EVAL_1814 = _RAND_150[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _EVAL_1827 = _RAND_151[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _EVAL_1831 = _RAND_152[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _EVAL_1832 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _EVAL_1835 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _EVAL_1844 = _RAND_155[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _EVAL_1847 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _EVAL_1851 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge dcache_clock_gate_out) begin
    if (_EVAL_336) begin
      _EVAL_155 <= _EVAL_1606;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_162 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_165 <= _EVAL_1594;
    end
    if (_EVAL_336) begin
      _EVAL_190 <= _EVAL_139;
    end
    if (_EVAL_336) begin
      _EVAL_204 <= _EVAL_135;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_211 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_239 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_16) begin
      if (_EVAL_1400) begin
        _EVAL_254 <= _EVAL_208;
      end else begin
        _EVAL_254 <= _EVAL_203;
      end
    end
    _EVAL_263 <= _EVAL_1602 == 1'h0;
    if (_EVAL_1616) begin
      _EVAL_277 <= _EVAL_258;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_280 <= _EVAL_1370;
        end
      end
    end
    if (_EVAL_591) begin
      _EVAL_291 <= _EVAL_1774;
    end
    if (_EVAL_374) begin
      _EVAL_293 <= _EVAL_962;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_300 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_374) begin
      if (_EVAL_1361) begin
        if (_EVAL_813) begin
          if (_EVAL_1609) begin
            if (_EVAL_722) begin
              _EVAL_320 <= _EVAL_277;
            end else begin
              _EVAL_320 <= _EVAL_1062;
            end
          end else begin
            _EVAL_320 <= _EVAL_1439;
          end
        end else begin
          _EVAL_320 <= _EVAL_258;
        end
      end else begin
        _EVAL_320 <= 4'h0;
      end
    end
    _EVAL_322 <= _EVAL_206 | _EVAL_591;
    if (_EVAL_18) begin
      _EVAL_332 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_1778) begin
                _EVAL_332 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_635) begin
              _EVAL_332 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_1778) begin
                    _EVAL_332 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_1778) begin
                  _EVAL_332 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_1778) begin
              _EVAL_332 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_336) begin
      _EVAL_341 <= _EVAL_1498;
    end
    _EVAL_356 <= _EVAL_643 & _EVAL_1567;
    if (_EVAL_18) begin
      _EVAL_357 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_1455) begin
                _EVAL_357 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_975) begin
              _EVAL_357 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_1455) begin
                    _EVAL_357 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_1455) begin
                  _EVAL_357 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_1455) begin
              _EVAL_357 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_374) begin
      _EVAL_359 <= _EVAL_1077;
    end
    if (_EVAL_374) begin
      _EVAL_367 <= _EVAL_458;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_375 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_376 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_377 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_387 <= _EVAL_1370;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_389 <= tlb__EVAL_38;
    end
    if (_EVAL_430) begin
      if (_EVAL_1542) begin
        _EVAL_393 <= _EVAL_77;
      end else begin
        _EVAL_393 <= _EVAL_1653;
      end
    end
    if (_EVAL_18) begin
      _EVAL_396 <= 3'h0;
    end else begin
      if (_EVAL_1416) begin
        _EVAL_396 <= 3'h0;
      end else begin
        if (_EVAL_1609) begin
          if (_EVAL_560) begin
            _EVAL_396 <= 3'h6;
          end else begin
            if (_EVAL_731) begin
              if (_EVAL_560) begin
                _EVAL_396 <= 3'h7;
              end else begin
                if (_EVAL_1865) begin
                  if (_EVAL_560) begin
                    _EVAL_396 <= 3'h7;
                  end else begin
                    if (_EVAL_720) begin
                      if (_EVAL_560) begin
                        _EVAL_396 <= 3'h0;
                      end else begin
                        if (_EVAL_403) begin
                          if (_EVAL_351) begin
                            _EVAL_396 <= 3'h0;
                          end else begin
                            if (_EVAL_1450) begin
                              if (_EVAL_1098) begin
                                _EVAL_396 <= 3'h2;
                              end else begin
                                if (_EVAL_1430) begin
                                  if (_EVAL_560) begin
                                    _EVAL_396 <= 3'h7;
                                  end else begin
                                    _EVAL_396 <= 3'h3;
                                  end
                                end else begin
                                  if (_EVAL_560) begin
                                    _EVAL_396 <= 3'h0;
                                  end else begin
                                    _EVAL_396 <= 3'h5;
                                  end
                                end
                              end
                            end else begin
                              if (_EVAL_1139) begin
                                if (_EVAL_668) begin
                                  _EVAL_396 <= 3'h1;
                                end else begin
                                  _EVAL_396 <= 3'h6;
                                end
                              end
                            end
                          end
                        end else begin
                          if (_EVAL_1450) begin
                            if (_EVAL_1098) begin
                              _EVAL_396 <= 3'h2;
                            end else begin
                              if (_EVAL_1430) begin
                                if (_EVAL_560) begin
                                  _EVAL_396 <= 3'h7;
                                end else begin
                                  _EVAL_396 <= 3'h3;
                                end
                              end else begin
                                if (_EVAL_560) begin
                                  _EVAL_396 <= 3'h0;
                                end else begin
                                  _EVAL_396 <= 3'h5;
                                end
                              end
                            end
                          end else begin
                            if (_EVAL_1139) begin
                              if (_EVAL_668) begin
                                _EVAL_396 <= 3'h1;
                              end else begin
                                _EVAL_396 <= 3'h6;
                              end
                            end
                          end
                        end
                      end
                    end else begin
                      if (_EVAL_403) begin
                        if (_EVAL_351) begin
                          _EVAL_396 <= 3'h0;
                        end else begin
                          if (_EVAL_1450) begin
                            if (_EVAL_1098) begin
                              _EVAL_396 <= 3'h2;
                            end else begin
                              if (_EVAL_1430) begin
                                if (_EVAL_560) begin
                                  _EVAL_396 <= 3'h7;
                                end else begin
                                  _EVAL_396 <= 3'h3;
                                end
                              end else begin
                                if (_EVAL_560) begin
                                  _EVAL_396 <= 3'h0;
                                end else begin
                                  _EVAL_396 <= 3'h5;
                                end
                              end
                            end
                          end else begin
                            if (_EVAL_1139) begin
                              if (_EVAL_668) begin
                                _EVAL_396 <= 3'h1;
                              end else begin
                                _EVAL_396 <= 3'h6;
                              end
                            end
                          end
                        end
                      end else begin
                        if (_EVAL_1450) begin
                          if (_EVAL_1098) begin
                            _EVAL_396 <= 3'h2;
                          end else begin
                            if (_EVAL_1430) begin
                              if (_EVAL_560) begin
                                _EVAL_396 <= 3'h7;
                              end else begin
                                _EVAL_396 <= 3'h3;
                              end
                            end else begin
                              if (_EVAL_560) begin
                                _EVAL_396 <= 3'h0;
                              end else begin
                                _EVAL_396 <= 3'h5;
                              end
                            end
                          end
                        end else begin
                          if (_EVAL_1139) begin
                            if (_EVAL_668) begin
                              _EVAL_396 <= 3'h1;
                            end else begin
                              _EVAL_396 <= 3'h6;
                            end
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_EVAL_720) begin
                    if (_EVAL_560) begin
                      _EVAL_396 <= 3'h0;
                    end else begin
                      if (_EVAL_403) begin
                        if (_EVAL_351) begin
                          _EVAL_396 <= 3'h0;
                        end else begin
                          _EVAL_396 <= _EVAL_1640;
                        end
                      end else begin
                        _EVAL_396 <= _EVAL_1640;
                      end
                    end
                  end else begin
                    if (_EVAL_403) begin
                      if (_EVAL_351) begin
                        _EVAL_396 <= 3'h0;
                      end else begin
                        _EVAL_396 <= _EVAL_1640;
                      end
                    end else begin
                      _EVAL_396 <= _EVAL_1640;
                    end
                  end
                end
              end
            end else begin
              if (_EVAL_1865) begin
                if (_EVAL_560) begin
                  _EVAL_396 <= 3'h7;
                end else begin
                  if (_EVAL_720) begin
                    if (_EVAL_560) begin
                      _EVAL_396 <= 3'h0;
                    end else begin
                      _EVAL_396 <= _EVAL_1150;
                    end
                  end else begin
                    _EVAL_396 <= _EVAL_1150;
                  end
                end
              end else begin
                if (_EVAL_720) begin
                  if (_EVAL_560) begin
                    _EVAL_396 <= 3'h0;
                  end else begin
                    _EVAL_396 <= _EVAL_1150;
                  end
                end else begin
                  _EVAL_396 <= _EVAL_1150;
                end
              end
            end
          end
        end else begin
          if (_EVAL_731) begin
            if (_EVAL_560) begin
              _EVAL_396 <= 3'h7;
            end else begin
              if (_EVAL_1865) begin
                if (_EVAL_560) begin
                  _EVAL_396 <= 3'h7;
                end else begin
                  _EVAL_396 <= _EVAL_1559;
                end
              end else begin
                _EVAL_396 <= _EVAL_1559;
              end
            end
          end else begin
            if (_EVAL_1865) begin
              if (_EVAL_560) begin
                _EVAL_396 <= 3'h7;
              end else begin
                _EVAL_396 <= _EVAL_1559;
              end
            end else begin
              _EVAL_396 <= _EVAL_1559;
            end
          end
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_401 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_374) begin
      _EVAL_433 <= _EVAL_534;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_451 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_591) begin
      _EVAL_461 <= _EVAL_831;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_477 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_487 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_502 <= 5'h0;
    end else begin
      if (_EVAL_531) begin
        if (_EVAL_682) begin
          if (_EVAL_605) begin
            _EVAL_502 <= _EVAL_908;
          end else begin
            _EVAL_502 <= 5'h0;
          end
        end else begin
          _EVAL_502 <= _EVAL_1526;
        end
      end
    end
    if (_EVAL_591) begin
      _EVAL_506 <= _EVAL_781;
    end
    if (_EVAL_1332) begin
      _EVAL_526 <= tlb__EVAL_23;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_541 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_1332) begin
      if (_EVAL_973) begin
        _EVAL_549 <= _EVAL_1418;
      end else begin
        if (_EVAL_1666) begin
          _EVAL_549 <= _EVAL_799;
        end else begin
          if (_EVAL_563) begin
            _EVAL_549 <= _EVAL_1218;
          end else begin
            _EVAL_549 <= _EVAL_545;
          end
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_559 <= 1'h0;
    end else begin
      if (_EVAL_1609) begin
        if (_EVAL_1085) begin
          _EVAL_559 <= 1'h1;
        end else begin
          if (_EVAL_1718) begin
            if (!(_EVAL_1564)) begin
              if (!(_EVAL_264)) begin
                if (_EVAL_1477) begin
                  _EVAL_559 <= 1'h0;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1718) begin
          if (!(_EVAL_1564)) begin
            if (!(_EVAL_264)) begin
              if (_EVAL_1477) begin
                _EVAL_559 <= 1'h0;
              end
            end
          end
        end
      end
    end
    _EVAL_588 <= tlb__EVAL_41 & _EVAL_1408;
    if (_EVAL_1139) begin
      _EVAL_598 <= 2'h0;
    end else begin
      if (_EVAL_974) begin
        _EVAL_598 <= _EVAL_773;
      end
    end
    if (_EVAL_1332) begin
      _EVAL_611 <= tlb__EVAL_58;
    end
    if (_EVAL_1332) begin
      _EVAL_612 <= tlb__EVAL_69;
    end
    if (_EVAL_18) begin
      _EVAL_613 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_331) begin
                _EVAL_613 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_176) begin
              _EVAL_613 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_331) begin
                    _EVAL_613 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_331) begin
                  _EVAL_613 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_331) begin
              _EVAL_613 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_614 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_629 <= _EVAL_1370;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_631 <= tlb__EVAL_9;
    end
    if (_EVAL_575) begin
      _EVAL_632 <= _EVAL_714;
    end
    if (_EVAL_18) begin
      _EVAL_655 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_661) begin
                _EVAL_655 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_807) begin
              _EVAL_655 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_661) begin
                    _EVAL_655 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_661) begin
                  _EVAL_655 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_661) begin
              _EVAL_655 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_659 <= 5'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1438) begin
          if (_EVAL_1738) begin
            _EVAL_659 <= _EVAL_462;
          end else begin
            _EVAL_659 <= 5'h0;
          end
        end else begin
          _EVAL_659 <= _EVAL_900;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_700 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_591) begin
      _EVAL_730 <= _EVAL_820;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_732 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_1332) begin
      if (_EVAL_1422) begin
        _EVAL_746 <= _EVAL_615;
      end else begin
        _EVAL_746 <= _EVAL_1556;
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_753 <= _EVAL_1370;
        end
      end
    end
    if (_EVAL_591) begin
      _EVAL_763 <= _EVAL_1030;
    end
    if (_EVAL_430) begin
      _EVAL_769 <= _EVAL_204;
    end
    if (_EVAL_18) begin
      _EVAL_800 <= 1'h0;
    end else begin
      if (_EVAL_800) begin
        if (_EVAL_881) begin
          _EVAL_800 <= 1'h0;
        end else begin
          if (_EVAL_1620) begin
            _EVAL_800 <= 1'h1;
          end
        end
      end else begin
        if (_EVAL_1620) begin
          _EVAL_800 <= 1'h1;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_801 <= _EVAL_389;
        end
      end
    end
    if (_EVAL_430) begin
      _EVAL_831 <= _EVAL_258;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_846 <= _EVAL_389;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_872 <= tlb__EVAL_68;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_874 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_893 <= 7'h0;
    end else begin
      if (_EVAL_926) begin
        _EVAL_893 <= 7'h0;
      end else begin
        if (_EVAL_1530) begin
          _EVAL_893 <= 7'h3;
        end else begin
          if (_EVAL_509) begin
            _EVAL_893 <= _EVAL_1652;
          end else begin
            if (_EVAL_575) begin
              if (_EVAL_1376) begin
                _EVAL_893 <= 7'h7f;
              end else begin
                _EVAL_893 <= 7'h0;
              end
            end
          end
        end
      end
    end
    _EVAL_907 <= _EVAL_42;
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_918 <= _EVAL_165;
        end
      end
    end
    _EVAL_924 <= _EVAL_876 & _EVAL_1766;
    if (_EVAL_18) begin
      _EVAL_926 <= 1'h0;
    end else begin
      if (_EVAL_403) begin
        if (_EVAL_351) begin
          _EVAL_926 <= 1'h1;
        end else begin
          _EVAL_926 <= _EVAL_974;
        end
      end else begin
        _EVAL_926 <= _EVAL_974;
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_937 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_951 <= _EVAL_793;
    end
    if (_EVAL_1332) begin
      _EVAL_981 <= _EVAL_1661;
    end
    if (_EVAL_1609) begin
      if (_EVAL_1085) begin
        _EVAL_982 <= _EVAL_1107;
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_1001 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1032 <= 3'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_553) begin
            _EVAL_1032 <= 3'h7;
          end else begin
            if (_EVAL_694) begin
              _EVAL_1032 <= _EVAL_1451;
            end
          end
        end else begin
          if (_EVAL_694) begin
            _EVAL_1032 <= _EVAL_1451;
          end
        end
      end else begin
        if (_EVAL_694) begin
          _EVAL_1032 <= _EVAL_1451;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_1049 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_685) begin
      if (_EVAL_1443) begin
        _EVAL_1058 <= _EVAL_981;
      end
    end
    if (_EVAL_18) begin
      _EVAL_1060 <= 8'hc0;
    end else begin
      _EVAL_1060 <= _EVAL_890[7:0];
    end
    if (_EVAL_430) begin
      _EVAL_1096 <= _EVAL_8;
    end
    if (_EVAL_18) begin
      _EVAL_1100 <= 1'h1;
    end else begin
      if (_EVAL_1422) begin
        if (_EVAL_1278) begin
          if (_EVAL_881) begin
            _EVAL_1100 <= 1'h1;
          end else begin
            if (_EVAL_961) begin
              _EVAL_1100 <= 1'h0;
            end
          end
        end else begin
          if (_EVAL_961) begin
            _EVAL_1100 <= 1'h0;
          end
        end
      end else begin
        if (_EVAL_961) begin
          _EVAL_1100 <= 1'h0;
        end
      end
    end
    _EVAL_1104 <= _EVAL_356 & _EVAL_959;
    if (_EVAL_1139) begin
      _EVAL_1107 <= _EVAL_628;
    end else begin
      if (_EVAL_974) begin
        _EVAL_1107 <= _EVAL_1476;
      end
    end
    if (_EVAL_18) begin
      _EVAL_1109 <= 1'h0;
    end else begin
      _EVAL_1109 <= _EVAL_1404;
    end
    if (_EVAL_591) begin
      _EVAL_1121 <= _EVAL_721;
    end
    if (_EVAL_18) begin
      _EVAL_1122 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_1110) begin
                _EVAL_1122 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_1668) begin
              _EVAL_1122 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_1110) begin
                    _EVAL_1122 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_1110) begin
                  _EVAL_1122 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_1110) begin
              _EVAL_1122 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_1134 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_1135 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_1140 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1172 <= _EVAL_389;
        end
      end
    end
    if (_EVAL_591) begin
      _EVAL_1195 <= _EVAL_839;
    end
    if (_EVAL_1332) begin
      if (_EVAL_973) begin
        _EVAL_1200 <= _EVAL_1561;
      end else begin
        if (_EVAL_1666) begin
          _EVAL_1200 <= _EVAL_313;
        end else begin
          if (_EVAL_563) begin
            _EVAL_1200 <= _EVAL_1264;
          end else begin
            _EVAL_1200 <= _EVAL_693;
          end
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_1213 <= _EVAL_1390;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1225 <= 5'h0;
    end else begin
      if (_EVAL_531) begin
        if (_EVAL_1426) begin
          if (_EVAL_605) begin
            _EVAL_1225 <= _EVAL_908;
          end else begin
            _EVAL_1225 <= 5'h0;
          end
        end else begin
          _EVAL_1225 <= _EVAL_371;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1240 <= _EVAL_1390;
        end
      end
    end
    _EVAL_1252 <= _EVAL_224 & _EVAL_1621;
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_1269 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1271 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_1046) begin
                _EVAL_1271 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_729) begin
              _EVAL_1271 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_1046) begin
                    _EVAL_1271 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_1046) begin
                  _EVAL_1271 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_1046) begin
              _EVAL_1271 <= 1'h1;
            end
          end
        end
      end
    end
    _EVAL_1278 <= _EVAL_1733;
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_1300 <= _EVAL_1390;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_1316 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1319 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_553) begin
            _EVAL_1319 <= 1'h0;
          end else begin
            _EVAL_1319 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1325 <= _EVAL_204;
    end
    if (_EVAL_18) begin
      _EVAL_1350 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_1658) begin
            if (_EVAL_1088) begin
              if (_EVAL_1673) begin
                _EVAL_1350 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_264) begin
            if (_EVAL_1624) begin
              _EVAL_1350 <= 1'h0;
            end else begin
              if (_EVAL_1658) begin
                if (_EVAL_1088) begin
                  if (_EVAL_1673) begin
                    _EVAL_1350 <= 1'h1;
                  end
                end
              end
            end
          end else begin
            if (_EVAL_1658) begin
              if (_EVAL_1088) begin
                if (_EVAL_1673) begin
                  _EVAL_1350 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (_EVAL_1088) begin
            if (_EVAL_1673) begin
              _EVAL_1350 <= 1'h1;
            end
          end
        end
      end
    end
    if (_EVAL_1139) begin
      _EVAL_1366 <= 4'h0;
    end else begin
      if (_EVAL_974) begin
        _EVAL_1366 <= _EVAL_931;
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1370 <= _EVAL_190;
    end
    if (_EVAL_926) begin
      _EVAL_1373 <= _EVAL_793;
    end
    if (_EVAL_336) begin
      if (_EVAL_1516) begin
        _EVAL_1374 <= 1'h1;
      end else begin
        _EVAL_1374 <= _EVAL_117;
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_1387 <= _EVAL_1390;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1390 <= _EVAL_1844;
    end
    if (_EVAL_1332) begin
      _EVAL_1417 <= _EVAL_155;
    end
    if (_EVAL_18) begin
      _EVAL_1422 <= 1'h0;
    end else begin
      if (_EVAL_1422) begin
        if (_EVAL_1491) begin
          _EVAL_1422 <= 1'h0;
        end else begin
          if (_EVAL_685) begin
            if (_EVAL_1443) begin
              _EVAL_1422 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_685) begin
          if (_EVAL_1443) begin
            _EVAL_1422 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_374) begin
      _EVAL_1431 <= _EVAL_600;
    end
    if (_EVAL_926) begin
      _EVAL_1439 <= _EVAL_258;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_1441 <= _EVAL_389;
        end
      end
    end
    _EVAL_1442 <= _EVAL_16;
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_1444 <= _EVAL_1370;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1450 <= 1'h0;
    end else begin
      _EVAL_1450 <= _EVAL_926;
    end
    if (_EVAL_430) begin
      _EVAL_1486 <= _EVAL_1568;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_1489 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1500 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_1139) begin
      _EVAL_1502 <= 3'h0;
    end else begin
      if (_EVAL_974) begin
        _EVAL_1502 <= _EVAL_1529;
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1506 <= tlb__EVAL_52;
    end
    if (_EVAL_374) begin
      _EVAL_1527 <= _EVAL_493;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_1541 <= _EVAL_1390;
        end
      end
    end
    if (_EVAL_336) begin
      _EVAL_1555 <= _EVAL_148;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_331) begin
          _EVAL_1569 <= _EVAL_981;
        end
      end
    end
    if (_EVAL_336) begin
      _EVAL_1594 <= _EVAL_104;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1110) begin
          _EVAL_1595 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_374) begin
      _EVAL_1619 <= _EVAL_1507;
    end
    _EVAL_1620 <= _EVAL_18;
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_1625 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_1626 <= _EVAL_389;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1650 <= _EVAL_1374;
    end
    if (_EVAL_336) begin
      _EVAL_1661 <= _EVAL_56;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1688 <= _EVAL_1370;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1697 <= 1'h0;
    end else begin
      _EVAL_1697 <= _EVAL_1456;
    end
    if (_EVAL_374) begin
      _EVAL_1709 <= _EVAL_1761;
    end
    if (_EVAL_1332) begin
      _EVAL_1716 <= tlb__EVAL_18;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_1724 <= _EVAL_389;
        end
      end
    end
    _EVAL_1733 <= _EVAL_627 & _EVAL_1611;
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1739 <= _EVAL_1650;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1740 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_1756 <= _EVAL_1325;
        end
      end
    end
    if (_EVAL_430) begin
      _EVAL_1774 <= _EVAL_155;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_1784 <= _EVAL_389;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1046) begin
          _EVAL_1800 <= _EVAL_1832;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1805 <= tlb__EVAL_64;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1673) begin
          _EVAL_1810 <= _EVAL_1390;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_1814 <= 5'h0;
    end else begin
      if (_EVAL_1658) begin
        if (_EVAL_879) begin
          if (_EVAL_716) begin
            _EVAL_1814 <= _EVAL_1681;
          end else begin
            _EVAL_1814 <= 5'h0;
          end
        end else begin
          _EVAL_1814 <= _EVAL_1055;
        end
      end
    end
    if (_EVAL_374) begin
      if (_EVAL_1190) begin
        if (_EVAL_813) begin
          if (_EVAL_1609) begin
            if (_EVAL_722) begin
              _EVAL_1827 <= _EVAL_277;
            end else begin
              _EVAL_1827 <= _EVAL_1062;
            end
          end else begin
            _EVAL_1827 <= _EVAL_1439;
          end
        end else begin
          _EVAL_1827 <= _EVAL_258;
        end
      end else begin
        _EVAL_1827 <= 4'h0;
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1455) begin
          _EVAL_1831 <= _EVAL_1390;
        end
      end
    end
    if (_EVAL_1332) begin
      _EVAL_1832 <= _EVAL_1555;
    end
    if (_EVAL_18) begin
      _EVAL_1835 <= 1'h0;
    end else begin
      if (_EVAL_1718) begin
        if (_EVAL_1564) begin
          if (_EVAL_553) begin
            _EVAL_1835 <= 1'h0;
          end else begin
            if (_EVAL_1658) begin
              if (!(_EVAL_1088)) begin
                _EVAL_1835 <= 1'h1;
              end
            end
          end
        end else begin
          if (_EVAL_1658) begin
            if (!(_EVAL_1088)) begin
              _EVAL_1835 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_1658) begin
          if (!(_EVAL_1088)) begin
            _EVAL_1835 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_336) begin
      _EVAL_1844 <= _EVAL_133;
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_661) begin
          _EVAL_1847 <= _EVAL_165;
        end
      end
    end
    if (_EVAL_1658) begin
      if (_EVAL_1088) begin
        if (_EVAL_1778) begin
          _EVAL_1851 <= _EVAL_1370;
        end
      end
    end
  end
  always @(posedge _EVAL_72) begin
    _EVAL_759 <= _EVAL_744 | _EVAL_694;
  end
endmodule
