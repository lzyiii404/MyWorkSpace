//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_64(
  output [31:0] _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  output        _EVAL_3,
  output [2:0]  _EVAL_4,
  input  [4:0]  _EVAL_5,
  output [31:0] _EVAL_6,
  input  [31:0] _EVAL_7,
  input  [2:0]  _EVAL_8,
  output        _EVAL_9,
  output [4:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  output        _EVAL_14,
  input  [3:0]  _EVAL_15,
  output [2:0]  _EVAL_16,
  input  [4:0]  _EVAL_17,
  output [1:0]  _EVAL_18,
  output [2:0]  _EVAL_19,
  input  [31:0] _EVAL_20,
  input         _EVAL_21,
  output [3:0]  _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  output [3:0]  _EVAL_26,
  output [4:0]  _EVAL_27,
  input         _EVAL_28,
  output        _EVAL_29,
  input  [2:0]  _EVAL_30,
  input         _EVAL_31,
  input  [3:0]  _EVAL_32,
  input  [3:0]  _EVAL_33,
  output [3:0]  _EVAL_34,
  output        _EVAL_35,
  output        _EVAL_36,
  output [31:0] _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40
);
  reg  _EVAL_41;
  reg [31:0] _RAND_0;
  reg  _EVAL_93;
  reg [31:0] _RAND_1;
  reg  _EVAL_97;
  reg [31:0] _RAND_2;
  reg  _EVAL_103;
  reg [31:0] _RAND_3;
  reg  _EVAL_107;
  reg [31:0] _RAND_4;
  reg  _EVAL_134;
  reg [31:0] _RAND_5;
  reg  _EVAL_137;
  reg [31:0] _RAND_6;
  reg  _EVAL_143;
  reg [31:0] _RAND_7;
  reg  _EVAL_152;
  reg [31:0] _RAND_8;
  reg  _EVAL_173;
  reg [31:0] _RAND_9;
  reg  _EVAL_174;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_176;
  reg [31:0] _RAND_11;
  reg  _EVAL_186;
  reg [31:0] _RAND_12;
  reg  _EVAL_191;
  reg [31:0] _RAND_13;
  reg  _EVAL_193;
  reg [31:0] _RAND_14;
  reg  _EVAL_210;
  reg [31:0] _RAND_15;
  reg  _EVAL_211;
  reg [31:0] _RAND_16;
  reg  _EVAL_214;
  reg [31:0] _RAND_17;
  reg  _EVAL_215;
  reg [31:0] _RAND_18;
  reg  _EVAL_217;
  reg [31:0] _RAND_19;
  reg  _EVAL_251;
  reg [31:0] _RAND_20;
  reg  _EVAL_252;
  reg [31:0] _RAND_21;
  reg [5:0] _EVAL_253;
  reg [31:0] _RAND_22;
  reg  _EVAL_256;
  reg [31:0] _RAND_23;
  reg  _EVAL_260;
  reg [31:0] _RAND_24;
  reg [1:0] _EVAL_263;
  reg [31:0] _RAND_25;
  reg  _EVAL_266;
  reg [31:0] _RAND_26;
  reg  _EVAL_273;
  reg [31:0] _RAND_27;
  reg  _EVAL_275;
  reg [31:0] _RAND_28;
  reg  _EVAL_276;
  reg [31:0] _RAND_29;
  reg  _EVAL_279;
  reg [31:0] _RAND_30;
  reg [1:0] _EVAL_283;
  reg [31:0] _RAND_31;
  reg  _EVAL_292;
  reg [31:0] _RAND_32;
  reg [5:0] _EVAL_315;
  reg [31:0] _RAND_33;
  reg  _EVAL_337;
  reg [31:0] _RAND_34;
  reg  _EVAL_338;
  reg [31:0] _RAND_35;
  reg  _EVAL_344;
  reg [31:0] _RAND_36;
  reg [1:0] _EVAL_346;
  reg [31:0] _RAND_37;
  wire  _EVAL_87;
  wire [22:0] _EVAL_85;
  wire [7:0] _EVAL_329;
  wire [7:0] _EVAL_320;
  wire [5:0] _EVAL_213;
  wire  _EVAL_319;
  wire [1:0] _EVAL_297;
  wire  _EVAL_246;
  wire  _EVAL_136;
  wire  _EVAL_177;
  wire  _EVAL_301;
  wire  _EVAL_146;
  wire  _EVAL_171;
  wire  _EVAL_285;
  wire  _EVAL_115;
  wire  _EVAL_96;
  wire  _EVAL_72;
  wire [31:0] _EVAL_99;
  wire [32:0] _EVAL_51;
  wire [32:0] _EVAL_64;
  wire [32:0] _EVAL_271;
  wire  _EVAL_183;
  wire [1:0] _EVAL_102;
  wire [32:0] _EVAL_314;
  wire [32:0] _EVAL_195;
  wire [32:0] _EVAL_43;
  wire  _EVAL_50;
  wire [1:0] _EVAL_294;
  wire [1:0] _EVAL_254;
  wire  _EVAL_262;
  wire  _EVAL_242;
  wire  _EVAL_240;
  wire  _EVAL_105;
  wire  _EVAL_59;
  wire  _EVAL_132;
  wire  _EVAL_83;
  wire  _EVAL_327;
  wire  _EVAL_264;
  wire  _EVAL_249;
  wire  _EVAL_175;
  wire  _EVAL_311;
  wire  _EVAL_159;
  wire  _EVAL_272;
  wire  _EVAL_244;
  wire  _EVAL_139;
  wire  _EVAL_68;
  wire  _EVAL_56;
  wire  _EVAL_239;
  wire  _EVAL_153;
  wire  _EVAL_91;
  wire  _EVAL_44;
  wire  _EVAL_208;
  wire  _EVAL_160;
  wire  _EVAL_336;
  wire  _EVAL_278;
  wire  _EVAL_126;
  wire  _EVAL_49;
  wire  _EVAL_268;
  wire  _EVAL_112;
  wire  _EVAL_258;
  wire  _EVAL_142;
  wire  _EVAL_117;
  wire  _EVAL_189;
  wire  _EVAL_89;
  wire  _EVAL_157;
  wire  _EVAL_151;
  wire  _EVAL_222;
  wire  _EVAL_150;
  wire  _EVAL_198;
  wire  _EVAL_168;
  wire  _EVAL_62;
  wire  _EVAL_116;
  wire  _EVAL_187;
  wire  _EVAL_84;
  wire  _EVAL_192;
  wire  _EVAL_236;
  wire  _EVAL_69;
  wire  _EVAL_55;
  wire  _EVAL_170;
  wire  _EVAL_330;
  wire  _EVAL_231;
  wire  _EVAL_156;
  wire  _EVAL_180;
  wire  _EVAL_288;
  wire  _EVAL_172;
  wire [22:0] _EVAL_281;
  wire [7:0] _EVAL_75;
  wire [7:0] _EVAL_114;
  wire [5:0] _EVAL_267;
  wire  _EVAL_135;
  wire [5:0] _EVAL_71;
  wire  _EVAL_110;
  wire  _EVAL_63;
  wire [5:0] _EVAL_141;
  wire  _EVAL_274;
  wire  _EVAL_212;
  assign _EVAL_87 = _EVAL_30[0];
  assign _EVAL_85 = 23'hff << _EVAL_33;
  assign _EVAL_329 = _EVAL_85[7:0];
  assign _EVAL_320 = ~ _EVAL_329;
  assign _EVAL_213 = _EVAL_320[7:2];
  assign _EVAL_319 = _EVAL_315 == 6'h0;
  assign _EVAL_297 = _EVAL_17[4:3];
  assign _EVAL_246 = _EVAL_297 == 2'h0;
  assign _EVAL_136 = _EVAL_246 & _EVAL_319;
  assign _EVAL_177 = _EVAL_134 | _EVAL_93;
  assign _EVAL_301 = _EVAL_177 | _EVAL_210;
  assign _EVAL_146 = _EVAL_301 | _EVAL_217;
  assign _EVAL_171 = _EVAL_146 | _EVAL_107;
  assign _EVAL_285 = _EVAL_171 | _EVAL_41;
  assign _EVAL_115 = _EVAL_285 | _EVAL_152;
  assign _EVAL_96 = _EVAL_115 | _EVAL_292;
  assign _EVAL_72 = _EVAL_136 & _EVAL_96;
  assign _EVAL_99 = _EVAL_20 ^ 32'h40000000;
  assign _EVAL_51 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_64 = $signed(_EVAL_51) & $signed(33'shc0000000);
  assign _EVAL_271 = $signed(_EVAL_64);
  assign _EVAL_183 = $signed(_EVAL_271) == $signed(33'sh0);
  assign _EVAL_102 = {{1'd0}, _EVAL_183};
  assign _EVAL_314 = {1'b0,$signed(_EVAL_20)};
  assign _EVAL_195 = $signed(_EVAL_314) & $signed(33'shc0000000);
  assign _EVAL_43 = $signed(_EVAL_195);
  assign _EVAL_50 = $signed(_EVAL_43) == $signed(33'sh0);
  assign _EVAL_294 = _EVAL_50 ? 2'h2 : 2'h0;
  assign _EVAL_254 = _EVAL_102 | _EVAL_294;
  assign _EVAL_262 = _EVAL_254 == 2'h0;
  assign _EVAL_242 = _EVAL_346 != _EVAL_254;
  assign _EVAL_240 = _EVAL_262 | _EVAL_242;
  assign _EVAL_105 = _EVAL_72 & _EVAL_240;
  assign _EVAL_59 = _EVAL_297 == 2'h1;
  assign _EVAL_132 = _EVAL_59 & _EVAL_319;
  assign _EVAL_83 = _EVAL_191 | _EVAL_174;
  assign _EVAL_327 = _EVAL_83 | _EVAL_344;
  assign _EVAL_264 = _EVAL_327 | _EVAL_266;
  assign _EVAL_249 = _EVAL_264 | _EVAL_193;
  assign _EVAL_175 = _EVAL_249 | _EVAL_338;
  assign _EVAL_311 = _EVAL_175 | _EVAL_279;
  assign _EVAL_159 = _EVAL_311 | _EVAL_276;
  assign _EVAL_272 = _EVAL_132 & _EVAL_159;
  assign _EVAL_244 = _EVAL_263 != _EVAL_254;
  assign _EVAL_139 = _EVAL_262 | _EVAL_244;
  assign _EVAL_68 = _EVAL_272 & _EVAL_139;
  assign _EVAL_56 = _EVAL_105 | _EVAL_68;
  assign _EVAL_239 = _EVAL_297 == 2'h2;
  assign _EVAL_153 = _EVAL_239 & _EVAL_319;
  assign _EVAL_91 = _EVAL_273 | _EVAL_97;
  assign _EVAL_44 = _EVAL_91 | _EVAL_137;
  assign _EVAL_208 = _EVAL_44 | _EVAL_173;
  assign _EVAL_160 = _EVAL_208 | _EVAL_275;
  assign _EVAL_336 = _EVAL_160 | _EVAL_252;
  assign _EVAL_278 = _EVAL_336 | _EVAL_211;
  assign _EVAL_126 = _EVAL_278 | _EVAL_186;
  assign _EVAL_49 = _EVAL_153 & _EVAL_126;
  assign _EVAL_268 = _EVAL_283 != _EVAL_254;
  assign _EVAL_112 = _EVAL_262 | _EVAL_268;
  assign _EVAL_258 = _EVAL_49 & _EVAL_112;
  assign _EVAL_142 = _EVAL_56 | _EVAL_258;
  assign _EVAL_117 = _EVAL_297 == 2'h3;
  assign _EVAL_189 = _EVAL_117 & _EVAL_319;
  assign _EVAL_89 = _EVAL_337 | _EVAL_103;
  assign _EVAL_157 = _EVAL_89 | _EVAL_251;
  assign _EVAL_151 = _EVAL_157 | _EVAL_215;
  assign _EVAL_222 = _EVAL_151 | _EVAL_260;
  assign _EVAL_150 = _EVAL_222 | _EVAL_143;
  assign _EVAL_198 = _EVAL_150 | _EVAL_214;
  assign _EVAL_168 = _EVAL_198 | _EVAL_256;
  assign _EVAL_62 = _EVAL_189 & _EVAL_168;
  assign _EVAL_116 = _EVAL_176 != _EVAL_254;
  assign _EVAL_187 = _EVAL_262 | _EVAL_116;
  assign _EVAL_84 = _EVAL_62 & _EVAL_187;
  assign _EVAL_192 = _EVAL_142 | _EVAL_84;
  assign _EVAL_236 = _EVAL_192 == 1'h0;
  assign _EVAL_69 = _EVAL_1 & _EVAL_236;
  assign _EVAL_55 = _EVAL_69 & _EVAL_39;
  assign _EVAL_170 = _EVAL_319 & _EVAL_55;
  assign _EVAL_330 = _EVAL_253 == 6'h0;
  assign _EVAL_231 = _EVAL_30 != 3'h6;
  assign _EVAL_156 = _EVAL_330 & _EVAL_231;
  assign _EVAL_180 = _EVAL_12 & _EVAL_31;
  assign _EVAL_288 = _EVAL_156 & _EVAL_180;
  assign _EVAL_172 = _EVAL_8[2];
  assign _EVAL_281 = 23'hff << _EVAL_15;
  assign _EVAL_75 = _EVAL_281[7:0];
  assign _EVAL_114 = ~ _EVAL_75;
  assign _EVAL_267 = _EVAL_114[7:2];
  assign _EVAL_135 = _EVAL_172 == 1'h0;
  assign _EVAL_71 = _EVAL_315 - 6'h1;
  assign _EVAL_110 = _EVAL_55 & _EVAL_246;
  assign _EVAL_63 = _EVAL_55 & _EVAL_117;
  assign _EVAL_141 = _EVAL_253 - 6'h1;
  assign _EVAL_274 = _EVAL_55 & _EVAL_59;
  assign _EVAL_212 = _EVAL_55 & _EVAL_239;
  assign _EVAL_25 = _EVAL_23;
  assign _EVAL = _EVAL_7;
  assign _EVAL_29 = _EVAL_11;
  assign _EVAL_35 = _EVAL_1 & _EVAL_236;
  assign _EVAL_6 = _EVAL_13;
  assign _EVAL_34 = _EVAL_33;
  assign _EVAL_4 = _EVAL_8;
  assign _EVAL_10 = _EVAL_5;
  assign _EVAL_14 = _EVAL_39 & _EVAL_236;
  assign _EVAL_16 = _EVAL_30;
  assign _EVAL_19 = _EVAL_0;
  assign _EVAL_24 = _EVAL_40;
  assign _EVAL_36 = _EVAL_38;
  assign _EVAL_37 = _EVAL_20;
  assign _EVAL_9 = _EVAL_31;
  assign _EVAL_22 = _EVAL_32;
  assign _EVAL_18 = _EVAL_2;
  assign _EVAL_3 = _EVAL_12;
  assign _EVAL_26 = _EVAL_15;
  assign _EVAL_27 = _EVAL_17;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_41 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_93 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_97 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_103 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_107 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_134 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_137 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_143 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_152 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_173 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_174 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_176 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_186 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_191 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_193 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_210 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_211 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_214 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_215 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_217 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_251 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_252 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_253 = _RAND_22[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_256 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_260 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_263 = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_266 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_273 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_275 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_276 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_279 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_283 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_292 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_315 = _RAND_33[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_337 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_338 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_344 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_346 = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_28) begin
    if (_EVAL_21) begin
      _EVAL_41 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h5 == _EVAL_5) begin
          _EVAL_41 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h5 == _EVAL_17) begin
              _EVAL_41 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h5 == _EVAL_17) begin
            _EVAL_41 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_93 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1 == _EVAL_5) begin
          _EVAL_93 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1 == _EVAL_17) begin
              _EVAL_93 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1 == _EVAL_17) begin
            _EVAL_93 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_97 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h11 == _EVAL_5) begin
          _EVAL_97 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h11 == _EVAL_17) begin
              _EVAL_97 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h11 == _EVAL_17) begin
            _EVAL_97 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_103 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h19 == _EVAL_5) begin
          _EVAL_103 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h19 == _EVAL_17) begin
              _EVAL_103 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h19 == _EVAL_17) begin
            _EVAL_103 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_107 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h4 == _EVAL_5) begin
          _EVAL_107 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h4 == _EVAL_17) begin
              _EVAL_107 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h4 == _EVAL_17) begin
            _EVAL_107 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_134 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h0 == _EVAL_5) begin
          _EVAL_134 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h0 == _EVAL_17) begin
              _EVAL_134 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h0 == _EVAL_17) begin
            _EVAL_134 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_137 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h12 == _EVAL_5) begin
          _EVAL_137 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h12 == _EVAL_17) begin
              _EVAL_137 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h12 == _EVAL_17) begin
            _EVAL_137 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_143 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1d == _EVAL_5) begin
          _EVAL_143 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1d == _EVAL_17) begin
              _EVAL_143 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1d == _EVAL_17) begin
            _EVAL_143 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_152 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h6 == _EVAL_5) begin
          _EVAL_152 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h6 == _EVAL_17) begin
              _EVAL_152 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h6 == _EVAL_17) begin
            _EVAL_152 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_173 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h13 == _EVAL_5) begin
          _EVAL_173 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h13 == _EVAL_17) begin
              _EVAL_173 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h13 == _EVAL_17) begin
            _EVAL_173 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_174 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h9 == _EVAL_5) begin
          _EVAL_174 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h9 == _EVAL_17) begin
              _EVAL_174 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h9 == _EVAL_17) begin
            _EVAL_174 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_176 <= _EVAL_254;
    end
    if (_EVAL_21) begin
      _EVAL_186 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h17 == _EVAL_5) begin
          _EVAL_186 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h17 == _EVAL_17) begin
              _EVAL_186 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h17 == _EVAL_17) begin
            _EVAL_186 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_191 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h8 == _EVAL_5) begin
          _EVAL_191 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h8 == _EVAL_17) begin
              _EVAL_191 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h8 == _EVAL_17) begin
            _EVAL_191 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_193 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'hc == _EVAL_5) begin
          _EVAL_193 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'hc == _EVAL_17) begin
              _EVAL_193 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'hc == _EVAL_17) begin
            _EVAL_193 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_210 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h2 == _EVAL_5) begin
          _EVAL_210 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h2 == _EVAL_17) begin
              _EVAL_210 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h2 == _EVAL_17) begin
            _EVAL_210 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_211 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h16 == _EVAL_5) begin
          _EVAL_211 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h16 == _EVAL_17) begin
              _EVAL_211 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h16 == _EVAL_17) begin
            _EVAL_211 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_214 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1e == _EVAL_5) begin
          _EVAL_214 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1e == _EVAL_17) begin
              _EVAL_214 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1e == _EVAL_17) begin
            _EVAL_214 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_215 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1b == _EVAL_5) begin
          _EVAL_215 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1b == _EVAL_17) begin
              _EVAL_215 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1b == _EVAL_17) begin
            _EVAL_215 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_217 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h3 == _EVAL_5) begin
          _EVAL_217 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h3 == _EVAL_17) begin
              _EVAL_217 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h3 == _EVAL_17) begin
            _EVAL_217 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_251 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1a == _EVAL_5) begin
          _EVAL_251 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1a == _EVAL_17) begin
              _EVAL_251 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1a == _EVAL_17) begin
            _EVAL_251 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_252 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h15 == _EVAL_5) begin
          _EVAL_252 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h15 == _EVAL_17) begin
              _EVAL_252 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h15 == _EVAL_17) begin
            _EVAL_252 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_253 <= 6'h0;
    end else begin
      if (_EVAL_180) begin
        if (_EVAL_330) begin
          if (_EVAL_87) begin
            _EVAL_253 <= _EVAL_213;
          end else begin
            _EVAL_253 <= 6'h0;
          end
        end else begin
          _EVAL_253 <= _EVAL_141;
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_256 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1f == _EVAL_5) begin
          _EVAL_256 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1f == _EVAL_17) begin
              _EVAL_256 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1f == _EVAL_17) begin
            _EVAL_256 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_260 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h1c == _EVAL_5) begin
          _EVAL_260 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h1c == _EVAL_17) begin
              _EVAL_260 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h1c == _EVAL_17) begin
            _EVAL_260 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_274) begin
      _EVAL_263 <= _EVAL_254;
    end
    if (_EVAL_21) begin
      _EVAL_266 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'hb == _EVAL_5) begin
          _EVAL_266 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'hb == _EVAL_17) begin
              _EVAL_266 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'hb == _EVAL_17) begin
            _EVAL_266 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_273 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h10 == _EVAL_5) begin
          _EVAL_273 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h10 == _EVAL_17) begin
              _EVAL_273 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h10 == _EVAL_17) begin
            _EVAL_273 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_275 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h14 == _EVAL_5) begin
          _EVAL_275 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h14 == _EVAL_17) begin
              _EVAL_275 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h14 == _EVAL_17) begin
            _EVAL_275 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_276 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'hf == _EVAL_5) begin
          _EVAL_276 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'hf == _EVAL_17) begin
              _EVAL_276 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'hf == _EVAL_17) begin
            _EVAL_276 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_279 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'he == _EVAL_5) begin
          _EVAL_279 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'he == _EVAL_17) begin
              _EVAL_279 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'he == _EVAL_17) begin
            _EVAL_279 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_212) begin
      _EVAL_283 <= _EVAL_254;
    end
    if (_EVAL_21) begin
      _EVAL_292 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h7 == _EVAL_5) begin
          _EVAL_292 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h7 == _EVAL_17) begin
              _EVAL_292 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h7 == _EVAL_17) begin
            _EVAL_292 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_315 <= 6'h0;
    end else begin
      if (_EVAL_55) begin
        if (_EVAL_319) begin
          if (_EVAL_135) begin
            _EVAL_315 <= _EVAL_267;
          end else begin
            _EVAL_315 <= 6'h0;
          end
        end else begin
          _EVAL_315 <= _EVAL_71;
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_337 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'h18 == _EVAL_5) begin
          _EVAL_337 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'h18 == _EVAL_17) begin
              _EVAL_337 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'h18 == _EVAL_17) begin
            _EVAL_337 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_338 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'hd == _EVAL_5) begin
          _EVAL_338 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'hd == _EVAL_17) begin
              _EVAL_338 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'hd == _EVAL_17) begin
            _EVAL_338 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_21) begin
      _EVAL_344 <= 1'h0;
    end else begin
      if (_EVAL_288) begin
        if (5'ha == _EVAL_5) begin
          _EVAL_344 <= 1'h0;
        end else begin
          if (_EVAL_170) begin
            if (5'ha == _EVAL_17) begin
              _EVAL_344 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_170) begin
          if (5'ha == _EVAL_17) begin
            _EVAL_344 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_110) begin
      _EVAL_346 <= _EVAL_254;
    end
  end
endmodule
