//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_277(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  input  [31:0] _EVAL_1,
  output        _EVAL_2,
  output [6:0]  _EVAL_3,
  output [31:0] _EVAL_4,
  output [2:0]  _EVAL_5,
  input  [6:0]  _EVAL_6,
  output        _EVAL_7,
  input  [31:0] _EVAL_8,
  input  [24:0] _EVAL_9,
  input  [1:0]  _EVAL_10,
  output [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  output [2:0]  _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  input  [24:0] _EVAL_22,
  output [2:0]  _EVAL_23,
  output [2:0]  _EVAL_24,
  output [31:0] _EVAL_25,
  output [24:0] _EVAL_26,
  input         _EVAL_27,
  output [6:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  output [3:0]  _EVAL_31,
  input  [1:0]  _EVAL_32,
  output        _EVAL_33,
  output [1:0]  _EVAL_34,
  input  [6:0]  _EVAL_35,
  output [1:0]  _EVAL_36,
  output [1:0]  _EVAL_37,
  output        _EVAL_38,
  input  [2:0]  _EVAL_39,
  input         _EVAL_40,
  input  [3:0]  _EVAL_41,
  input  [6:0]  _EVAL_42,
  input  [3:0]  _EVAL_43,
  output        _EVAL_44,
  output [31:0] _EVAL_45,
  input  [2:0]  _EVAL_46,
  input         _EVAL_47,
  output [1:0]  _EVAL_48,
  input  [2:0]  _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input  [2:0]  _EVAL_52,
  output        _EVAL_53,
  output [2:0]  _EVAL_54,
  output [6:0]  _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  input  [2:0]  _EVAL_60
);
  wire [24:0] RationalCrossingSink__EVAL;
  wire [2:0] RationalCrossingSink__EVAL_0;
  wire [1:0] RationalCrossingSink__EVAL_1;
  wire [2:0] RationalCrossingSink__EVAL_2;
  wire  RationalCrossingSink__EVAL_3;
  wire  RationalCrossingSink__EVAL_4;
  wire [2:0] RationalCrossingSink__EVAL_5;
  wire [31:0] RationalCrossingSink__EVAL_6;
  wire [2:0] RationalCrossingSink__EVAL_7;
  wire [3:0] RationalCrossingSink__EVAL_8;
  wire  RationalCrossingSink__EVAL_9;
  wire [2:0] RationalCrossingSink__EVAL_10;
  wire [24:0] RationalCrossingSink__EVAL_11;
  wire [6:0] RationalCrossingSink__EVAL_12;
  wire  RationalCrossingSink__EVAL_13;
  wire [2:0] RationalCrossingSink__EVAL_14;
  wire [31:0] RationalCrossingSink__EVAL_15;
  wire  RationalCrossingSink__EVAL_16;
  wire [24:0] RationalCrossingSink__EVAL_17;
  wire [31:0] RationalCrossingSink__EVAL_18;
  wire [6:0] RationalCrossingSink__EVAL_19;
  wire [3:0] RationalCrossingSink__EVAL_20;
  wire [2:0] RationalCrossingSink__EVAL_21;
  wire  RationalCrossingSink__EVAL_22;
  wire  RationalCrossingSink__EVAL_23;
  wire [6:0] RationalCrossingSink__EVAL_24;
  wire [2:0] RationalCrossingSink__EVAL_25;
  wire [2:0] RationalCrossingSink__EVAL_26;
  wire  RationalCrossingSink__EVAL_27;
  wire  RationalCrossingSink__EVAL_28;
  wire [1:0] RationalCrossingSink__EVAL_29;
  wire [3:0] RationalCrossingSink__EVAL_30;
  wire  RationalCrossingSource__EVAL;
  wire  RationalCrossingSource__EVAL_0;
  wire  RationalCrossingSource__EVAL_1;
  wire [2:0] RationalCrossingSource__EVAL_2;
  wire [6:0] RationalCrossingSource__EVAL_3;
  wire  RationalCrossingSource__EVAL_4;
  wire [2:0] RationalCrossingSource__EVAL_5;
  wire [31:0] RationalCrossingSource__EVAL_6;
  wire [6:0] RationalCrossingSource__EVAL_7;
  wire [1:0] RationalCrossingSource__EVAL_8;
  wire  RationalCrossingSource__EVAL_9;
  wire  RationalCrossingSource__EVAL_10;
  wire  RationalCrossingSource__EVAL_11;
  wire [1:0] RationalCrossingSource__EVAL_12;
  wire  RationalCrossingSource__EVAL_13;
  wire  RationalCrossingSource__EVAL_14;
  wire [31:0] RationalCrossingSource__EVAL_15;
  wire  RationalCrossingSource__EVAL_16;
  wire [2:0] RationalCrossingSource__EVAL_17;
  wire [6:0] RationalCrossingSource__EVAL_18;
  wire [1:0] RationalCrossingSource__EVAL_19;
  wire [2:0] RationalCrossingSource__EVAL_20;
  wire  RationalCrossingSource__EVAL_21;
  wire [31:0] RationalCrossingSource__EVAL_22;
  wire [1:0] RationalCrossingSource__EVAL_23;
  wire  RationalCrossingSource__EVAL_24;
  wire [1:0] RationalCrossingSource__EVAL_25;
  wire  RationalCrossingSource__EVAL_26;
  wire [2:0] RationalCrossingSource__EVAL_27;
  wire  RationalCrossingSource__EVAL_28;
  wire  RationalCrossingSource__EVAL_29;
  wire [2:0] RationalCrossingSource__EVAL_30;
  SiFive__EVAL_275 RationalCrossingSink (
    ._EVAL(RationalCrossingSink__EVAL),
    ._EVAL_0(RationalCrossingSink__EVAL_0),
    ._EVAL_1(RationalCrossingSink__EVAL_1),
    ._EVAL_2(RationalCrossingSink__EVAL_2),
    ._EVAL_3(RationalCrossingSink__EVAL_3),
    ._EVAL_4(RationalCrossingSink__EVAL_4),
    ._EVAL_5(RationalCrossingSink__EVAL_5),
    ._EVAL_6(RationalCrossingSink__EVAL_6),
    ._EVAL_7(RationalCrossingSink__EVAL_7),
    ._EVAL_8(RationalCrossingSink__EVAL_8),
    ._EVAL_9(RationalCrossingSink__EVAL_9),
    ._EVAL_10(RationalCrossingSink__EVAL_10),
    ._EVAL_11(RationalCrossingSink__EVAL_11),
    ._EVAL_12(RationalCrossingSink__EVAL_12),
    ._EVAL_13(RationalCrossingSink__EVAL_13),
    ._EVAL_14(RationalCrossingSink__EVAL_14),
    ._EVAL_15(RationalCrossingSink__EVAL_15),
    ._EVAL_16(RationalCrossingSink__EVAL_16),
    ._EVAL_17(RationalCrossingSink__EVAL_17),
    ._EVAL_18(RationalCrossingSink__EVAL_18),
    ._EVAL_19(RationalCrossingSink__EVAL_19),
    ._EVAL_20(RationalCrossingSink__EVAL_20),
    ._EVAL_21(RationalCrossingSink__EVAL_21),
    ._EVAL_22(RationalCrossingSink__EVAL_22),
    ._EVAL_23(RationalCrossingSink__EVAL_23),
    ._EVAL_24(RationalCrossingSink__EVAL_24),
    ._EVAL_25(RationalCrossingSink__EVAL_25),
    ._EVAL_26(RationalCrossingSink__EVAL_26),
    ._EVAL_27(RationalCrossingSink__EVAL_27),
    ._EVAL_28(RationalCrossingSink__EVAL_28),
    ._EVAL_29(RationalCrossingSink__EVAL_29),
    ._EVAL_30(RationalCrossingSink__EVAL_30)
  );
  SiFive__EVAL_276 RationalCrossingSource (
    ._EVAL(RationalCrossingSource__EVAL),
    ._EVAL_0(RationalCrossingSource__EVAL_0),
    ._EVAL_1(RationalCrossingSource__EVAL_1),
    ._EVAL_2(RationalCrossingSource__EVAL_2),
    ._EVAL_3(RationalCrossingSource__EVAL_3),
    ._EVAL_4(RationalCrossingSource__EVAL_4),
    ._EVAL_5(RationalCrossingSource__EVAL_5),
    ._EVAL_6(RationalCrossingSource__EVAL_6),
    ._EVAL_7(RationalCrossingSource__EVAL_7),
    ._EVAL_8(RationalCrossingSource__EVAL_8),
    ._EVAL_9(RationalCrossingSource__EVAL_9),
    ._EVAL_10(RationalCrossingSource__EVAL_10),
    ._EVAL_11(RationalCrossingSource__EVAL_11),
    ._EVAL_12(RationalCrossingSource__EVAL_12),
    ._EVAL_13(RationalCrossingSource__EVAL_13),
    ._EVAL_14(RationalCrossingSource__EVAL_14),
    ._EVAL_15(RationalCrossingSource__EVAL_15),
    ._EVAL_16(RationalCrossingSource__EVAL_16),
    ._EVAL_17(RationalCrossingSource__EVAL_17),
    ._EVAL_18(RationalCrossingSource__EVAL_18),
    ._EVAL_19(RationalCrossingSource__EVAL_19),
    ._EVAL_20(RationalCrossingSource__EVAL_20),
    ._EVAL_21(RationalCrossingSource__EVAL_21),
    ._EVAL_22(RationalCrossingSource__EVAL_22),
    ._EVAL_23(RationalCrossingSource__EVAL_23),
    ._EVAL_24(RationalCrossingSource__EVAL_24),
    ._EVAL_25(RationalCrossingSource__EVAL_25),
    ._EVAL_26(RationalCrossingSource__EVAL_26),
    ._EVAL_27(RationalCrossingSource__EVAL_27),
    ._EVAL_28(RationalCrossingSource__EVAL_28),
    ._EVAL_29(RationalCrossingSource__EVAL_29),
    ._EVAL_30(RationalCrossingSource__EVAL_30)
  );
  assign RationalCrossingSink__EVAL_19 = _EVAL_35;
  assign RationalCrossingSink__EVAL_4 = _EVAL_58;
  assign _EVAL_11 = RationalCrossingSink__EVAL_10;
  assign _EVAL_2 = RationalCrossingSource__EVAL;
  assign RationalCrossingSource__EVAL_1 = _EVAL_21;
  assign RationalCrossingSink__EVAL_24 = _EVAL_42;
  assign RationalCrossingSink__EVAL_2 = _EVAL_46;
  assign RationalCrossingSink__EVAL_22 = _EVAL_27;
  assign RationalCrossingSource__EVAL_25 = _EVAL_32;
  assign RationalCrossingSink__EVAL_5 = _EVAL_12;
  assign _EVAL_18 = RationalCrossingSource__EVAL_26;
  assign _EVAL_5 = RationalCrossingSink__EVAL_14;
  assign RationalCrossingSink__EVAL_11 = _EVAL_9;
  assign _EVAL_37 = RationalCrossingSource__EVAL_8;
  assign RationalCrossingSource__EVAL_22 = _EVAL_8;
  assign RationalCrossingSource__EVAL_11 = _EVAL_27;
  assign _EVAL_3 = RationalCrossingSource__EVAL_3;
  assign _EVAL_30 = RationalCrossingSource__EVAL_30;
  assign _EVAL_38 = RationalCrossingSource__EVAL_4;
  assign RationalCrossingSource__EVAL_20 = _EVAL_60;
  assign _EVAL_7 = RationalCrossingSource__EVAL_9;
  assign RationalCrossingSource__EVAL_19 = _EVAL_10;
  assign RationalCrossingSource__EVAL_2 = _EVAL_15;
  assign RationalCrossingSink__EVAL_16 = _EVAL_14;
  assign RationalCrossingSource__EVAL_18 = _EVAL_6;
  assign RationalCrossingSink__EVAL_0 = _EVAL_52;
  assign RationalCrossingSink__EVAL_15 = _EVAL_0;
  assign RationalCrossingSink__EVAL_23 = _EVAL_40;
  assign RationalCrossingSource__EVAL_0 = _EVAL_57;
  assign _EVAL = RationalCrossingSource__EVAL_16;
  assign _EVAL_33 = RationalCrossingSource__EVAL_24;
  assign _EVAL_45 = RationalCrossingSink__EVAL_6;
  assign RationalCrossingSource__EVAL_14 = _EVAL_59;
  assign _EVAL_24 = RationalCrossingSource__EVAL_17;
  assign RationalCrossingSink__EVAL_9 = _EVAL_21;
  assign RationalCrossingSource__EVAL_29 = _EVAL_51;
  assign RationalCrossingSource__EVAL_28 = _EVAL_56;
  assign _EVAL_53 = RationalCrossingSource__EVAL_10;
  assign _EVAL_19 = RationalCrossingSink__EVAL_25;
  assign RationalCrossingSink__EVAL_26 = _EVAL_49;
  assign _EVAL_36 = RationalCrossingSink__EVAL_1;
  assign _EVAL_44 = RationalCrossingSink__EVAL_27;
  assign RationalCrossingSink__EVAL_18 = _EVAL_1;
  assign RationalCrossingSink__EVAL_17 = _EVAL_22;
  assign RationalCrossingSink__EVAL_28 = _EVAL_47;
  assign _EVAL_31 = RationalCrossingSink__EVAL_30;
  assign _EVAL_20 = RationalCrossingSink__EVAL_3;
  assign _EVAL_16 = RationalCrossingSink__EVAL_13;
  assign _EVAL_4 = RationalCrossingSource__EVAL_6;
  assign RationalCrossingSink__EVAL_7 = _EVAL_29;
  assign _EVAL_54 = RationalCrossingSource__EVAL_5;
  assign RationalCrossingSink__EVAL_20 = _EVAL_43;
  assign _EVAL_25 = RationalCrossingSource__EVAL_15;
  assign RationalCrossingSink__EVAL_8 = _EVAL_41;
  assign RationalCrossingSink__EVAL_29 = _EVAL_13;
  assign _EVAL_23 = RationalCrossingSource__EVAL_27;
  assign _EVAL_34 = RationalCrossingSource__EVAL_12;
  assign _EVAL_28 = RationalCrossingSink__EVAL_12;
  assign _EVAL_55 = RationalCrossingSource__EVAL_7;
  assign _EVAL_26 = RationalCrossingSink__EVAL;
  assign _EVAL_48 = RationalCrossingSource__EVAL_23;
  assign RationalCrossingSource__EVAL_13 = _EVAL_50;
  assign RationalCrossingSink__EVAL_21 = _EVAL_39;
  assign _EVAL_17 = RationalCrossingSource__EVAL_21;
endmodule
