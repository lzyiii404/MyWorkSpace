//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_314_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [3:0]  _EVAL_5,
  input         _EVAL_6,
  input  [14:0] _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [11:0] _EVAL_12,
  input         _EVAL_13,
  input  [11:0] _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_58;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_59;
  reg [31:0] _RAND_1;
  reg  _EVAL_71;
  reg [31:0] _RAND_2;
  reg [11:0] _EVAL_72;
  reg [31:0] _RAND_3;
  reg [2335:0] _EVAL_99;
  reg [2335:0] _RAND_4;
  reg [14:0] _EVAL_104;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_107;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_115;
  reg [31:0] _RAND_7;
  reg  _EVAL_131;
  reg [31:0] _RAND_8;
  reg  _EVAL_136;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_171;
  reg [31:0] _RAND_10;
  reg  _EVAL_215;
  reg [31:0] _RAND_11;
  reg [1:0] _EVAL_223;
  reg [31:0] _RAND_12;
  reg [11:0] _EVAL_227;
  reg [31:0] _RAND_13;
  wire  _EVAL_137;
  wire [2335:0] _EVAL_160;
  wire  _EVAL_24;
  wire  _EVAL_98;
  wire [1:0] _EVAL_105;
  wire [1:0] _EVAL_158;
  wire  _EVAL_41;
  wire  _EVAL_82;
  wire  _EVAL_151;
  wire  _EVAL_91;
  wire  _EVAL_166;
  wire  _EVAL_159;
  wire  _EVAL_172;
  wire  _EVAL_139;
  wire  _EVAL_126;
  wire  _EVAL_185;
  wire  _EVAL_117;
  wire  _EVAL_89;
  wire  _EVAL_182;
  wire  _EVAL_38;
  wire  _EVAL_141;
  wire  _EVAL_175;
  wire  _EVAL_23;
  wire  _EVAL_102;
  wire  _EVAL_130;
  wire  _EVAL_236;
  wire  _EVAL_147;
  wire  _EVAL_208;
  wire [3:0] _EVAL_93;
  wire  _EVAL_20;
  wire  _EVAL_17;
  wire  _EVAL_103;
  wire [4:0] _EVAL_46;
  wire [1:0] _EVAL_210;
  wire  _EVAL_177;
  wire [14:0] _EVAL_212;
  wire  _EVAL_194;
  wire  _EVAL_149;
  wire  _EVAL_76;
  wire  _EVAL_123;
  wire  _EVAL_198;
  wire  _EVAL_178;
  wire  _EVAL_180;
  wire  _EVAL_87;
  wire  _EVAL_85;
  wire  _EVAL_183;
  wire  _EVAL_196;
  wire  _EVAL_135;
  wire  _EVAL_233;
  wire  _EVAL_36;
  wire  _EVAL_129;
  wire  _EVAL_232;
  wire [4095:0] _EVAL_86;
  wire [4095:0] _EVAL_106;
  wire [2335:0] _EVAL_118;
  wire  _EVAL_51;
  wire  _EVAL_235;
  wire  _EVAL_18;
  wire  _EVAL_67;
  wire  _EVAL_95;
  wire [2335:0] _EVAL_174;
  wire  _EVAL_56;
  wire  _EVAL_32;
  wire  _EVAL_22;
  wire  _EVAL_199;
  wire  _EVAL_202;
  wire  _EVAL_146;
  wire  _EVAL_33;
  wire  _EVAL_148;
  wire  _EVAL_111;
  wire  _EVAL_203;
  wire  _EVAL_61;
  wire  _EVAL_84;
  wire  _EVAL_28;
  wire  _EVAL_64;
  wire  _EVAL_200;
  wire [4095:0] _EVAL_228;
  wire [4095:0] _EVAL_220;
  wire [2335:0] _EVAL_21;
  wire  _EVAL_15;
  wire  _EVAL_37;
  wire  _EVAL_65;
  wire  _EVAL_77;
  wire  _EVAL_122;
  wire  _EVAL_119;
  wire  _EVAL_150;
  wire  _EVAL_54;
  wire  _EVAL_140;
  wire  _EVAL_164;
  wire [1:0] _EVAL_189;
  wire [14:0] _EVAL_218;
  wire [14:0] _EVAL_176;
  wire  _EVAL_48;
  wire [15:0] _EVAL_214;
  wire [15:0] _EVAL_19;
  wire [15:0] _EVAL_193;
  wire  _EVAL_43;
  wire  _EVAL_50;
  wire  _EVAL_35;
  wire  _EVAL_133;
  wire [2335:0] _EVAL_121;
  wire [2335:0] _EVAL_101;
  wire  _EVAL_204;
  wire  _EVAL_112;
  wire  _EVAL_234;
  wire  _EVAL_230;
  wire  _EVAL_187;
  wire  _EVAL_197;
  wire  _EVAL_231;
  wire  _EVAL_219;
  wire  _EVAL_209;
  wire  _EVAL_152;
  wire  _EVAL_206;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_201;
  wire  _EVAL_173;
  wire  _EVAL_57;
  wire  _EVAL_134;
  wire  _EVAL_161;
  wire  _EVAL_26;
  wire  _EVAL_114;
  wire  _EVAL_83;
  wire  _EVAL_125;
  wire  _EVAL_109;
  wire  _EVAL_155;
  wire  _EVAL_55;
  wire  _EVAL_124;
  wire  _EVAL_188;
  wire  _EVAL_45;
  wire  _EVAL_132;
  wire  _EVAL_211;
  wire  _EVAL_225;
  wire [3:0] _EVAL_217;
  wire [3:0] _EVAL_157;
  wire [3:0] _EVAL_31;
  wire  _EVAL_68;
  wire  _EVAL_184;
  wire  _EVAL_213;
  wire  _EVAL_169;
  wire  _EVAL_145;
  wire  _EVAL_110;
  wire  _EVAL_224;
  wire  _EVAL_78;
  wire  _EVAL_40;
  wire  _EVAL_53;
  wire [31:0] _EVAL_60;
  wire  _EVAL_165;
  wire  _EVAL_92;
  wire  _EVAL_108;
  wire  _EVAL_100;
  wire  _EVAL_156;
  wire  _EVAL_153;
  wire  _EVAL_181;
  wire  _EVAL_30;
  wire  _EVAL_229;
  wire  _EVAL_222;
  wire  _EVAL_63;
  wire  _EVAL_138;
  wire  _EVAL_195;
  wire  _EVAL_27;
  wire  _EVAL_29;
  wire  _EVAL_127;
  wire  _EVAL_154;
  wire [2335:0] _EVAL_79;
  wire [2335:0] _EVAL_80;
  wire  _EVAL_120;
  wire  _EVAL_128;
  wire  _EVAL_216;
  wire  _EVAL_25;
  wire  _EVAL_167;
  wire  _EVAL_163;
  wire  _EVAL_116;
  wire  _EVAL_47;
  wire  _EVAL_226;
  wire  _EVAL_44;
  wire  _EVAL_75;
  wire  _EVAL_88;
  wire  _EVAL_90;
  wire  _EVAL_39;
  wire  _EVAL_66;
  wire  _EVAL_97;
  wire  _EVAL_81;
  wire  _EVAL_221;
  wire  _EVAL_192;
  wire  _EVAL_42;
  wire  _EVAL_74;
  wire  _EVAL_34;
  wire  _EVAL_207;
  wire  _EVAL_96;
  wire  _EVAL_62;
  wire  _EVAL_52;
  wire  _EVAL_205;
  wire  _EVAL_162;
  wire  _EVAL_94;
  wire  _EVAL_190;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_137 = _EVAL_10 <= 3'h2;
  assign _EVAL_160 = _EVAL_99 >> _EVAL_12;
  assign _EVAL_24 = _EVAL_11 >= 2'h2;
  assign _EVAL_98 = _EVAL_11[0];
  assign _EVAL_105 = 2'h1 << _EVAL_98;
  assign _EVAL_158 = _EVAL_105 | 2'h1;
  assign _EVAL_41 = _EVAL_158[1];
  assign _EVAL_82 = _EVAL_7[1];
  assign _EVAL_151 = _EVAL_41 & _EVAL_82;
  assign _EVAL_91 = _EVAL_24 | _EVAL_151;
  assign _EVAL_166 = _EVAL_158[0];
  assign _EVAL_159 = _EVAL_7[0];
  assign _EVAL_172 = _EVAL_82 & _EVAL_159;
  assign _EVAL_139 = _EVAL_166 & _EVAL_172;
  assign _EVAL_126 = _EVAL_91 | _EVAL_139;
  assign _EVAL_185 = _EVAL_159 == 1'h0;
  assign _EVAL_117 = _EVAL_82 & _EVAL_185;
  assign _EVAL_89 = _EVAL_166 & _EVAL_117;
  assign _EVAL_182 = _EVAL_91 | _EVAL_89;
  assign _EVAL_38 = _EVAL_82 == 1'h0;
  assign _EVAL_141 = _EVAL_41 & _EVAL_38;
  assign _EVAL_175 = _EVAL_24 | _EVAL_141;
  assign _EVAL_23 = _EVAL_38 & _EVAL_159;
  assign _EVAL_102 = _EVAL_166 & _EVAL_23;
  assign _EVAL_130 = _EVAL_175 | _EVAL_102;
  assign _EVAL_236 = _EVAL_38 & _EVAL_185;
  assign _EVAL_147 = _EVAL_166 & _EVAL_236;
  assign _EVAL_208 = _EVAL_175 | _EVAL_147;
  assign _EVAL_93 = {_EVAL_126,_EVAL_182,_EVAL_130,_EVAL_208};
  assign _EVAL_20 = _EVAL_5 == _EVAL_93;
  assign _EVAL_17 = _EVAL_20 | _EVAL_13;
  assign _EVAL_103 = _EVAL_17 == 1'h0;
  assign _EVAL_46 = 5'h3 << _EVAL_11;
  assign _EVAL_210 = _EVAL_46[1:0];
  assign _EVAL_177 = _EVAL_9 == 3'h5;
  assign _EVAL_212 = _EVAL_7 ^ 15'h4000;
  assign _EVAL_194 = _EVAL_215 == 1'h0;
  assign _EVAL_149 = _EVAL_194 == 1'h0;
  assign _EVAL_76 = _EVAL_1 & _EVAL_149;
  assign _EVAL_123 = _EVAL_8 == 3'h2;
  assign _EVAL_198 = _EVAL & _EVAL_123;
  assign _EVAL_178 = _EVAL_71 - 1'h1;
  assign _EVAL_180 = _EVAL_8 == 3'h3;
  assign _EVAL_87 = _EVAL & _EVAL_180;
  assign _EVAL_85 = _EVAL_1 & _EVAL_177;
  assign _EVAL_183 = _EVAL_0 & _EVAL;
  assign _EVAL_196 = _EVAL_6 & _EVAL_1;
  assign _EVAL_135 = _EVAL_131 == 1'h0;
  assign _EVAL_233 = _EVAL_196 & _EVAL_135;
  assign _EVAL_36 = _EVAL_9 == 3'h6;
  assign _EVAL_129 = _EVAL_36 == 1'h0;
  assign _EVAL_232 = _EVAL_233 & _EVAL_129;
  assign _EVAL_86 = 4096'h1 << _EVAL_14;
  assign _EVAL_106 = _EVAL_232 ? _EVAL_86 : 4096'h0;
  assign _EVAL_118 = _EVAL_106[2335:0];
  assign _EVAL_51 = _EVAL_14 <= 12'h91f;
  assign _EVAL_235 = _EVAL_196 & _EVAL_194;
  assign _EVAL_18 = _EVAL_71 == 1'h0;
  assign _EVAL_67 = _EVAL_9 == _EVAL_107;
  assign _EVAL_95 = _EVAL_67 | _EVAL_13;
  assign _EVAL_174 = ~ _EVAL_118;
  assign _EVAL_56 = _EVAL_99 != 2336'h0;
  assign _EVAL_32 = _EVAL_56 == 1'h0;
  assign _EVAL_22 = plusarg_reader_out == 32'h0;
  assign _EVAL_199 = _EVAL_32 | _EVAL_22;
  assign _EVAL_202 = _EVAL_59 < plusarg_reader_out;
  assign _EVAL_146 = _EVAL_199 | _EVAL_202;
  assign _EVAL_33 = _EVAL_146 | _EVAL_13;
  assign _EVAL_148 = _EVAL_33 == 1'h0;
  assign _EVAL_111 = _EVAL_12 <= 12'h91f;
  assign _EVAL_203 = _EVAL_111 | _EVAL_13;
  assign _EVAL_61 = _EVAL_203 == 1'h0;
  assign _EVAL_84 = _EVAL_9 == 3'h2;
  assign _EVAL_28 = _EVAL_1 & _EVAL_84;
  assign _EVAL_64 = _EVAL_136 == 1'h0;
  assign _EVAL_200 = _EVAL_183 & _EVAL_64;
  assign _EVAL_228 = 4096'h1 << _EVAL_12;
  assign _EVAL_220 = _EVAL_200 ? _EVAL_228 : 4096'h0;
  assign _EVAL_21 = _EVAL_220[2335:0];
  assign _EVAL_15 = _EVAL_21 != _EVAL_118;
  assign _EVAL_37 = _EVAL_21 != 2336'h0;
  assign _EVAL_65 = _EVAL_37 == 1'h0;
  assign _EVAL_77 = _EVAL_15 | _EVAL_65;
  assign _EVAL_122 = _EVAL_77 | _EVAL_13;
  assign _EVAL_119 = _EVAL_122 == 1'h0;
  assign _EVAL_150 = _EVAL_24 | _EVAL_13;
  assign _EVAL_54 = _EVAL_150 == 1'h0;
  assign _EVAL_140 = _EVAL_8 == 3'h6;
  assign _EVAL_164 = _EVAL & _EVAL_140;
  assign _EVAL_189 = ~ _EVAL_210;
  assign _EVAL_218 = {{13'd0}, _EVAL_189};
  assign _EVAL_176 = _EVAL_7 & _EVAL_218;
  assign _EVAL_48 = _EVAL_11 <= 2'h2;
  assign _EVAL_214 = {1'b0,$signed(_EVAL_212)};
  assign _EVAL_19 = $signed(_EVAL_214) & $signed(-16'sh1000);
  assign _EVAL_193 = $signed(_EVAL_19);
  assign _EVAL_43 = $signed(_EVAL_193) == $signed(16'sh0);
  assign _EVAL_50 = _EVAL_48 & _EVAL_43;
  assign _EVAL_35 = _EVAL_50 | _EVAL_13;
  assign _EVAL_133 = _EVAL_35 == 1'h0;
  assign _EVAL_121 = _EVAL_21 | _EVAL_99;
  assign _EVAL_101 = _EVAL_121 >> _EVAL_14;
  assign _EVAL_204 = _EVAL_101[0];
  assign _EVAL_112 = _EVAL_204 | _EVAL_13;
  assign _EVAL_234 = _EVAL_112 == 1'h0;
  assign _EVAL_230 = _EVAL_2 >= 2'h2;
  assign _EVAL_187 = _EVAL_51 | _EVAL_13;
  assign _EVAL_197 = _EVAL_187 == 1'h0;
  assign _EVAL_231 = _EVAL_2 == _EVAL_223;
  assign _EVAL_219 = _EVAL_231 | _EVAL_13;
  assign _EVAL_209 = _EVAL_219 == 1'h0;
  assign _EVAL_152 = _EVAL_4 == 1'h0;
  assign _EVAL_206 = _EVAL_8 == 3'h7;
  assign _EVAL_237 = _EVAL & _EVAL_206;
  assign _EVAL_238 = _EVAL_10 == 3'h0;
  assign _EVAL_201 = _EVAL_238 | _EVAL_13;
  assign _EVAL_173 = _EVAL_10 != 3'h0;
  assign _EVAL_57 = _EVAL_173 | _EVAL_13;
  assign _EVAL_134 = _EVAL_57 == 1'h0;
  assign _EVAL_161 = _EVAL_8 == 3'h4;
  assign _EVAL_26 = _EVAL & _EVAL_161;
  assign _EVAL_114 = _EVAL_131 - 1'h1;
  assign _EVAL_83 = _EVAL_10 <= 3'h3;
  assign _EVAL_125 = _EVAL_83 | _EVAL_13;
  assign _EVAL_109 = _EVAL_125 == 1'h0;
  assign _EVAL_155 = _EVAL_8 == 3'h0;
  assign _EVAL_55 = _EVAL_1 & _EVAL_36;
  assign _EVAL_124 = _EVAL_9 <= 3'h6;
  assign _EVAL_188 = _EVAL_124 | _EVAL_13;
  assign _EVAL_45 = _EVAL_14 == _EVAL_227;
  assign _EVAL_132 = _EVAL_13 == 1'h0;
  assign _EVAL_211 = _EVAL_8 == 3'h5;
  assign _EVAL_225 = _EVAL & _EVAL_211;
  assign _EVAL_217 = ~ _EVAL_93;
  assign _EVAL_157 = _EVAL_5 & _EVAL_217;
  assign _EVAL_31 = ~ _EVAL_5;
  assign _EVAL_68 = _EVAL_31 == 4'h0;
  assign _EVAL_184 = _EVAL_68 | _EVAL_13;
  assign _EVAL_213 = _EVAL_184 == 1'h0;
  assign _EVAL_169 = _EVAL_176 == 15'h0;
  assign _EVAL_145 = _EVAL_169 | _EVAL_13;
  assign _EVAL_110 = _EVAL_136 - 1'h1;
  assign _EVAL_224 = _EVAL_10 <= 3'h4;
  assign _EVAL_78 = _EVAL_45 | _EVAL_13;
  assign _EVAL_40 = _EVAL_78 == 1'h0;
  assign _EVAL_53 = _EVAL_183 | _EVAL_196;
  assign _EVAL_60 = _EVAL_59 + 32'h1;
  assign _EVAL_165 = _EVAL_152 | _EVAL_13;
  assign _EVAL_92 = _EVAL_165 == 1'h0;
  assign _EVAL_108 = _EVAL_137 | _EVAL_13;
  assign _EVAL_100 = _EVAL_108 == 1'h0;
  assign _EVAL_156 = _EVAL_9 == 3'h4;
  assign _EVAL_153 = _EVAL_1 & _EVAL_156;
  assign _EVAL_181 = _EVAL_160[0];
  assign _EVAL_30 = _EVAL_181 == 1'h0;
  assign _EVAL_229 = _EVAL_30 | _EVAL_13;
  assign _EVAL_222 = _EVAL_229 == 1'h0;
  assign _EVAL_63 = _EVAL_10 == _EVAL_115;
  assign _EVAL_138 = _EVAL_63 | _EVAL_13;
  assign _EVAL_195 = _EVAL_230 | _EVAL_13;
  assign _EVAL_27 = _EVAL_224 | _EVAL_13;
  assign _EVAL_29 = _EVAL_27 == 1'h0;
  assign _EVAL_127 = _EVAL_215 - 1'h1;
  assign _EVAL_154 = _EVAL_12 == _EVAL_72;
  assign _EVAL_79 = _EVAL_99 | _EVAL_21;
  assign _EVAL_80 = _EVAL_79 & _EVAL_174;
  assign _EVAL_120 = _EVAL_154 | _EVAL_13;
  assign _EVAL_128 = _EVAL_120 == 1'h0;
  assign _EVAL_216 = _EVAL_8 == 3'h1;
  assign _EVAL_25 = _EVAL & _EVAL_216;
  assign _EVAL_167 = _EVAL_18 == 1'h0;
  assign _EVAL_163 = _EVAL & _EVAL_167;
  assign _EVAL_116 = _EVAL_8 == _EVAL_58;
  assign _EVAL_47 = _EVAL_145 == 1'h0;
  assign _EVAL_226 = _EVAL_116 | _EVAL_13;
  assign _EVAL_44 = _EVAL_226 == 1'h0;
  assign _EVAL_75 = _EVAL_7 == _EVAL_104;
  assign _EVAL_88 = _EVAL_188 == 1'h0;
  assign _EVAL_90 = _EVAL_75 | _EVAL_13;
  assign _EVAL_39 = _EVAL_195 == 1'h0;
  assign _EVAL_66 = _EVAL_9 == 3'h0;
  assign _EVAL_97 = _EVAL_11 == _EVAL_171;
  assign _EVAL_81 = _EVAL_97 | _EVAL_13;
  assign _EVAL_221 = _EVAL_90 == 1'h0;
  assign _EVAL_192 = _EVAL_9 == 3'h1;
  assign _EVAL_42 = _EVAL_157 == 4'h0;
  assign _EVAL_74 = _EVAL_81 == 1'h0;
  assign _EVAL_34 = _EVAL_138 == 1'h0;
  assign _EVAL_207 = _EVAL_1 & _EVAL_192;
  assign _EVAL_96 = _EVAL_183 & _EVAL_18;
  assign _EVAL_62 = _EVAL_42 | _EVAL_13;
  assign _EVAL_52 = _EVAL_62 == 1'h0;
  assign _EVAL_205 = _EVAL_1 & _EVAL_66;
  assign _EVAL_162 = _EVAL_201 == 1'h0;
  assign _EVAL_94 = _EVAL_95 == 1'h0;
  assign _EVAL_190 = _EVAL & _EVAL_155;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_58 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_59 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_71 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_72 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {73{`RANDOM}};
  _EVAL_99 = _RAND_4[2335:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_104 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_107 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_115 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_131 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_136 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_171 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_215 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_223 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_227 = _RAND_13[11:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_96) begin
      _EVAL_58 <= _EVAL_8;
    end
    if (_EVAL_13) begin
      _EVAL_59 <= 32'h0;
    end else begin
      if (_EVAL_53) begin
        _EVAL_59 <= 32'h0;
      end else begin
        _EVAL_59 <= _EVAL_60;
      end
    end
    if (_EVAL_13) begin
      _EVAL_71 <= 1'h0;
    end else begin
      if (_EVAL_183) begin
        if (_EVAL_18) begin
          _EVAL_71 <= 1'h0;
        end else begin
          _EVAL_71 <= _EVAL_178;
        end
      end
    end
    if (_EVAL_96) begin
      _EVAL_72 <= _EVAL_12;
    end
    if (_EVAL_13) begin
      _EVAL_99 <= 2336'h0;
    end else begin
      _EVAL_99 <= _EVAL_80;
    end
    if (_EVAL_96) begin
      _EVAL_104 <= _EVAL_7;
    end
    if (_EVAL_235) begin
      _EVAL_107 <= _EVAL_9;
    end
    if (_EVAL_96) begin
      _EVAL_115 <= _EVAL_10;
    end
    if (_EVAL_13) begin
      _EVAL_131 <= 1'h0;
    end else begin
      if (_EVAL_196) begin
        if (_EVAL_135) begin
          _EVAL_131 <= 1'h0;
        end else begin
          _EVAL_131 <= _EVAL_114;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_136 <= 1'h0;
    end else begin
      if (_EVAL_183) begin
        if (_EVAL_64) begin
          _EVAL_136 <= 1'h0;
        end else begin
          _EVAL_136 <= _EVAL_110;
        end
      end
    end
    if (_EVAL_96) begin
      _EVAL_171 <= _EVAL_11;
    end
    if (_EVAL_13) begin
      _EVAL_215 <= 1'h0;
    end else begin
      if (_EVAL_196) begin
        if (_EVAL_194) begin
          _EVAL_215 <= 1'h0;
        end else begin
          _EVAL_215 <= _EVAL_127;
        end
      end
    end
    if (_EVAL_235) begin
      _EVAL_223 <= _EVAL_2;
    end
    if (_EVAL_235) begin
      _EVAL_227 <= _EVAL_14;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf9925e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19602c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae8b84db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea95ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b03b1ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9817991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19018510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb96d4bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a862eb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5f9d6c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(200415a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61b1fc54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79d91f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4196f9ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2eb311c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca76bcab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bddf239)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb473fef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33873282)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f0684c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf1d82c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31908dd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e35df6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82cf291b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5e59717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aefe180f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7de7288c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d828a416)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e35e5e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8edc821)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f2d746c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccd2bcb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f3b5520)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b0d2de4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf66ce67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b13b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c719695b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb1c749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbc6fcaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ad58fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30d40d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2c3c631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25cce22e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a0f91ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de60b4b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e679fbfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6786ba22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7935cf94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f215a32e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb0c3065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6bc7fe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d37cc6e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98c955fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fc1c20e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffd2a09d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(147f55b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1840a173)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df9b0213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10eecbaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6db5bf11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e37cbfe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3849315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf58451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b62bc31e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6070b9c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1809643b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee9ed123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5649fbd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46bd5adc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d71f4482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60540a4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3287683)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
