//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_259_assert(
  input        _EVAL_1,
  input        _EVAL_18,
  input        _EVAL_42,
  input  [3:0] _EVAL_77,
  input        _EVAL_332,
  input        _EVAL_357,
  input        _EVAL_559,
  input        _EVAL_613,
  input        _EVAL_655,
  input        _EVAL_1122,
  input        _EVAL_1271,
  input        _EVAL_1278,
  input        _EVAL_1350,
  input        _EVAL_1422,
  input        _EVAL_1442,
  input        _EVAL_1486,
  input        _EVAL_1835,
  input  [3:0] _EVAL_1653,
  input        _EVAL_209,
  input        _EVAL_153,
  input        _EVAL_1564,
  input        _EVAL_1542,
  input        _EVAL_838,
  input        _EVAL_699,
  input        _EVAL_583,
  input        _EVAL_1438,
  input        _EVAL_1757,
  input        _EVAL_1016,
  input        _EVAL_1221,
  input        _EVAL_1718,
  input        _EVAL_1524,
  input        _EVAL_276,
  input        _EVAL_264,
  input        _EVAL_176,
  input        _EVAL_406,
  input        _EVAL_497,
  input        _EVAL_1315,
  input        _EVAL_1624,
  input        _EVAL_807,
  input        _EVAL_1519,
  input        _EVAL_1139,
  input        _EVAL_1786,
  input        _EVAL_1403,
  input        _EVAL_1477,
  input        _EVAL_975,
  input        _EVAL_729,
  input        _EVAL_635,
  input        _EVAL_665,
  input        _EVAL_325,
  input        _EVAL_1668,
  input        dcache_clock_gate_out
);
  wire  _EVAL_1802;
  wire  _EVAL_1035;
  wire  _EVAL_372;
  wire  _EVAL_181;
  wire  _EVAL_408;
  wire  _EVAL_221;
  wire [3:0] _EVAL_1558;
  wire  _EVAL_1690;
  wire  _EVAL_1677;
  wire  _EVAL_1501;
  wire  _EVAL_933;
  wire  _EVAL_543;
  wire  _EVAL_1057;
  wire  _EVAL_472;
  wire  _EVAL_215;
  wire  _EVAL_538;
  wire  _EVAL_1482;
  wire  _EVAL_474;
  wire  _EVAL_1796;
  wire [3:0] _EVAL_1801;
  wire  _EVAL_1490;
  wire  _EVAL_1047;
  wire  _EVAL_503;
  wire  _EVAL_519;
  wire  _EVAL_1590;
  wire  _EVAL_1285;
  wire  _EVAL_989;
  wire  _EVAL_1870;
  wire  _EVAL_1101;
  wire  _EVAL_943;
  wire  _EVAL_1051;
  wire  _EVAL_1470;
  wire  _EVAL_1544;
  wire  _EVAL_1513;
  wire  _EVAL_1266;
  wire  _EVAL_582;
  wire  _EVAL_766;
  wire  _EVAL_953;
  wire  _EVAL_1079;
  wire  _EVAL_1816;
  wire  _EVAL_1310;
  wire  _EVAL_1598;
  wire  _EVAL_1375;
  wire  _EVAL_1634;
  wire  _EVAL_1203;
  wire  _EVAL_573;
  wire  _EVAL_1286;
  wire  _EVAL_1492;
  wire  _EVAL_152;
  wire  _EVAL_938;
  wire  _EVAL_480;
  wire  _EVAL_1356;
  wire  _EVAL_1875;
  wire  _EVAL_1171;
  wire  _EVAL_1324;
  wire  _EVAL_1852;
  wire  _EVAL_1767;
  wire  _EVAL_1234;
  wire  _EVAL_1755;
  wire  _EVAL_1472;
  wire  _EVAL_1804;
  wire  _EVAL_289;
  wire  _EVAL_786;
  wire  _EVAL_1275;
  wire  _EVAL_1013;
  wire  _EVAL_645;
  wire  _EVAL_853;
  wire  _EVAL_1678;
  wire  _EVAL_1167;
  wire  _EVAL_1365;
  wire  _EVAL_485;
  wire  _EVAL_915;
  wire  _EVAL_703;
  wire  _EVAL_488;
  wire  _EVAL_514;
  wire  _EVAL_1731;
  wire  _EVAL_1147;
  wire  _EVAL_1238;
  wire  _EVAL_265;
  wire  _EVAL_1742;
  wire  _EVAL_1090;
  wire  _EVAL_1044;
  wire  _EVAL_1033;
  assign _EVAL_1802 = _EVAL_209 == _EVAL_153;
  assign _EVAL_1035 = _EVAL_1486 | _EVAL_1802;
  assign _EVAL_372 = _EVAL_1035 | _EVAL_18;
  assign _EVAL_181 = _EVAL_372 == 1'h0;
  assign _EVAL_408 = _EVAL_357 | _EVAL_18;
  assign _EVAL_221 = _EVAL_408 == 1'h0;
  assign _EVAL_1558 = ~ _EVAL_77;
  assign _EVAL_1690 = 1'h0;
  assign _EVAL_1677 = _EVAL_1690;
  assign _EVAL_1501 = _EVAL_1422 & _EVAL_1677;
  assign _EVAL_933 = _EVAL_406 & _EVAL_1501;
  assign _EVAL_543 = _EVAL_1564 == 1'h0;
  assign _EVAL_1057 = _EVAL_1718 & _EVAL_543;
  assign _EVAL_472 = _EVAL_1057 & _EVAL_264;
  assign _EVAL_215 = _EVAL_472 & _EVAL_807;
  assign _EVAL_538 = _EVAL_1122 | _EVAL_18;
  assign _EVAL_1482 = _EVAL_538 == 1'h0;
  assign _EVAL_474 = _EVAL_1315 & _EVAL_1542;
  assign _EVAL_1796 = _EVAL_474 == 1'h0;
  assign _EVAL_1801 = _EVAL_1653 | _EVAL_1558;
  assign _EVAL_1490 = _EVAL_1801 == 4'hf;
  assign _EVAL_1047 = _EVAL_1796 | _EVAL_1490;
  assign _EVAL_503 = _EVAL_1519 | _EVAL_1278;
  assign _EVAL_519 = _EVAL_503 | _EVAL_42;
  assign _EVAL_1590 = _EVAL_153 & _EVAL_583;
  assign _EVAL_1285 = _EVAL_1690 == 1'h0;
  assign _EVAL_989 = _EVAL_1422 & _EVAL_1285;
  assign _EVAL_1870 = _EVAL_497 & _EVAL_989;
  assign _EVAL_1101 = _EVAL_472 & _EVAL_729;
  assign _EVAL_943 = _EVAL_1757 & _EVAL_276;
  assign _EVAL_1051 = _EVAL_1786 & _EVAL_1677;
  assign _EVAL_1470 = _EVAL_406 & _EVAL_1051;
  assign _EVAL_1544 = _EVAL_1403 == 1'h0;
  assign _EVAL_1513 = _EVAL_1718 & _EVAL_1438;
  assign _EVAL_1266 = _EVAL_1513 & _EVAL_1564;
  assign _EVAL_582 = _EVAL_1786 & _EVAL_1285;
  assign _EVAL_766 = _EVAL_406 & _EVAL_582;
  assign _EVAL_953 = _EVAL_1271 | _EVAL_18;
  assign _EVAL_1079 = _EVAL_497 & _EVAL_1051;
  assign _EVAL_1816 = _EVAL_613 | _EVAL_18;
  assign _EVAL_1310 = _EVAL_1816 == 1'h0;
  assign _EVAL_1598 = _EVAL_519 | _EVAL_18;
  assign _EVAL_1375 = _EVAL_1598 == 1'h0;
  assign _EVAL_1634 = _EVAL_1 & _EVAL_1564;
  assign _EVAL_1203 = _EVAL_264 == 1'h0;
  assign _EVAL_573 = _EVAL_1047 | _EVAL_18;
  assign _EVAL_1286 = _EVAL_1835 | _EVAL_18;
  assign _EVAL_1492 = _EVAL_1286 == 1'h0;
  assign _EVAL_152 = _EVAL_1524 & _EVAL_1544;
  assign _EVAL_938 = _EVAL_472 & _EVAL_176;
  assign _EVAL_480 = _EVAL_559 | _EVAL_18;
  assign _EVAL_1356 = _EVAL_943 == _EVAL_1266;
  assign _EVAL_1875 = _EVAL_665 | _EVAL_18;
  assign _EVAL_1171 = _EVAL_325 == 1'h0;
  assign _EVAL_1324 = _EVAL_573 == 1'h0;
  assign _EVAL_1852 = _EVAL_406 & _EVAL_989;
  assign _EVAL_1767 = _EVAL_1356 | _EVAL_18;
  assign _EVAL_1234 = _EVAL_1016 == 1'h0;
  assign _EVAL_1755 = _EVAL_1171 | _EVAL_699;
  assign _EVAL_1472 = _EVAL_1767 == 1'h0;
  assign _EVAL_1804 = _EVAL_18 == 1'h0;
  assign _EVAL_289 = _EVAL_1350 | _EVAL_18;
  assign _EVAL_786 = _EVAL_472 & _EVAL_635;
  assign _EVAL_1275 = _EVAL_1755 | _EVAL_18;
  assign _EVAL_1013 = _EVAL_1275 == 1'h0;
  assign _EVAL_645 = _EVAL_472 & _EVAL_975;
  assign _EVAL_853 = _EVAL_497 & _EVAL_1501;
  assign _EVAL_1678 = _EVAL_655 | _EVAL_18;
  assign _EVAL_1167 = _EVAL_1678 == 1'h0;
  assign _EVAL_1365 = _EVAL_480 == 1'h0;
  assign _EVAL_485 = _EVAL_332 | _EVAL_18;
  assign _EVAL_915 = _EVAL_953 == 1'h0;
  assign _EVAL_703 = _EVAL_1718 & _EVAL_1564;
  assign _EVAL_488 = _EVAL_472 & _EVAL_1668;
  assign _EVAL_514 = _EVAL_1 & _EVAL_543;
  assign _EVAL_1731 = _EVAL_1057 & _EVAL_1203;
  assign _EVAL_1147 = _EVAL_1221 & _EVAL_1234;
  assign _EVAL_1238 = _EVAL_472 & _EVAL_1624;
  assign _EVAL_265 = _EVAL_289 == 1'h0;
  assign _EVAL_1742 = _EVAL_1731 & _EVAL_1477;
  assign _EVAL_1090 = _EVAL_485 == 1'h0;
  assign _EVAL_1044 = _EVAL_497 & _EVAL_582;
  assign _EVAL_1033 = _EVAL_1875 == 1'h0;
  always @(posedge dcache_clock_gate_out) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_838 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a0f52cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1238 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1013) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9493fc4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1147 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a52624)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1101 & _EVAL_915) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fac9748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1870 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ab001bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_1482) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1472) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43d0e9c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d18f1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1139 & _EVAL_1375) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(386131ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_1167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_1310) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_1033) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80d137d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_703 & _EVAL_1492) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ead9bfb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1742 & _EVAL_1365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d01cc4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1139 & _EVAL_1375) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_1482) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_514 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b56b10ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfbcb13c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1590 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4740af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1238 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1472) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1079 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3045bc85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_1310) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1101 & _EVAL_915) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_1167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ae93070)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_1033) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1013) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1852 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb3637e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1634 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d8cbf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1742 & _EVAL_1365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_1090) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1013) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d43039a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_703 & _EVAL_1492) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1044 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb8c5a23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1013) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d43039a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1470 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f10025eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_1090) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0dcc8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_933 & _EVAL_1804) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43afd797)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
