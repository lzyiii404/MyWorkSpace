//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_288(
  input  [32:0] _EVAL,
  output        _EVAL_0,
  output [23:0] _EVAL_1,
  output [25:0] _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input  [32:0] _EVAL_6,
  output        _EVAL_7,
  output [4:0]  _EVAL_8,
  output        _EVAL_9,
  output [23:0] _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output [47:0] _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  input  [32:0] _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  output [9:0]  _EVAL_20
);
  wire [22:0] _EVAL_143;
  wire  _EVAL_47;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_48;
  wire  _EVAL_110;
  wire [8:0] _EVAL_98;
  wire [2:0] _EVAL_138;
  wire  _EVAL_63;
  wire  _EVAL_94;
  wire [22:0] _EVAL_67;
  wire [24:0] _EVAL_37;
  wire [24:0] _EVAL_112;
  wire [24:0] _EVAL_117;
  wire [52:0] _EVAL_72;
  wire [77:0] _EVAL_34;
  wire [8:0] _EVAL_36;
  wire  _EVAL_127;
  wire  _EVAL_114;
  wire [2:0] _EVAL_26;
  wire  _EVAL_77;
  wire  _EVAL_91;
  wire [8:0] _EVAL_57;
  wire [2:0] _EVAL_134;
  wire  _EVAL_59;
  wire  _EVAL_109;
  wire [9:0] _EVAL_44;
  wire [9:0] _EVAL_132;
  wire [10:0] _EVAL_88;
  wire [10:0] _EVAL_41;
  wire [10:0] _EVAL_76;
  wire [9:0] _EVAL_71;
  wire [10:0] _EVAL_65;
  wire [10:0] _EVAL_29;
  wire [10:0] _EVAL_70;
  wire  _EVAL_60;
  wire  _EVAL_136;
  wire [9:0] _EVAL_118;
  wire  _EVAL_139;
  wire [6:0] _EVAL_113;
  wire [6:0] _EVAL_100;
  wire [6:0] _EVAL_142;
  wire [4:0] _EVAL_64;
  wire [32:0] _EVAL_101;
  wire  _EVAL_43;
  wire  _EVAL_49;
  wire  _EVAL_75;
  wire [10:0] _EVAL_22;
  wire [10:0] _EVAL_92;
  wire [10:0] _EVAL_93;
  wire [77:0] _EVAL_58;
  wire [77:0] _EVAL_21;
  wire [74:0] _EVAL_69;
  wire [74:0] _EVAL_123;
  wire [2:0] _EVAL_27;
  wire  _EVAL_84;
  wire [26:0] _EVAL_53;
  wire [2:0] _EVAL_31;
  wire  _EVAL_56;
  wire [3:0] _EVAL_55;
  wire  _EVAL_39;
  wire [3:0] _EVAL_80;
  wire  _EVAL_50;
  wire [3:0] _EVAL_129;
  wire  _EVAL_68;
  wire [3:0] _EVAL_120;
  wire  _EVAL_125;
  wire [3:0] _EVAL_73;
  wire  _EVAL_51;
  wire [3:0] _EVAL_131;
  wire  _EVAL_96;
  wire [6:0] _EVAL_89;
  wire [5:0] _EVAL_52;
  wire [3:0] _EVAL_102;
  wire [1:0] _EVAL_116;
  wire  _EVAL_133;
  wire  _EVAL_126;
  wire [1:0] _EVAL_104;
  wire  _EVAL_90;
  wire  _EVAL_86;
  wire [1:0] _EVAL_25;
  wire  _EVAL_82;
  wire  _EVAL_74;
  wire [5:0] _EVAL_23;
  wire [6:0] _EVAL_66;
  wire [6:0] _EVAL_128;
  wire  _EVAL_137;
  wire  _EVAL_54;
  wire  _EVAL_124;
  wire  _EVAL_107;
  wire  _EVAL_106;
  wire  _EVAL_78;
  wire [75:0] _EVAL_85;
  wire  _EVAL_135;
  wire  _EVAL_122;
  wire [1:0] _EVAL_81;
  wire [1:0] _EVAL_115;
  wire  _EVAL_24;
  wire  _EVAL_140;
  wire [22:0] _EVAL_97;
  wire [24:0] _EVAL_42;
  wire  _EVAL_40;
  wire  _EVAL_105;
  wire  _EVAL_103;
  wire  _EVAL_61;
  wire [24:0] _EVAL_111;
  wire  _EVAL_95;
  wire  _EVAL_46;
  wire [1:0] _EVAL_130;
  wire  _EVAL_83;
  wire  _EVAL_87;
  wire  _EVAL_30;
  wire  _EVAL_108;
  wire  _EVAL_121;
  wire  _EVAL_119;
  wire  _EVAL_38;
  wire  _EVAL_35;
  wire  _EVAL_28;
  wire [9:0] _EVAL_62;
  wire  _EVAL_141;
  wire  _EVAL_45;
  assign _EVAL_143 = _EVAL[22:0];
  assign _EVAL_47 = _EVAL[32];
  assign _EVAL_32 = _EVAL_17[32];
  assign _EVAL_33 = _EVAL_47 ^ _EVAL_32;
  assign _EVAL_48 = _EVAL_6[32];
  assign _EVAL_110 = _EVAL_33 ^ _EVAL_48;
  assign _EVAL_98 = _EVAL_6[31:23];
  assign _EVAL_138 = _EVAL_98[8:6];
  assign _EVAL_63 = _EVAL_138 == 3'h0;
  assign _EVAL_94 = _EVAL_63 == 1'h0;
  assign _EVAL_67 = _EVAL_6[22:0];
  assign _EVAL_37 = {1'h0,_EVAL_94,_EVAL_67};
  assign _EVAL_112 = ~ _EVAL_37;
  assign _EVAL_117 = _EVAL_110 ? _EVAL_112 : _EVAL_37;
  assign _EVAL_72 = _EVAL_110 ? 53'h1fffffffffffff : 53'h0;
  assign _EVAL_34 = {_EVAL_117,_EVAL_72};
  assign _EVAL_36 = _EVAL_17[31:23];
  assign _EVAL_127 = _EVAL_36[6];
  assign _EVAL_114 = _EVAL_127 == 1'h0;
  assign _EVAL_26 = _EVAL_36[8:6];
  assign _EVAL_77 = _EVAL_26 == 3'h0;
  assign _EVAL_91 = _EVAL_77 == 1'h0;
  assign _EVAL_57 = _EVAL[31:23];
  assign _EVAL_134 = _EVAL_57[8:6];
  assign _EVAL_59 = _EVAL_134 == 3'h0;
  assign _EVAL_109 = _EVAL_59 | _EVAL_77;
  assign _EVAL_44 = {1'b0,$signed(_EVAL_57)};
  assign _EVAL_132 = {1'b0,$signed(_EVAL_36)};
  assign _EVAL_88 = $signed(_EVAL_44) + $signed(_EVAL_132);
  assign _EVAL_41 = $signed(_EVAL_88) + $signed(-11'she5);
  assign _EVAL_76 = $signed(_EVAL_41);
  assign _EVAL_71 = {1'b0,$signed(_EVAL_98)};
  assign _EVAL_65 = {{1{_EVAL_71[9]}},_EVAL_71};
  assign _EVAL_29 = $signed(_EVAL_76) - $signed(_EVAL_65);
  assign _EVAL_70 = $signed(_EVAL_29);
  assign _EVAL_60 = $signed(_EVAL_70) < $signed(11'sh0);
  assign _EVAL_136 = _EVAL_109 | _EVAL_60;
  assign _EVAL_118 = _EVAL_70[9:0];
  assign _EVAL_139 = _EVAL_118 < 10'h4a;
  assign _EVAL_113 = _EVAL_118[6:0];
  assign _EVAL_100 = _EVAL_139 ? _EVAL_113 : 7'h4a;
  assign _EVAL_142 = _EVAL_136 ? 7'h0 : _EVAL_100;
  assign _EVAL_64 = _EVAL_142[6:2];
  assign _EVAL_101 = $signed(-33'sh100000000) >>> _EVAL_64;
  assign _EVAL_43 = _EVAL_118 <= 10'h18;
  assign _EVAL_49 = _EVAL_136 | _EVAL_43;
  assign _EVAL_75 = _EVAL_94 & _EVAL_49;
  assign _EVAL_22 = $signed(_EVAL_76) - $signed(11'sh18);
  assign _EVAL_92 = $signed(_EVAL_22);
  assign _EVAL_93 = _EVAL_75 ? $signed({{1{_EVAL_71[9]}},_EVAL_71}) : $signed(_EVAL_92);
  assign _EVAL_58 = $signed(_EVAL_34);
  assign _EVAL_21 = $signed(_EVAL_58) >>> _EVAL_142;
  assign _EVAL_69 = _EVAL_21[77:3];
  assign _EVAL_123 = $unsigned(_EVAL_69);
  assign _EVAL_27 = _EVAL_21[2:0];
  assign _EVAL_84 = _EVAL_27 == 3'h7;
  assign _EVAL_53 = {_EVAL_37, 2'h0};
  assign _EVAL_31 = _EVAL_53[26:24];
  assign _EVAL_56 = _EVAL_31 != 3'h0;
  assign _EVAL_55 = _EVAL_53[23:20];
  assign _EVAL_39 = _EVAL_55 != 4'h0;
  assign _EVAL_80 = _EVAL_53[19:16];
  assign _EVAL_50 = _EVAL_80 != 4'h0;
  assign _EVAL_129 = _EVAL_53[15:12];
  assign _EVAL_68 = _EVAL_129 != 4'h0;
  assign _EVAL_120 = _EVAL_53[11:8];
  assign _EVAL_125 = _EVAL_120 != 4'h0;
  assign _EVAL_73 = _EVAL_53[7:4];
  assign _EVAL_51 = _EVAL_73 != 4'h0;
  assign _EVAL_131 = _EVAL_53[3:0];
  assign _EVAL_96 = _EVAL_131 != 4'h0;
  assign _EVAL_89 = {_EVAL_56,_EVAL_39,_EVAL_50,_EVAL_68,_EVAL_125,_EVAL_51,_EVAL_96};
  assign _EVAL_52 = _EVAL_101[19:14];
  assign _EVAL_102 = _EVAL_52[3:0];
  assign _EVAL_116 = _EVAL_102[1:0];
  assign _EVAL_133 = _EVAL_116[0];
  assign _EVAL_126 = _EVAL_116[1];
  assign _EVAL_104 = _EVAL_102[3:2];
  assign _EVAL_90 = _EVAL_104[0];
  assign _EVAL_86 = _EVAL_104[1];
  assign _EVAL_25 = _EVAL_52[5:4];
  assign _EVAL_82 = _EVAL_25[0];
  assign _EVAL_74 = _EVAL_25[1];
  assign _EVAL_23 = {_EVAL_133,_EVAL_126,_EVAL_90,_EVAL_86,_EVAL_82,_EVAL_74};
  assign _EVAL_66 = {{1'd0}, _EVAL_23};
  assign _EVAL_128 = _EVAL_89 & _EVAL_66;
  assign _EVAL_137 = _EVAL_128 != 7'h0;
  assign _EVAL_54 = _EVAL_137 == 1'h0;
  assign _EVAL_124 = _EVAL_84 & _EVAL_54;
  assign _EVAL_107 = _EVAL_27 != 3'h0;
  assign _EVAL_106 = _EVAL_107 | _EVAL_137;
  assign _EVAL_78 = _EVAL_110 ? _EVAL_124 : _EVAL_106;
  assign _EVAL_85 = {_EVAL_123,_EVAL_78};
  assign _EVAL_135 = _EVAL_37[22];
  assign _EVAL_122 = _EVAL_135 == 1'h0;
  assign _EVAL_81 = _EVAL_98[8:7];
  assign _EVAL_115 = _EVAL_36[8:7];
  assign _EVAL_24 = _EVAL_115 == 2'h3;
  assign _EVAL_140 = _EVAL_24 & _EVAL_127;
  assign _EVAL_97 = _EVAL_17[22:0];
  assign _EVAL_42 = {1'h0,_EVAL_91,_EVAL_97};
  assign _EVAL_40 = _EVAL_42[22];
  assign _EVAL_105 = _EVAL_40 == 1'h0;
  assign _EVAL_103 = _EVAL_140 & _EVAL_105;
  assign _EVAL_61 = _EVAL_59 == 1'h0;
  assign _EVAL_111 = {1'h0,_EVAL_61,_EVAL_143};
  assign _EVAL_95 = _EVAL_111[22];
  assign _EVAL_46 = _EVAL_95 == 1'h0;
  assign _EVAL_130 = _EVAL_57[8:7];
  assign _EVAL_83 = _EVAL_130 == 2'h3;
  assign _EVAL_87 = _EVAL_57[6];
  assign _EVAL_30 = _EVAL_83 & _EVAL_87;
  assign _EVAL_108 = _EVAL_30 & _EVAL_46;
  assign _EVAL_121 = _EVAL_98[6];
  assign _EVAL_119 = _EVAL_121 == 1'h0;
  assign _EVAL_38 = _EVAL_87 == 1'h0;
  assign _EVAL_35 = _EVAL_81 == 2'h3;
  assign _EVAL_28 = _EVAL_35 & _EVAL_121;
  assign _EVAL_62 = _EVAL_93[9:0];
  assign _EVAL_141 = _EVAL_108 | _EVAL_103;
  assign _EVAL_45 = _EVAL_28 & _EVAL_122;
  assign _EVAL_18 = _EVAL_35 & _EVAL_121;
  assign _EVAL_19 = _EVAL_141 | _EVAL_45;
  assign _EVAL_8 = _EVAL_142[4:0];
  assign _EVAL_13 = _EVAL_85[48:1];
  assign _EVAL_20 = $signed(_EVAL_62);
  assign _EVAL_11 = _EVAL_33 ^ _EVAL_48;
  assign _EVAL_12 = _EVAL_26 == 3'h0;
  assign _EVAL_0 = _EVAL_85[0];
  assign _EVAL_7 = _EVAL_24 & _EVAL_114;
  assign _EVAL_5 = _EVAL_83 & _EVAL_38;
  assign _EVAL_3 = _EVAL_94 & _EVAL_49;
  assign _EVAL_10 = _EVAL_42[23:0];
  assign _EVAL_4 = _EVAL_30 | _EVAL_140;
  assign _EVAL_16 = _EVAL_47 ^ _EVAL_32;
  assign _EVAL_14 = _EVAL_134 == 3'h0;
  assign _EVAL_2 = _EVAL_85[74:49];
  assign _EVAL_9 = _EVAL_138 == 3'h0;
  assign _EVAL_1 = _EVAL_111[23:0];
  assign _EVAL_15 = _EVAL_35 & _EVAL_119;
endmodule
