//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive_CoreIPSubsystem(
  input          clock,
  input          reset,
  input          debug_psd_test_mode,
  input          debug_psd_test_mode_reset,
  input          debug_systemjtag_jtag_TCK,
  input          debug_systemjtag_jtag_TMS,
  input          debug_systemjtag_jtag_TDI,
  output         debug_systemjtag_jtag_TDO_data,
  output         debug_systemjtag_jtag_TDO_driven,
  input          debug_systemjtag_reset,
  input  [10:0]  debug_systemjtag_mfr_id,
  output         debug_ndreset,
  output         debug_dmactive,
  input          core_clock_0,
  input  [31:0]  reset_vector_0,
  input          rtc_toggle,
  input  [126:0] global_interrupts,
  input          mem_port_axi4_0_aw_ready,
  output         mem_port_axi4_0_aw_valid,
  output [3:0]   mem_port_axi4_0_aw_bits_id,
  output [31:0]  mem_port_axi4_0_aw_bits_addr,
  output [7:0]   mem_port_axi4_0_aw_bits_len,
  output [2:0]   mem_port_axi4_0_aw_bits_size,
  output [1:0]   mem_port_axi4_0_aw_bits_burst,
  output         mem_port_axi4_0_aw_bits_lock,
  output [3:0]   mem_port_axi4_0_aw_bits_cache,
  output [2:0]   mem_port_axi4_0_aw_bits_prot,
  output [3:0]   mem_port_axi4_0_aw_bits_qos,
  input          mem_port_axi4_0_w_ready,
  output         mem_port_axi4_0_w_valid,
  output [63:0]  mem_port_axi4_0_w_bits_data,
  output [7:0]   mem_port_axi4_0_w_bits_strb,
  output         mem_port_axi4_0_w_bits_last,
  output         mem_port_axi4_0_w_bits_corrupt,
  output         mem_port_axi4_0_b_ready,
  input          mem_port_axi4_0_b_valid,
  input  [3:0]   mem_port_axi4_0_b_bits_id,
  input  [1:0]   mem_port_axi4_0_b_bits_resp,
  input          mem_port_axi4_0_ar_ready,
  output         mem_port_axi4_0_ar_valid,
  output [3:0]   mem_port_axi4_0_ar_bits_id,
  output [31:0]  mem_port_axi4_0_ar_bits_addr,
  output [7:0]   mem_port_axi4_0_ar_bits_len,
  output [2:0]   mem_port_axi4_0_ar_bits_size,
  output [1:0]   mem_port_axi4_0_ar_bits_burst,
  output         mem_port_axi4_0_ar_bits_lock,
  output [3:0]   mem_port_axi4_0_ar_bits_cache,
  output [2:0]   mem_port_axi4_0_ar_bits_prot,
  output [3:0]   mem_port_axi4_0_ar_bits_qos,
  output         mem_port_axi4_0_r_ready,
  input          mem_port_axi4_0_r_valid,
  input  [3:0]   mem_port_axi4_0_r_bits_id,
  input  [63:0]  mem_port_axi4_0_r_bits_data,
  input  [1:0]   mem_port_axi4_0_r_bits_resp,
  input          mem_port_axi4_0_r_bits_last,
  input          sys_port_axi4_0_aw_ready,
  output         sys_port_axi4_0_aw_valid,
  output [3:0]   sys_port_axi4_0_aw_bits_id,
  output [30:0]  sys_port_axi4_0_aw_bits_addr,
  output [7:0]   sys_port_axi4_0_aw_bits_len,
  output [2:0]   sys_port_axi4_0_aw_bits_size,
  output [1:0]   sys_port_axi4_0_aw_bits_burst,
  output         sys_port_axi4_0_aw_bits_lock,
  output [3:0]   sys_port_axi4_0_aw_bits_cache,
  output [2:0]   sys_port_axi4_0_aw_bits_prot,
  output [3:0]   sys_port_axi4_0_aw_bits_qos,
  input          sys_port_axi4_0_w_ready,
  output         sys_port_axi4_0_w_valid,
  output [31:0]  sys_port_axi4_0_w_bits_data,
  output [3:0]   sys_port_axi4_0_w_bits_strb,
  output         sys_port_axi4_0_w_bits_last,
  output         sys_port_axi4_0_b_ready,
  input          sys_port_axi4_0_b_valid,
  input  [3:0]   sys_port_axi4_0_b_bits_id,
  input  [1:0]   sys_port_axi4_0_b_bits_resp,
  input          sys_port_axi4_0_ar_ready,
  output         sys_port_axi4_0_ar_valid,
  output [3:0]   sys_port_axi4_0_ar_bits_id,
  output [30:0]  sys_port_axi4_0_ar_bits_addr,
  output [7:0]   sys_port_axi4_0_ar_bits_len,
  output [2:0]   sys_port_axi4_0_ar_bits_size,
  output [1:0]   sys_port_axi4_0_ar_bits_burst,
  output         sys_port_axi4_0_ar_bits_lock,
  output [3:0]   sys_port_axi4_0_ar_bits_cache,
  output [2:0]   sys_port_axi4_0_ar_bits_prot,
  output [3:0]   sys_port_axi4_0_ar_bits_qos,
  output         sys_port_axi4_0_r_ready,
  input          sys_port_axi4_0_r_valid,
  input  [3:0]   sys_port_axi4_0_r_bits_id,
  input  [31:0]  sys_port_axi4_0_r_bits_data,
  input  [1:0]   sys_port_axi4_0_r_bits_resp,
  input          sys_port_axi4_0_r_bits_last,
  input          periph_port_axi4_0_aw_ready,
  output         periph_port_axi4_0_aw_valid,
  output         periph_port_axi4_0_aw_bits_id,
  output [29:0]  periph_port_axi4_0_aw_bits_addr,
  output [7:0]   periph_port_axi4_0_aw_bits_len,
  output [2:0]   periph_port_axi4_0_aw_bits_size,
  output [1:0]   periph_port_axi4_0_aw_bits_burst,
  output         periph_port_axi4_0_aw_bits_lock,
  output [3:0]   periph_port_axi4_0_aw_bits_cache,
  output [2:0]   periph_port_axi4_0_aw_bits_prot,
  output [3:0]   periph_port_axi4_0_aw_bits_qos,
  input          periph_port_axi4_0_w_ready,
  output         periph_port_axi4_0_w_valid,
  output [31:0]  periph_port_axi4_0_w_bits_data,
  output [3:0]   periph_port_axi4_0_w_bits_strb,
  output         periph_port_axi4_0_w_bits_last,
  output         periph_port_axi4_0_b_ready,
  input          periph_port_axi4_0_b_valid,
  input          periph_port_axi4_0_b_bits_id,
  input  [1:0]   periph_port_axi4_0_b_bits_resp,
  input          periph_port_axi4_0_ar_ready,
  output         periph_port_axi4_0_ar_valid,
  output         periph_port_axi4_0_ar_bits_id,
  output [29:0]  periph_port_axi4_0_ar_bits_addr,
  output [7:0]   periph_port_axi4_0_ar_bits_len,
  output [2:0]   periph_port_axi4_0_ar_bits_size,
  output [1:0]   periph_port_axi4_0_ar_bits_burst,
  output         periph_port_axi4_0_ar_bits_lock,
  output [3:0]   periph_port_axi4_0_ar_bits_cache,
  output [2:0]   periph_port_axi4_0_ar_bits_prot,
  output [3:0]   periph_port_axi4_0_ar_bits_qos,
  output         periph_port_axi4_0_r_ready,
  input          periph_port_axi4_0_r_valid,
  input          periph_port_axi4_0_r_bits_id,
  input  [31:0]  periph_port_axi4_0_r_bits_data,
  input  [1:0]   periph_port_axi4_0_r_bits_resp,
  input          periph_port_axi4_0_r_bits_last,
  output         front_port_axi4_0_aw_ready,
  input          front_port_axi4_0_aw_valid,
  input  [7:0]   front_port_axi4_0_aw_bits_id,
  input  [31:0]  front_port_axi4_0_aw_bits_addr,
  input  [7:0]   front_port_axi4_0_aw_bits_len,
  input  [2:0]   front_port_axi4_0_aw_bits_size,
  input  [1:0]   front_port_axi4_0_aw_bits_burst,
  input          front_port_axi4_0_aw_bits_lock,
  input  [3:0]   front_port_axi4_0_aw_bits_cache,
  input  [2:0]   front_port_axi4_0_aw_bits_prot,
  input  [3:0]   front_port_axi4_0_aw_bits_qos,
  output         front_port_axi4_0_w_ready,
  input          front_port_axi4_0_w_valid,
  input  [31:0]  front_port_axi4_0_w_bits_data,
  input  [3:0]   front_port_axi4_0_w_bits_strb,
  input          front_port_axi4_0_w_bits_last,
  input          front_port_axi4_0_b_ready,
  output         front_port_axi4_0_b_valid,
  output [7:0]   front_port_axi4_0_b_bits_id,
  output [1:0]   front_port_axi4_0_b_bits_resp,
  output         front_port_axi4_0_ar_ready,
  input          front_port_axi4_0_ar_valid,
  input  [7:0]   front_port_axi4_0_ar_bits_id,
  input  [31:0]  front_port_axi4_0_ar_bits_addr,
  input  [7:0]   front_port_axi4_0_ar_bits_len,
  input  [2:0]   front_port_axi4_0_ar_bits_size,
  input  [1:0]   front_port_axi4_0_ar_bits_burst,
  input          front_port_axi4_0_ar_bits_lock,
  input  [3:0]   front_port_axi4_0_ar_bits_cache,
  input  [2:0]   front_port_axi4_0_ar_bits_prot,
  input  [3:0]   front_port_axi4_0_ar_bits_qos,
  input          front_port_axi4_0_r_ready,
  output         front_port_axi4_0_r_valid,
  output [7:0]   front_port_axi4_0_r_bits_id,
  output [31:0]  front_port_axi4_0_r_bits_data,
  output [1:0]   front_port_axi4_0_r_bits_resp,
  output         front_port_axi4_0_r_bits_last
);
  wire  SynchronizerShiftReg_w1_d3__EVAL;
  wire  SynchronizerShiftReg_w1_d3__EVAL_0;
  wire  SynchronizerShiftReg_w1_d3__EVAL_1;
  wire  dmiResetCatch__EVAL;
  wire  dmiResetCatch__EVAL_0;
  wire  dmiResetCatch__EVAL_1;
  wire  dmiResetCatch__EVAL_2;
  wire  dmiResetCatch__EVAL_3;
  wire [63:0] sagesafety__EVAL;
  wire  sagesafety__EVAL_0;
  wire [3:0] sagesafety__EVAL_1;
  wire [6:0] sagesafety__EVAL_2;
  wire  sagesafety__EVAL_3;
  wire [29:0] sagesafety__EVAL_4;
  wire [6:0] sagesafety__EVAL_5;
  wire [3:0] sagesafety__EVAL_6;
  wire [3:0] sagesafety__EVAL_7;
  wire [2:0] sagesafety__EVAL_8;
  wire [63:0] sagesafety__EVAL_9;
  wire [3:0] sagesafety__EVAL_10;
  wire [1:0] sagesafety__EVAL_11;
  wire [29:0] sagesafety__EVAL_12;
  wire [2:0] sagesafety__EVAL_13;
  wire  sagesafety__EVAL_14;
  wire  sagesafety__EVAL_15;
  wire [1:0] sagesafety__EVAL_16;
  wire  sagesafety__EVAL_17;
  wire  sagesafety__EVAL_18;
  wire [6:0] sagesafety__EVAL_19;
  wire  sagesafety__EVAL_20;
  wire [6:0] sagesafety__EVAL_21;
  wire  sagesafety__EVAL_22;
  wire  sagesafety__EVAL_23;
  wire [63:0] sagesafety__EVAL_24;
  wire [2:0] sagesafety__EVAL_25;
  wire  sagesafety__EVAL_26;
  wire [2:0] sagesafety__EVAL_27;
  wire  sagesafety__EVAL_28;
  wire  sagesafety__EVAL_29;
  wire  sagesafety__EVAL_30;
  wire  sagesafety__EVAL_31;
  wire [2:0] sagesafety__EVAL_32;
  wire [7:0] sagesafety__EVAL_33;
  wire  sagesafety__EVAL_34;
  wire  sagesafety__EVAL_35;
  wire [7:0] sagesafety__EVAL_36;
  wire [63:0] sagesafety__EVAL_37;
  wire  sagesafety__EVAL_38;
  wire [2:0] sagesafety__EVAL_39;
  wire  sagesafety__EVAL_40;
  wire  dtm__EVAL;
  wire  dtm__EVAL_0;
  wire  dtm__EVAL_1;
  wire  dtm__EVAL_2;
  wire  dtm__EVAL_3;
  wire  dtm__EVAL_4;
  wire  dtm__EVAL_5;
  wire [10:0] dtm__EVAL_6;
  wire  dtm__EVAL_7;
  wire [31:0] dtm__EVAL_8;
  wire [31:0] dtm__EVAL_9;
  wire  dtm__EVAL_10;
  wire  dtm__EVAL_11;
  wire [1:0] dtm__EVAL_12;
  wire [1:0] dtm__EVAL_13;
  wire  dtm__EVAL_14;
  wire [6:0] dtm__EVAL_15;
  wire  dtm__EVAL_16;
  wire [31:0] tile__EVAL;
  wire  tile__EVAL_0;
  wire [31:0] tile__EVAL_1;
  wire  tile__EVAL_2;
  wire [63:0] tile__EVAL_3;
  wire [2:0] tile__EVAL_4;
  wire [6:0] tile__EVAL_5;
  wire [2:0] tile__EVAL_6;
  wire [3:0] tile__EVAL_7;
  wire [1:0] tile__EVAL_8;
  wire  tile__EVAL_9;
  wire [1:0] tile__EVAL_10;
  wire [3:0] tile__EVAL_11;
  wire [2:0] tile__EVAL_12;
  wire  tile__EVAL_13;
  wire [1:0] tile__EVAL_14;
  wire  tile__EVAL_15;
  wire [7:0] tile__EVAL_16;
  wire  tile__EVAL_17;
  wire [3:0] tile__EVAL_18;
  wire [1:0] tile__EVAL_19;
  wire  tile__EVAL_20;
  wire [1:0] tile__EVAL_21;
  wire [31:0] tile__EVAL_22;
  wire  tile__EVAL_23;
  wire  tile__EVAL_24;
  wire [7:0] tile__EVAL_25;
  wire [31:0] tile__EVAL_26;
  wire [31:0] tile__EVAL_27;
  wire [2:0] tile__EVAL_28;
  wire [3:0] tile__EVAL_29;
  wire [1:0] tile__EVAL_30;
  wire  tile__EVAL_31;
  wire  tile__EVAL_32;
  wire [2:0] tile__EVAL_33;
  wire [2:0] tile__EVAL_34;
  wire  tile__EVAL_35;
  wire [2:0] tile__EVAL_36;
  wire [2:0] tile__EVAL_37;
  wire [31:0] tile__EVAL_38;
  wire [31:0] tile__EVAL_39;
  wire [2:0] tile__EVAL_40;
  wire [3:0] tile__EVAL_41;
  wire  tile__EVAL_42;
  wire [1:0] tile__EVAL_43;
  wire  tile__EVAL_44;
  wire [63:0] tile__EVAL_45;
  wire [3:0] tile__EVAL_46;
  wire  tile__EVAL_47;
  wire [6:0] tile__EVAL_48;
  wire [31:0] tile__EVAL_49;
  wire [31:0] tile__EVAL_50;
  wire [1:0] tile__EVAL_51;
  wire [1:0] tile__EVAL_52;
  wire  tile__EVAL_53;
  wire [1:0] tile__EVAL_54;
  wire [2:0] tile__EVAL_55;
  wire [1:0] tile__EVAL_56;
  wire [3:0] tile__EVAL_57;
  wire [2:0] tile__EVAL_58;
  wire [6:0] tile__EVAL_59;
  wire [1:0] tile__EVAL_60;
  wire [1:0] tile__EVAL_61;
  wire [3:0] tile__EVAL_62;
  wire [3:0] tile__EVAL_63;
  wire  tile__EVAL_64;
  wire  tile__EVAL_65;
  wire  tile__EVAL_66;
  wire  tile__EVAL_67;
  wire  tile__EVAL_68;
  wire  tile__EVAL_69;
  wire [1:0] tile__EVAL_70;
  wire [1:0] tile__EVAL_71;
  wire  tile__EVAL_72;
  wire [2:0] tile__EVAL_73;
  wire  tile__EVAL_74;
  wire  tile__EVAL_75;
  wire  tile__EVAL_76;
  wire [2:0] tile__EVAL_77;
  wire [63:0] tile__EVAL_78;
  wire [2:0] tile__EVAL_79;
  wire  tile__EVAL_80;
  wire [1:0] tile__EVAL_81;
  wire [31:0] tile__EVAL_82;
  wire  tile__EVAL_83;
  wire [2:0] tile__EVAL_84;
  wire [6:0] tile__EVAL_85;
  wire [1:0] tile__EVAL_86;
  wire  tile__EVAL_87;
  wire [31:0] tile__EVAL_88;
  wire  tile__EVAL_89;
  wire [24:0] tile__EVAL_90;
  wire [3:0] tile__EVAL_91;
  wire  tile__EVAL_92;
  wire [3:0] tile__EVAL_93;
  wire [2:0] tile__EVAL_94;
  wire  tile__EVAL_95;
  wire [2:0] tile__EVAL_96;
  wire [2:0] tile__EVAL_97;
  wire [24:0] tile__EVAL_98;
  wire [3:0] tile__EVAL_99;
  wire  tile__EVAL_100;
  wire  tile__EVAL_101;
  wire  tile__EVAL_102;
  wire [63:0] tile__EVAL_103;
  wire [3:0] tile__EVAL_104;
  wire  tile__EVAL_105;
  wire [63:0] tile__EVAL_106;
  wire [3:0] tile__EVAL_107;
  wire [1:0] tile__EVAL_108;
  wire  tile__EVAL_109;
  wire [1:0] tile__EVAL_110;
  wire [1:0] tile__EVAL_111;
  wire  tile__EVAL_112;
  wire  tile__EVAL_113;
  wire [2:0] tile__EVAL_114;
  wire [2:0] tile__EVAL_115;
  wire [63:0] tile__EVAL_116;
  wire  tile__EVAL_117;
  wire  tile__EVAL_118;
  wire [11:0] plic__EVAL;
  wire  plic__EVAL_0;
  wire  plic__EVAL_1;
  wire  plic__EVAL_2;
  wire  plic__EVAL_3;
  wire  plic__EVAL_4;
  wire  plic__EVAL_5;
  wire  plic__EVAL_6;
  wire  plic__EVAL_7;
  wire  plic__EVAL_8;
  wire  plic__EVAL_9;
  wire  plic__EVAL_10;
  wire  plic__EVAL_11;
  wire  plic__EVAL_12;
  wire  plic__EVAL_13;
  wire  plic__EVAL_14;
  wire  plic__EVAL_15;
  wire  plic__EVAL_16;
  wire  plic__EVAL_17;
  wire  plic__EVAL_18;
  wire  plic__EVAL_19;
  wire [11:0] plic__EVAL_20;
  wire  plic__EVAL_21;
  wire  plic__EVAL_22;
  wire  plic__EVAL_23;
  wire  plic__EVAL_24;
  wire  plic__EVAL_25;
  wire  plic__EVAL_26;
  wire  plic__EVAL_27;
  wire  plic__EVAL_28;
  wire  plic__EVAL_29;
  wire  plic__EVAL_30;
  wire  plic__EVAL_31;
  wire  plic__EVAL_32;
  wire  plic__EVAL_33;
  wire  plic__EVAL_34;
  wire  plic__EVAL_35;
  wire  plic__EVAL_36;
  wire  plic__EVAL_37;
  wire [2:0] plic__EVAL_38;
  wire  plic__EVAL_39;
  wire  plic__EVAL_40;
  wire  plic__EVAL_41;
  wire  plic__EVAL_42;
  wire  plic__EVAL_43;
  wire  plic__EVAL_44;
  wire  plic__EVAL_45;
  wire  plic__EVAL_46;
  wire  plic__EVAL_47;
  wire  plic__EVAL_48;
  wire  plic__EVAL_49;
  wire  plic__EVAL_50;
  wire [27:0] plic__EVAL_51;
  wire  plic__EVAL_52;
  wire  plic__EVAL_53;
  wire  plic__EVAL_54;
  wire  plic__EVAL_55;
  wire  plic__EVAL_56;
  wire  plic__EVAL_57;
  wire  plic__EVAL_58;
  wire  plic__EVAL_59;
  wire  plic__EVAL_60;
  wire  plic__EVAL_61;
  wire [1:0] plic__EVAL_62;
  wire  plic__EVAL_63;
  wire  plic__EVAL_64;
  wire  plic__EVAL_65;
  wire  plic__EVAL_66;
  wire  plic__EVAL_67;
  wire  plic__EVAL_68;
  wire [3:0] plic__EVAL_69;
  wire  plic__EVAL_70;
  wire  plic__EVAL_71;
  wire  plic__EVAL_72;
  wire  plic__EVAL_73;
  wire  plic__EVAL_74;
  wire  plic__EVAL_75;
  wire  plic__EVAL_76;
  wire  plic__EVAL_77;
  wire  plic__EVAL_78;
  wire [1:0] plic__EVAL_79;
  wire  plic__EVAL_80;
  wire  plic__EVAL_81;
  wire  plic__EVAL_82;
  wire  plic__EVAL_83;
  wire [31:0] plic__EVAL_84;
  wire  plic__EVAL_85;
  wire [2:0] plic__EVAL_86;
  wire  plic__EVAL_87;
  wire  plic__EVAL_88;
  wire  plic__EVAL_89;
  wire  plic__EVAL_90;
  wire  plic__EVAL_91;
  wire  plic__EVAL_92;
  wire  plic__EVAL_93;
  wire  plic__EVAL_94;
  wire  plic__EVAL_95;
  wire  plic__EVAL_96;
  wire  plic__EVAL_97;
  wire  plic__EVAL_98;
  wire  plic__EVAL_99;
  wire  plic__EVAL_100;
  wire  plic__EVAL_101;
  wire  plic__EVAL_102;
  wire  plic__EVAL_103;
  wire  plic__EVAL_104;
  wire  plic__EVAL_105;
  wire  plic__EVAL_106;
  wire  plic__EVAL_107;
  wire  plic__EVAL_108;
  wire  plic__EVAL_109;
  wire  plic__EVAL_110;
  wire  plic__EVAL_111;
  wire  plic__EVAL_112;
  wire  plic__EVAL_113;
  wire  plic__EVAL_114;
  wire  plic__EVAL_115;
  wire  plic__EVAL_116;
  wire  plic__EVAL_117;
  wire  plic__EVAL_118;
  wire  plic__EVAL_119;
  wire  plic__EVAL_120;
  wire  plic__EVAL_121;
  wire  plic__EVAL_122;
  wire  plic__EVAL_123;
  wire  plic__EVAL_124;
  wire  plic__EVAL_125;
  wire  plic__EVAL_126;
  wire  plic__EVAL_127;
  wire  plic__EVAL_128;
  wire  plic__EVAL_129;
  wire [31:0] plic__EVAL_130;
  wire  plic__EVAL_131;
  wire  plic__EVAL_132;
  wire  plic__EVAL_133;
  wire  plic__EVAL_134;
  wire  plic__EVAL_135;
  wire  plic__EVAL_136;
  wire  plic__EVAL_137;
  wire  plic__EVAL_138;
  wire  plic__EVAL_139;
  wire  plic__EVAL_140;
  wire  plic__EVAL_141;
  wire  plic__EVAL_142;
  wire [2:0] plic__EVAL_143;
  wire  plic__EVAL_144;
  wire [8:0] ww__EVAL;
  wire [8:0] ww__EVAL_0;
  wire [8:0] ww__EVAL_1;
  wire [7:0] ww__EVAL_2;
  wire [8:0] ww__EVAL_3;
  wire  ww__EVAL_4;
  wire [2:0] ww__EVAL_5;
  wire  ww__EVAL_6;
  wire [2:0] ww__EVAL_7;
  wire [31:0] ww__EVAL_8;
  wire  ww__EVAL_9;
  wire [63:0] ww__EVAL_10;
  wire  ww__EVAL_11;
  wire [2:0] ww__EVAL_12;
  wire  ww__EVAL_13;
  wire [63:0] ww__EVAL_14;
  wire  ww__EVAL_15;
  wire  ww__EVAL_16;
  wire [2:0] ww__EVAL_17;
  wire [2:0] ww__EVAL_18;
  wire [2:0] ww__EVAL_19;
  wire  ww__EVAL_20;
  wire  ww__EVAL_21;
  wire  ww__EVAL_22;
  wire [63:0] ww__EVAL_23;
  wire [2:0] ww__EVAL_24;
  wire [7:0] ww__EVAL_25;
  wire [2:0] ww__EVAL_26;
  wire [2:0] ww__EVAL_27;
  wire  ww__EVAL_28;
  wire [63:0] ww__EVAL_29;
  wire  ww__EVAL_30;
  wire  ww__EVAL_31;
  wire  ww__EVAL_32;
  wire  ww__EVAL_33;
  wire [2:0] ww__EVAL_34;
  wire [31:0] ww__EVAL_35;
  wire  ww__EVAL_36;
  wire  sbus__EVAL;
  wire [3:0] sbus__EVAL_0;
  wire [1:0] sbus__EVAL_1;
  wire [7:0] sbus__EVAL_2;
  wire [2:0] sbus__EVAL_3;
  wire [63:0] sbus__EVAL_4;
  wire  sbus__EVAL_5;
  wire  sbus__EVAL_6;
  wire  sbus__EVAL_7;
  wire [3:0] sbus__EVAL_8;
  wire [63:0] sbus__EVAL_9;
  wire [1:0] sbus__EVAL_10;
  wire [31:0] sbus__EVAL_11;
  wire [3:0] sbus__EVAL_12;
  wire [1:0] sbus__EVAL_13;
  wire  sbus__EVAL_14;
  wire [7:0] sbus__EVAL_15;
  wire [31:0] sbus__EVAL_16;
  wire  sbus__EVAL_17;
  wire [2:0] sbus__EVAL_18;
  wire  sbus__EVAL_19;
  wire [2:0] sbus__EVAL_20;
  wire [1:0] sbus__EVAL_21;
  wire [1:0] sbus__EVAL_22;
  wire [2:0] sbus__EVAL_23;
  wire [1:0] sbus__EVAL_24;
  wire [6:0] sbus__EVAL_25;
  wire [3:0] sbus__EVAL_26;
  wire  sbus__EVAL_27;
  wire [2:0] sbus__EVAL_28;
  wire [3:0] sbus__EVAL_29;
  wire [30:0] sbus__EVAL_30;
  wire  sbus__EVAL_31;
  wire  sbus__EVAL_32;
  wire  sbus__EVAL_33;
  wire [3:0] sbus__EVAL_34;
  wire [2:0] sbus__EVAL_35;
  wire [3:0] sbus__EVAL_36;
  wire [2:0] sbus__EVAL_37;
  wire [3:0] sbus__EVAL_38;
  wire [2:0] sbus__EVAL_39;
  wire [2:0] sbus__EVAL_40;
  wire  sbus__EVAL_41;
  wire [2:0] sbus__EVAL_42;
  wire  sbus__EVAL_43;
  wire [5:0] sbus__EVAL_44;
  wire [1:0] sbus__EVAL_45;
  wire  sbus__EVAL_46;
  wire [3:0] sbus__EVAL_47;
  wire [31:0] sbus__EVAL_48;
  wire [2:0] sbus__EVAL_49;
  wire  sbus__EVAL_50;
  wire [1:0] sbus__EVAL_51;
  wire  sbus__EVAL_52;
  wire  sbus__EVAL_53;
  wire [1:0] sbus__EVAL_54;
  wire [3:0] sbus__EVAL_55;
  wire  sbus__EVAL_56;
  wire  sbus__EVAL_57;
  wire  sbus__EVAL_58;
  wire [1:0] sbus__EVAL_59;
  wire [2:0] sbus__EVAL_60;
  wire  sbus__EVAL_61;
  wire [31:0] sbus__EVAL_62;
  wire  sbus__EVAL_63;
  wire [6:0] sbus__EVAL_64;
  wire [2:0] sbus__EVAL_65;
  wire [31:0] sbus__EVAL_66;
  wire  sbus__EVAL_67;
  wire [1:0] sbus__EVAL_68;
  wire  sbus__EVAL_69;
  wire [63:0] sbus__EVAL_70;
  wire [63:0] sbus__EVAL_71;
  wire [30:0] sbus__EVAL_72;
  wire [63:0] sbus__EVAL_73;
  wire [63:0] sbus__EVAL_74;
  wire [31:0] sbus__EVAL_75;
  wire  sbus__EVAL_76;
  wire [1:0] sbus__EVAL_77;
  wire [2:0] sbus__EVAL_78;
  wire [3:0] sbus__EVAL_79;
  wire [6:0] sbus__EVAL_80;
  wire [3:0] sbus__EVAL_81;
  wire  sbus__EVAL_82;
  wire  sbus__EVAL_83;
  wire [31:0] sbus__EVAL_84;
  wire [2:0] sbus__EVAL_85;
  wire [2:0] sbus__EVAL_86;
  wire [1:0] sbus__EVAL_87;
  wire [6:0] sbus__EVAL_88;
  wire [31:0] sbus__EVAL_89;
  wire  sbus__EVAL_90;
  wire  sbus__EVAL_91;
  wire [31:0] sbus__EVAL_92;
  wire [31:0] sbus__EVAL_93;
  wire [1:0] sbus__EVAL_94;
  wire [2:0] sbus__EVAL_95;
  wire [31:0] sbus__EVAL_96;
  wire [1:0] sbus__EVAL_97;
  wire  sbus__EVAL_98;
  wire [3:0] sbus__EVAL_99;
  wire [1:0] sbus__EVAL_100;
  wire  sbus__EVAL_101;
  wire [7:0] sbus__EVAL_102;
  wire  sbus__EVAL_103;
  wire  sbus__EVAL_104;
  wire [63:0] sbus__EVAL_105;
  wire  sbus__EVAL_106;
  wire [3:0] sbus__EVAL_107;
  wire [1:0] sbus__EVAL_108;
  wire [3:0] sbus__EVAL_109;
  wire  sbus__EVAL_110;
  wire [2:0] sbus__EVAL_111;
  wire [2:0] sbus__EVAL_112;
  wire  sbus__EVAL_113;
  wire  sbus__EVAL_114;
  wire  sbus__EVAL_115;
  wire [6:0] sbus__EVAL_116;
  wire [3:0] sbus__EVAL_117;
  wire [3:0] sbus__EVAL_118;
  wire [6:0] sbus__EVAL_119;
  wire [3:0] sbus__EVAL_120;
  wire  sbus__EVAL_121;
  wire  sbus__EVAL_122;
  wire [1:0] sbus__EVAL_123;
  wire  sbus__EVAL_124;
  wire [29:0] sbus__EVAL_125;
  wire  sbus__EVAL_126;
  wire  sbus__EVAL_127;
  wire [6:0] sbus__EVAL_128;
  wire  sbus__EVAL_129;
  wire [2:0] sbus__EVAL_130;
  wire [3:0] sbus__EVAL_131;
  wire [2:0] sbus__EVAL_132;
  wire  sbus__EVAL_133;
  wire  sbus__EVAL_134;
  wire  sbus__EVAL_135;
  wire  sbus__EVAL_136;
  wire  sbus__EVAL_137;
  wire [3:0] sbus__EVAL_138;
  wire  sbus__EVAL_139;
  wire [2:0] sbus__EVAL_140;
  wire  sbus__EVAL_141;
  wire [7:0] sbus__EVAL_142;
  wire [63:0] sbus__EVAL_143;
  wire  sbus__EVAL_144;
  wire [31:0] sbus__EVAL_145;
  wire  sbus__EVAL_146;
  wire  sbus__EVAL_147;
  wire  sbus__EVAL_148;
  wire  sbus__EVAL_149;
  wire  sbus__EVAL_150;
  wire [3:0] sbus__EVAL_151;
  wire [6:0] sbus__EVAL_152;
  wire  sbus__EVAL_153;
  wire  sbus__EVAL_154;
  wire [2:0] sbus__EVAL_155;
  wire  sbus__EVAL_156;
  wire [2:0] sbus__EVAL_157;
  wire [2:0] sbus__EVAL_158;
  wire  sbus__EVAL_159;
  wire  sbus__EVAL_160;
  wire [1:0] sbus__EVAL_161;
  wire [2:0] sbus__EVAL_162;
  wire [3:0] sbus__EVAL_163;
  wire  sbus__EVAL_164;
  wire  sbus__EVAL_165;
  wire  sbus__EVAL_166;
  wire  sbus__EVAL_167;
  wire [7:0] sbus__EVAL_168;
  wire  sbus__EVAL_169;
  wire  sbus__EVAL_170;
  wire  sbus__EVAL_171;
  wire [31:0] sbus__EVAL_172;
  wire [3:0] sbus__EVAL_173;
  wire [1:0] sbus__EVAL_174;
  wire [3:0] sbus__EVAL_175;
  wire [3:0] sbus__EVAL_176;
  wire [31:0] sbus__EVAL_177;
  wire  sbus__EVAL_178;
  wire [3:0] sbus__EVAL_179;
  wire [31:0] sbus__EVAL_180;
  wire [29:0] sbus__EVAL_181;
  wire [3:0] sbus__EVAL_182;
  wire  sbus__EVAL_183;
  wire [63:0] sbus__EVAL_184;
  wire [7:0] sbus__EVAL_185;
  wire [2:0] sbus__EVAL_186;
  wire [31:0] sbus__EVAL_187;
  wire [5:0] sbus__EVAL_188;
  wire [2:0] sbus__EVAL_189;
  wire [63:0] sbus__EVAL_190;
  wire [2:0] sbus__EVAL_191;
  wire [6:0] sbus__EVAL_192;
  wire [63:0] sbus__EVAL_193;
  wire [2:0] sbus__EVAL_194;
  wire  sbus__EVAL_195;
  wire [3:0] sbus__EVAL_196;
  wire [63:0] sbus__EVAL_197;
  wire [1:0] sbus__EVAL_198;
  wire [29:0] sbus__EVAL_199;
  wire [63:0] sbus__EVAL_200;
  wire [3:0] sbus__EVAL_201;
  wire  sbus__EVAL_202;
  wire  sbus__EVAL_203;
  wire [1:0] sbus__EVAL_204;
  wire  sbus__EVAL_205;
  wire [2:0] sbus__EVAL_206;
  wire  sbus__EVAL_207;
  wire [1:0] sbus__EVAL_208;
  wire [2:0] sbus__EVAL_209;
  wire [7:0] sbus__EVAL_210;
  wire  sbus__EVAL_211;
  wire  sbus__EVAL_212;
  wire  sbus__EVAL_213;
  wire  sbus__EVAL_214;
  wire [1:0] sbus__EVAL_215;
  wire  sbus__EVAL_216;
  wire [2:0] sbus__EVAL_217;
  wire  sbus__EVAL_218;
  wire  sbus__EVAL_219;
  wire  sbus__EVAL_220;
  wire [3:0] sbus__EVAL_221;
  wire  sbus__EVAL_222;
  wire [3:0] sbus__EVAL_223;
  wire [2:0] sbus__EVAL_224;
  wire  int_bus__EVAL;
  wire  int_bus__EVAL_0;
  wire  int_bus__EVAL_1;
  wire  int_bus__EVAL_2;
  wire  int_bus__EVAL_3;
  wire  int_bus__EVAL_4;
  wire  int_bus__EVAL_5;
  wire  int_bus__EVAL_6;
  wire  int_bus__EVAL_7;
  wire  int_bus__EVAL_8;
  wire  int_bus__EVAL_9;
  wire  int_bus__EVAL_10;
  wire  int_bus__EVAL_11;
  wire  int_bus__EVAL_12;
  wire  int_bus__EVAL_13;
  wire  int_bus__EVAL_14;
  wire  int_bus__EVAL_15;
  wire  int_bus__EVAL_16;
  wire  int_bus__EVAL_17;
  wire  int_bus__EVAL_18;
  wire  int_bus__EVAL_19;
  wire  int_bus__EVAL_20;
  wire  int_bus__EVAL_21;
  wire  int_bus__EVAL_22;
  wire  int_bus__EVAL_23;
  wire  int_bus__EVAL_24;
  wire  int_bus__EVAL_25;
  wire  int_bus__EVAL_26;
  wire  int_bus__EVAL_27;
  wire  int_bus__EVAL_28;
  wire  int_bus__EVAL_29;
  wire  int_bus__EVAL_30;
  wire  int_bus__EVAL_31;
  wire  int_bus__EVAL_32;
  wire  int_bus__EVAL_33;
  wire  int_bus__EVAL_34;
  wire  int_bus__EVAL_35;
  wire  int_bus__EVAL_36;
  wire  int_bus__EVAL_37;
  wire  int_bus__EVAL_38;
  wire  int_bus__EVAL_39;
  wire  int_bus__EVAL_40;
  wire  int_bus__EVAL_41;
  wire  int_bus__EVAL_42;
  wire  int_bus__EVAL_43;
  wire  int_bus__EVAL_44;
  wire  int_bus__EVAL_45;
  wire  int_bus__EVAL_46;
  wire  int_bus__EVAL_47;
  wire  int_bus__EVAL_48;
  wire  int_bus__EVAL_49;
  wire  int_bus__EVAL_50;
  wire  int_bus__EVAL_51;
  wire  int_bus__EVAL_52;
  wire  int_bus__EVAL_53;
  wire  int_bus__EVAL_54;
  wire  int_bus__EVAL_55;
  wire  int_bus__EVAL_56;
  wire  int_bus__EVAL_57;
  wire  int_bus__EVAL_58;
  wire  int_bus__EVAL_59;
  wire  int_bus__EVAL_60;
  wire  int_bus__EVAL_61;
  wire  int_bus__EVAL_62;
  wire  int_bus__EVAL_63;
  wire  int_bus__EVAL_64;
  wire  int_bus__EVAL_65;
  wire  int_bus__EVAL_66;
  wire  int_bus__EVAL_67;
  wire  int_bus__EVAL_68;
  wire  int_bus__EVAL_69;
  wire  int_bus__EVAL_70;
  wire  int_bus__EVAL_71;
  wire  int_bus__EVAL_72;
  wire  int_bus__EVAL_73;
  wire  int_bus__EVAL_74;
  wire  int_bus__EVAL_75;
  wire  int_bus__EVAL_76;
  wire  int_bus__EVAL_77;
  wire  int_bus__EVAL_78;
  wire  int_bus__EVAL_79;
  wire  int_bus__EVAL_80;
  wire  int_bus__EVAL_81;
  wire  int_bus__EVAL_82;
  wire  int_bus__EVAL_83;
  wire  int_bus__EVAL_84;
  wire  int_bus__EVAL_85;
  wire  int_bus__EVAL_86;
  wire  int_bus__EVAL_87;
  wire  int_bus__EVAL_88;
  wire  int_bus__EVAL_89;
  wire  int_bus__EVAL_90;
  wire  int_bus__EVAL_91;
  wire  int_bus__EVAL_92;
  wire  int_bus__EVAL_93;
  wire  int_bus__EVAL_94;
  wire  int_bus__EVAL_95;
  wire  int_bus__EVAL_96;
  wire  int_bus__EVAL_97;
  wire  int_bus__EVAL_98;
  wire  int_bus__EVAL_99;
  wire  int_bus__EVAL_100;
  wire  int_bus__EVAL_101;
  wire  int_bus__EVAL_102;
  wire  int_bus__EVAL_103;
  wire  int_bus__EVAL_104;
  wire  int_bus__EVAL_105;
  wire  int_bus__EVAL_106;
  wire  int_bus__EVAL_107;
  wire  int_bus__EVAL_108;
  wire  int_bus__EVAL_109;
  wire  int_bus__EVAL_110;
  wire  int_bus__EVAL_111;
  wire  int_bus__EVAL_112;
  wire  int_bus__EVAL_113;
  wire  int_bus__EVAL_114;
  wire  int_bus__EVAL_115;
  wire  int_bus__EVAL_116;
  wire  int_bus__EVAL_117;
  wire  int_bus__EVAL_118;
  wire  int_bus__EVAL_119;
  wire  int_bus__EVAL_120;
  wire  int_bus__EVAL_121;
  wire  int_bus__EVAL_122;
  wire  int_bus__EVAL_123;
  wire  int_bus__EVAL_124;
  wire  int_bus__EVAL_125;
  wire  int_bus__EVAL_126;
  wire  int_bus__EVAL_127;
  wire  int_bus__EVAL_128;
  wire  int_bus__EVAL_129;
  wire  int_bus__EVAL_130;
  wire  int_bus__EVAL_131;
  wire  int_bus__EVAL_132;
  wire  int_bus__EVAL_133;
  wire  int_bus__EVAL_134;
  wire  int_bus__EVAL_135;
  wire  int_bus__EVAL_136;
  wire  int_bus__EVAL_137;
  wire  int_bus__EVAL_138;
  wire  int_bus__EVAL_139;
  wire  int_bus__EVAL_140;
  wire  int_bus__EVAL_141;
  wire  int_bus__EVAL_142;
  wire  int_bus__EVAL_143;
  wire  int_bus__EVAL_144;
  wire  int_bus__EVAL_145;
  wire  int_bus__EVAL_146;
  wire  int_bus__EVAL_147;
  wire  int_bus__EVAL_148;
  wire  int_bus__EVAL_149;
  wire  int_bus__EVAL_150;
  wire  int_bus__EVAL_151;
  wire  int_bus__EVAL_152;
  wire  int_bus__EVAL_153;
  wire  int_bus__EVAL_154;
  wire  int_bus__EVAL_155;
  wire  int_bus__EVAL_156;
  wire  int_bus__EVAL_157;
  wire  int_bus__EVAL_158;
  wire  int_bus__EVAL_159;
  wire  int_bus__EVAL_160;
  wire  int_bus__EVAL_161;
  wire  int_bus__EVAL_162;
  wire  int_bus__EVAL_163;
  wire  int_bus__EVAL_164;
  wire  int_bus__EVAL_165;
  wire  int_bus__EVAL_166;
  wire  int_bus__EVAL_167;
  wire  int_bus__EVAL_168;
  wire  int_bus__EVAL_169;
  wire  int_bus__EVAL_170;
  wire  int_bus__EVAL_171;
  wire  int_bus__EVAL_172;
  wire  int_bus__EVAL_173;
  wire  int_bus__EVAL_174;
  wire  int_bus__EVAL_175;
  wire  int_bus__EVAL_176;
  wire  int_bus__EVAL_177;
  wire  int_bus__EVAL_178;
  wire  int_bus__EVAL_179;
  wire  int_bus__EVAL_180;
  wire  int_bus__EVAL_181;
  wire  int_bus__EVAL_182;
  wire  int_bus__EVAL_183;
  wire  int_bus__EVAL_184;
  wire  int_bus__EVAL_185;
  wire  int_bus__EVAL_186;
  wire  int_bus__EVAL_187;
  wire  int_bus__EVAL_188;
  wire  int_bus__EVAL_189;
  wire  int_bus__EVAL_190;
  wire  int_bus__EVAL_191;
  wire  int_bus__EVAL_192;
  wire  int_bus__EVAL_193;
  wire  int_bus__EVAL_194;
  wire  int_bus__EVAL_195;
  wire  int_bus__EVAL_196;
  wire  int_bus__EVAL_197;
  wire  int_bus__EVAL_198;
  wire  int_bus__EVAL_199;
  wire  int_bus__EVAL_200;
  wire  int_bus__EVAL_201;
  wire  int_bus__EVAL_202;
  wire  int_bus__EVAL_203;
  wire  int_bus__EVAL_204;
  wire  int_bus__EVAL_205;
  wire  int_bus__EVAL_206;
  wire  int_bus__EVAL_207;
  wire  int_bus__EVAL_208;
  wire  int_bus__EVAL_209;
  wire  int_bus__EVAL_210;
  wire  int_bus__EVAL_211;
  wire  int_bus__EVAL_212;
  wire  int_bus__EVAL_213;
  wire  int_bus__EVAL_214;
  wire  int_bus__EVAL_215;
  wire  int_bus__EVAL_216;
  wire  int_bus__EVAL_217;
  wire  int_bus__EVAL_218;
  wire  int_bus__EVAL_219;
  wire  int_bus__EVAL_220;
  wire  int_bus__EVAL_221;
  wire  int_bus__EVAL_222;
  wire  int_bus__EVAL_223;
  wire  int_bus__EVAL_224;
  wire  int_bus__EVAL_225;
  wire  int_bus__EVAL_226;
  wire  int_bus__EVAL_227;
  wire  int_bus__EVAL_228;
  wire  int_bus__EVAL_229;
  wire  int_bus__EVAL_230;
  wire  int_bus__EVAL_231;
  wire  int_bus__EVAL_232;
  wire  int_bus__EVAL_233;
  wire  int_bus__EVAL_234;
  wire  int_bus__EVAL_235;
  wire  int_bus__EVAL_236;
  wire  int_bus__EVAL_237;
  wire  int_bus__EVAL_238;
  wire  int_bus__EVAL_239;
  wire  int_bus__EVAL_240;
  wire  int_bus__EVAL_241;
  wire  int_bus__EVAL_242;
  wire  int_bus__EVAL_243;
  wire  int_bus__EVAL_244;
  wire  int_bus__EVAL_245;
  wire  int_bus__EVAL_246;
  wire  int_bus__EVAL_247;
  wire  int_bus__EVAL_248;
  wire  int_bus__EVAL_249;
  wire  int_bus__EVAL_250;
  wire  int_bus__EVAL_251;
  wire  int_bus__EVAL_252;
  wire  intsource__EVAL;
  wire  intsource__EVAL_0;
  wire  intsource__EVAL_1;
  wire  intsource__EVAL_2;
  wire  intsource__EVAL_3;
  wire  intsource__EVAL_4;
  wire [5:0] fbus__EVAL;
  wire  fbus__EVAL_0;
  wire [7:0] fbus__EVAL_1;
  wire  fbus__EVAL_2;
  wire  fbus__EVAL_3;
  wire  fbus__EVAL_4;
  wire [31:0] fbus__EVAL_5;
  wire [7:0] fbus__EVAL_6;
  wire  fbus__EVAL_7;
  wire [31:0] fbus__EVAL_8;
  wire  fbus__EVAL_9;
  wire [7:0] fbus__EVAL_10;
  wire [2:0] fbus__EVAL_11;
  wire [2:0] fbus__EVAL_12;
  wire [31:0] fbus__EVAL_13;
  wire [2:0] fbus__EVAL_14;
  wire  fbus__EVAL_15;
  wire [2:0] fbus__EVAL_16;
  wire [7:0] fbus__EVAL_17;
  wire [1:0] fbus__EVAL_18;
  wire  fbus__EVAL_19;
  wire [3:0] fbus__EVAL_20;
  wire  fbus__EVAL_21;
  wire  fbus__EVAL_22;
  wire [31:0] fbus__EVAL_23;
  wire  fbus__EVAL_24;
  wire  fbus__EVAL_25;
  wire [31:0] fbus__EVAL_26;
  wire  fbus__EVAL_27;
  wire [7:0] fbus__EVAL_28;
  wire [1:0] fbus__EVAL_29;
  wire  fbus__EVAL_30;
  wire [7:0] fbus__EVAL_31;
  wire [1:0] fbus__EVAL_32;
  wire [7:0] fbus__EVAL_33;
  wire [1:0] fbus__EVAL_34;
  wire [2:0] fbus__EVAL_35;
  wire  fbus__EVAL_36;
  wire  fbus__EVAL_37;
  wire  fbus__EVAL_38;
  wire  fbus__EVAL_39;
  wire [5:0] fbus__EVAL_40;
  wire [7:0] fbus__EVAL_41;
  wire  fbus__EVAL_42;
  wire  fbus__EVAL_43;
  wire  fbus__EVAL_44;
  wire [3:0] fbus__EVAL_45;
  wire [31:0] fbus__EVAL_46;
  wire [3:0] fbus__EVAL_47;
  wire [2:0] fbus__EVAL_48;
  wire  fbus__EVAL_49;
  wire [31:0] fbus__EVAL_50;
  wire  fbus__EVAL_51;
  wire [3:0] fbus__EVAL_52;
  wire  fbus__EVAL_53;
  wire  fbus__EVAL_54;
  wire  fbus__EVAL_55;
  wire [3:0] fbus__EVAL_56;
  wire  fbus__EVAL_57;
  wire [31:0] fbus__EVAL_58;
  wire [1:0] fbus__EVAL_59;
  wire  fbus__EVAL_60;
  wire [1:0] debug_1__EVAL;
  wire  debug_1__EVAL_0;
  wire [2:0] debug_1__EVAL_1;
  wire [11:0] debug_1__EVAL_2;
  wire  debug_1__EVAL_3;
  wire [1:0] debug_1__EVAL_4;
  wire  debug_1__EVAL_5;
  wire [11:0] debug_1__EVAL_6;
  wire  debug_1__EVAL_7;
  wire  debug_1__EVAL_8;
  wire  debug_1__EVAL_9;
  wire [1:0] debug_1__EVAL_10;
  wire [31:0] debug_1__EVAL_11;
  wire  debug_1__EVAL_12;
  wire [31:0] debug_1__EVAL_13;
  wire [7:0] debug_1__EVAL_14;
  wire [2:0] debug_1__EVAL_15;
  wire [3:0] debug_1__EVAL_16;
  wire [2:0] debug_1__EVAL_17;
  wire [1:0] debug_1__EVAL_18;
  wire  debug_1__EVAL_19;
  wire  debug_1__EVAL_20;
  wire  debug_1__EVAL_21;
  wire  debug_1__EVAL_22;
  wire  debug_1__EVAL_23;
  wire  debug_1__EVAL_24;
  wire [31:0] debug_1__EVAL_25;
  wire [2:0] debug_1__EVAL_26;
  wire [31:0] debug_1__EVAL_27;
  wire  debug_1__EVAL_28;
  wire  debug_1__EVAL_29;
  wire  debug_1__EVAL_30;
  wire  debug_1__EVAL_31;
  wire [7:0] debug_1__EVAL_32;
  wire [31:0] debug_1__EVAL_33;
  wire  debug_1__EVAL_34;
  wire [6:0] debug_1__EVAL_35;
  wire  debug_1__EVAL_36;
  wire  debug_1__EVAL_37;
  wire  debug_1__EVAL_38;
  wire  debug_1__EVAL_39;
  wire  debug_1__EVAL_40;
  wire [3:0] debug_1__EVAL_41;
  wire [11:0] debug_1__EVAL_42;
  wire  debug_1__EVAL_43;
  wire [2:0] cbus__EVAL;
  wire  cbus__EVAL_0;
  wire [1:0] cbus__EVAL_1;
  wire [1:0] cbus__EVAL_2;
  wire [2:0] cbus__EVAL_3;
  wire [3:0] cbus__EVAL_4;
  wire  cbus__EVAL_5;
  wire  cbus__EVAL_6;
  wire [3:0] cbus__EVAL_7;
  wire [31:0] cbus__EVAL_8;
  wire [27:0] cbus__EVAL_9;
  wire [1:0] cbus__EVAL_10;
  wire  cbus__EVAL_11;
  wire  cbus__EVAL_12;
  wire [31:0] cbus__EVAL_13;
  wire [1:0] cbus__EVAL_14;
  wire [31:0] cbus__EVAL_15;
  wire [6:0] cbus__EVAL_16;
  wire [31:0] cbus__EVAL_17;
  wire [29:0] cbus__EVAL_18;
  wire [31:0] cbus__EVAL_19;
  wire [2:0] cbus__EVAL_20;
  wire [2:0] cbus__EVAL_21;
  wire  cbus__EVAL_22;
  wire [29:0] cbus__EVAL_23;
  wire [1:0] cbus__EVAL_24;
  wire  cbus__EVAL_25;
  wire [2:0] cbus__EVAL_26;
  wire [1:0] cbus__EVAL_27;
  wire [6:0] cbus__EVAL_28;
  wire [6:0] cbus__EVAL_29;
  wire  cbus__EVAL_30;
  wire [2:0] cbus__EVAL_31;
  wire [3:0] cbus__EVAL_32;
  wire [1:0] cbus__EVAL_33;
  wire [3:0] cbus__EVAL_34;
  wire [2:0] cbus__EVAL_35;
  wire  cbus__EVAL_36;
  wire [3:0] cbus__EVAL_37;
  wire  cbus__EVAL_38;
  wire [1:0] cbus__EVAL_39;
  wire [2:0] cbus__EVAL_40;
  wire [1:0] cbus__EVAL_41;
  wire [31:0] cbus__EVAL_42;
  wire  cbus__EVAL_43;
  wire  cbus__EVAL_44;
  wire [2:0] cbus__EVAL_45;
  wire [31:0] cbus__EVAL_46;
  wire [7:0] cbus__EVAL_47;
  wire  cbus__EVAL_48;
  wire [31:0] cbus__EVAL_49;
  wire [2:0] cbus__EVAL_50;
  wire  cbus__EVAL_51;
  wire [1:0] cbus__EVAL_52;
  wire  cbus__EVAL_53;
  wire [31:0] cbus__EVAL_54;
  wire [2:0] cbus__EVAL_55;
  wire [3:0] cbus__EVAL_56;
  wire [31:0] cbus__EVAL_57;
  wire  cbus__EVAL_58;
  wire [31:0] cbus__EVAL_59;
  wire [1:0] cbus__EVAL_60;
  wire [1:0] cbus__EVAL_61;
  wire [1:0] cbus__EVAL_62;
  wire  cbus__EVAL_63;
  wire [2:0] cbus__EVAL_64;
  wire  cbus__EVAL_65;
  wire [2:0] cbus__EVAL_66;
  wire [2:0] cbus__EVAL_67;
  wire [2:0] cbus__EVAL_68;
  wire  cbus__EVAL_69;
  wire [24:0] cbus__EVAL_70;
  wire  cbus__EVAL_71;
  wire [11:0] cbus__EVAL_72;
  wire [1:0] cbus__EVAL_73;
  wire [2:0] cbus__EVAL_74;
  wire [11:0] cbus__EVAL_75;
  wire [3:0] cbus__EVAL_76;
  wire [2:0] cbus__EVAL_77;
  wire [14:0] cbus__EVAL_78;
  wire [7:0] cbus__EVAL_79;
  wire [2:0] cbus__EVAL_80;
  wire [11:0] cbus__EVAL_81;
  wire  cbus__EVAL_82;
  wire [11:0] cbus__EVAL_83;
  wire  cbus__EVAL_84;
  wire  cbus__EVAL_85;
  wire  cbus__EVAL_86;
  wire [31:0] cbus__EVAL_87;
  wire  cbus__EVAL_88;
  wire [6:0] cbus__EVAL_89;
  wire  cbus__EVAL_90;
  wire [25:0] cbus__EVAL_91;
  wire  cbus__EVAL_92;
  wire [2:0] cbus__EVAL_93;
  wire [2:0] cbus__EVAL_94;
  wire  cbus__EVAL_95;
  wire  cbus__EVAL_96;
  wire [11:0] cbus__EVAL_97;
  wire  cbus__EVAL_98;
  wire [3:0] cbus__EVAL_99;
  wire [29:0] cbus__EVAL_100;
  wire [2:0] cbus__EVAL_101;
  wire [2:0] cbus__EVAL_102;
  wire  cbus__EVAL_103;
  wire  cbus__EVAL_104;
  wire [1:0] cbus__EVAL_105;
  wire  cbus__EVAL_106;
  wire  cbus__EVAL_107;
  wire [24:0] cbus__EVAL_108;
  wire [1:0] cbus__EVAL_109;
  wire  cbus__EVAL_110;
  wire  cbus__EVAL_111;
  wire [3:0] cbus__EVAL_112;
  wire [11:0] cbus__EVAL_113;
  wire [2:0] cbus__EVAL_114;
  wire [6:0] cbus__EVAL_115;
  wire  cbus__EVAL_116;
  wire  cbus__EVAL_117;
  wire [3:0] cbus__EVAL_118;
  wire  cbus__EVAL_119;
  wire [31:0] cbus__EVAL_120;
  wire  cbus__EVAL_121;
  wire  cbus__EVAL_122;
  wire [3:0] cbus__EVAL_123;
  wire  cbus__EVAL_124;
  wire [2:0] cbus__EVAL_125;
  wire [2:0] cbus__EVAL_126;
  wire [1:0] cbus__EVAL_127;
  wire  cbus__EVAL_128;
  wire  cbus__EVAL_129;
  wire  cbus__EVAL_130;
  wire  cbus__EVAL_131;
  wire [2:0] cbus__EVAL_132;
  wire [31:0] cbus__EVAL_133;
  wire [11:0] cbus__EVAL_134;
  wire  cbus__EVAL_135;
  wire  cbus__EVAL_136;
  wire [31:0] cbus__EVAL_137;
  wire [11:0] cbus__EVAL_138;
  wire  cbus__EVAL_139;
  wire [6:0] cbus__EVAL_140;
  wire [11:0] cbus__EVAL_141;
  wire  cbus__EVAL_142;
  wire  cbus__EVAL_143;
  wire [3:0] cbus__EVAL_144;
  wire [1:0] cbus__EVAL_145;
  wire  cbus__EVAL_146;
  wire [31:0] cbus__EVAL_147;
  wire [3:0] cbus__EVAL_148;
  wire  cbus__EVAL_149;
  wire  cbus__EVAL_150;
  wire  cbus__EVAL_151;
  wire [1:0] cbus__EVAL_152;
  wire  cbus__EVAL_153;
  wire  cbus__EVAL_154;
  wire [2:0] cbus__EVAL_155;
  wire [2:0] cbus__EVAL_156;
  wire [3:0] cbus__EVAL_157;
  wire  cbus__EVAL_158;
  wire [2:0] cbus__EVAL_159;
  wire [2:0] clint__EVAL;
  wire  clint__EVAL_0;
  wire [11:0] clint__EVAL_1;
  wire  clint__EVAL_2;
  wire  clint__EVAL_3;
  wire  clint__EVAL_4;
  wire [11:0] clint__EVAL_5;
  wire [1:0] clint__EVAL_6;
  wire  clint__EVAL_7;
  wire  clint__EVAL_8;
  wire [2:0] clint__EVAL_9;
  wire  clint__EVAL_10;
  wire  clint__EVAL_11;
  wire  clint__EVAL_12;
  wire [31:0] clint__EVAL_13;
  wire [31:0] clint__EVAL_14;
  wire [25:0] clint__EVAL_15;
  wire [2:0] clint__EVAL_16;
  wire [1:0] clint__EVAL_17;
  wire  clint__EVAL_18;
  wire [3:0] clint__EVAL_19;
  wire [2:0] shrinker__EVAL;
  wire [2:0] shrinker__EVAL_0;
  wire [2:0] shrinker__EVAL_1;
  wire  shrinker__EVAL_2;
  wire  shrinker__EVAL_3;
  wire  shrinker__EVAL_4;
  wire  shrinker__EVAL_5;
  wire  shrinker__EVAL_6;
  wire [8:0] shrinker__EVAL_7;
  wire  shrinker__EVAL_8;
  wire [7:0] shrinker__EVAL_9;
  wire [8:0] shrinker__EVAL_10;
  wire [63:0] shrinker__EVAL_11;
  wire [2:0] shrinker__EVAL_12;
  wire [2:0] shrinker__EVAL_13;
  wire  shrinker__EVAL_14;
  wire  shrinker__EVAL_15;
  wire  shrinker__EVAL_16;
  wire  shrinker__EVAL_17;
  wire [2:0] shrinker__EVAL_18;
  wire [63:0] shrinker__EVAL_19;
  wire [31:0] shrinker__EVAL_20;
  wire  shrinker__EVAL_21;
  wire [2:0] shrinker__EVAL_22;
  wire  shrinker__EVAL_23;
  wire  shrinker__EVAL_24;
  wire [2:0] shrinker__EVAL_25;
  wire [63:0] shrinker__EVAL_26;
  wire  shrinker__EVAL_27;
  wire [7:0] shrinker__EVAL_28;
  wire [63:0] shrinker__EVAL_29;
  wire [31:0] shrinker__EVAL_30;
  wire [2:0] shrinker__EVAL_31;
  wire [2:0] shrinker__EVAL_32;
  wire  shrinker__EVAL_33;
  wire  shrinker__EVAL_34;
  wire  shrinker__EVAL_35;
  wire  shrinker__EVAL_36;
  wire  testIndicator_clock;
  wire  testIndicator_reset;
  wire  testIndicator_auto_in_a_ready;
  wire  testIndicator_auto_in_a_valid;
  wire [2:0] testIndicator_auto_in_a_bits_opcode;
  wire [2:0] testIndicator_auto_in_a_bits_param;
  wire [1:0] testIndicator_auto_in_a_bits_size;
  wire [11:0] testIndicator_auto_in_a_bits_source;
  wire [14:0] testIndicator_auto_in_a_bits_address;
  wire [3:0] testIndicator_auto_in_a_bits_mask;
  wire [31:0] testIndicator_auto_in_a_bits_data;
  wire  testIndicator_auto_in_a_bits_corrupt;
  wire  testIndicator_auto_in_d_ready;
  wire  testIndicator_auto_in_d_valid;
  wire [2:0] testIndicator_auto_in_d_bits_opcode;
  wire [1:0] testIndicator_auto_in_d_bits_size;
  wire [11:0] testIndicator_auto_in_d_bits_source;
  wire [31:0] testIndicator_auto_in_d_bits_data;
  wire  intsource_1__EVAL;
  wire  intsource_1__EVAL_0;
  wire  intsource_1__EVAL_1;
  wire  intsource_1__EVAL_2;
  wire [63:0] bh__EVAL;
  wire  bh__EVAL_0;
  wire [31:0] bh__EVAL_1;
  wire [6:0] bh__EVAL_2;
  wire  bh__EVAL_3;
  wire [2:0] bh__EVAL_4;
  wire  bh__EVAL_5;
  wire [2:0] bh__EVAL_6;
  wire [63:0] bh__EVAL_7;
  wire [31:0] bh__EVAL_8;
  wire [8:0] bh__EVAL_9;
  wire  bh__EVAL_10;
  wire [2:0] bh__EVAL_11;
  wire [2:0] bh__EVAL_12;
  wire  bh__EVAL_13;
  wire [2:0] bh__EVAL_14;
  wire [2:0] bh__EVAL_15;
  wire  bh__EVAL_16;
  wire [2:0] bh__EVAL_17;
  wire  bh__EVAL_18;
  wire  bh__EVAL_19;
  wire [2:0] bh__EVAL_20;
  wire [6:0] bh__EVAL_21;
  wire  bh__EVAL_22;
  wire [2:0] bh__EVAL_23;
  wire  bh__EVAL_24;
  wire  bh__EVAL_25;
  wire [1:0] bh__EVAL_26;
  wire [63:0] bh__EVAL_27;
  wire [63:0] bh__EVAL_28;
  wire  bh__EVAL_29;
  wire [2:0] bh__EVAL_30;
  wire [31:0] bh__EVAL_31;
  wire [8:0] bh__EVAL_32;
  wire  bh__EVAL_33;
  wire  bh__EVAL_34;
  wire [2:0] bh__EVAL_35;
  wire [7:0] bh__EVAL_36;
  wire [2:0] bh__EVAL_37;
  wire  bh__EVAL_38;
  wire  bh__EVAL_39;
  wire  bh__EVAL_40;
  wire  bh__EVAL_41;
  wire  bh__EVAL_42;
  wire  bh__EVAL_43;
  wire [1:0] bh__EVAL_44;
  wire  bh__EVAL_45;
  wire [6:0] bh__EVAL_46;
  wire  bh__EVAL_47;
  wire [2:0] bh__EVAL_48;
  wire [7:0] bh__EVAL_49;
  wire [63:0] bh__EVAL_50;
  wire [31:0] bh__EVAL_51;
  wire  bh__EVAL_52;
  wire  bh__EVAL_53;
  wire  mbus__EVAL;
  wire  mbus__EVAL_0;
  wire  mbus__EVAL_1;
  wire  mbus__EVAL_2;
  wire [3:0] mbus__EVAL_3;
  wire [2:0] mbus__EVAL_4;
  wire [3:0] mbus__EVAL_5;
  wire  mbus__EVAL_6;
  wire  mbus__EVAL_7;
  wire  mbus__EVAL_8;
  wire  mbus__EVAL_9;
  wire [2:0] mbus__EVAL_10;
  wire [31:0] mbus__EVAL_11;
  wire  mbus__EVAL_12;
  wire [2:0] mbus__EVAL_13;
  wire  mbus__EVAL_14;
  wire [63:0] mbus__EVAL_15;
  wire [7:0] mbus__EVAL_16;
  wire [31:0] mbus__EVAL_17;
  wire  mbus__EVAL_18;
  wire [63:0] mbus__EVAL_19;
  wire [2:0] mbus__EVAL_20;
  wire  mbus__EVAL_21;
  wire [63:0] mbus__EVAL_22;
  wire [31:0] mbus__EVAL_23;
  wire [2:0] mbus__EVAL_24;
  wire  mbus__EVAL_25;
  wire  mbus__EVAL_26;
  wire [2:0] mbus__EVAL_27;
  wire [1:0] mbus__EVAL_28;
  wire [2:0] mbus__EVAL_29;
  wire [3:0] mbus__EVAL_30;
  wire  mbus__EVAL_31;
  wire [1:0] mbus__EVAL_32;
  wire  mbus__EVAL_33;
  wire  mbus__EVAL_34;
  wire  mbus__EVAL_35;
  wire [7:0] mbus__EVAL_36;
  wire  mbus__EVAL_37;
  wire [63:0] mbus__EVAL_38;
  wire  mbus__EVAL_39;
  wire [3:0] mbus__EVAL_40;
  wire [1:0] mbus__EVAL_41;
  wire [3:0] mbus__EVAL_42;
  wire [3:0] mbus__EVAL_43;
  wire [3:0] mbus__EVAL_44;
  wire  mbus__EVAL_45;
  wire  mbus__EVAL_46;
  wire  mbus__EVAL_47;
  wire [7:0] mbus__EVAL_48;
  wire [3:0] mbus__EVAL_49;
  wire [1:0] mbus__EVAL_50;
  wire [7:0] mbus__EVAL_51;
  wire  mbus__EVAL_52;
  wire  mbus__EVAL_53;
  wire [2:0] mbus__EVAL_54;
  wire [2:0] mbus__EVAL_55;
  wire  mbus__EVAL_56;
  reg  _EVAL_1;
  reg [31:0] _RAND_0;
  reg  _EVAL_4;
  reg [31:0] _RAND_1;
  wire  _EVAL_2;
  wire  _EVAL_3;
  wire  _EVAL;
  wire [1:0] _EVAL_0;
  SiFive__EVAL_278 SynchronizerShiftReg_w1_d3 (
    ._EVAL(SynchronizerShiftReg_w1_d3__EVAL),
    ._EVAL_0(SynchronizerShiftReg_w1_d3__EVAL_0),
    ._EVAL_1(SynchronizerShiftReg_w1_d3__EVAL_1)
  );
  SiFive__EVAL_218 dmiResetCatch (
    ._EVAL(dmiResetCatch__EVAL),
    ._EVAL_0(dmiResetCatch__EVAL_0),
    ._EVAL_1(dmiResetCatch__EVAL_1),
    ._EVAL_2(dmiResetCatch__EVAL_2),
    ._EVAL_3(dmiResetCatch__EVAL_3)
  );
  SiFive__EVAL_326 sagesafety (
    ._EVAL(sagesafety__EVAL),
    ._EVAL_0(sagesafety__EVAL_0),
    ._EVAL_1(sagesafety__EVAL_1),
    ._EVAL_2(sagesafety__EVAL_2),
    ._EVAL_3(sagesafety__EVAL_3),
    ._EVAL_4(sagesafety__EVAL_4),
    ._EVAL_5(sagesafety__EVAL_5),
    ._EVAL_6(sagesafety__EVAL_6),
    ._EVAL_7(sagesafety__EVAL_7),
    ._EVAL_8(sagesafety__EVAL_8),
    ._EVAL_9(sagesafety__EVAL_9),
    ._EVAL_10(sagesafety__EVAL_10),
    ._EVAL_11(sagesafety__EVAL_11),
    ._EVAL_12(sagesafety__EVAL_12),
    ._EVAL_13(sagesafety__EVAL_13),
    ._EVAL_14(sagesafety__EVAL_14),
    ._EVAL_15(sagesafety__EVAL_15),
    ._EVAL_16(sagesafety__EVAL_16),
    ._EVAL_17(sagesafety__EVAL_17),
    ._EVAL_18(sagesafety__EVAL_18),
    ._EVAL_19(sagesafety__EVAL_19),
    ._EVAL_20(sagesafety__EVAL_20),
    ._EVAL_21(sagesafety__EVAL_21),
    ._EVAL_22(sagesafety__EVAL_22),
    ._EVAL_23(sagesafety__EVAL_23),
    ._EVAL_24(sagesafety__EVAL_24),
    ._EVAL_25(sagesafety__EVAL_25),
    ._EVAL_26(sagesafety__EVAL_26),
    ._EVAL_27(sagesafety__EVAL_27),
    ._EVAL_28(sagesafety__EVAL_28),
    ._EVAL_29(sagesafety__EVAL_29),
    ._EVAL_30(sagesafety__EVAL_30),
    ._EVAL_31(sagesafety__EVAL_31),
    ._EVAL_32(sagesafety__EVAL_32),
    ._EVAL_33(sagesafety__EVAL_33),
    ._EVAL_34(sagesafety__EVAL_34),
    ._EVAL_35(sagesafety__EVAL_35),
    ._EVAL_36(sagesafety__EVAL_36),
    ._EVAL_37(sagesafety__EVAL_37),
    ._EVAL_38(sagesafety__EVAL_38),
    ._EVAL_39(sagesafety__EVAL_39),
    ._EVAL_40(sagesafety__EVAL_40)
  );
  SiFive__EVAL_335 dtm (
    ._EVAL(dtm__EVAL),
    ._EVAL_0(dtm__EVAL_0),
    ._EVAL_1(dtm__EVAL_1),
    ._EVAL_2(dtm__EVAL_2),
    ._EVAL_3(dtm__EVAL_3),
    ._EVAL_4(dtm__EVAL_4),
    ._EVAL_5(dtm__EVAL_5),
    ._EVAL_6(dtm__EVAL_6),
    ._EVAL_7(dtm__EVAL_7),
    ._EVAL_8(dtm__EVAL_8),
    ._EVAL_9(dtm__EVAL_9),
    ._EVAL_10(dtm__EVAL_10),
    ._EVAL_11(dtm__EVAL_11),
    ._EVAL_12(dtm__EVAL_12),
    ._EVAL_13(dtm__EVAL_13),
    ._EVAL_14(dtm__EVAL_14),
    ._EVAL_15(dtm__EVAL_15),
    ._EVAL_16(dtm__EVAL_16)
  );
  SiFive__EVAL_310 tile (
    ._EVAL(tile__EVAL),
    ._EVAL_0(tile__EVAL_0),
    ._EVAL_1(tile__EVAL_1),
    ._EVAL_2(tile__EVAL_2),
    ._EVAL_3(tile__EVAL_3),
    ._EVAL_4(tile__EVAL_4),
    ._EVAL_5(tile__EVAL_5),
    ._EVAL_6(tile__EVAL_6),
    ._EVAL_7(tile__EVAL_7),
    ._EVAL_8(tile__EVAL_8),
    ._EVAL_9(tile__EVAL_9),
    ._EVAL_10(tile__EVAL_10),
    ._EVAL_11(tile__EVAL_11),
    ._EVAL_12(tile__EVAL_12),
    ._EVAL_13(tile__EVAL_13),
    ._EVAL_14(tile__EVAL_14),
    ._EVAL_15(tile__EVAL_15),
    ._EVAL_16(tile__EVAL_16),
    ._EVAL_17(tile__EVAL_17),
    ._EVAL_18(tile__EVAL_18),
    ._EVAL_19(tile__EVAL_19),
    ._EVAL_20(tile__EVAL_20),
    ._EVAL_21(tile__EVAL_21),
    ._EVAL_22(tile__EVAL_22),
    ._EVAL_23(tile__EVAL_23),
    ._EVAL_24(tile__EVAL_24),
    ._EVAL_25(tile__EVAL_25),
    ._EVAL_26(tile__EVAL_26),
    ._EVAL_27(tile__EVAL_27),
    ._EVAL_28(tile__EVAL_28),
    ._EVAL_29(tile__EVAL_29),
    ._EVAL_30(tile__EVAL_30),
    ._EVAL_31(tile__EVAL_31),
    ._EVAL_32(tile__EVAL_32),
    ._EVAL_33(tile__EVAL_33),
    ._EVAL_34(tile__EVAL_34),
    ._EVAL_35(tile__EVAL_35),
    ._EVAL_36(tile__EVAL_36),
    ._EVAL_37(tile__EVAL_37),
    ._EVAL_38(tile__EVAL_38),
    ._EVAL_39(tile__EVAL_39),
    ._EVAL_40(tile__EVAL_40),
    ._EVAL_41(tile__EVAL_41),
    ._EVAL_42(tile__EVAL_42),
    ._EVAL_43(tile__EVAL_43),
    ._EVAL_44(tile__EVAL_44),
    ._EVAL_45(tile__EVAL_45),
    ._EVAL_46(tile__EVAL_46),
    ._EVAL_47(tile__EVAL_47),
    ._EVAL_48(tile__EVAL_48),
    ._EVAL_49(tile__EVAL_49),
    ._EVAL_50(tile__EVAL_50),
    ._EVAL_51(tile__EVAL_51),
    ._EVAL_52(tile__EVAL_52),
    ._EVAL_53(tile__EVAL_53),
    ._EVAL_54(tile__EVAL_54),
    ._EVAL_55(tile__EVAL_55),
    ._EVAL_56(tile__EVAL_56),
    ._EVAL_57(tile__EVAL_57),
    ._EVAL_58(tile__EVAL_58),
    ._EVAL_59(tile__EVAL_59),
    ._EVAL_60(tile__EVAL_60),
    ._EVAL_61(tile__EVAL_61),
    ._EVAL_62(tile__EVAL_62),
    ._EVAL_63(tile__EVAL_63),
    ._EVAL_64(tile__EVAL_64),
    ._EVAL_65(tile__EVAL_65),
    ._EVAL_66(tile__EVAL_66),
    ._EVAL_67(tile__EVAL_67),
    ._EVAL_68(tile__EVAL_68),
    ._EVAL_69(tile__EVAL_69),
    ._EVAL_70(tile__EVAL_70),
    ._EVAL_71(tile__EVAL_71),
    ._EVAL_72(tile__EVAL_72),
    ._EVAL_73(tile__EVAL_73),
    ._EVAL_74(tile__EVAL_74),
    ._EVAL_75(tile__EVAL_75),
    ._EVAL_76(tile__EVAL_76),
    ._EVAL_77(tile__EVAL_77),
    ._EVAL_78(tile__EVAL_78),
    ._EVAL_79(tile__EVAL_79),
    ._EVAL_80(tile__EVAL_80),
    ._EVAL_81(tile__EVAL_81),
    ._EVAL_82(tile__EVAL_82),
    ._EVAL_83(tile__EVAL_83),
    ._EVAL_84(tile__EVAL_84),
    ._EVAL_85(tile__EVAL_85),
    ._EVAL_86(tile__EVAL_86),
    ._EVAL_87(tile__EVAL_87),
    ._EVAL_88(tile__EVAL_88),
    ._EVAL_89(tile__EVAL_89),
    ._EVAL_90(tile__EVAL_90),
    ._EVAL_91(tile__EVAL_91),
    ._EVAL_92(tile__EVAL_92),
    ._EVAL_93(tile__EVAL_93),
    ._EVAL_94(tile__EVAL_94),
    ._EVAL_95(tile__EVAL_95),
    ._EVAL_96(tile__EVAL_96),
    ._EVAL_97(tile__EVAL_97),
    ._EVAL_98(tile__EVAL_98),
    ._EVAL_99(tile__EVAL_99),
    ._EVAL_100(tile__EVAL_100),
    ._EVAL_101(tile__EVAL_101),
    ._EVAL_102(tile__EVAL_102),
    ._EVAL_103(tile__EVAL_103),
    ._EVAL_104(tile__EVAL_104),
    ._EVAL_105(tile__EVAL_105),
    ._EVAL_106(tile__EVAL_106),
    ._EVAL_107(tile__EVAL_107),
    ._EVAL_108(tile__EVAL_108),
    ._EVAL_109(tile__EVAL_109),
    ._EVAL_110(tile__EVAL_110),
    ._EVAL_111(tile__EVAL_111),
    ._EVAL_112(tile__EVAL_112),
    ._EVAL_113(tile__EVAL_113),
    ._EVAL_114(tile__EVAL_114),
    ._EVAL_115(tile__EVAL_115),
    ._EVAL_116(tile__EVAL_116),
    ._EVAL_117(tile__EVAL_117),
    ._EVAL_118(tile__EVAL_118)
  );
  SiFive__EVAL_185 plic (
    ._EVAL(plic__EVAL),
    ._EVAL_0(plic__EVAL_0),
    ._EVAL_1(plic__EVAL_1),
    ._EVAL_2(plic__EVAL_2),
    ._EVAL_3(plic__EVAL_3),
    ._EVAL_4(plic__EVAL_4),
    ._EVAL_5(plic__EVAL_5),
    ._EVAL_6(plic__EVAL_6),
    ._EVAL_7(plic__EVAL_7),
    ._EVAL_8(plic__EVAL_8),
    ._EVAL_9(plic__EVAL_9),
    ._EVAL_10(plic__EVAL_10),
    ._EVAL_11(plic__EVAL_11),
    ._EVAL_12(plic__EVAL_12),
    ._EVAL_13(plic__EVAL_13),
    ._EVAL_14(plic__EVAL_14),
    ._EVAL_15(plic__EVAL_15),
    ._EVAL_16(plic__EVAL_16),
    ._EVAL_17(plic__EVAL_17),
    ._EVAL_18(plic__EVAL_18),
    ._EVAL_19(plic__EVAL_19),
    ._EVAL_20(plic__EVAL_20),
    ._EVAL_21(plic__EVAL_21),
    ._EVAL_22(plic__EVAL_22),
    ._EVAL_23(plic__EVAL_23),
    ._EVAL_24(plic__EVAL_24),
    ._EVAL_25(plic__EVAL_25),
    ._EVAL_26(plic__EVAL_26),
    ._EVAL_27(plic__EVAL_27),
    ._EVAL_28(plic__EVAL_28),
    ._EVAL_29(plic__EVAL_29),
    ._EVAL_30(plic__EVAL_30),
    ._EVAL_31(plic__EVAL_31),
    ._EVAL_32(plic__EVAL_32),
    ._EVAL_33(plic__EVAL_33),
    ._EVAL_34(plic__EVAL_34),
    ._EVAL_35(plic__EVAL_35),
    ._EVAL_36(plic__EVAL_36),
    ._EVAL_37(plic__EVAL_37),
    ._EVAL_38(plic__EVAL_38),
    ._EVAL_39(plic__EVAL_39),
    ._EVAL_40(plic__EVAL_40),
    ._EVAL_41(plic__EVAL_41),
    ._EVAL_42(plic__EVAL_42),
    ._EVAL_43(plic__EVAL_43),
    ._EVAL_44(plic__EVAL_44),
    ._EVAL_45(plic__EVAL_45),
    ._EVAL_46(plic__EVAL_46),
    ._EVAL_47(plic__EVAL_47),
    ._EVAL_48(plic__EVAL_48),
    ._EVAL_49(plic__EVAL_49),
    ._EVAL_50(plic__EVAL_50),
    ._EVAL_51(plic__EVAL_51),
    ._EVAL_52(plic__EVAL_52),
    ._EVAL_53(plic__EVAL_53),
    ._EVAL_54(plic__EVAL_54),
    ._EVAL_55(plic__EVAL_55),
    ._EVAL_56(plic__EVAL_56),
    ._EVAL_57(plic__EVAL_57),
    ._EVAL_58(plic__EVAL_58),
    ._EVAL_59(plic__EVAL_59),
    ._EVAL_60(plic__EVAL_60),
    ._EVAL_61(plic__EVAL_61),
    ._EVAL_62(plic__EVAL_62),
    ._EVAL_63(plic__EVAL_63),
    ._EVAL_64(plic__EVAL_64),
    ._EVAL_65(plic__EVAL_65),
    ._EVAL_66(plic__EVAL_66),
    ._EVAL_67(plic__EVAL_67),
    ._EVAL_68(plic__EVAL_68),
    ._EVAL_69(plic__EVAL_69),
    ._EVAL_70(plic__EVAL_70),
    ._EVAL_71(plic__EVAL_71),
    ._EVAL_72(plic__EVAL_72),
    ._EVAL_73(plic__EVAL_73),
    ._EVAL_74(plic__EVAL_74),
    ._EVAL_75(plic__EVAL_75),
    ._EVAL_76(plic__EVAL_76),
    ._EVAL_77(plic__EVAL_77),
    ._EVAL_78(plic__EVAL_78),
    ._EVAL_79(plic__EVAL_79),
    ._EVAL_80(plic__EVAL_80),
    ._EVAL_81(plic__EVAL_81),
    ._EVAL_82(plic__EVAL_82),
    ._EVAL_83(plic__EVAL_83),
    ._EVAL_84(plic__EVAL_84),
    ._EVAL_85(plic__EVAL_85),
    ._EVAL_86(plic__EVAL_86),
    ._EVAL_87(plic__EVAL_87),
    ._EVAL_88(plic__EVAL_88),
    ._EVAL_89(plic__EVAL_89),
    ._EVAL_90(plic__EVAL_90),
    ._EVAL_91(plic__EVAL_91),
    ._EVAL_92(plic__EVAL_92),
    ._EVAL_93(plic__EVAL_93),
    ._EVAL_94(plic__EVAL_94),
    ._EVAL_95(plic__EVAL_95),
    ._EVAL_96(plic__EVAL_96),
    ._EVAL_97(plic__EVAL_97),
    ._EVAL_98(plic__EVAL_98),
    ._EVAL_99(plic__EVAL_99),
    ._EVAL_100(plic__EVAL_100),
    ._EVAL_101(plic__EVAL_101),
    ._EVAL_102(plic__EVAL_102),
    ._EVAL_103(plic__EVAL_103),
    ._EVAL_104(plic__EVAL_104),
    ._EVAL_105(plic__EVAL_105),
    ._EVAL_106(plic__EVAL_106),
    ._EVAL_107(plic__EVAL_107),
    ._EVAL_108(plic__EVAL_108),
    ._EVAL_109(plic__EVAL_109),
    ._EVAL_110(plic__EVAL_110),
    ._EVAL_111(plic__EVAL_111),
    ._EVAL_112(plic__EVAL_112),
    ._EVAL_113(plic__EVAL_113),
    ._EVAL_114(plic__EVAL_114),
    ._EVAL_115(plic__EVAL_115),
    ._EVAL_116(plic__EVAL_116),
    ._EVAL_117(plic__EVAL_117),
    ._EVAL_118(plic__EVAL_118),
    ._EVAL_119(plic__EVAL_119),
    ._EVAL_120(plic__EVAL_120),
    ._EVAL_121(plic__EVAL_121),
    ._EVAL_122(plic__EVAL_122),
    ._EVAL_123(plic__EVAL_123),
    ._EVAL_124(plic__EVAL_124),
    ._EVAL_125(plic__EVAL_125),
    ._EVAL_126(plic__EVAL_126),
    ._EVAL_127(plic__EVAL_127),
    ._EVAL_128(plic__EVAL_128),
    ._EVAL_129(plic__EVAL_129),
    ._EVAL_130(plic__EVAL_130),
    ._EVAL_131(plic__EVAL_131),
    ._EVAL_132(plic__EVAL_132),
    ._EVAL_133(plic__EVAL_133),
    ._EVAL_134(plic__EVAL_134),
    ._EVAL_135(plic__EVAL_135),
    ._EVAL_136(plic__EVAL_136),
    ._EVAL_137(plic__EVAL_137),
    ._EVAL_138(plic__EVAL_138),
    ._EVAL_139(plic__EVAL_139),
    ._EVAL_140(plic__EVAL_140),
    ._EVAL_141(plic__EVAL_141),
    ._EVAL_142(plic__EVAL_142),
    ._EVAL_143(plic__EVAL_143),
    ._EVAL_144(plic__EVAL_144)
  );
  SiFive__EVAL_322 ww (
    ._EVAL(ww__EVAL),
    ._EVAL_0(ww__EVAL_0),
    ._EVAL_1(ww__EVAL_1),
    ._EVAL_2(ww__EVAL_2),
    ._EVAL_3(ww__EVAL_3),
    ._EVAL_4(ww__EVAL_4),
    ._EVAL_5(ww__EVAL_5),
    ._EVAL_6(ww__EVAL_6),
    ._EVAL_7(ww__EVAL_7),
    ._EVAL_8(ww__EVAL_8),
    ._EVAL_9(ww__EVAL_9),
    ._EVAL_10(ww__EVAL_10),
    ._EVAL_11(ww__EVAL_11),
    ._EVAL_12(ww__EVAL_12),
    ._EVAL_13(ww__EVAL_13),
    ._EVAL_14(ww__EVAL_14),
    ._EVAL_15(ww__EVAL_15),
    ._EVAL_16(ww__EVAL_16),
    ._EVAL_17(ww__EVAL_17),
    ._EVAL_18(ww__EVAL_18),
    ._EVAL_19(ww__EVAL_19),
    ._EVAL_20(ww__EVAL_20),
    ._EVAL_21(ww__EVAL_21),
    ._EVAL_22(ww__EVAL_22),
    ._EVAL_23(ww__EVAL_23),
    ._EVAL_24(ww__EVAL_24),
    ._EVAL_25(ww__EVAL_25),
    ._EVAL_26(ww__EVAL_26),
    ._EVAL_27(ww__EVAL_27),
    ._EVAL_28(ww__EVAL_28),
    ._EVAL_29(ww__EVAL_29),
    ._EVAL_30(ww__EVAL_30),
    ._EVAL_31(ww__EVAL_31),
    ._EVAL_32(ww__EVAL_32),
    ._EVAL_33(ww__EVAL_33),
    ._EVAL_34(ww__EVAL_34),
    ._EVAL_35(ww__EVAL_35),
    ._EVAL_36(ww__EVAL_36)
  );
  SiFive__EVAL_49 sbus (
    ._EVAL(sbus__EVAL),
    ._EVAL_0(sbus__EVAL_0),
    ._EVAL_1(sbus__EVAL_1),
    ._EVAL_2(sbus__EVAL_2),
    ._EVAL_3(sbus__EVAL_3),
    ._EVAL_4(sbus__EVAL_4),
    ._EVAL_5(sbus__EVAL_5),
    ._EVAL_6(sbus__EVAL_6),
    ._EVAL_7(sbus__EVAL_7),
    ._EVAL_8(sbus__EVAL_8),
    ._EVAL_9(sbus__EVAL_9),
    ._EVAL_10(sbus__EVAL_10),
    ._EVAL_11(sbus__EVAL_11),
    ._EVAL_12(sbus__EVAL_12),
    ._EVAL_13(sbus__EVAL_13),
    ._EVAL_14(sbus__EVAL_14),
    ._EVAL_15(sbus__EVAL_15),
    ._EVAL_16(sbus__EVAL_16),
    ._EVAL_17(sbus__EVAL_17),
    ._EVAL_18(sbus__EVAL_18),
    ._EVAL_19(sbus__EVAL_19),
    ._EVAL_20(sbus__EVAL_20),
    ._EVAL_21(sbus__EVAL_21),
    ._EVAL_22(sbus__EVAL_22),
    ._EVAL_23(sbus__EVAL_23),
    ._EVAL_24(sbus__EVAL_24),
    ._EVAL_25(sbus__EVAL_25),
    ._EVAL_26(sbus__EVAL_26),
    ._EVAL_27(sbus__EVAL_27),
    ._EVAL_28(sbus__EVAL_28),
    ._EVAL_29(sbus__EVAL_29),
    ._EVAL_30(sbus__EVAL_30),
    ._EVAL_31(sbus__EVAL_31),
    ._EVAL_32(sbus__EVAL_32),
    ._EVAL_33(sbus__EVAL_33),
    ._EVAL_34(sbus__EVAL_34),
    ._EVAL_35(sbus__EVAL_35),
    ._EVAL_36(sbus__EVAL_36),
    ._EVAL_37(sbus__EVAL_37),
    ._EVAL_38(sbus__EVAL_38),
    ._EVAL_39(sbus__EVAL_39),
    ._EVAL_40(sbus__EVAL_40),
    ._EVAL_41(sbus__EVAL_41),
    ._EVAL_42(sbus__EVAL_42),
    ._EVAL_43(sbus__EVAL_43),
    ._EVAL_44(sbus__EVAL_44),
    ._EVAL_45(sbus__EVAL_45),
    ._EVAL_46(sbus__EVAL_46),
    ._EVAL_47(sbus__EVAL_47),
    ._EVAL_48(sbus__EVAL_48),
    ._EVAL_49(sbus__EVAL_49),
    ._EVAL_50(sbus__EVAL_50),
    ._EVAL_51(sbus__EVAL_51),
    ._EVAL_52(sbus__EVAL_52),
    ._EVAL_53(sbus__EVAL_53),
    ._EVAL_54(sbus__EVAL_54),
    ._EVAL_55(sbus__EVAL_55),
    ._EVAL_56(sbus__EVAL_56),
    ._EVAL_57(sbus__EVAL_57),
    ._EVAL_58(sbus__EVAL_58),
    ._EVAL_59(sbus__EVAL_59),
    ._EVAL_60(sbus__EVAL_60),
    ._EVAL_61(sbus__EVAL_61),
    ._EVAL_62(sbus__EVAL_62),
    ._EVAL_63(sbus__EVAL_63),
    ._EVAL_64(sbus__EVAL_64),
    ._EVAL_65(sbus__EVAL_65),
    ._EVAL_66(sbus__EVAL_66),
    ._EVAL_67(sbus__EVAL_67),
    ._EVAL_68(sbus__EVAL_68),
    ._EVAL_69(sbus__EVAL_69),
    ._EVAL_70(sbus__EVAL_70),
    ._EVAL_71(sbus__EVAL_71),
    ._EVAL_72(sbus__EVAL_72),
    ._EVAL_73(sbus__EVAL_73),
    ._EVAL_74(sbus__EVAL_74),
    ._EVAL_75(sbus__EVAL_75),
    ._EVAL_76(sbus__EVAL_76),
    ._EVAL_77(sbus__EVAL_77),
    ._EVAL_78(sbus__EVAL_78),
    ._EVAL_79(sbus__EVAL_79),
    ._EVAL_80(sbus__EVAL_80),
    ._EVAL_81(sbus__EVAL_81),
    ._EVAL_82(sbus__EVAL_82),
    ._EVAL_83(sbus__EVAL_83),
    ._EVAL_84(sbus__EVAL_84),
    ._EVAL_85(sbus__EVAL_85),
    ._EVAL_86(sbus__EVAL_86),
    ._EVAL_87(sbus__EVAL_87),
    ._EVAL_88(sbus__EVAL_88),
    ._EVAL_89(sbus__EVAL_89),
    ._EVAL_90(sbus__EVAL_90),
    ._EVAL_91(sbus__EVAL_91),
    ._EVAL_92(sbus__EVAL_92),
    ._EVAL_93(sbus__EVAL_93),
    ._EVAL_94(sbus__EVAL_94),
    ._EVAL_95(sbus__EVAL_95),
    ._EVAL_96(sbus__EVAL_96),
    ._EVAL_97(sbus__EVAL_97),
    ._EVAL_98(sbus__EVAL_98),
    ._EVAL_99(sbus__EVAL_99),
    ._EVAL_100(sbus__EVAL_100),
    ._EVAL_101(sbus__EVAL_101),
    ._EVAL_102(sbus__EVAL_102),
    ._EVAL_103(sbus__EVAL_103),
    ._EVAL_104(sbus__EVAL_104),
    ._EVAL_105(sbus__EVAL_105),
    ._EVAL_106(sbus__EVAL_106),
    ._EVAL_107(sbus__EVAL_107),
    ._EVAL_108(sbus__EVAL_108),
    ._EVAL_109(sbus__EVAL_109),
    ._EVAL_110(sbus__EVAL_110),
    ._EVAL_111(sbus__EVAL_111),
    ._EVAL_112(sbus__EVAL_112),
    ._EVAL_113(sbus__EVAL_113),
    ._EVAL_114(sbus__EVAL_114),
    ._EVAL_115(sbus__EVAL_115),
    ._EVAL_116(sbus__EVAL_116),
    ._EVAL_117(sbus__EVAL_117),
    ._EVAL_118(sbus__EVAL_118),
    ._EVAL_119(sbus__EVAL_119),
    ._EVAL_120(sbus__EVAL_120),
    ._EVAL_121(sbus__EVAL_121),
    ._EVAL_122(sbus__EVAL_122),
    ._EVAL_123(sbus__EVAL_123),
    ._EVAL_124(sbus__EVAL_124),
    ._EVAL_125(sbus__EVAL_125),
    ._EVAL_126(sbus__EVAL_126),
    ._EVAL_127(sbus__EVAL_127),
    ._EVAL_128(sbus__EVAL_128),
    ._EVAL_129(sbus__EVAL_129),
    ._EVAL_130(sbus__EVAL_130),
    ._EVAL_131(sbus__EVAL_131),
    ._EVAL_132(sbus__EVAL_132),
    ._EVAL_133(sbus__EVAL_133),
    ._EVAL_134(sbus__EVAL_134),
    ._EVAL_135(sbus__EVAL_135),
    ._EVAL_136(sbus__EVAL_136),
    ._EVAL_137(sbus__EVAL_137),
    ._EVAL_138(sbus__EVAL_138),
    ._EVAL_139(sbus__EVAL_139),
    ._EVAL_140(sbus__EVAL_140),
    ._EVAL_141(sbus__EVAL_141),
    ._EVAL_142(sbus__EVAL_142),
    ._EVAL_143(sbus__EVAL_143),
    ._EVAL_144(sbus__EVAL_144),
    ._EVAL_145(sbus__EVAL_145),
    ._EVAL_146(sbus__EVAL_146),
    ._EVAL_147(sbus__EVAL_147),
    ._EVAL_148(sbus__EVAL_148),
    ._EVAL_149(sbus__EVAL_149),
    ._EVAL_150(sbus__EVAL_150),
    ._EVAL_151(sbus__EVAL_151),
    ._EVAL_152(sbus__EVAL_152),
    ._EVAL_153(sbus__EVAL_153),
    ._EVAL_154(sbus__EVAL_154),
    ._EVAL_155(sbus__EVAL_155),
    ._EVAL_156(sbus__EVAL_156),
    ._EVAL_157(sbus__EVAL_157),
    ._EVAL_158(sbus__EVAL_158),
    ._EVAL_159(sbus__EVAL_159),
    ._EVAL_160(sbus__EVAL_160),
    ._EVAL_161(sbus__EVAL_161),
    ._EVAL_162(sbus__EVAL_162),
    ._EVAL_163(sbus__EVAL_163),
    ._EVAL_164(sbus__EVAL_164),
    ._EVAL_165(sbus__EVAL_165),
    ._EVAL_166(sbus__EVAL_166),
    ._EVAL_167(sbus__EVAL_167),
    ._EVAL_168(sbus__EVAL_168),
    ._EVAL_169(sbus__EVAL_169),
    ._EVAL_170(sbus__EVAL_170),
    ._EVAL_171(sbus__EVAL_171),
    ._EVAL_172(sbus__EVAL_172),
    ._EVAL_173(sbus__EVAL_173),
    ._EVAL_174(sbus__EVAL_174),
    ._EVAL_175(sbus__EVAL_175),
    ._EVAL_176(sbus__EVAL_176),
    ._EVAL_177(sbus__EVAL_177),
    ._EVAL_178(sbus__EVAL_178),
    ._EVAL_179(sbus__EVAL_179),
    ._EVAL_180(sbus__EVAL_180),
    ._EVAL_181(sbus__EVAL_181),
    ._EVAL_182(sbus__EVAL_182),
    ._EVAL_183(sbus__EVAL_183),
    ._EVAL_184(sbus__EVAL_184),
    ._EVAL_185(sbus__EVAL_185),
    ._EVAL_186(sbus__EVAL_186),
    ._EVAL_187(sbus__EVAL_187),
    ._EVAL_188(sbus__EVAL_188),
    ._EVAL_189(sbus__EVAL_189),
    ._EVAL_190(sbus__EVAL_190),
    ._EVAL_191(sbus__EVAL_191),
    ._EVAL_192(sbus__EVAL_192),
    ._EVAL_193(sbus__EVAL_193),
    ._EVAL_194(sbus__EVAL_194),
    ._EVAL_195(sbus__EVAL_195),
    ._EVAL_196(sbus__EVAL_196),
    ._EVAL_197(sbus__EVAL_197),
    ._EVAL_198(sbus__EVAL_198),
    ._EVAL_199(sbus__EVAL_199),
    ._EVAL_200(sbus__EVAL_200),
    ._EVAL_201(sbus__EVAL_201),
    ._EVAL_202(sbus__EVAL_202),
    ._EVAL_203(sbus__EVAL_203),
    ._EVAL_204(sbus__EVAL_204),
    ._EVAL_205(sbus__EVAL_205),
    ._EVAL_206(sbus__EVAL_206),
    ._EVAL_207(sbus__EVAL_207),
    ._EVAL_208(sbus__EVAL_208),
    ._EVAL_209(sbus__EVAL_209),
    ._EVAL_210(sbus__EVAL_210),
    ._EVAL_211(sbus__EVAL_211),
    ._EVAL_212(sbus__EVAL_212),
    ._EVAL_213(sbus__EVAL_213),
    ._EVAL_214(sbus__EVAL_214),
    ._EVAL_215(sbus__EVAL_215),
    ._EVAL_216(sbus__EVAL_216),
    ._EVAL_217(sbus__EVAL_217),
    ._EVAL_218(sbus__EVAL_218),
    ._EVAL_219(sbus__EVAL_219),
    ._EVAL_220(sbus__EVAL_220),
    ._EVAL_221(sbus__EVAL_221),
    ._EVAL_222(sbus__EVAL_222),
    ._EVAL_223(sbus__EVAL_223),
    ._EVAL_224(sbus__EVAL_224)
  );
  SiFive__EVAL int_bus (
    ._EVAL(int_bus__EVAL),
    ._EVAL_0(int_bus__EVAL_0),
    ._EVAL_1(int_bus__EVAL_1),
    ._EVAL_2(int_bus__EVAL_2),
    ._EVAL_3(int_bus__EVAL_3),
    ._EVAL_4(int_bus__EVAL_4),
    ._EVAL_5(int_bus__EVAL_5),
    ._EVAL_6(int_bus__EVAL_6),
    ._EVAL_7(int_bus__EVAL_7),
    ._EVAL_8(int_bus__EVAL_8),
    ._EVAL_9(int_bus__EVAL_9),
    ._EVAL_10(int_bus__EVAL_10),
    ._EVAL_11(int_bus__EVAL_11),
    ._EVAL_12(int_bus__EVAL_12),
    ._EVAL_13(int_bus__EVAL_13),
    ._EVAL_14(int_bus__EVAL_14),
    ._EVAL_15(int_bus__EVAL_15),
    ._EVAL_16(int_bus__EVAL_16),
    ._EVAL_17(int_bus__EVAL_17),
    ._EVAL_18(int_bus__EVAL_18),
    ._EVAL_19(int_bus__EVAL_19),
    ._EVAL_20(int_bus__EVAL_20),
    ._EVAL_21(int_bus__EVAL_21),
    ._EVAL_22(int_bus__EVAL_22),
    ._EVAL_23(int_bus__EVAL_23),
    ._EVAL_24(int_bus__EVAL_24),
    ._EVAL_25(int_bus__EVAL_25),
    ._EVAL_26(int_bus__EVAL_26),
    ._EVAL_27(int_bus__EVAL_27),
    ._EVAL_28(int_bus__EVAL_28),
    ._EVAL_29(int_bus__EVAL_29),
    ._EVAL_30(int_bus__EVAL_30),
    ._EVAL_31(int_bus__EVAL_31),
    ._EVAL_32(int_bus__EVAL_32),
    ._EVAL_33(int_bus__EVAL_33),
    ._EVAL_34(int_bus__EVAL_34),
    ._EVAL_35(int_bus__EVAL_35),
    ._EVAL_36(int_bus__EVAL_36),
    ._EVAL_37(int_bus__EVAL_37),
    ._EVAL_38(int_bus__EVAL_38),
    ._EVAL_39(int_bus__EVAL_39),
    ._EVAL_40(int_bus__EVAL_40),
    ._EVAL_41(int_bus__EVAL_41),
    ._EVAL_42(int_bus__EVAL_42),
    ._EVAL_43(int_bus__EVAL_43),
    ._EVAL_44(int_bus__EVAL_44),
    ._EVAL_45(int_bus__EVAL_45),
    ._EVAL_46(int_bus__EVAL_46),
    ._EVAL_47(int_bus__EVAL_47),
    ._EVAL_48(int_bus__EVAL_48),
    ._EVAL_49(int_bus__EVAL_49),
    ._EVAL_50(int_bus__EVAL_50),
    ._EVAL_51(int_bus__EVAL_51),
    ._EVAL_52(int_bus__EVAL_52),
    ._EVAL_53(int_bus__EVAL_53),
    ._EVAL_54(int_bus__EVAL_54),
    ._EVAL_55(int_bus__EVAL_55),
    ._EVAL_56(int_bus__EVAL_56),
    ._EVAL_57(int_bus__EVAL_57),
    ._EVAL_58(int_bus__EVAL_58),
    ._EVAL_59(int_bus__EVAL_59),
    ._EVAL_60(int_bus__EVAL_60),
    ._EVAL_61(int_bus__EVAL_61),
    ._EVAL_62(int_bus__EVAL_62),
    ._EVAL_63(int_bus__EVAL_63),
    ._EVAL_64(int_bus__EVAL_64),
    ._EVAL_65(int_bus__EVAL_65),
    ._EVAL_66(int_bus__EVAL_66),
    ._EVAL_67(int_bus__EVAL_67),
    ._EVAL_68(int_bus__EVAL_68),
    ._EVAL_69(int_bus__EVAL_69),
    ._EVAL_70(int_bus__EVAL_70),
    ._EVAL_71(int_bus__EVAL_71),
    ._EVAL_72(int_bus__EVAL_72),
    ._EVAL_73(int_bus__EVAL_73),
    ._EVAL_74(int_bus__EVAL_74),
    ._EVAL_75(int_bus__EVAL_75),
    ._EVAL_76(int_bus__EVAL_76),
    ._EVAL_77(int_bus__EVAL_77),
    ._EVAL_78(int_bus__EVAL_78),
    ._EVAL_79(int_bus__EVAL_79),
    ._EVAL_80(int_bus__EVAL_80),
    ._EVAL_81(int_bus__EVAL_81),
    ._EVAL_82(int_bus__EVAL_82),
    ._EVAL_83(int_bus__EVAL_83),
    ._EVAL_84(int_bus__EVAL_84),
    ._EVAL_85(int_bus__EVAL_85),
    ._EVAL_86(int_bus__EVAL_86),
    ._EVAL_87(int_bus__EVAL_87),
    ._EVAL_88(int_bus__EVAL_88),
    ._EVAL_89(int_bus__EVAL_89),
    ._EVAL_90(int_bus__EVAL_90),
    ._EVAL_91(int_bus__EVAL_91),
    ._EVAL_92(int_bus__EVAL_92),
    ._EVAL_93(int_bus__EVAL_93),
    ._EVAL_94(int_bus__EVAL_94),
    ._EVAL_95(int_bus__EVAL_95),
    ._EVAL_96(int_bus__EVAL_96),
    ._EVAL_97(int_bus__EVAL_97),
    ._EVAL_98(int_bus__EVAL_98),
    ._EVAL_99(int_bus__EVAL_99),
    ._EVAL_100(int_bus__EVAL_100),
    ._EVAL_101(int_bus__EVAL_101),
    ._EVAL_102(int_bus__EVAL_102),
    ._EVAL_103(int_bus__EVAL_103),
    ._EVAL_104(int_bus__EVAL_104),
    ._EVAL_105(int_bus__EVAL_105),
    ._EVAL_106(int_bus__EVAL_106),
    ._EVAL_107(int_bus__EVAL_107),
    ._EVAL_108(int_bus__EVAL_108),
    ._EVAL_109(int_bus__EVAL_109),
    ._EVAL_110(int_bus__EVAL_110),
    ._EVAL_111(int_bus__EVAL_111),
    ._EVAL_112(int_bus__EVAL_112),
    ._EVAL_113(int_bus__EVAL_113),
    ._EVAL_114(int_bus__EVAL_114),
    ._EVAL_115(int_bus__EVAL_115),
    ._EVAL_116(int_bus__EVAL_116),
    ._EVAL_117(int_bus__EVAL_117),
    ._EVAL_118(int_bus__EVAL_118),
    ._EVAL_119(int_bus__EVAL_119),
    ._EVAL_120(int_bus__EVAL_120),
    ._EVAL_121(int_bus__EVAL_121),
    ._EVAL_122(int_bus__EVAL_122),
    ._EVAL_123(int_bus__EVAL_123),
    ._EVAL_124(int_bus__EVAL_124),
    ._EVAL_125(int_bus__EVAL_125),
    ._EVAL_126(int_bus__EVAL_126),
    ._EVAL_127(int_bus__EVAL_127),
    ._EVAL_128(int_bus__EVAL_128),
    ._EVAL_129(int_bus__EVAL_129),
    ._EVAL_130(int_bus__EVAL_130),
    ._EVAL_131(int_bus__EVAL_131),
    ._EVAL_132(int_bus__EVAL_132),
    ._EVAL_133(int_bus__EVAL_133),
    ._EVAL_134(int_bus__EVAL_134),
    ._EVAL_135(int_bus__EVAL_135),
    ._EVAL_136(int_bus__EVAL_136),
    ._EVAL_137(int_bus__EVAL_137),
    ._EVAL_138(int_bus__EVAL_138),
    ._EVAL_139(int_bus__EVAL_139),
    ._EVAL_140(int_bus__EVAL_140),
    ._EVAL_141(int_bus__EVAL_141),
    ._EVAL_142(int_bus__EVAL_142),
    ._EVAL_143(int_bus__EVAL_143),
    ._EVAL_144(int_bus__EVAL_144),
    ._EVAL_145(int_bus__EVAL_145),
    ._EVAL_146(int_bus__EVAL_146),
    ._EVAL_147(int_bus__EVAL_147),
    ._EVAL_148(int_bus__EVAL_148),
    ._EVAL_149(int_bus__EVAL_149),
    ._EVAL_150(int_bus__EVAL_150),
    ._EVAL_151(int_bus__EVAL_151),
    ._EVAL_152(int_bus__EVAL_152),
    ._EVAL_153(int_bus__EVAL_153),
    ._EVAL_154(int_bus__EVAL_154),
    ._EVAL_155(int_bus__EVAL_155),
    ._EVAL_156(int_bus__EVAL_156),
    ._EVAL_157(int_bus__EVAL_157),
    ._EVAL_158(int_bus__EVAL_158),
    ._EVAL_159(int_bus__EVAL_159),
    ._EVAL_160(int_bus__EVAL_160),
    ._EVAL_161(int_bus__EVAL_161),
    ._EVAL_162(int_bus__EVAL_162),
    ._EVAL_163(int_bus__EVAL_163),
    ._EVAL_164(int_bus__EVAL_164),
    ._EVAL_165(int_bus__EVAL_165),
    ._EVAL_166(int_bus__EVAL_166),
    ._EVAL_167(int_bus__EVAL_167),
    ._EVAL_168(int_bus__EVAL_168),
    ._EVAL_169(int_bus__EVAL_169),
    ._EVAL_170(int_bus__EVAL_170),
    ._EVAL_171(int_bus__EVAL_171),
    ._EVAL_172(int_bus__EVAL_172),
    ._EVAL_173(int_bus__EVAL_173),
    ._EVAL_174(int_bus__EVAL_174),
    ._EVAL_175(int_bus__EVAL_175),
    ._EVAL_176(int_bus__EVAL_176),
    ._EVAL_177(int_bus__EVAL_177),
    ._EVAL_178(int_bus__EVAL_178),
    ._EVAL_179(int_bus__EVAL_179),
    ._EVAL_180(int_bus__EVAL_180),
    ._EVAL_181(int_bus__EVAL_181),
    ._EVAL_182(int_bus__EVAL_182),
    ._EVAL_183(int_bus__EVAL_183),
    ._EVAL_184(int_bus__EVAL_184),
    ._EVAL_185(int_bus__EVAL_185),
    ._EVAL_186(int_bus__EVAL_186),
    ._EVAL_187(int_bus__EVAL_187),
    ._EVAL_188(int_bus__EVAL_188),
    ._EVAL_189(int_bus__EVAL_189),
    ._EVAL_190(int_bus__EVAL_190),
    ._EVAL_191(int_bus__EVAL_191),
    ._EVAL_192(int_bus__EVAL_192),
    ._EVAL_193(int_bus__EVAL_193),
    ._EVAL_194(int_bus__EVAL_194),
    ._EVAL_195(int_bus__EVAL_195),
    ._EVAL_196(int_bus__EVAL_196),
    ._EVAL_197(int_bus__EVAL_197),
    ._EVAL_198(int_bus__EVAL_198),
    ._EVAL_199(int_bus__EVAL_199),
    ._EVAL_200(int_bus__EVAL_200),
    ._EVAL_201(int_bus__EVAL_201),
    ._EVAL_202(int_bus__EVAL_202),
    ._EVAL_203(int_bus__EVAL_203),
    ._EVAL_204(int_bus__EVAL_204),
    ._EVAL_205(int_bus__EVAL_205),
    ._EVAL_206(int_bus__EVAL_206),
    ._EVAL_207(int_bus__EVAL_207),
    ._EVAL_208(int_bus__EVAL_208),
    ._EVAL_209(int_bus__EVAL_209),
    ._EVAL_210(int_bus__EVAL_210),
    ._EVAL_211(int_bus__EVAL_211),
    ._EVAL_212(int_bus__EVAL_212),
    ._EVAL_213(int_bus__EVAL_213),
    ._EVAL_214(int_bus__EVAL_214),
    ._EVAL_215(int_bus__EVAL_215),
    ._EVAL_216(int_bus__EVAL_216),
    ._EVAL_217(int_bus__EVAL_217),
    ._EVAL_218(int_bus__EVAL_218),
    ._EVAL_219(int_bus__EVAL_219),
    ._EVAL_220(int_bus__EVAL_220),
    ._EVAL_221(int_bus__EVAL_221),
    ._EVAL_222(int_bus__EVAL_222),
    ._EVAL_223(int_bus__EVAL_223),
    ._EVAL_224(int_bus__EVAL_224),
    ._EVAL_225(int_bus__EVAL_225),
    ._EVAL_226(int_bus__EVAL_226),
    ._EVAL_227(int_bus__EVAL_227),
    ._EVAL_228(int_bus__EVAL_228),
    ._EVAL_229(int_bus__EVAL_229),
    ._EVAL_230(int_bus__EVAL_230),
    ._EVAL_231(int_bus__EVAL_231),
    ._EVAL_232(int_bus__EVAL_232),
    ._EVAL_233(int_bus__EVAL_233),
    ._EVAL_234(int_bus__EVAL_234),
    ._EVAL_235(int_bus__EVAL_235),
    ._EVAL_236(int_bus__EVAL_236),
    ._EVAL_237(int_bus__EVAL_237),
    ._EVAL_238(int_bus__EVAL_238),
    ._EVAL_239(int_bus__EVAL_239),
    ._EVAL_240(int_bus__EVAL_240),
    ._EVAL_241(int_bus__EVAL_241),
    ._EVAL_242(int_bus__EVAL_242),
    ._EVAL_243(int_bus__EVAL_243),
    ._EVAL_244(int_bus__EVAL_244),
    ._EVAL_245(int_bus__EVAL_245),
    ._EVAL_246(int_bus__EVAL_246),
    ._EVAL_247(int_bus__EVAL_247),
    ._EVAL_248(int_bus__EVAL_248),
    ._EVAL_249(int_bus__EVAL_249),
    ._EVAL_250(int_bus__EVAL_250),
    ._EVAL_251(int_bus__EVAL_251),
    ._EVAL_252(int_bus__EVAL_252)
  );
  SiFive__EVAL_312 intsource (
    ._EVAL(intsource__EVAL),
    ._EVAL_0(intsource__EVAL_0),
    ._EVAL_1(intsource__EVAL_1),
    ._EVAL_2(intsource__EVAL_2),
    ._EVAL_3(intsource__EVAL_3),
    ._EVAL_4(intsource__EVAL_4)
  );
  SiFive__EVAL_85 fbus (
    ._EVAL(fbus__EVAL),
    ._EVAL_0(fbus__EVAL_0),
    ._EVAL_1(fbus__EVAL_1),
    ._EVAL_2(fbus__EVAL_2),
    ._EVAL_3(fbus__EVAL_3),
    ._EVAL_4(fbus__EVAL_4),
    ._EVAL_5(fbus__EVAL_5),
    ._EVAL_6(fbus__EVAL_6),
    ._EVAL_7(fbus__EVAL_7),
    ._EVAL_8(fbus__EVAL_8),
    ._EVAL_9(fbus__EVAL_9),
    ._EVAL_10(fbus__EVAL_10),
    ._EVAL_11(fbus__EVAL_11),
    ._EVAL_12(fbus__EVAL_12),
    ._EVAL_13(fbus__EVAL_13),
    ._EVAL_14(fbus__EVAL_14),
    ._EVAL_15(fbus__EVAL_15),
    ._EVAL_16(fbus__EVAL_16),
    ._EVAL_17(fbus__EVAL_17),
    ._EVAL_18(fbus__EVAL_18),
    ._EVAL_19(fbus__EVAL_19),
    ._EVAL_20(fbus__EVAL_20),
    ._EVAL_21(fbus__EVAL_21),
    ._EVAL_22(fbus__EVAL_22),
    ._EVAL_23(fbus__EVAL_23),
    ._EVAL_24(fbus__EVAL_24),
    ._EVAL_25(fbus__EVAL_25),
    ._EVAL_26(fbus__EVAL_26),
    ._EVAL_27(fbus__EVAL_27),
    ._EVAL_28(fbus__EVAL_28),
    ._EVAL_29(fbus__EVAL_29),
    ._EVAL_30(fbus__EVAL_30),
    ._EVAL_31(fbus__EVAL_31),
    ._EVAL_32(fbus__EVAL_32),
    ._EVAL_33(fbus__EVAL_33),
    ._EVAL_34(fbus__EVAL_34),
    ._EVAL_35(fbus__EVAL_35),
    ._EVAL_36(fbus__EVAL_36),
    ._EVAL_37(fbus__EVAL_37),
    ._EVAL_38(fbus__EVAL_38),
    ._EVAL_39(fbus__EVAL_39),
    ._EVAL_40(fbus__EVAL_40),
    ._EVAL_41(fbus__EVAL_41),
    ._EVAL_42(fbus__EVAL_42),
    ._EVAL_43(fbus__EVAL_43),
    ._EVAL_44(fbus__EVAL_44),
    ._EVAL_45(fbus__EVAL_45),
    ._EVAL_46(fbus__EVAL_46),
    ._EVAL_47(fbus__EVAL_47),
    ._EVAL_48(fbus__EVAL_48),
    ._EVAL_49(fbus__EVAL_49),
    ._EVAL_50(fbus__EVAL_50),
    ._EVAL_51(fbus__EVAL_51),
    ._EVAL_52(fbus__EVAL_52),
    ._EVAL_53(fbus__EVAL_53),
    ._EVAL_54(fbus__EVAL_54),
    ._EVAL_55(fbus__EVAL_55),
    ._EVAL_56(fbus__EVAL_56),
    ._EVAL_57(fbus__EVAL_57),
    ._EVAL_58(fbus__EVAL_58),
    ._EVAL_59(fbus__EVAL_59),
    ._EVAL_60(fbus__EVAL_60)
  );
  SiFive__EVAL_222 debug_1 (
    ._EVAL(debug_1__EVAL),
    ._EVAL_0(debug_1__EVAL_0),
    ._EVAL_1(debug_1__EVAL_1),
    ._EVAL_2(debug_1__EVAL_2),
    ._EVAL_3(debug_1__EVAL_3),
    ._EVAL_4(debug_1__EVAL_4),
    ._EVAL_5(debug_1__EVAL_5),
    ._EVAL_6(debug_1__EVAL_6),
    ._EVAL_7(debug_1__EVAL_7),
    ._EVAL_8(debug_1__EVAL_8),
    ._EVAL_9(debug_1__EVAL_9),
    ._EVAL_10(debug_1__EVAL_10),
    ._EVAL_11(debug_1__EVAL_11),
    ._EVAL_12(debug_1__EVAL_12),
    ._EVAL_13(debug_1__EVAL_13),
    ._EVAL_14(debug_1__EVAL_14),
    ._EVAL_15(debug_1__EVAL_15),
    ._EVAL_16(debug_1__EVAL_16),
    ._EVAL_17(debug_1__EVAL_17),
    ._EVAL_18(debug_1__EVAL_18),
    ._EVAL_19(debug_1__EVAL_19),
    ._EVAL_20(debug_1__EVAL_20),
    ._EVAL_21(debug_1__EVAL_21),
    ._EVAL_22(debug_1__EVAL_22),
    ._EVAL_23(debug_1__EVAL_23),
    ._EVAL_24(debug_1__EVAL_24),
    ._EVAL_25(debug_1__EVAL_25),
    ._EVAL_26(debug_1__EVAL_26),
    ._EVAL_27(debug_1__EVAL_27),
    ._EVAL_28(debug_1__EVAL_28),
    ._EVAL_29(debug_1__EVAL_29),
    ._EVAL_30(debug_1__EVAL_30),
    ._EVAL_31(debug_1__EVAL_31),
    ._EVAL_32(debug_1__EVAL_32),
    ._EVAL_33(debug_1__EVAL_33),
    ._EVAL_34(debug_1__EVAL_34),
    ._EVAL_35(debug_1__EVAL_35),
    ._EVAL_36(debug_1__EVAL_36),
    ._EVAL_37(debug_1__EVAL_37),
    ._EVAL_38(debug_1__EVAL_38),
    ._EVAL_39(debug_1__EVAL_39),
    ._EVAL_40(debug_1__EVAL_40),
    ._EVAL_41(debug_1__EVAL_41),
    ._EVAL_42(debug_1__EVAL_42),
    ._EVAL_43(debug_1__EVAL_43)
  );
  SiFive__EVAL_180 cbus (
    ._EVAL(cbus__EVAL),
    ._EVAL_0(cbus__EVAL_0),
    ._EVAL_1(cbus__EVAL_1),
    ._EVAL_2(cbus__EVAL_2),
    ._EVAL_3(cbus__EVAL_3),
    ._EVAL_4(cbus__EVAL_4),
    ._EVAL_5(cbus__EVAL_5),
    ._EVAL_6(cbus__EVAL_6),
    ._EVAL_7(cbus__EVAL_7),
    ._EVAL_8(cbus__EVAL_8),
    ._EVAL_9(cbus__EVAL_9),
    ._EVAL_10(cbus__EVAL_10),
    ._EVAL_11(cbus__EVAL_11),
    ._EVAL_12(cbus__EVAL_12),
    ._EVAL_13(cbus__EVAL_13),
    ._EVAL_14(cbus__EVAL_14),
    ._EVAL_15(cbus__EVAL_15),
    ._EVAL_16(cbus__EVAL_16),
    ._EVAL_17(cbus__EVAL_17),
    ._EVAL_18(cbus__EVAL_18),
    ._EVAL_19(cbus__EVAL_19),
    ._EVAL_20(cbus__EVAL_20),
    ._EVAL_21(cbus__EVAL_21),
    ._EVAL_22(cbus__EVAL_22),
    ._EVAL_23(cbus__EVAL_23),
    ._EVAL_24(cbus__EVAL_24),
    ._EVAL_25(cbus__EVAL_25),
    ._EVAL_26(cbus__EVAL_26),
    ._EVAL_27(cbus__EVAL_27),
    ._EVAL_28(cbus__EVAL_28),
    ._EVAL_29(cbus__EVAL_29),
    ._EVAL_30(cbus__EVAL_30),
    ._EVAL_31(cbus__EVAL_31),
    ._EVAL_32(cbus__EVAL_32),
    ._EVAL_33(cbus__EVAL_33),
    ._EVAL_34(cbus__EVAL_34),
    ._EVAL_35(cbus__EVAL_35),
    ._EVAL_36(cbus__EVAL_36),
    ._EVAL_37(cbus__EVAL_37),
    ._EVAL_38(cbus__EVAL_38),
    ._EVAL_39(cbus__EVAL_39),
    ._EVAL_40(cbus__EVAL_40),
    ._EVAL_41(cbus__EVAL_41),
    ._EVAL_42(cbus__EVAL_42),
    ._EVAL_43(cbus__EVAL_43),
    ._EVAL_44(cbus__EVAL_44),
    ._EVAL_45(cbus__EVAL_45),
    ._EVAL_46(cbus__EVAL_46),
    ._EVAL_47(cbus__EVAL_47),
    ._EVAL_48(cbus__EVAL_48),
    ._EVAL_49(cbus__EVAL_49),
    ._EVAL_50(cbus__EVAL_50),
    ._EVAL_51(cbus__EVAL_51),
    ._EVAL_52(cbus__EVAL_52),
    ._EVAL_53(cbus__EVAL_53),
    ._EVAL_54(cbus__EVAL_54),
    ._EVAL_55(cbus__EVAL_55),
    ._EVAL_56(cbus__EVAL_56),
    ._EVAL_57(cbus__EVAL_57),
    ._EVAL_58(cbus__EVAL_58),
    ._EVAL_59(cbus__EVAL_59),
    ._EVAL_60(cbus__EVAL_60),
    ._EVAL_61(cbus__EVAL_61),
    ._EVAL_62(cbus__EVAL_62),
    ._EVAL_63(cbus__EVAL_63),
    ._EVAL_64(cbus__EVAL_64),
    ._EVAL_65(cbus__EVAL_65),
    ._EVAL_66(cbus__EVAL_66),
    ._EVAL_67(cbus__EVAL_67),
    ._EVAL_68(cbus__EVAL_68),
    ._EVAL_69(cbus__EVAL_69),
    ._EVAL_70(cbus__EVAL_70),
    ._EVAL_71(cbus__EVAL_71),
    ._EVAL_72(cbus__EVAL_72),
    ._EVAL_73(cbus__EVAL_73),
    ._EVAL_74(cbus__EVAL_74),
    ._EVAL_75(cbus__EVAL_75),
    ._EVAL_76(cbus__EVAL_76),
    ._EVAL_77(cbus__EVAL_77),
    ._EVAL_78(cbus__EVAL_78),
    ._EVAL_79(cbus__EVAL_79),
    ._EVAL_80(cbus__EVAL_80),
    ._EVAL_81(cbus__EVAL_81),
    ._EVAL_82(cbus__EVAL_82),
    ._EVAL_83(cbus__EVAL_83),
    ._EVAL_84(cbus__EVAL_84),
    ._EVAL_85(cbus__EVAL_85),
    ._EVAL_86(cbus__EVAL_86),
    ._EVAL_87(cbus__EVAL_87),
    ._EVAL_88(cbus__EVAL_88),
    ._EVAL_89(cbus__EVAL_89),
    ._EVAL_90(cbus__EVAL_90),
    ._EVAL_91(cbus__EVAL_91),
    ._EVAL_92(cbus__EVAL_92),
    ._EVAL_93(cbus__EVAL_93),
    ._EVAL_94(cbus__EVAL_94),
    ._EVAL_95(cbus__EVAL_95),
    ._EVAL_96(cbus__EVAL_96),
    ._EVAL_97(cbus__EVAL_97),
    ._EVAL_98(cbus__EVAL_98),
    ._EVAL_99(cbus__EVAL_99),
    ._EVAL_100(cbus__EVAL_100),
    ._EVAL_101(cbus__EVAL_101),
    ._EVAL_102(cbus__EVAL_102),
    ._EVAL_103(cbus__EVAL_103),
    ._EVAL_104(cbus__EVAL_104),
    ._EVAL_105(cbus__EVAL_105),
    ._EVAL_106(cbus__EVAL_106),
    ._EVAL_107(cbus__EVAL_107),
    ._EVAL_108(cbus__EVAL_108),
    ._EVAL_109(cbus__EVAL_109),
    ._EVAL_110(cbus__EVAL_110),
    ._EVAL_111(cbus__EVAL_111),
    ._EVAL_112(cbus__EVAL_112),
    ._EVAL_113(cbus__EVAL_113),
    ._EVAL_114(cbus__EVAL_114),
    ._EVAL_115(cbus__EVAL_115),
    ._EVAL_116(cbus__EVAL_116),
    ._EVAL_117(cbus__EVAL_117),
    ._EVAL_118(cbus__EVAL_118),
    ._EVAL_119(cbus__EVAL_119),
    ._EVAL_120(cbus__EVAL_120),
    ._EVAL_121(cbus__EVAL_121),
    ._EVAL_122(cbus__EVAL_122),
    ._EVAL_123(cbus__EVAL_123),
    ._EVAL_124(cbus__EVAL_124),
    ._EVAL_125(cbus__EVAL_125),
    ._EVAL_126(cbus__EVAL_126),
    ._EVAL_127(cbus__EVAL_127),
    ._EVAL_128(cbus__EVAL_128),
    ._EVAL_129(cbus__EVAL_129),
    ._EVAL_130(cbus__EVAL_130),
    ._EVAL_131(cbus__EVAL_131),
    ._EVAL_132(cbus__EVAL_132),
    ._EVAL_133(cbus__EVAL_133),
    ._EVAL_134(cbus__EVAL_134),
    ._EVAL_135(cbus__EVAL_135),
    ._EVAL_136(cbus__EVAL_136),
    ._EVAL_137(cbus__EVAL_137),
    ._EVAL_138(cbus__EVAL_138),
    ._EVAL_139(cbus__EVAL_139),
    ._EVAL_140(cbus__EVAL_140),
    ._EVAL_141(cbus__EVAL_141),
    ._EVAL_142(cbus__EVAL_142),
    ._EVAL_143(cbus__EVAL_143),
    ._EVAL_144(cbus__EVAL_144),
    ._EVAL_145(cbus__EVAL_145),
    ._EVAL_146(cbus__EVAL_146),
    ._EVAL_147(cbus__EVAL_147),
    ._EVAL_148(cbus__EVAL_148),
    ._EVAL_149(cbus__EVAL_149),
    ._EVAL_150(cbus__EVAL_150),
    ._EVAL_151(cbus__EVAL_151),
    ._EVAL_152(cbus__EVAL_152),
    ._EVAL_153(cbus__EVAL_153),
    ._EVAL_154(cbus__EVAL_154),
    ._EVAL_155(cbus__EVAL_155),
    ._EVAL_156(cbus__EVAL_156),
    ._EVAL_157(cbus__EVAL_157),
    ._EVAL_158(cbus__EVAL_158),
    ._EVAL_159(cbus__EVAL_159)
  );
  SiFive__EVAL_187 clint (
    ._EVAL(clint__EVAL),
    ._EVAL_0(clint__EVAL_0),
    ._EVAL_1(clint__EVAL_1),
    ._EVAL_2(clint__EVAL_2),
    ._EVAL_3(clint__EVAL_3),
    ._EVAL_4(clint__EVAL_4),
    ._EVAL_5(clint__EVAL_5),
    ._EVAL_6(clint__EVAL_6),
    ._EVAL_7(clint__EVAL_7),
    ._EVAL_8(clint__EVAL_8),
    ._EVAL_9(clint__EVAL_9),
    ._EVAL_10(clint__EVAL_10),
    ._EVAL_11(clint__EVAL_11),
    ._EVAL_12(clint__EVAL_12),
    ._EVAL_13(clint__EVAL_13),
    ._EVAL_14(clint__EVAL_14),
    ._EVAL_15(clint__EVAL_15),
    ._EVAL_16(clint__EVAL_16),
    ._EVAL_17(clint__EVAL_17),
    ._EVAL_18(clint__EVAL_18),
    ._EVAL_19(clint__EVAL_19)
  );
  SiFive__EVAL_324 shrinker (
    ._EVAL(shrinker__EVAL),
    ._EVAL_0(shrinker__EVAL_0),
    ._EVAL_1(shrinker__EVAL_1),
    ._EVAL_2(shrinker__EVAL_2),
    ._EVAL_3(shrinker__EVAL_3),
    ._EVAL_4(shrinker__EVAL_4),
    ._EVAL_5(shrinker__EVAL_5),
    ._EVAL_6(shrinker__EVAL_6),
    ._EVAL_7(shrinker__EVAL_7),
    ._EVAL_8(shrinker__EVAL_8),
    ._EVAL_9(shrinker__EVAL_9),
    ._EVAL_10(shrinker__EVAL_10),
    ._EVAL_11(shrinker__EVAL_11),
    ._EVAL_12(shrinker__EVAL_12),
    ._EVAL_13(shrinker__EVAL_13),
    ._EVAL_14(shrinker__EVAL_14),
    ._EVAL_15(shrinker__EVAL_15),
    ._EVAL_16(shrinker__EVAL_16),
    ._EVAL_17(shrinker__EVAL_17),
    ._EVAL_18(shrinker__EVAL_18),
    ._EVAL_19(shrinker__EVAL_19),
    ._EVAL_20(shrinker__EVAL_20),
    ._EVAL_21(shrinker__EVAL_21),
    ._EVAL_22(shrinker__EVAL_22),
    ._EVAL_23(shrinker__EVAL_23),
    ._EVAL_24(shrinker__EVAL_24),
    ._EVAL_25(shrinker__EVAL_25),
    ._EVAL_26(shrinker__EVAL_26),
    ._EVAL_27(shrinker__EVAL_27),
    ._EVAL_28(shrinker__EVAL_28),
    ._EVAL_29(shrinker__EVAL_29),
    ._EVAL_30(shrinker__EVAL_30),
    ._EVAL_31(shrinker__EVAL_31),
    ._EVAL_32(shrinker__EVAL_32),
    ._EVAL_33(shrinker__EVAL_33),
    ._EVAL_34(shrinker__EVAL_34),
    ._EVAL_35(shrinker__EVAL_35),
    ._EVAL_36(shrinker__EVAL_36)
  );
  SiFive_TLTestIndicator testIndicator (
    .clock(testIndicator_clock),
    .reset(testIndicator_reset),
    .auto_in_a_ready(testIndicator_auto_in_a_ready),
    .auto_in_a_valid(testIndicator_auto_in_a_valid),
    .auto_in_a_bits_opcode(testIndicator_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(testIndicator_auto_in_a_bits_param),
    .auto_in_a_bits_size(testIndicator_auto_in_a_bits_size),
    .auto_in_a_bits_source(testIndicator_auto_in_a_bits_source),
    .auto_in_a_bits_address(testIndicator_auto_in_a_bits_address),
    .auto_in_a_bits_mask(testIndicator_auto_in_a_bits_mask),
    .auto_in_a_bits_data(testIndicator_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(testIndicator_auto_in_a_bits_corrupt),
    .auto_in_d_ready(testIndicator_auto_in_d_ready),
    .auto_in_d_valid(testIndicator_auto_in_d_valid),
    .auto_in_d_bits_opcode(testIndicator_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(testIndicator_auto_in_d_bits_size),
    .auto_in_d_bits_source(testIndicator_auto_in_d_bits_source),
    .auto_in_d_bits_data(testIndicator_auto_in_d_bits_data)
  );
  SiFive__EVAL_313 intsource_1 (
    ._EVAL(intsource_1__EVAL),
    ._EVAL_0(intsource_1__EVAL_0),
    ._EVAL_1(intsource_1__EVAL_1),
    ._EVAL_2(intsource_1__EVAL_2)
  );
  SiFive__EVAL_320 bh (
    ._EVAL(bh__EVAL),
    ._EVAL_0(bh__EVAL_0),
    ._EVAL_1(bh__EVAL_1),
    ._EVAL_2(bh__EVAL_2),
    ._EVAL_3(bh__EVAL_3),
    ._EVAL_4(bh__EVAL_4),
    ._EVAL_5(bh__EVAL_5),
    ._EVAL_6(bh__EVAL_6),
    ._EVAL_7(bh__EVAL_7),
    ._EVAL_8(bh__EVAL_8),
    ._EVAL_9(bh__EVAL_9),
    ._EVAL_10(bh__EVAL_10),
    ._EVAL_11(bh__EVAL_11),
    ._EVAL_12(bh__EVAL_12),
    ._EVAL_13(bh__EVAL_13),
    ._EVAL_14(bh__EVAL_14),
    ._EVAL_15(bh__EVAL_15),
    ._EVAL_16(bh__EVAL_16),
    ._EVAL_17(bh__EVAL_17),
    ._EVAL_18(bh__EVAL_18),
    ._EVAL_19(bh__EVAL_19),
    ._EVAL_20(bh__EVAL_20),
    ._EVAL_21(bh__EVAL_21),
    ._EVAL_22(bh__EVAL_22),
    ._EVAL_23(bh__EVAL_23),
    ._EVAL_24(bh__EVAL_24),
    ._EVAL_25(bh__EVAL_25),
    ._EVAL_26(bh__EVAL_26),
    ._EVAL_27(bh__EVAL_27),
    ._EVAL_28(bh__EVAL_28),
    ._EVAL_29(bh__EVAL_29),
    ._EVAL_30(bh__EVAL_30),
    ._EVAL_31(bh__EVAL_31),
    ._EVAL_32(bh__EVAL_32),
    ._EVAL_33(bh__EVAL_33),
    ._EVAL_34(bh__EVAL_34),
    ._EVAL_35(bh__EVAL_35),
    ._EVAL_36(bh__EVAL_36),
    ._EVAL_37(bh__EVAL_37),
    ._EVAL_38(bh__EVAL_38),
    ._EVAL_39(bh__EVAL_39),
    ._EVAL_40(bh__EVAL_40),
    ._EVAL_41(bh__EVAL_41),
    ._EVAL_42(bh__EVAL_42),
    ._EVAL_43(bh__EVAL_43),
    ._EVAL_44(bh__EVAL_44),
    ._EVAL_45(bh__EVAL_45),
    ._EVAL_46(bh__EVAL_46),
    ._EVAL_47(bh__EVAL_47),
    ._EVAL_48(bh__EVAL_48),
    ._EVAL_49(bh__EVAL_49),
    ._EVAL_50(bh__EVAL_50),
    ._EVAL_51(bh__EVAL_51),
    ._EVAL_52(bh__EVAL_52),
    ._EVAL_53(bh__EVAL_53)
  );
  SiFive__EVAL_110 mbus (
    ._EVAL(mbus__EVAL),
    ._EVAL_0(mbus__EVAL_0),
    ._EVAL_1(mbus__EVAL_1),
    ._EVAL_2(mbus__EVAL_2),
    ._EVAL_3(mbus__EVAL_3),
    ._EVAL_4(mbus__EVAL_4),
    ._EVAL_5(mbus__EVAL_5),
    ._EVAL_6(mbus__EVAL_6),
    ._EVAL_7(mbus__EVAL_7),
    ._EVAL_8(mbus__EVAL_8),
    ._EVAL_9(mbus__EVAL_9),
    ._EVAL_10(mbus__EVAL_10),
    ._EVAL_11(mbus__EVAL_11),
    ._EVAL_12(mbus__EVAL_12),
    ._EVAL_13(mbus__EVAL_13),
    ._EVAL_14(mbus__EVAL_14),
    ._EVAL_15(mbus__EVAL_15),
    ._EVAL_16(mbus__EVAL_16),
    ._EVAL_17(mbus__EVAL_17),
    ._EVAL_18(mbus__EVAL_18),
    ._EVAL_19(mbus__EVAL_19),
    ._EVAL_20(mbus__EVAL_20),
    ._EVAL_21(mbus__EVAL_21),
    ._EVAL_22(mbus__EVAL_22),
    ._EVAL_23(mbus__EVAL_23),
    ._EVAL_24(mbus__EVAL_24),
    ._EVAL_25(mbus__EVAL_25),
    ._EVAL_26(mbus__EVAL_26),
    ._EVAL_27(mbus__EVAL_27),
    ._EVAL_28(mbus__EVAL_28),
    ._EVAL_29(mbus__EVAL_29),
    ._EVAL_30(mbus__EVAL_30),
    ._EVAL_31(mbus__EVAL_31),
    ._EVAL_32(mbus__EVAL_32),
    ._EVAL_33(mbus__EVAL_33),
    ._EVAL_34(mbus__EVAL_34),
    ._EVAL_35(mbus__EVAL_35),
    ._EVAL_36(mbus__EVAL_36),
    ._EVAL_37(mbus__EVAL_37),
    ._EVAL_38(mbus__EVAL_38),
    ._EVAL_39(mbus__EVAL_39),
    ._EVAL_40(mbus__EVAL_40),
    ._EVAL_41(mbus__EVAL_41),
    ._EVAL_42(mbus__EVAL_42),
    ._EVAL_43(mbus__EVAL_43),
    ._EVAL_44(mbus__EVAL_44),
    ._EVAL_45(mbus__EVAL_45),
    ._EVAL_46(mbus__EVAL_46),
    ._EVAL_47(mbus__EVAL_47),
    ._EVAL_48(mbus__EVAL_48),
    ._EVAL_49(mbus__EVAL_49),
    ._EVAL_50(mbus__EVAL_50),
    ._EVAL_51(mbus__EVAL_51),
    ._EVAL_52(mbus__EVAL_52),
    ._EVAL_53(mbus__EVAL_53),
    ._EVAL_54(mbus__EVAL_54),
    ._EVAL_55(mbus__EVAL_55),
    ._EVAL_56(mbus__EVAL_56)
  );
  assign _EVAL_2 = SynchronizerShiftReg_w1_d3__EVAL_0;
  assign _EVAL_3 = ~ _EVAL_1;
  assign _EVAL = _EVAL_2 & _EVAL_3;
  assign _EVAL_0 = 2'h0;
  assign tile__EVAL_61 = sbus__EVAL_198;
  assign int_bus__EVAL_64 = global_interrupts[116];
  assign sbus__EVAL_97 = tile__EVAL_71;
  assign sbus__EVAL_179 = tile__EVAL_11;
  assign mem_port_axi4_0_ar_bits_prot = mbus__EVAL_24;
  assign fbus__EVAL_2 = debug_1__EVAL_24;
  assign sbus__EVAL_192 = sagesafety__EVAL_19;
  assign bh__EVAL_16 = ww__EVAL_28;
  assign fbus__EVAL_52 = debug_1__EVAL_16;
  assign int_bus__EVAL_89 = global_interrupts[62];
  assign sys_port_axi4_0_aw_bits_len = sbus__EVAL_142;
  assign sys_port_axi4_0_r_ready = sbus__EVAL_167;
  assign sbus__EVAL_116 = bh__EVAL_2;
  assign int_bus__EVAL_103 = global_interrupts[89];
  assign fbus__EVAL_8 = front_port_axi4_0_aw_bits_addr;
  assign plic__EVAL_115 = int_bus__EVAL_46;
  assign int_bus__EVAL_209 = global_interrupts[30];
  assign plic__EVAL_21 = int_bus__EVAL_242;
  assign tile__EVAL_51 = sbus__EVAL_68;
  assign fbus__EVAL_30 = front_port_axi4_0_ar_valid;
  assign plic__EVAL_118 = int_bus__EVAL_76;
  assign int_bus__EVAL_212 = global_interrupts[51];
  assign shrinker__EVAL_15 = mbus__EVAL_39;
  assign plic__EVAL_75 = int_bus__EVAL_202;
  assign int_bus__EVAL_68 = global_interrupts[76];
  assign sbus__EVAL_112 = tile__EVAL_34;
  assign plic__EVAL_51 = cbus__EVAL_9;
  assign mem_port_axi4_0_aw_bits_len = mbus__EVAL_48;
  assign testIndicator_auto_in_a_bits_address = cbus__EVAL_78;
  assign plic__EVAL_39 = int_bus__EVAL_170;
  assign ww__EVAL_26 = bh__EVAL_15;
  assign sbus__EVAL_120 = tile__EVAL_57;
  assign debug_1__EVAL_17 = cbus__EVAL_132;
  assign shrinker__EVAL_32 = ww__EVAL_24;
  assign int_bus__EVAL_116 = global_interrupts[59];
  assign int_bus__EVAL_17 = global_interrupts[79];
  assign periph_port_axi4_0_r_ready = cbus__EVAL_150;
  assign fbus__EVAL_32 = front_port_axi4_0_aw_bits_burst;
  assign tile__EVAL_21 = sbus__EVAL_100;
  assign ww__EVAL_19 = bh__EVAL_48;
  assign sys_port_axi4_0_ar_bits_lock = sbus__EVAL_122;
  assign plic__EVAL_132 = int_bus__EVAL_63;
  assign tile__EVAL_53 = cbus__EVAL_149;
  assign sbus__EVAL_85 = tile__EVAL_79;
  assign mbus__EVAL_55 = shrinker__EVAL_31;
  assign sbus__EVAL_37 = sagesafety__EVAL_39;
  assign sbus__EVAL_69 = cbus__EVAL_48;
  assign cbus__EVAL_84 = periph_port_axi4_0_r_valid;
  assign sbus__EVAL_106 = tile__EVAL_66;
  assign cbus__EVAL_144 = sbus__EVAL_26;
  assign sbus__EVAL_1 = bh__EVAL_26;
  assign tile__EVAL_59 = cbus__EVAL_28;
  assign bh__EVAL_40 = ww__EVAL_11;
  assign mbus__EVAL_15 = mem_port_axi4_0_r_bits_data;
  assign shrinker__EVAL = ww__EVAL_34;
  assign periph_port_axi4_0_aw_bits_size = cbus__EVAL_125;
  assign sys_port_axi4_0_aw_bits_burst = sbus__EVAL_22;
  assign int_bus__EVAL_79 = global_interrupts[32];
  assign mbus__EVAL_22 = shrinker__EVAL_29;
  assign sbus__EVAL_157 = sagesafety__EVAL_8;
  assign int_bus__EVAL_124 = global_interrupts[3];
  assign bh__EVAL_21 = sbus__EVAL_64;
  assign mbus__EVAL_51 = shrinker__EVAL_28;
  assign sys_port_axi4_0_ar_bits_prot = sbus__EVAL_42;
  assign plic__EVAL_35 = int_bus__EVAL_78;
  assign ww__EVAL_23 = shrinker__EVAL_11;
  assign plic__EVAL_84 = cbus__EVAL_17;
  assign cbus__EVAL_141 = debug_1__EVAL_42;
  assign plic__EVAL_17 = int_bus__EVAL_144;
  assign mem_port_axi4_0_aw_bits_qos = mbus__EVAL_30;
  assign tile__EVAL_72 = sbus__EVAL_147;
  assign ww__EVAL_17 = shrinker__EVAL_22;
  assign plic__EVAL_86 = cbus__EVAL_21;
  assign plic__EVAL_110 = int_bus__EVAL_208;
  assign bh__EVAL_39 = sbus__EVAL_129;
  assign plic__EVAL_19 = int_bus__EVAL_44;
  assign debug_1__EVAL_34 = cbus__EVAL_65;
  assign int_bus__EVAL_166 = global_interrupts[57];
  assign int_bus__EVAL_122 = global_interrupts[5];
  assign plic__EVAL_124 = int_bus__EVAL_127;
  assign sys_port_axi4_0_aw_bits_cache = sbus__EVAL_201;
  assign cbus__EVAL_83 = plic__EVAL;
  assign ww__EVAL = shrinker__EVAL_7;
  assign sbus__EVAL_93 = fbus__EVAL_13;
  assign int_bus__EVAL_225 = global_interrupts[1];
  assign sbus__EVAL_59 = sys_port_axi4_0_r_bits_resp;
  assign int_bus__EVAL_81 = global_interrupts[29];
  assign periph_port_axi4_0_w_valid = cbus__EVAL_95;
  assign fbus__EVAL_44 = front_port_axi4_0_b_ready;
  assign plic__EVAL_69 = cbus__EVAL_4;
  assign plic__EVAL_93 = int_bus__EVAL_159;
  assign shrinker__EVAL_23 = ww__EVAL_13;
  assign sbus__EVAL_66 = sys_port_axi4_0_r_bits_data;
  assign int_bus__EVAL_204 = global_interrupts[56];
  assign tile__EVAL_39 = cbus__EVAL_87;
  assign fbus__EVAL_10 = front_port_axi4_0_ar_bits_len;
  assign cbus__EVAL_57 = periph_port_axi4_0_r_bits_data;
  assign int_bus__EVAL_98 = global_interrupts[80];
  assign int_bus__EVAL_229 = global_interrupts[69];
  assign sbus__EVAL_54 = sys_port_axi4_0_b_bits_resp;
  assign fbus__EVAL_45 = sbus__EVAL_12;
  assign mbus__EVAL_2 = reset;
  assign shrinker__EVAL_36 = ww__EVAL_22;
  assign sbus__EVAL_134 = sys_port_axi4_0_aw_ready;
  assign tile__EVAL_6 = cbus__EVAL_40;
  assign sbus__EVAL_131 = tile__EVAL_29;
  assign mem_port_axi4_0_aw_bits_id = mbus__EVAL_43;
  assign plic__EVAL_7 = int_bus__EVAL_160;
  assign plic__EVAL_56 = int_bus__EVAL_91;
  assign int_bus__EVAL_214 = global_interrupts[58];
  assign sbus__EVAL_14 = sagesafety__EVAL_34;
  assign int_bus__EVAL_136 = global_interrupts[72];
  assign int_bus__EVAL_18 = global_interrupts[97];
  assign sbus__EVAL_158 = fbus__EVAL_12;
  assign debug_1__EVAL_37 = debug_psd_test_mode_reset;
  assign plic__EVAL_1 = int_bus__EVAL_118;
  assign plic__EVAL_104 = int_bus__EVAL_16;
  assign fbus__EVAL_48 = debug_1__EVAL_1;
  assign shrinker__EVAL_21 = ww__EVAL_20;
  assign plic__EVAL_70 = int_bus__EVAL_58;
  assign int_bus__EVAL_13 = global_interrupts[114];
  assign int_bus__EVAL_161 = global_interrupts[28];
  assign int_bus__EVAL_233 = global_interrupts[92];
  assign plic__EVAL_137 = int_bus__EVAL_59;
  assign plic__EVAL_87 = int_bus__EVAL_192;
  assign sbus__EVAL_153 = sagesafety__EVAL_28;
  assign mem_port_axi4_0_ar_bits_lock = mbus__EVAL_25;
  assign mem_port_axi4_0_aw_bits_size = mbus__EVAL_13;
  assign plic__EVAL_59 = cbus__EVAL_151;
  assign sbus__EVAL_74 = sagesafety__EVAL;
  assign sbus__EVAL_105 = tile__EVAL_103;
  assign cbus__EVAL_15 = sbus__EVAL_96;
  assign plic__EVAL_91 = int_bus__EVAL_231;
  assign sys_port_axi4_0_b_ready = sbus__EVAL_216;
  assign mbus__EVAL_45 = mem_port_axi4_0_r_bits_last;
  assign plic__EVAL_2 = int_bus__EVAL_201;
  assign sbus__EVAL_127 = tile__EVAL_15;
  assign sbus__EVAL_70 = tile__EVAL_116;
  assign plic__EVAL_114 = int_bus__EVAL_143;
  assign cbus__EVAL_8 = debug_1__EVAL_11;
  assign front_port_axi4_0_b_bits_id = fbus__EVAL_1;
  assign sbus__EVAL_40 = tile__EVAL_40;
  assign sbus__EVAL_221 = tile__EVAL_99;
  assign cbus__EVAL_86 = debug_1__EVAL_7;
  assign shrinker__EVAL_16 = mbus__EVAL_21;
  assign shrinker__EVAL_30 = ww__EVAL_35;
  assign fbus__EVAL_37 = front_port_axi4_0_aw_valid;
  assign plic__EVAL_108 = int_bus__EVAL_47;
  assign dtm__EVAL_2 = debug_1__EVAL_30;
  assign int_bus__EVAL_65 = global_interrupts[112];
  assign sbus__EVAL_56 = bh__EVAL_38;
  assign tile__EVAL_19 = sbus__EVAL_94;
  assign shrinker__EVAL_8 = mbus__EVAL_26;
  assign int_bus__EVAL_142 = global_interrupts[22];
  assign plic__EVAL_23 = int_bus__EVAL_74;
  assign bh__EVAL_51 = sbus__EVAL_92;
  assign int_bus__EVAL_37 = global_interrupts[18];
  assign plic__EVAL_12 = int_bus__EVAL_88;
  assign debug_1__EVAL_32 = fbus__EVAL_6;
  assign sbus__EVAL_166 = bh__EVAL_34;
  assign cbus__EVAL_54 = plic__EVAL_130;
  assign mbus__EVAL_11 = shrinker__EVAL_20;
  assign fbus__EVAL_11 = front_port_axi4_0_ar_bits_size;
  assign sagesafety__EVAL_18 = reset;
  assign int_bus__EVAL_211 = global_interrupts[109];
  assign mem_port_axi4_0_aw_bits_prot = mbus__EVAL_4;
  assign int_bus__EVAL_27 = global_interrupts[37];
  assign periph_port_axi4_0_b_ready = cbus__EVAL_36;
  assign sbus__EVAL_48 = fbus__EVAL_5;
  assign mem_port_axi4_0_ar_bits_burst = mbus__EVAL_32;
  assign mem_port_axi4_0_ar_valid = mbus__EVAL_47;
  assign sbus__EVAL_138 = sys_port_axi4_0_r_bits_id;
  assign debug_1__EVAL_22 = clock;
  assign int_bus__EVAL_4 = global_interrupts[9];
  assign sbus__EVAL_186 = cbus__EVAL_68;
  assign sys_port_axi4_0_aw_bits_qos = sbus__EVAL_117;
  assign sbus__EVAL_6 = sagesafety__EVAL_30;
  assign int_bus__EVAL_193 = global_interrupts[126];
  assign int_bus__EVAL_2 = global_interrupts[0];
  assign plic__EVAL_83 = int_bus__EVAL_6;
  assign sbus__EVAL_79 = tile__EVAL_18;
  assign plic__EVAL_55 = int_bus__EVAL_31;
  assign ww__EVAL_9 = clock;
  assign int_bus__EVAL_163 = global_interrupts[86];
  assign mem_port_axi4_0_aw_bits_addr = mbus__EVAL_23;
  assign int_bus__EVAL_11 = global_interrupts[25];
  assign front_port_axi4_0_ar_ready = fbus__EVAL_42;
  assign int_bus__EVAL_216 = global_interrupts[35];
  assign fbus__EVAL_33 = debug_1__EVAL_14;
  assign bh__EVAL_8 = sbus__EVAL_11;
  assign cbus__EVAL_147 = testIndicator_auto_in_d_bits_data;
  assign testIndicator_auto_in_a_bits_data = cbus__EVAL_49;
  assign plic__EVAL_88 = int_bus__EVAL_129;
  assign tile__EVAL_94 = sbus__EVAL_162;
  assign cbus__EVAL_116 = periph_port_axi4_0_r_bits_last;
  assign mem_port_axi4_0_ar_bits_addr = mbus__EVAL_17;
  assign tile__EVAL_70 = cbus__EVAL_2;
  assign fbus__EVAL_22 = debug_1__EVAL_28;
  assign fbus__EVAL_56 = front_port_axi4_0_w_bits_strb;
  assign plic__EVAL_133 = int_bus__EVAL_104;
  assign periph_port_axi4_0_w_bits_data = cbus__EVAL_59;
  assign plic__EVAL_33 = int_bus__EVAL_26;
  assign mem_port_axi4_0_b_ready = mbus__EVAL_7;
  assign sys_port_axi4_0_aw_valid = sbus__EVAL_61;
  assign clint__EVAL_3 = cbus__EVAL_136;
  assign tile__EVAL_112 = sbus__EVAL_220;
  assign fbus__EVAL_41 = front_port_axi4_0_aw_bits_id;
  assign int_bus__EVAL_244 = global_interrupts[64];
  assign plic__EVAL_31 = int_bus__EVAL_220;
  assign bh__EVAL_28 = sbus__EVAL_73;
  assign mem_port_axi4_0_aw_valid = mbus__EVAL_37;
  assign sys_port_axi4_0_w_bits_data = sbus__EVAL_75;
  assign periph_port_axi4_0_aw_bits_prot = cbus__EVAL_64;
  assign tile__EVAL_26 = sbus__EVAL_177;
  assign tile__EVAL_111 = sbus__EVAL_77;
  assign sagesafety__EVAL_25 = sbus__EVAL_18;
  assign mem_port_axi4_0_w_valid = mbus__EVAL_34;
  assign plic__EVAL_26 = int_bus__EVAL_99;
  assign sbus__EVAL_204 = tile__EVAL_10;
  assign cbus__EVAL_13 = clint__EVAL_14;
  assign cbus__EVAL_52 = tile__EVAL_110;
  assign sbus__EVAL_137 = clock;
  assign sagesafety__EVAL_3 = sbus__EVAL_170;
  assign debug_1__EVAL_6 = cbus__EVAL_81;
  assign plic__EVAL_28 = int_bus__EVAL_195;
  assign tile__EVAL_7 = sbus__EVAL_223;
  assign int_bus__EVAL_146 = global_interrupts[102];
  assign plic__EVAL_29 = int_bus__EVAL_112;
  assign sbus__EVAL_62 = cbus__EVAL_120;
  assign plic__EVAL_143 = cbus__EVAL_66;
  assign periph_port_axi4_0_aw_valid = cbus__EVAL_110;
  assign plic__EVAL_72 = int_bus__EVAL_57;
  assign front_port_axi4_0_aw_ready = fbus__EVAL_21;
  assign mbus__EVAL_54 = shrinker__EVAL_25;
  assign sbus__EVAL_21 = tile__EVAL_108;
  assign plic__EVAL_73 = int_bus__EVAL_239;
  assign sys_port_axi4_0_ar_bits_cache = sbus__EVAL_8;
  assign mbus__EVAL_35 = mem_port_axi4_0_w_ready;
  assign cbus__EVAL_131 = plic__EVAL_15;
  assign plic__EVAL_67 = int_bus__EVAL_138;
  assign front_port_axi4_0_w_ready = fbus__EVAL_36;
  assign sbus__EVAL_0 = tile__EVAL_46;
  assign plic__EVAL_36 = int_bus__EVAL_177;
  assign ww__EVAL_2 = bh__EVAL_36;
  assign dtm__EVAL_16 = debug_systemjtag_jtag_TDI;
  assign front_port_axi4_0_r_bits_id = fbus__EVAL_17;
  assign int_bus__EVAL_217 = global_interrupts[71];
  assign shrinker__EVAL_24 = reset;
  assign mem_port_axi4_0_w_bits_last = mbus__EVAL_9;
  assign cbus__EVAL_80 = testIndicator_auto_in_d_bits_opcode;
  assign sbus__EVAL_163 = cbus__EVAL_118;
  assign sys_port_axi4_0_w_valid = sbus__EVAL_218;
  assign cbus__EVAL_85 = plic__EVAL_3;
  assign ww__EVAL_36 = shrinker__EVAL_4;
  assign plic__EVAL_46 = int_bus__EVAL_167;
  assign int_bus__EVAL_121 = global_interrupts[40];
  assign debug_1__EVAL_20 = fbus__EVAL_38;
  assign plic__EVAL_144 = int_bus__EVAL_190;
  assign clint__EVAL_16 = cbus__EVAL_114;
  assign sbus__EVAL_98 = sys_port_axi4_0_r_valid;
  assign plic__EVAL_43 = int_bus__EVAL_140;
  assign int_bus__EVAL_72 = global_interrupts[49];
  assign tile__EVAL_31 = sbus__EVAL;
  assign debug_1__EVAL_40 = dtm__EVAL_3;
  assign cbus__EVAL_117 = sbus__EVAL_33;
  assign sys_port_axi4_0_w_bits_last = sbus__EVAL_82;
  assign sbus__EVAL_44 = fbus__EVAL;
  assign shrinker__EVAL_9 = ww__EVAL_25;
  assign bh__EVAL_0 = sbus__EVAL_103;
  assign periph_port_axi4_0_aw_bits_qos = cbus__EVAL_76;
  assign plic__EVAL_81 = int_bus__EVAL_12;
  assign tile__EVAL_67 = _EVAL_0[0];
  assign plic__EVAL_103 = int_bus__EVAL_45;
  assign sagesafety__EVAL_9 = sbus__EVAL_193;
  assign plic__EVAL_74 = int_bus__EVAL_111;
  assign plic__EVAL_95 = int_bus__EVAL_241;
  assign shrinker__EVAL_26 = ww__EVAL_10;
  assign front_port_axi4_0_b_bits_resp = fbus__EVAL_59;
  assign dtm__EVAL_5 = debug_systemjtag_jtag_TMS;
  assign plic__EVAL_140 = int_bus__EVAL_87;
  assign mbus__EVAL_12 = mem_port_axi4_0_b_valid;
  assign int_bus__EVAL_120 = global_interrupts[52];
  assign sbus__EVAL_168 = tile__EVAL_25;
  assign testIndicator_auto_in_a_bits_mask = cbus__EVAL_123;
  assign int_bus__EVAL_134 = global_interrupts[53];
  assign sbus__EVAL_178 = bh__EVAL_25;
  assign int_bus__EVAL_251 = global_interrupts[77];
  assign cbus__EVAL_41 = periph_port_axi4_0_r_bits_resp;
  assign front_port_axi4_0_r_bits_data = fbus__EVAL_26;
  assign dtm__EVAL_12 = debug_1__EVAL_10;
  assign sys_port_axi4_0_aw_bits_addr = sbus__EVAL_72;
  assign sbus__EVAL_161 = bh__EVAL_44;
  assign cbus__EVAL_44 = periph_port_axi4_0_aw_ready;
  assign cbus__EVAL_128 = periph_port_axi4_0_ar_ready;
  assign plic__EVAL_42 = int_bus__EVAL_151;
  assign fbus__EVAL_28 = front_port_axi4_0_aw_bits_len;
  assign cbus__EVAL_33 = clint__EVAL_6;
  assign debug_1__EVAL_5 = fbus__EVAL_43;
  assign cbus__EVAL_7 = sbus__EVAL_38;
  assign shrinker__EVAL_27 = mbus__EVAL_8;
  assign cbus__EVAL_102 = sbus__EVAL_60;
  assign debug_1__EVAL_2 = cbus__EVAL_75;
  assign testIndicator_auto_in_a_bits_corrupt = cbus__EVAL_5;
  assign int_bus__EVAL_182 = global_interrupts[122];
  assign sbus__EVAL_45 = sagesafety__EVAL_11;
  assign cbus__EVAL_27 = tile__EVAL_56;
  assign sbus__EVAL_50 = cbus__EVAL_103;
  assign int_bus__EVAL_82 = global_interrupts[88];
  assign plic__EVAL_65 = int_bus__EVAL_10;
  assign sbus__EVAL_101 = sagesafety__EVAL_23;
  assign intsource__EVAL = reset;
  assign shrinker__EVAL_1 = ww__EVAL_18;
  assign debug_1__EVAL_18 = cbus__EVAL_60;
  assign sbus__EVAL_123 = tile__EVAL_52;
  assign int_bus__EVAL_131 = global_interrupts[106];
  assign sbus__EVAL_46 = sys_port_axi4_0_b_valid;
  assign int_bus__EVAL_83 = global_interrupts[13];
  assign ww__EVAL_30 = bh__EVAL_45;
  assign sagesafety__EVAL_35 = sbus__EVAL_202;
  assign tile__EVAL_83 = cbus__EVAL_111;
  assign sbus__EVAL_41 = tile__EVAL_20;
  assign int_bus__EVAL_171 = global_interrupts[125];
  assign plic__EVAL_80 = int_bus__EVAL_125;
  assign sbus__EVAL_10 = tile__EVAL_81;
  assign sagesafety__EVAL_33 = sbus__EVAL_185;
  assign sagesafety__EVAL_7 = sbus__EVAL_29;
  assign sbus__EVAL_90 = sagesafety__EVAL_22;
  assign testIndicator_auto_in_a_bits_param = cbus__EVAL_126;
  assign int_bus__EVAL_123 = global_interrupts[119];
  assign testIndicator_auto_in_a_bits_opcode = cbus__EVAL_155;
  assign plic__EVAL_60 = int_bus__EVAL_22;
  assign int_bus__EVAL_178 = global_interrupts[60];
  assign front_port_axi4_0_r_valid = fbus__EVAL_25;
  assign mem_port_axi4_0_w_bits_data = mbus__EVAL_19;
  assign plic__EVAL_120 = int_bus__EVAL_148;
  assign clint__EVAL_1 = cbus__EVAL_134;
  assign cbus__EVAL_1 = testIndicator_auto_in_d_bits_size;
  assign periph_port_axi4_0_ar_bits_lock = cbus__EVAL_11;
  assign debug_1__EVAL_3 = fbus__EVAL_54;
  assign sys_port_axi4_0_ar_bits_burst = sbus__EVAL_215;
  assign sbus__EVAL_143 = tile__EVAL_106;
  assign cbus__EVAL_127 = plic__EVAL_62;
  assign plic__EVAL_119 = int_bus__EVAL_185;
  assign testIndicator_auto_in_a_bits_source = cbus__EVAL_113;
  assign int_bus__EVAL_40 = global_interrupts[26];
  assign tile__EVAL_38 = reset_vector_0;
  assign tile__EVAL_8 = cbus__EVAL_14;
  assign int_bus__EVAL_238 = global_interrupts[110];
  assign sagesafety__EVAL_2 = sbus__EVAL_80;
  assign bh__EVAL_52 = sbus__EVAL_154;
  assign fbus__EVAL_58 = front_port_axi4_0_w_bits_data;
  assign int_bus__EVAL_30 = global_interrupts[46];
  assign debug_1__EVAL_4 = dtm__EVAL_13;
  assign plic__EVAL_48 = int_bus__EVAL_66;
  assign cbus__EVAL_77 = clint__EVAL_9;
  assign int_bus__EVAL_250 = global_interrupts[91];
  assign tile__EVAL_74 = sbus__EVAL_83;
  assign sbus__EVAL_151 = tile__EVAL_62;
  assign testIndicator_reset = reset;
  assign fbus__EVAL_46 = debug_1__EVAL_25;
  assign sbus__EVAL_67 = cbus__EVAL_119;
  assign sbus__EVAL_89 = tile__EVAL_88;
  assign mem_port_axi4_0_aw_bits_burst = mbus__EVAL_41;
  assign cbus__EVAL_98 = sbus__EVAL_139;
  assign plic__EVAL_16 = int_bus__EVAL_75;
  assign plic__EVAL_109 = int_bus__EVAL_247;
  assign fbus__EVAL_9 = clock;
  assign int_bus__EVAL_36 = global_interrupts[123];
  assign SynchronizerShiftReg_w1_d3__EVAL_1 = clock;
  assign debug_1__EVAL_0 = debug_systemjtag_jtag_TCK;
  assign mbus__EVAL_0 = shrinker__EVAL_14;
  assign sagesafety__EVAL_40 = sbus__EVAL_58;
  assign tile__EVAL_30 = sbus__EVAL_174;
  assign mem_port_axi4_0_w_bits_corrupt = mbus__EVAL_18;
  assign sbus__EVAL_209 = tile__EVAL_96;
  assign bh__EVAL_33 = clock;
  assign plic__EVAL_85 = int_bus__EVAL_172;
  assign plic__EVAL_116 = int_bus__EVAL_133;
  assign cbus__EVAL_45 = sbus__EVAL_217;
  assign mem_port_axi4_0_ar_bits_size = mbus__EVAL_29;
  assign plic__EVAL_68 = int_bus__EVAL_219;
  assign sbus__EVAL_28 = sagesafety__EVAL_13;
  assign periph_port_axi4_0_aw_bits_cache = cbus__EVAL_148;
  assign sbus__EVAL_7 = tile__EVAL_105;
  assign sagesafety__EVAL_38 = sbus__EVAL_63;
  assign sbus__EVAL_173 = fbus__EVAL_47;
  assign plic__EVAL_0 = int_bus__EVAL_109;
  assign int_bus__EVAL_43 = global_interrupts[4];
  assign int_bus__EVAL_110 = global_interrupts[87];
  assign bh__EVAL_11 = ww__EVAL_7;
  assign sbus__EVAL_114 = bh__EVAL_29;
  assign cbus__EVAL_107 = debug_1__EVAL_23;
  assign sbus__EVAL_91 = tile__EVAL_87;
  assign cbus__EVAL_159 = tile__EVAL_77;
  assign clint__EVAL_13 = cbus__EVAL_19;
  assign int_bus__EVAL_246 = global_interrupts[74];
  assign sagesafety__EVAL_6 = sbus__EVAL_81;
  assign sbus__EVAL_159 = reset;
  assign int_bus__EVAL_184 = global_interrupts[99];
  assign cbus__EVAL_94 = tile__EVAL_114;
  assign debug_1__EVAL_19 = cbus__EVAL_154;
  assign periph_port_axi4_0_aw_bits_burst = cbus__EVAL_24;
  assign ww__EVAL_21 = shrinker__EVAL_3;
  assign plic__EVAL_99 = int_bus__EVAL_203;
  assign sbus__EVAL_88 = sagesafety__EVAL_21;
  assign plic__EVAL_30 = int_bus__EVAL_145;
  assign plic__EVAL_9 = int_bus__EVAL_196;
  assign mbus__EVAL_14 = shrinker__EVAL_5;
  assign fbus__EVAL_40 = sbus__EVAL_188;
  assign tile__EVAL_28 = cbus__EVAL_74;
  assign plic__EVAL_105 = reset;
  assign bh__EVAL_23 = sbus__EVAL_140;
  assign int_bus__EVAL_149 = global_interrupts[108];
  assign int_bus__EVAL_194 = global_interrupts[68];
  assign int_bus__EVAL_73 = global_interrupts[27];
  assign sbus__EVAL_189 = tile__EVAL_4;
  assign tile__EVAL_78 = sbus__EVAL_71;
  assign plic__EVAL_41 = int_bus__EVAL_152;
  assign dtm__EVAL_6 = debug_systemjtag_mfr_id;
  assign clint__EVAL_18 = cbus__EVAL_135;
  assign int_bus__EVAL_221 = global_interrupts[117];
  assign plic__EVAL_136 = int_bus__EVAL_141;
  assign sbus__EVAL_150 = sys_port_axi4_0_w_ready;
  assign int_bus__EVAL_228 = global_interrupts[101];
  assign plic__EVAL_47 = int_bus__EVAL_119;
  assign int_bus__EVAL_29 = global_interrupts[45];
  assign fbus__EVAL_55 = front_port_axi4_0_r_ready;
  assign sbus__EVAL_169 = cbus__EVAL_129;
  assign plic__EVAL_126 = int_bus__EVAL_71;
  assign tile__EVAL_9 = intsource__EVAL_4;
  assign plic__EVAL_45 = int_bus__EVAL_232;
  assign int_bus__EVAL_9 = global_interrupts[70];
  assign tile__EVAL_32 = reset;
  assign plic__EVAL_92 = int_bus__EVAL_15;
  assign dtm__EVAL_8 = debug_1__EVAL_13;
  assign bh__EVAL_4 = ww__EVAL_27;
  assign shrinker__EVAL_10 = ww__EVAL_3;
  assign dmiResetCatch__EVAL = debug_systemjtag_reset;
  assign sagesafety__EVAL_4 = sbus__EVAL_125;
  assign sbus__EVAL_149 = sys_port_axi4_0_ar_ready;
  assign shrinker__EVAL_12 = mbus__EVAL_10;
  assign int_bus__EVAL_197 = global_interrupts[44];
  assign mem_port_axi4_0_aw_bits_lock = mbus__EVAL;
  assign cbus__EVAL_89 = tile__EVAL_85;
  assign plic__EVAL_117 = int_bus__EVAL_200;
  assign intsource__EVAL_3 = clint__EVAL_0;
  assign int_bus__EVAL_226 = global_interrupts[20];
  assign mem_port_axi4_0_ar_bits_cache = mbus__EVAL_3;
  assign cbus__EVAL_50 = plic__EVAL_38;
  assign cbus__EVAL_145 = debug_1__EVAL;
  assign cbus__EVAL_122 = testIndicator_auto_in_d_valid;
  assign sys_port_axi4_0_ar_bits_qos = sbus__EVAL_109;
  assign int_bus__EVAL_69 = global_interrupts[39];
  assign ww__EVAL_32 = bh__EVAL_43;
  assign tile__EVAL_42 = sbus__EVAL_113;
  assign tile__EVAL_41 = sbus__EVAL_176;
  assign ww__EVAL_12 = shrinker__EVAL_18;
  assign testIndicator_clock = clock;
  assign cbus__EVAL_72 = clint__EVAL_5;
  assign ww__EVAL_15 = reset;
  assign debug_1__EVAL_35 = dtm__EVAL_15;
  assign bh__EVAL_46 = sbus__EVAL_25;
  assign sbus__EVAL_35 = tile__EVAL_73;
  assign int_bus__EVAL_55 = global_interrupts[83];
  assign plic__EVAL_20 = cbus__EVAL_97;
  assign tile__EVAL_75 = sbus__EVAL_214;
  assign plic__EVAL_97 = int_bus__EVAL_90;
  assign cbus__EVAL_29 = tile__EVAL_5;
  assign sys_port_axi4_0_aw_bits_size = sbus__EVAL_224;
  assign tile__EVAL_80 = debug_1__EVAL_43;
  assign int_bus__EVAL_19 = global_interrupts[78];
  assign plic__EVAL_57 = int_bus__EVAL_179;
  assign cbus__EVAL_82 = clock;
  assign mbus__EVAL_27 = shrinker__EVAL_13;
  assign sbus__EVAL_187 = tile__EVAL_82;
  assign sbus__EVAL_144 = tile__EVAL_69;
  assign int_bus__EVAL_173 = global_interrupts[36];
  assign plic__EVAL_131 = cbus__EVAL_88;
  assign plic__EVAL_6 = int_bus__EVAL_51;
  assign bh__EVAL = sbus__EVAL_200;
  assign plic__EVAL_49 = int_bus__EVAL_180;
  assign int_bus__EVAL_33 = global_interrupts[120];
  assign cbus__EVAL_140 = sbus__EVAL_119;
  assign int_bus__EVAL_227 = global_interrupts[115];
  assign periph_port_axi4_0_ar_bits_burst = cbus__EVAL_73;
  assign int_bus__EVAL_54 = global_interrupts[85];
  assign sbus__EVAL_199 = sagesafety__EVAL_12;
  assign int_bus__EVAL_49 = global_interrupts[90];
  assign sbus__EVAL_207 = bh__EVAL_42;
  assign sbus__EVAL_190 = sagesafety__EVAL_37;
  assign tile__EVAL_12 = cbus__EVAL_101;
  assign int_bus__EVAL_222 = global_interrupts[2];
  assign sbus__EVAL_211 = sagesafety__EVAL_14;
  assign ww__EVAL_14 = bh__EVAL_50;
  assign sbus__EVAL_31 = sys_port_axi4_0_r_bits_last;
  assign int_bus__EVAL_95 = global_interrupts[15];
  assign sbus__EVAL_191 = tile__EVAL_33;
  assign debug_1__EVAL_21 = debug_psd_test_mode;
  assign front_port_axi4_0_b_valid = fbus__EVAL_39;
  assign bh__EVAL_47 = sbus__EVAL_121;
  assign periph_port_axi4_0_ar_valid = cbus__EVAL_143;
  assign int_bus__EVAL_70 = global_interrupts[8];
  assign sagesafety__EVAL_29 = sbus__EVAL_183;
  assign fbus__EVAL_24 = sbus__EVAL_53;
  assign debug_1__EVAL_12 = fbus__EVAL_27;
  assign cbus__EVAL_146 = testIndicator_auto_in_a_ready;
  assign bh__EVAL_53 = sbus__EVAL_136;
  assign dmiResetCatch__EVAL_2 = debug_psd_test_mode_reset;
  assign cbus__EVAL_0 = tile__EVAL_117;
  assign debug_systemjtag_jtag_TDO_driven = dtm__EVAL_10;
  assign sagesafety__EVAL_31 = sbus__EVAL_57;
  assign shrinker__EVAL_17 = clock;
  assign debug_systemjtag_jtag_TDO_data = dtm__EVAL_4;
  assign plic__EVAL_34 = int_bus__EVAL_102;
  assign int_bus__EVAL_28 = global_interrupts[105];
  assign int_bus__EVAL_168 = global_interrupts[63];
  assign plic__EVAL_71 = int_bus__EVAL_80;
  assign tile__EVAL_36 = cbus__EVAL_26;
  assign mbus__EVAL_52 = mem_port_axi4_0_r_valid;
  assign sagesafety__EVAL_32 = sbus__EVAL_111;
  assign fbus__EVAL_3 = front_port_axi4_0_w_bits_last;
  assign plic__EVAL_40 = int_bus__EVAL_156;
  assign fbus__EVAL_60 = sbus__EVAL_205;
  assign bh__EVAL_37 = sbus__EVAL_78;
  assign plic__EVAL_90 = int_bus__EVAL_106;
  assign periph_port_axi4_0_ar_bits_qos = cbus__EVAL_34;
  assign sbus__EVAL_104 = fbus__EVAL_0;
  assign sbus__EVAL_172 = bh__EVAL_31;
  assign cbus__EVAL_109 = periph_port_axi4_0_b_bits_resp;
  assign sys_port_axi4_0_aw_bits_prot = sbus__EVAL_49;
  assign sbus__EVAL_34 = tile__EVAL_93;
  assign shrinker__EVAL_0 = mbus__EVAL_20;
  assign plic__EVAL_11 = int_bus__EVAL_187;
  assign plic__EVAL_22 = int_bus__EVAL_86;
  assign sbus__EVAL_2 = sagesafety__EVAL_36;
  assign sbus__EVAL_17 = tile__EVAL_17;
  assign sbus__EVAL_76 = fbus__EVAL_19;
  assign sbus__EVAL_95 = tile__EVAL_37;
  assign mem_port_axi4_0_r_ready = mbus__EVAL_31;
  assign sbus__EVAL_135 = cbus__EVAL_71;
  assign tile__EVAL_98 = cbus__EVAL_70;
  assign sbus__EVAL_4 = bh__EVAL_27;
  assign int_bus__EVAL_92 = global_interrupts[31];
  assign int_bus__EVAL_96 = global_interrupts[75];
  assign sbus__EVAL_126 = bh__EVAL_5;
  assign periph_port_axi4_0_w_bits_last = cbus__EVAL_43;
  assign tile__EVAL_107 = sbus__EVAL_107;
  assign tile__EVAL_0 = sbus__EVAL_164;
  assign debug_1__EVAL_38 = cbus__EVAL_22;
  assign int_bus__EVAL_215 = global_interrupts[113];
  assign int_bus__EVAL_1 = global_interrupts[10];
  assign int_bus__EVAL_139 = global_interrupts[55];
  assign int_bus__EVAL_130 = global_interrupts[84];
  assign plic__EVAL_4 = int_bus__EVAL_188;
  assign tile__EVAL_47 = intsource__EVAL_1;
  assign int_bus__EVAL_3 = global_interrupts[14];
  assign clint__EVAL_19 = cbus__EVAL_157;
  assign bh__EVAL_24 = sbus__EVAL_160;
  assign sbus__EVAL_43 = bh__EVAL_41;
  assign periph_port_axi4_0_ar_bits_len = cbus__EVAL_79;
  assign plic__EVAL_52 = int_bus__EVAL_84;
  assign int_bus__EVAL_7 = global_interrupts[42];
  assign int_bus__EVAL_245 = global_interrupts[104];
  assign plic__EVAL_121 = int_bus__EVAL_191;
  assign sagesafety__EVAL_20 = sbus__EVAL_156;
  assign plic__EVAL_112 = int_bus__EVAL_94;
  assign debug_1__EVAL_27 = cbus__EVAL_46;
  assign int_bus__EVAL_21 = global_interrupts[38];
  assign fbus__EVAL_35 = front_port_axi4_0_aw_bits_size;
  assign mbus__EVAL_50 = mem_port_axi4_0_r_bits_resp;
  assign mbus__EVAL_28 = mem_port_axi4_0_b_bits_resp;
  assign tile__EVAL_89 = cbus__EVAL_69;
  assign plic__EVAL_50 = int_bus__EVAL_108;
  assign bh__EVAL_19 = reset;
  assign cbus__EVAL_63 = tile__EVAL_92;
  assign plic__EVAL_141 = int_bus__EVAL_135;
  assign sbus__EVAL_110 = tile__EVAL_13;
  assign cbus__EVAL_12 = periph_port_axi4_0_b_valid;
  assign tile__EVAL_55 = cbus__EVAL_3;
  assign bh__EVAL_17 = sbus__EVAL_155;
  assign mem_port_axi4_0_ar_bits_id = mbus__EVAL_49;
  assign int_bus__EVAL_41 = global_interrupts[19];
  assign plic__EVAL_82 = int_bus__EVAL_115;
  assign bh__EVAL_13 = ww__EVAL_31;
  assign int_bus__EVAL_189 = global_interrupts[103];
  assign plic__EVAL_122 = int_bus__EVAL_249;
  assign clint__EVAL_10 = clock;
  assign plic__EVAL_61 = int_bus__EVAL_234;
  assign dtm__EVAL_14 = debug_systemjtag_jtag_TCK;
  assign cbus__EVAL_53 = sbus__EVAL_32;
  assign cbus__EVAL_30 = tile__EVAL_95;
  assign sagesafety__EVAL_16 = sbus__EVAL_87;
  assign sbus__EVAL_182 = sagesafety__EVAL_1;
  assign int_bus__EVAL_153 = global_interrupts[100];
  assign plic__EVAL_77 = int_bus__EVAL_164;
  assign debug_1__EVAL_39 = dmiResetCatch__EVAL_0;
  assign testIndicator_auto_in_a_bits_size = cbus__EVAL_39;
  assign int_bus__EVAL_199 = global_interrupts[41];
  assign dtm__EVAL_1 = debug_1__EVAL_36;
  assign plic__EVAL_13 = int_bus__EVAL_97;
  assign sbus__EVAL_222 = tile__EVAL_109;
  assign sbus__EVAL_99 = sagesafety__EVAL_10;
  assign plic__EVAL_37 = int_bus__EVAL_107;
  assign sys_port_axi4_0_w_bits_strb = sbus__EVAL_196;
  assign plic__EVAL_78 = int_bus__EVAL_183;
  assign int_bus__EVAL_67 = global_interrupts[82];
  assign int_bus__EVAL_132 = global_interrupts[34];
  assign int_bus__EVAL_158 = global_interrupts[23];
  assign sbus__EVAL_145 = tile__EVAL_27;
  assign tile__EVAL_90 = cbus__EVAL_108;
  assign cbus__EVAL_67 = tile__EVAL_97;
  assign sbus__EVAL_108 = cbus__EVAL_10;
  assign plic__EVAL_98 = int_bus__EVAL_174;
  assign int_bus__EVAL_50 = global_interrupts[98];
  assign ww__EVAL_4 = shrinker__EVAL_2;
  assign debug_1__EVAL_41 = cbus__EVAL_112;
  assign periph_port_axi4_0_ar_bits_prot = cbus__EVAL_35;
  assign fbus__EVAL_50 = sbus__EVAL_84;
  assign testIndicator_auto_in_d_ready = cbus__EVAL_6;
  assign tile__EVAL_115 = sbus__EVAL_206;
  assign mem_port_axi4_0_aw_bits_cache = mbus__EVAL_5;
  assign int_bus__EVAL_61 = global_interrupts[7];
  assign int_bus__EVAL_114 = global_interrupts[21];
  assign tile__EVAL_45 = sbus__EVAL_184;
  assign fbus__EVAL_23 = front_port_axi4_0_ar_bits_addr;
  assign shrinker__EVAL_33 = mbus__EVAL_46;
  assign clint__EVAL_15 = cbus__EVAL_91;
  assign SynchronizerShiftReg_w1_d3__EVAL = rtc_toggle;
  assign bh__EVAL_30 = sbus__EVAL_39;
  assign int_bus__EVAL_25 = global_interrupts[48];
  assign cbus__EVAL_62 = tile__EVAL_43;
  assign sbus__EVAL_115 = tile__EVAL_76;
  assign testIndicator_auto_in_a_valid = cbus__EVAL_38;
  assign int_bus__EVAL_23 = global_interrupts[6];
  assign int_bus__EVAL_105 = global_interrupts[111];
  assign debug_1__EVAL_33 = dtm__EVAL_9;
  assign sbus__EVAL_203 = sagesafety__EVAL_17;
  assign sys_port_axi4_0_aw_bits_id = sbus__EVAL_36;
  assign int_bus__EVAL = global_interrupts[66];
  assign debug_1__EVAL_31 = reset;
  assign tile__EVAL_84 = cbus__EVAL_156;
  assign sbus__EVAL_130 = bh__EVAL_35;
  assign plic__EVAL_66 = int_bus__EVAL_150;
  assign periph_port_axi4_0_aw_bits_lock = cbus__EVAL_158;
  assign sys_port_axi4_0_aw_bits_lock = sbus__EVAL_52;
  assign bh__EVAL_12 = sbus__EVAL_3;
  assign mbus__EVAL_56 = mem_port_axi4_0_aw_ready;
  assign sagesafety__EVAL_26 = sbus__EVAL_171;
  assign cbus__EVAL_42 = tile__EVAL_1;
  assign sbus__EVAL_5 = sagesafety__EVAL_15;
  assign plic__EVAL_100 = int_bus__EVAL_218;
  assign front_port_axi4_0_r_bits_resp = fbus__EVAL_29;
  assign ww__EVAL_33 = bh__EVAL_18;
  assign sys_port_axi4_0_ar_bits_len = sbus__EVAL_15;
  assign periph_port_axi4_0_ar_bits_cache = cbus__EVAL_56;
  assign int_bus__EVAL_77 = global_interrupts[50];
  assign int_bus__EVAL_162 = global_interrupts[96];
  assign ww__EVAL_5 = bh__EVAL_14;
  assign sbus__EVAL_27 = fbus__EVAL_15;
  assign cbus__EVAL_138 = testIndicator_auto_in_d_bits_source;
  assign cbus__EVAL_20 = debug_1__EVAL_26;
  assign plic__EVAL_10 = int_bus__EVAL_213;
  assign tile__EVAL_86 = sbus__EVAL_51;
  assign cbus__EVAL_25 = tile__EVAL_113;
  assign sagesafety__EVAL_5 = sbus__EVAL_152;
  assign fbus__EVAL_31 = front_port_axi4_0_ar_bits_id;
  assign plic__EVAL_89 = int_bus__EVAL_165;
  assign clint__EVAL = cbus__EVAL_55;
  assign cbus__EVAL_130 = periph_port_axi4_0_w_ready;
  assign bh__EVAL_22 = ww__EVAL_16;
  assign sbus__EVAL_197 = tile__EVAL_3;
  assign fbus__EVAL_51 = sbus__EVAL_141;
  assign int_bus__EVAL_205 = global_interrupts[81];
  assign intsource__EVAL_2 = clint__EVAL_12;
  assign plic__EVAL_128 = int_bus__EVAL_240;
  assign int_bus__EVAL_56 = global_interrupts[11];
  assign int_bus__EVAL_48 = global_interrupts[43];
  assign plic__EVAL_63 = int_bus__EVAL_147;
  assign int_bus__EVAL_24 = global_interrupts[24];
  assign plic__EVAL_123 = int_bus__EVAL_128;
  assign plic__EVAL_142 = clock;
  assign cbus__EVAL_137 = tile__EVAL_49;
  assign mbus__EVAL_6 = mem_port_axi4_0_ar_ready;
  assign debug_ndreset = debug_1__EVAL_8;
  assign plic__EVAL_27 = int_bus__EVAL_34;
  assign periph_port_axi4_0_ar_bits_addr = cbus__EVAL_18;
  assign mbus__EVAL_33 = shrinker__EVAL_6;
  assign periph_port_axi4_0_ar_bits_size = cbus__EVAL_93;
  assign cbus__EVAL_51 = tile__EVAL_65;
  assign intsource_1__EVAL_2 = plic__EVAL_138;
  assign cbus__EVAL_124 = clint__EVAL_4;
  assign clint__EVAL_17 = cbus__EVAL_61;
  assign clint__EVAL_11 = reset;
  assign intsource_1__EVAL_1 = reset;
  assign cbus__EVAL_90 = reset;
  assign cbus__EVAL_31 = tile__EVAL_58;
  assign cbus__EVAL_23 = sbus__EVAL_181;
  assign int_bus__EVAL_100 = global_interrupts[107];
  assign shrinker__EVAL_19 = mbus__EVAL_38;
  assign mem_port_axi4_0_w_bits_strb = mbus__EVAL_36;
  assign plic__EVAL_101 = int_bus__EVAL_85;
  assign mem_port_axi4_0_ar_bits_len = mbus__EVAL_16;
  assign int_bus__EVAL_248 = global_interrupts[67];
  assign plic__EVAL_134 = int_bus__EVAL_32;
  assign tile__EVAL_14 = sbus__EVAL_13;
  assign cbus__EVAL_58 = clint__EVAL_8;
  assign tile__EVAL_2 = sbus__EVAL_146;
  assign sagesafety__EVAL_0 = clock;
  assign int_bus__EVAL_210 = global_interrupts[121];
  assign mbus__EVAL_53 = clock;
  assign plic__EVAL_139 = int_bus__EVAL_237;
  assign sbus__EVAL_133 = tile__EVAL_35;
  assign periph_port_axi4_0_w_bits_strb = cbus__EVAL_99;
  assign plic__EVAL_58 = cbus__EVAL_96;
  assign plic__EVAL_129 = int_bus__EVAL_230;
  assign sagesafety__EVAL_24 = sbus__EVAL_9;
  assign fbus__EVAL_4 = front_port_axi4_0_w_valid;
  assign sys_port_axi4_0_ar_bits_size = sbus__EVAL_23;
  assign plic__EVAL_14 = int_bus__EVAL_157;
  assign int_bus__EVAL_53 = global_interrupts[94];
  assign int_bus__EVAL_62 = global_interrupts[93];
  assign tile__EVAL_102 = sbus__EVAL_213;
  assign intsource_1__EVAL = clock;
  assign int_bus__EVAL_5 = global_interrupts[33];
  assign intsource__EVAL_0 = clock;
  assign periph_port_axi4_0_ar_bits_id = cbus__EVAL_142;
  assign tile__EVAL_68 = sbus__EVAL_19;
  assign mbus__EVAL_40 = mem_port_axi4_0_b_bits_id;
  assign plic__EVAL_135 = int_bus__EVAL_169;
  assign clint__EVAL_7 = _EVAL_4;
  assign int_bus__EVAL_8 = global_interrupts[118];
  assign tile__EVAL_100 = core_clock_0;
  assign tile__EVAL_91 = sbus__EVAL_55;
  assign tile__EVAL_104 = cbus__EVAL_32;
  assign cbus__EVAL_121 = tile__EVAL_118;
  assign fbus__EVAL_34 = front_port_axi4_0_ar_bits_burst;
  assign bh__EVAL_3 = sbus__EVAL_148;
  assign plic__EVAL_44 = int_bus__EVAL_186;
  assign plic__EVAL_64 = int_bus__EVAL_154;
  assign dtm__EVAL = debug_systemjtag_reset;
  assign int_bus__EVAL_235 = global_interrupts[12];
  assign sys_port_axi4_0_ar_valid = sbus__EVAL_219;
  assign clint__EVAL_2 = cbus__EVAL_92;
  assign bh__EVAL_20 = sbus__EVAL_65;
  assign dmiResetCatch__EVAL_1 = debug_systemjtag_jtag_TCK;
  assign front_port_axi4_0_r_bits_last = fbus__EVAL_53;
  assign plic__EVAL_24 = int_bus__EVAL_155;
  assign plic__EVAL_107 = int_bus__EVAL_35;
  assign int_bus__EVAL_101 = global_interrupts[54];
  assign debug_1__EVAL_15 = cbus__EVAL;
  assign mbus__EVAL_1 = shrinker__EVAL_35;
  assign plic__EVAL_96 = int_bus__EVAL_252;
  assign bh__EVAL_32 = ww__EVAL_0;
  assign periph_port_axi4_0_aw_bits_addr = cbus__EVAL_100;
  assign int_bus__EVAL_52 = global_interrupts[124];
  assign tile__EVAL_50 = sbus__EVAL_180;
  assign plic__EVAL_102 = int_bus__EVAL_39;
  assign int_bus__EVAL_14 = global_interrupts[73];
  assign mem_port_axi4_0_ar_bits_qos = mbus__EVAL_44;
  assign sbus__EVAL_128 = cbus__EVAL_115;
  assign plic__EVAL_76 = int_bus__EVAL_126;
  assign sys_port_axi4_0_ar_bits_id = sbus__EVAL_175;
  assign tile__EVAL_64 = sbus__EVAL_124;
  assign ww__EVAL_6 = shrinker__EVAL_34;
  assign plic__EVAL_113 = int_bus__EVAL_38;
  assign plic__EVAL_127 = int_bus__EVAL_243;
  assign plic__EVAL_94 = int_bus__EVAL_236;
  assign plic__EVAL_111 = int_bus__EVAL_176;
  assign plic__EVAL_5 = int_bus__EVAL_0;
  assign fbus__EVAL_49 = sbus__EVAL_195;
  assign debug_1__EVAL_9 = dtm__EVAL_7;
  assign ww__EVAL_1 = bh__EVAL_9;
  assign int_bus__EVAL_20 = global_interrupts[16];
  assign sbus__EVAL_118 = fbus__EVAL_20;
  assign dtm__EVAL_0 = dtm__EVAL_11;
  assign int_bus__EVAL_60 = global_interrupts[61];
  assign sbus__EVAL_194 = fbus__EVAL_14;
  assign cbus__EVAL_153 = tile__EVAL_44;
  assign plic__EVAL_53 = int_bus__EVAL_93;
  assign sagesafety__EVAL_27 = sbus__EVAL_20;
  assign sbus__EVAL_86 = bh__EVAL_6;
  assign plic__EVAL_106 = int_bus__EVAL_206;
  assign sbus__EVAL_210 = tile__EVAL_16;
  assign plic__EVAL_18 = int_bus__EVAL_181;
  assign plic__EVAL_79 = cbus__EVAL_152;
  assign plic__EVAL_25 = int_bus__EVAL_113;
  assign cbus__EVAL_104 = tile__EVAL_23;
  assign periph_port_axi4_0_aw_bits_len = cbus__EVAL_47;
  assign int_bus__EVAL_207 = global_interrupts[17];
  assign cbus__EVAL_105 = tile__EVAL_60;
  assign fbus__EVAL_16 = sbus__EVAL_132;
  assign tile__EVAL_24 = intsource_1__EVAL_0;
  assign plic__EVAL_54 = int_bus__EVAL_198;
  assign mbus__EVAL_42 = mem_port_axi4_0_r_bits_id;
  assign bh__EVAL_49 = sbus__EVAL_102;
  assign dmiResetCatch__EVAL_3 = debug_psd_test_mode;
  assign sys_port_axi4_0_ar_bits_addr = sbus__EVAL_30;
  assign plic__EVAL_8 = int_bus__EVAL_224;
  assign tile__EVAL_101 = cbus__EVAL_139;
  assign fbus__EVAL_18 = sbus__EVAL_208;
  assign bh__EVAL_10 = sbus__EVAL_212;
  assign tile__EVAL_22 = cbus__EVAL_133;
  assign fbus__EVAL_57 = sbus__EVAL_165;
  assign tile__EVAL_48 = cbus__EVAL_16;
  assign periph_port_axi4_0_aw_bits_id = cbus__EVAL_106;
  assign int_bus__EVAL_42 = global_interrupts[65];
  assign debug_dmactive = debug_1__EVAL_29;
  assign tile__EVAL_54 = sbus__EVAL_24;
  assign tile__EVAL_63 = cbus__EVAL_37;
  assign sbus__EVAL_16 = tile__EVAL;
  assign plic__EVAL_125 = int_bus__EVAL_223;
  assign sbus__EVAL_47 = sys_port_axi4_0_b_bits_id;
  assign bh__EVAL_7 = ww__EVAL_29;
  assign fbus__EVAL_7 = reset;
  assign ww__EVAL_8 = bh__EVAL_1;
  assign plic__EVAL_32 = int_bus__EVAL_137;
  assign int_bus__EVAL_175 = global_interrupts[47];
  assign int_bus__EVAL_117 = global_interrupts[95];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _EVAL_1 <= 1'h0;
    end else begin
      _EVAL_1 <= _EVAL_2;
    end
    if (reset) begin
      _EVAL_4 <= 1'h0;
    end else begin
      _EVAL_4 <= _EVAL;
    end
  end
endmodule
