//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_50_assert(
  input  [3:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [31:0] _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [5:0] _EVAL_29;
  reg [31:0] _RAND_0;
  reg [5:0] _EVAL_32;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_54;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_64;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_98;
  reg [31:0] _RAND_4;
  reg [1:0] _EVAL_105;
  reg [31:0] _RAND_5;
  reg  _EVAL_115;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_182;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_196;
  reg [31:0] _RAND_8;
  reg  _EVAL_208;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_258;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_259;
  reg [31:0] _RAND_11;
  reg  _EVAL_271;
  reg [31:0] _RAND_12;
  reg [3:0] _EVAL_276;
  reg [31:0] _RAND_13;
  wire [22:0] _EVAL_267;
  wire [7:0] _EVAL_163;
  wire [7:0] _EVAL_207;
  wire [31:0] _EVAL_217;
  wire [31:0] _EVAL_225;
  wire  _EVAL_265;
  wire  _EVAL_165;
  wire  _EVAL_19;
  wire [1:0] _EVAL_281;
  wire [1:0] _EVAL_286;
  wire  _EVAL_173;
  wire  _EVAL_209;
  wire  _EVAL_223;
  wire  _EVAL_190;
  wire  _EVAL_268;
  wire  _EVAL_184;
  wire  _EVAL_224;
  wire  _EVAL_49;
  wire  _EVAL_180;
  wire  _EVAL_23;
  wire  _EVAL_38;
  wire  _EVAL_44;
  wire  _EVAL_272;
  wire  _EVAL_28;
  wire  _EVAL_245;
  wire  _EVAL_31;
  wire  _EVAL_251;
  wire  _EVAL_123;
  wire  _EVAL_171;
  wire  _EVAL_97;
  wire  _EVAL_290;
  wire  _EVAL_253;
  wire [3:0] _EVAL_132;
  wire  _EVAL_140;
  wire  _EVAL_73;
  wire  _EVAL_229;
  wire  _EVAL_294;
  wire  _EVAL_128;
  wire [31:0] _EVAL_81;
  wire [32:0] _EVAL_242;
  wire [32:0] _EVAL_134;
  wire [32:0] _EVAL_186;
  wire  _EVAL_43;
  wire [31:0] _EVAL_187;
  wire [32:0] _EVAL_278;
  wire [32:0] _EVAL_269;
  wire [32:0] _EVAL_131;
  wire  _EVAL_66;
  wire  _EVAL_198;
  wire [31:0] _EVAL_84;
  wire [32:0] _EVAL_144;
  wire [32:0] _EVAL_289;
  wire [32:0] _EVAL_154;
  wire  _EVAL_254;
  wire  _EVAL_185;
  wire [31:0] _EVAL_26;
  wire [32:0] _EVAL_106;
  wire [32:0] _EVAL_239;
  wire [32:0] _EVAL_107;
  wire  _EVAL_136;
  wire  _EVAL_275;
  wire [32:0] _EVAL_55;
  wire [32:0] _EVAL_176;
  wire [32:0] _EVAL_193;
  wire  _EVAL_197;
  wire  _EVAL_141;
  wire [31:0] _EVAL_104;
  wire [32:0] _EVAL_243;
  wire [32:0] _EVAL_148;
  wire [32:0] _EVAL_47;
  wire  _EVAL_158;
  wire  _EVAL_287;
  wire  _EVAL_215;
  wire  _EVAL_279;
  wire  _EVAL_75;
  wire  _EVAL_74;
  wire  _EVAL_255;
  wire  _EVAL_175;
  wire  _EVAL_152;
  wire [1:0] _EVAL_210;
  wire  _EVAL_233;
  wire  _EVAL_129;
  wire  _EVAL_248;
  wire [5:0] _EVAL_189;
  wire  _EVAL_130;
  wire  _EVAL_153;
  wire  _EVAL_95;
  wire  _EVAL_234;
  wire  _EVAL_199;
  wire  _EVAL_249;
  wire  _EVAL_42;
  wire  _EVAL_204;
  wire  _EVAL_192;
  wire  _EVAL_201;
  wire [31:0] _EVAL_220;
  wire [32:0] _EVAL_113;
  wire [32:0] _EVAL_70;
  wire [32:0] _EVAL_69;
  wire  _EVAL_15;
  wire  _EVAL_45;
  wire [31:0] _EVAL_206;
  wire [32:0] _EVAL_33;
  wire [32:0] _EVAL_40;
  wire [32:0] _EVAL_147;
  wire  _EVAL_59;
  wire  _EVAL_296;
  wire  _EVAL_92;
  wire  _EVAL_82;
  wire  _EVAL_18;
  wire [31:0] _EVAL_178;
  wire [32:0] _EVAL_36;
  wire [32:0] _EVAL_120;
  wire [32:0] _EVAL_247;
  wire  _EVAL_86;
  wire  _EVAL_159;
  wire  _EVAL_266;
  wire  _EVAL_65;
  wire  _EVAL_91;
  wire  _EVAL_89;
  wire  _EVAL_126;
  wire  _EVAL_39;
  wire  _EVAL_149;
  wire  _EVAL_90;
  wire  _EVAL_241;
  wire  _EVAL_292;
  wire  _EVAL_218;
  wire [1:0] _EVAL_30;
  wire  _EVAL_121;
  wire  _EVAL_67;
  wire  _EVAL_211;
  wire  _EVAL_77;
  wire  _EVAL_219;
  wire  _EVAL_168;
  wire  _EVAL_116;
  wire  _EVAL_50;
  wire  _EVAL_53;
  wire  _EVAL_188;
  wire  _EVAL_122;
  wire  _EVAL_57;
  wire  _EVAL_135;
  wire  _EVAL_291;
  wire  _EVAL_203;
  wire  _EVAL_119;
  wire  _EVAL_227;
  wire [22:0] _EVAL_263;
  wire [7:0] _EVAL_112;
  wire [7:0] _EVAL_160;
  wire [5:0] _EVAL_257;
  wire [5:0] _EVAL_48;
  wire  _EVAL_34;
  wire  _EVAL_284;
  wire  _EVAL_195;
  wire  _EVAL_250;
  wire  _EVAL_191;
  wire [31:0] _EVAL_222;
  wire  _EVAL_143;
  wire  _EVAL_146;
  wire  _EVAL_183;
  wire  _EVAL_114;
  wire  _EVAL_238;
  wire  _EVAL_60;
  wire  _EVAL_221;
  wire  _EVAL_101;
  wire  _EVAL_200;
  wire  _EVAL_295;
  wire  _EVAL_63;
  wire  _EVAL_51;
  wire  _EVAL_216;
  wire [5:0] _EVAL_150;
  wire [5:0] _EVAL_181;
  wire  _EVAL_61;
  wire  _EVAL_80;
  wire [3:0] _EVAL_213;
  wire [3:0] _EVAL_274;
  wire  _EVAL_230;
  wire  _EVAL_280;
  wire  _EVAL_172;
  wire  _EVAL_85;
  wire  _EVAL_179;
  wire  _EVAL_205;
  wire  _EVAL_24;
  wire  _EVAL_137;
  wire  _EVAL_232;
  wire  _EVAL_293;
  wire  _EVAL_124;
  wire [5:0] _EVAL_283;
  wire  _EVAL_277;
  wire  _EVAL_273;
  wire  _EVAL_177;
  wire  _EVAL_164;
  wire [3:0] _EVAL_262;
  wire  _EVAL_68;
  wire  _EVAL_78;
  wire  _EVAL_118;
  wire  _EVAL_235;
  wire  _EVAL_155;
  wire  _EVAL_174;
  wire  _EVAL_151;
  wire  _EVAL_108;
  wire  _EVAL_297;
  wire  _EVAL_162;
  wire  _EVAL_261;
  wire  _EVAL_252;
  wire  _EVAL_41;
  wire  _EVAL_169;
  wire  _EVAL_288;
  wire  _EVAL_142;
  wire  _EVAL_46;
  wire  _EVAL_282;
  wire  _EVAL_35;
  wire  _EVAL_72;
  wire  _EVAL_37;
  wire  _EVAL_236;
  wire  _EVAL_56;
  wire  _EVAL_138;
  wire  _EVAL_170;
  wire  _EVAL_214;
  wire  _EVAL_167;
  wire  _EVAL_285;
  wire  _EVAL_260;
  wire  _EVAL_228;
  wire  _EVAL_157;
  wire  _EVAL_17;
  wire  _EVAL_83;
  wire  _EVAL_194;
  wire  _EVAL_87;
  wire  _EVAL_21;
  wire  _EVAL_212;
  wire  _EVAL_22;
  wire  _EVAL_240;
  wire  _EVAL_25;
  wire  _EVAL_161;
  wire  _EVAL_111;
  wire  _EVAL_99;
  wire  _EVAL_103;
  wire  _EVAL_226;
  wire  _EVAL_76;
  wire  _EVAL_133;
  wire  _EVAL_88;
  wire  _EVAL_117;
  wire  _EVAL_246;
  wire  _EVAL_100;
  wire  _EVAL_231;
  wire  _EVAL_145;
  wire  _EVAL_20;
  wire  _EVAL_264;
  wire  _EVAL_110;
  wire  _EVAL_109;
  wire  _EVAL_79;
  wire  _EVAL_102;
  wire  _EVAL_125;
  wire  _EVAL_62;
  wire  _EVAL_256;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_267 = 23'hff << _EVAL_4;
  assign _EVAL_163 = _EVAL_267[7:0];
  assign _EVAL_207 = ~ _EVAL_163;
  assign _EVAL_217 = {{24'd0}, _EVAL_207};
  assign _EVAL_225 = _EVAL_6 & _EVAL_217;
  assign _EVAL_265 = _EVAL_225 == 32'h0;
  assign _EVAL_165 = _EVAL_4 >= 4'h2;
  assign _EVAL_19 = _EVAL_4[0];
  assign _EVAL_281 = 2'h1 << _EVAL_19;
  assign _EVAL_286 = _EVAL_281 | 2'h1;
  assign _EVAL_173 = _EVAL_286[1];
  assign _EVAL_209 = _EVAL_6[1];
  assign _EVAL_223 = _EVAL_173 & _EVAL_209;
  assign _EVAL_190 = _EVAL_165 | _EVAL_223;
  assign _EVAL_268 = _EVAL_286[0];
  assign _EVAL_184 = _EVAL_6[0];
  assign _EVAL_224 = _EVAL_209 & _EVAL_184;
  assign _EVAL_49 = _EVAL_268 & _EVAL_224;
  assign _EVAL_180 = _EVAL_190 | _EVAL_49;
  assign _EVAL_23 = _EVAL_184 == 1'h0;
  assign _EVAL_38 = _EVAL_209 & _EVAL_23;
  assign _EVAL_44 = _EVAL_268 & _EVAL_38;
  assign _EVAL_272 = _EVAL_190 | _EVAL_44;
  assign _EVAL_28 = _EVAL_209 == 1'h0;
  assign _EVAL_245 = _EVAL_173 & _EVAL_28;
  assign _EVAL_31 = _EVAL_165 | _EVAL_245;
  assign _EVAL_251 = _EVAL_28 & _EVAL_184;
  assign _EVAL_123 = _EVAL_268 & _EVAL_251;
  assign _EVAL_171 = _EVAL_31 | _EVAL_123;
  assign _EVAL_97 = _EVAL_28 & _EVAL_23;
  assign _EVAL_290 = _EVAL_268 & _EVAL_97;
  assign _EVAL_253 = _EVAL_31 | _EVAL_290;
  assign _EVAL_132 = {_EVAL_180,_EVAL_272,_EVAL_171,_EVAL_253};
  assign _EVAL_140 = _EVAL_0 == _EVAL_132;
  assign _EVAL_73 = _EVAL_140 | _EVAL_11;
  assign _EVAL_229 = _EVAL_73 == 1'h0;
  assign _EVAL_294 = _EVAL_12 == 1'h0;
  assign _EVAL_128 = _EVAL_294 | _EVAL_11;
  assign _EVAL_81 = _EVAL_6 ^ 32'h40000000;
  assign _EVAL_242 = {1'b0,$signed(_EVAL_81)};
  assign _EVAL_134 = $signed(_EVAL_242) & $signed(-33'sh2000);
  assign _EVAL_186 = $signed(_EVAL_134);
  assign _EVAL_43 = $signed(_EVAL_186) == $signed(33'sh0);
  assign _EVAL_187 = _EVAL_6 ^ 32'h80000000;
  assign _EVAL_278 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_269 = $signed(_EVAL_278) & $signed(-33'sh20000);
  assign _EVAL_131 = $signed(_EVAL_269);
  assign _EVAL_66 = $signed(_EVAL_131) == $signed(33'sh0);
  assign _EVAL_198 = _EVAL_43 | _EVAL_66;
  assign _EVAL_84 = _EVAL_6 ^ 32'hc000000;
  assign _EVAL_144 = {1'b0,$signed(_EVAL_84)};
  assign _EVAL_289 = $signed(_EVAL_144) & $signed(-33'sh4000000);
  assign _EVAL_154 = $signed(_EVAL_289);
  assign _EVAL_254 = $signed(_EVAL_154) == $signed(33'sh0);
  assign _EVAL_185 = _EVAL_198 | _EVAL_254;
  assign _EVAL_26 = _EVAL_6 ^ 32'h2000000;
  assign _EVAL_106 = {1'b0,$signed(_EVAL_26)};
  assign _EVAL_239 = $signed(_EVAL_106) & $signed(-33'sh10000);
  assign _EVAL_107 = $signed(_EVAL_239);
  assign _EVAL_136 = $signed(_EVAL_107) == $signed(33'sh0);
  assign _EVAL_275 = _EVAL_185 | _EVAL_136;
  assign _EVAL_55 = {1'b0,$signed(_EVAL_6)};
  assign _EVAL_176 = $signed(_EVAL_55) & $signed(-33'sh5000);
  assign _EVAL_193 = $signed(_EVAL_176);
  assign _EVAL_197 = $signed(_EVAL_193) == $signed(33'sh0);
  assign _EVAL_141 = _EVAL_275 | _EVAL_197;
  assign _EVAL_104 = _EVAL_6 ^ 32'h1800000;
  assign _EVAL_243 = {1'b0,$signed(_EVAL_104)};
  assign _EVAL_148 = $signed(_EVAL_243) & $signed(-33'sh8000);
  assign _EVAL_47 = $signed(_EVAL_148);
  assign _EVAL_158 = $signed(_EVAL_47) == $signed(33'sh0);
  assign _EVAL_287 = _EVAL_141 | _EVAL_158;
  assign _EVAL_215 = _EVAL_1 != 2'h2;
  assign _EVAL_279 = _EVAL_215 | _EVAL_11;
  assign _EVAL_75 = _EVAL_279 == 1'h0;
  assign _EVAL_74 = _EVAL_4 <= 4'h2;
  assign _EVAL_255 = _EVAL_10 & _EVAL_5;
  assign _EVAL_175 = _EVAL_54 == 6'h0;
  assign _EVAL_152 = _EVAL_255 & _EVAL_175;
  assign _EVAL_210 = _EVAL_152 ? 2'h1 : 2'h0;
  assign _EVAL_233 = _EVAL_210[0];
  assign _EVAL_129 = _EVAL_233 | _EVAL_208;
  assign _EVAL_248 = _EVAL_129 | _EVAL_11;
  assign _EVAL_189 = _EVAL_54 - 6'h1;
  assign _EVAL_130 = _EVAL_6 == _EVAL_182;
  assign _EVAL_153 = _EVAL_130 | _EVAL_11;
  assign _EVAL_95 = _EVAL_2 & _EVAL_13;
  assign _EVAL_234 = _EVAL_32 == 6'h0;
  assign _EVAL_199 = _EVAL_95 & _EVAL_234;
  assign _EVAL_249 = _EVAL_3 == 3'h6;
  assign _EVAL_42 = _EVAL_249 == 1'h0;
  assign _EVAL_204 = _EVAL_199 & _EVAL_42;
  assign _EVAL_192 = _EVAL_7 == 3'h2;
  assign _EVAL_201 = _EVAL_4 <= 4'h6;
  assign _EVAL_220 = _EVAL_6 ^ 32'h1900000;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_220)};
  assign _EVAL_70 = $signed(_EVAL_113) & $signed(-33'sh2000);
  assign _EVAL_69 = $signed(_EVAL_70);
  assign _EVAL_15 = $signed(_EVAL_69) == $signed(33'sh0);
  assign _EVAL_45 = _EVAL_287 | _EVAL_15;
  assign _EVAL_206 = _EVAL_6 ^ 32'h20000000;
  assign _EVAL_33 = {1'b0,$signed(_EVAL_206)};
  assign _EVAL_40 = $signed(_EVAL_33) & $signed(-33'sh2000);
  assign _EVAL_147 = $signed(_EVAL_40);
  assign _EVAL_59 = $signed(_EVAL_147) == $signed(33'sh0);
  assign _EVAL_296 = _EVAL_45 | _EVAL_59;
  assign _EVAL_92 = _EVAL_201 & _EVAL_296;
  assign _EVAL_82 = plusarg_reader_out == 32'h0;
  assign _EVAL_18 = _EVAL_4 <= 4'h8;
  assign _EVAL_178 = _EVAL_6 ^ 32'h3000;
  assign _EVAL_36 = {1'b0,$signed(_EVAL_178)};
  assign _EVAL_120 = $signed(_EVAL_36) & $signed(-33'sh1000);
  assign _EVAL_247 = $signed(_EVAL_120);
  assign _EVAL_86 = $signed(_EVAL_247) == $signed(33'sh0);
  assign _EVAL_159 = _EVAL_18 & _EVAL_86;
  assign _EVAL_266 = _EVAL_159 | _EVAL_11;
  assign _EVAL_65 = _EVAL_258 == 6'h0;
  assign _EVAL_91 = _EVAL_92 | _EVAL_159;
  assign _EVAL_89 = _EVAL_86 | _EVAL_254;
  assign _EVAL_126 = _EVAL_89 | _EVAL_136;
  assign _EVAL_39 = _EVAL_126 | _EVAL_197;
  assign _EVAL_149 = _EVAL_39 | _EVAL_158;
  assign _EVAL_90 = _EVAL_149 | _EVAL_15;
  assign _EVAL_241 = _EVAL_90 | _EVAL_59;
  assign _EVAL_292 = _EVAL_74 & _EVAL_241;
  assign _EVAL_218 = _EVAL_292 | _EVAL_11;
  assign _EVAL_30 = _EVAL_204 ? 2'h1 : 2'h0;
  assign _EVAL_121 = _EVAL_30[0];
  assign _EVAL_67 = ~ _EVAL_121;
  assign _EVAL_211 = _EVAL_128 == 1'h0;
  assign _EVAL_77 = _EVAL_208 | _EVAL_233;
  assign _EVAL_219 = _EVAL_77 & _EVAL_67;
  assign _EVAL_168 = _EVAL_233 != _EVAL_121;
  assign _EVAL_116 = _EVAL_208 == 1'h0;
  assign _EVAL_50 = _EVAL_116 | _EVAL_82;
  assign _EVAL_53 = _EVAL_233 == 1'h0;
  assign _EVAL_188 = _EVAL_168 | _EVAL_53;
  assign _EVAL_122 = _EVAL_188 | _EVAL_11;
  assign _EVAL_57 = _EVAL_122 == 1'h0;
  assign _EVAL_135 = _EVAL_3 <= 3'h6;
  assign _EVAL_291 = _EVAL_135 | _EVAL_11;
  assign _EVAL_203 = _EVAL_201 & _EVAL_66;
  assign _EVAL_119 = _EVAL_12 == _EVAL_115;
  assign _EVAL_227 = _EVAL_3[0];
  assign _EVAL_263 = 23'hff << _EVAL;
  assign _EVAL_112 = _EVAL_263[7:0];
  assign _EVAL_160 = ~ _EVAL_112;
  assign _EVAL_257 = _EVAL_160[7:2];
  assign _EVAL_48 = _EVAL_32 - 6'h1;
  assign _EVAL_34 = _EVAL_65 == 1'h0;
  assign _EVAL_284 = _EVAL_13 & _EVAL_34;
  assign _EVAL_195 = _EVAL_165 | _EVAL_11;
  assign _EVAL_250 = _EVAL_203 | _EVAL_11;
  assign _EVAL_191 = _EVAL_255 | _EVAL_95;
  assign _EVAL_222 = _EVAL_98 + 32'h1;
  assign _EVAL_143 = _EVAL_7 == 3'h1;
  assign _EVAL_146 = _EVAL_9 == _EVAL_271;
  assign _EVAL_183 = _EVAL_146 | _EVAL_11;
  assign _EVAL_114 = _EVAL_183 == 1'h0;
  assign _EVAL_238 = _EVAL_294 | _EVAL_8;
  assign _EVAL_60 = _EVAL_238 | _EVAL_11;
  assign _EVAL_221 = _EVAL_60 == 1'h0;
  assign _EVAL_101 = _EVAL_7 == 3'h0;
  assign _EVAL_200 = _EVAL_3 == 3'h5;
  assign _EVAL_295 = _EVAL_13 & _EVAL_200;
  assign _EVAL_63 = _EVAL_29 == 6'h0;
  assign _EVAL_51 = _EVAL_7[2];
  assign _EVAL_216 = _EVAL_51 == 1'h0;
  assign _EVAL_150 = _EVAL_207[7:2];
  assign _EVAL_181 = _EVAL_29 - 6'h1;
  assign _EVAL_61 = _EVAL_1 == 2'h0;
  assign _EVAL_80 = _EVAL_61 | _EVAL_11;
  assign _EVAL_213 = ~ _EVAL_132;
  assign _EVAL_274 = _EVAL_0 & _EVAL_213;
  assign _EVAL_230 = _EVAL_91 | _EVAL_11;
  assign _EVAL_280 = _EVAL_7 == 3'h5;
  assign _EVAL_172 = _EVAL == _EVAL_276;
  assign _EVAL_85 = _EVAL_172 | _EVAL_11;
  assign _EVAL_179 = _EVAL_85 == 1'h0;
  assign _EVAL_205 = _EVAL >= 4'h2;
  assign _EVAL_24 = _EVAL_205 | _EVAL_11;
  assign _EVAL_137 = _EVAL_153 == 1'h0;
  assign _EVAL_232 = _EVAL_195 == 1'h0;
  assign _EVAL_293 = _EVAL_3 == 3'h0;
  assign _EVAL_124 = _EVAL_250 == 1'h0;
  assign _EVAL_283 = _EVAL_258 - 6'h1;
  assign _EVAL_277 = _EVAL_266 == 1'h0;
  assign _EVAL_273 = _EVAL_11 == 1'h0;
  assign _EVAL_177 = _EVAL_1 <= 2'h2;
  assign _EVAL_164 = _EVAL_177 | _EVAL_11;
  assign _EVAL_262 = ~ _EVAL_0;
  assign _EVAL_68 = _EVAL_7 == 3'h3;
  assign _EVAL_78 = _EVAL_5 & _EVAL_143;
  assign _EVAL_118 = _EVAL_265 | _EVAL_11;
  assign _EVAL_235 = _EVAL_118 == 1'h0;
  assign _EVAL_155 = _EVAL_262 == 4'h0;
  assign _EVAL_174 = _EVAL_255 & _EVAL_63;
  assign _EVAL_151 = _EVAL_155 | _EVAL_11;
  assign _EVAL_108 = _EVAL_151 == 1'h0;
  assign _EVAL_297 = _EVAL_7 == 3'h4;
  assign _EVAL_162 = _EVAL_5 & _EVAL_297;
  assign _EVAL_261 = _EVAL_248 == 1'h0;
  assign _EVAL_252 = _EVAL_230 == 1'h0;
  assign _EVAL_41 = _EVAL_63 == 1'h0;
  assign _EVAL_169 = _EVAL_5 & _EVAL_41;
  assign _EVAL_288 = _EVAL_7 == _EVAL_196;
  assign _EVAL_142 = _EVAL_288 | _EVAL_11;
  assign _EVAL_46 = _EVAL_142 == 1'h0;
  assign _EVAL_282 = _EVAL_3 == _EVAL_64;
  assign _EVAL_35 = _EVAL_282 | _EVAL_11;
  assign _EVAL_72 = _EVAL_35 == 1'h0;
  assign _EVAL_37 = _EVAL_7 == 3'h7;
  assign _EVAL_236 = _EVAL_5 & _EVAL_37;
  assign _EVAL_56 = _EVAL_98 < plusarg_reader_out;
  assign _EVAL_138 = _EVAL_50 | _EVAL_56;
  assign _EVAL_170 = _EVAL_138 | _EVAL_11;
  assign _EVAL_214 = _EVAL_3 == 3'h2;
  assign _EVAL_167 = _EVAL_13 & _EVAL_214;
  assign _EVAL_285 = _EVAL_8 == 1'h0;
  assign _EVAL_260 = _EVAL_291 == 1'h0;
  assign _EVAL_228 = _EVAL_95 & _EVAL_65;
  assign _EVAL_157 = _EVAL_5 & _EVAL_68;
  assign _EVAL_17 = _EVAL_164 == 1'h0;
  assign _EVAL_83 = _EVAL_119 | _EVAL_11;
  assign _EVAL_194 = _EVAL_274 == 4'h0;
  assign _EVAL_87 = _EVAL_194 | _EVAL_11;
  assign _EVAL_21 = _EVAL_218 == 1'h0;
  assign _EVAL_212 = _EVAL_5 & _EVAL_101;
  assign _EVAL_22 = _EVAL_1 == _EVAL_105;
  assign _EVAL_240 = _EVAL_285 | _EVAL_11;
  assign _EVAL_25 = _EVAL_240 == 1'h0;
  assign _EVAL_161 = _EVAL_5 & _EVAL_192;
  assign _EVAL_111 = _EVAL_3 == 3'h4;
  assign _EVAL_99 = _EVAL_13 & _EVAL_111;
  assign _EVAL_103 = _EVAL_22 | _EVAL_11;
  assign _EVAL_226 = _EVAL_116 | _EVAL_11;
  assign _EVAL_76 = _EVAL_226 == 1'h0;
  assign _EVAL_133 = _EVAL_7 == 3'h6;
  assign _EVAL_88 = _EVAL_5 & _EVAL_280;
  assign _EVAL_117 = _EVAL_170 == 1'h0;
  assign _EVAL_246 = _EVAL_13 & _EVAL_249;
  assign _EVAL_100 = _EVAL_24 == 1'h0;
  assign _EVAL_231 = _EVAL_4 == _EVAL_259;
  assign _EVAL_145 = _EVAL_80 == 1'h0;
  assign _EVAL_20 = _EVAL_13 & _EVAL_293;
  assign _EVAL_264 = _EVAL_231 | _EVAL_11;
  assign _EVAL_110 = _EVAL_83 == 1'h0;
  assign _EVAL_109 = _EVAL_5 & _EVAL_133;
  assign _EVAL_79 = _EVAL_3 == 3'h1;
  assign _EVAL_102 = _EVAL_13 & _EVAL_79;
  assign _EVAL_125 = _EVAL_87 == 1'h0;
  assign _EVAL_62 = _EVAL_103 == 1'h0;
  assign _EVAL_256 = _EVAL_264 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_29 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_32 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_54 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_64 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_98 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_105 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_115 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_182 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_196 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_208 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_258 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_259 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_271 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_276 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL_11) begin
      _EVAL_29 <= 6'h0;
    end else begin
      if (_EVAL_255) begin
        if (_EVAL_63) begin
          if (_EVAL_216) begin
            _EVAL_29 <= _EVAL_150;
          end else begin
            _EVAL_29 <= 6'h0;
          end
        end else begin
          _EVAL_29 <= _EVAL_181;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_32 <= 6'h0;
    end else begin
      if (_EVAL_95) begin
        if (_EVAL_234) begin
          if (_EVAL_227) begin
            _EVAL_32 <= _EVAL_257;
          end else begin
            _EVAL_32 <= 6'h0;
          end
        end else begin
          _EVAL_32 <= _EVAL_48;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_54 <= 6'h0;
    end else begin
      if (_EVAL_255) begin
        if (_EVAL_175) begin
          if (_EVAL_216) begin
            _EVAL_54 <= _EVAL_150;
          end else begin
            _EVAL_54 <= 6'h0;
          end
        end else begin
          _EVAL_54 <= _EVAL_189;
        end
      end
    end
    if (_EVAL_228) begin
      _EVAL_64 <= _EVAL_3;
    end
    if (_EVAL_11) begin
      _EVAL_98 <= 32'h0;
    end else begin
      if (_EVAL_191) begin
        _EVAL_98 <= 32'h0;
      end else begin
        _EVAL_98 <= _EVAL_222;
      end
    end
    if (_EVAL_228) begin
      _EVAL_105 <= _EVAL_1;
    end
    if (_EVAL_228) begin
      _EVAL_115 <= _EVAL_12;
    end
    if (_EVAL_174) begin
      _EVAL_182 <= _EVAL_6;
    end
    if (_EVAL_174) begin
      _EVAL_196 <= _EVAL_7;
    end
    if (_EVAL_11) begin
      _EVAL_208 <= 1'h0;
    end else begin
      _EVAL_208 <= _EVAL_219;
    end
    if (_EVAL_11) begin
      _EVAL_258 <= 6'h0;
    end else begin
      if (_EVAL_95) begin
        if (_EVAL_65) begin
          if (_EVAL_227) begin
            _EVAL_258 <= _EVAL_257;
          end else begin
            _EVAL_258 <= 6'h0;
          end
        end else begin
          _EVAL_258 <= _EVAL_283;
        end
      end
    end
    if (_EVAL_174) begin
      _EVAL_259 <= _EVAL_4;
    end
    if (_EVAL_228) begin
      _EVAL_271 <= _EVAL_9;
    end
    if (_EVAL_228) begin
      _EVAL_276 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf4d8e1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(985396ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ae02060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1f23288)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c474004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(823e028c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69b79593)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(621b5ca7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee732923)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb3abd59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27053cb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(335510a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f461f869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1bb6728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1ae1d6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b0eb700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c20d4ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2de87ad0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f54b100)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d883d4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11d1df28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2892221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(709d7c4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d121f16f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a63a9cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c28874d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f45b7c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e7e2052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9420ab2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d9b955)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eca14be9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(911085bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b8798d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed356e99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cabce42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32cc9f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3a149b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e7d8644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12d369aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ce5474)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67d489f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c2e4213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c2154ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd763aad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23c38dff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99c13d41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec3f5f2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae3ff6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4877920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c13e4523)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12b1bb67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(777d1771)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58b9b7a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ad724c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14b64b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dc815ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a39fa6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2c81bc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a863234)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebfae418)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
