//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_294(
  output        _EVAL,
  input         _EVAL_0,
  input  [32:0] _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  output [2:0]  _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output [26:0] _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input  [32:0] _EVAL_15,
  output [9:0]  _EVAL_16,
  input  [2:0]  _EVAL_17
);
  reg [22:0] _EVAL_57;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_59;
  reg [31:0] _RAND_1;
  reg  _EVAL_81;
  reg [31:0] _RAND_2;
  reg [9:0] _EVAL_83;
  reg [31:0] _RAND_3;
  reg  _EVAL_86;
  reg [31:0] _RAND_4;
  reg  _EVAL_107;
  reg [31:0] _RAND_5;
  reg  _EVAL_110;
  reg [31:0] _RAND_6;
  reg [25:0] _EVAL_117;
  reg [31:0] _RAND_7;
  reg  _EVAL_161;
  reg [31:0] _RAND_8;
  reg  _EVAL_168;
  reg [31:0] _RAND_9;
  reg  _EVAL_170;
  reg [31:0] _RAND_10;
  reg [25:0] _EVAL_199;
  reg [31:0] _RAND_11;
  reg [4:0] _EVAL_224;
  reg [31:0] _RAND_12;
  wire [26:0] _EVAL_204;
  wire  _EVAL_137;
  wire [8:0] _EVAL_133;
  wire [9:0] _EVAL_210;
  wire  _EVAL_219;
  wire  _EVAL_169;
  wire  _EVAL_152;
  wire  _EVAL_88;
  wire  _EVAL_36;
  wire  _EVAL_217;
  wire [2:0] _EVAL_30;
  wire  _EVAL_94;
  wire  _EVAL_89;
  wire [22:0] _EVAL_200;
  wire [24:0] _EVAL_102;
  wire [25:0] _EVAL_188;
  wire [25:0] _EVAL_25;
  wire [26:0] _EVAL_130;
  wire  _EVAL_84;
  wire [1:0] _EVAL_21;
  wire [1:0] _EVAL_174;
  wire [21:0] _EVAL_85;
  wire [24:0] _EVAL_190;
  wire [26:0] _EVAL_99;
  wire [26:0] _EVAL_126;
  wire [26:0] _EVAL_31;
  wire  _EVAL_27;
  wire [26:0] _EVAL_51;
  wire [26:0] _EVAL_131;
  wire [27:0] _EVAL_118;
  wire [30:0] _EVAL_29;
  wire [8:0] _EVAL_40;
  wire [2:0] _EVAL_48;
  wire  _EVAL_106;
  wire  _EVAL_119;
  wire [22:0] _EVAL_147;
  wire [24:0] _EVAL_164;
  wire [25:0] _EVAL_105;
  wire [25:0] _EVAL_53;
  wire  _EVAL_39;
  wire  _EVAL_146;
  wire  _EVAL_90;
  wire [24:0] _EVAL_187;
  wire [25:0] _EVAL_139;
  wire [25:0] _EVAL_167;
  wire [25:0] _EVAL_45;
  wire [25:0] _EVAL_124;
  wire  _EVAL_171;
  wire  _EVAL_35;
  wire [23:0] _EVAL_43;
  wire [24:0] _EVAL_132;
  wire [24:0] _EVAL_140;
  wire [25:0] _EVAL_172;
  wire [25:0] _EVAL_144;
  wire [29:0] _EVAL_34;
  wire  _EVAL_122;
  wire [26:0] _EVAL_120;
  wire [29:0] _EVAL_20;
  wire [31:0] _EVAL_37;
  wire [29:0] _EVAL_63;
  wire [29:0] _EVAL_205;
  wire [29:0] _EVAL_101;
  wire [29:0] _EVAL_121;
  wire [30:0] _EVAL_129;
  wire [30:0] _EVAL_165;
  wire [30:0] _EVAL_173;
  wire  _EVAL_71;
  wire [25:0] _EVAL_215;
  wire [25:0] _EVAL_23;
  wire  _EVAL_42;
  wire [24:0] _EVAL_26;
  wire [25:0] _EVAL_149;
  wire [25:0] _EVAL_65;
  wire [30:0] _EVAL_100;
  wire [1:0] _EVAL_163;
  wire  _EVAL_186;
  wire  _EVAL_95;
  wire  _EVAL_66;
  wire  _EVAL_177;
  wire [1:0] _EVAL_159;
  wire  _EVAL_47;
  wire  _EVAL_72;
  wire  _EVAL_151;
  wire  _EVAL_211;
  wire  _EVAL_221;
  wire [4:0] _EVAL_92;
  wire [4:0] _EVAL_202;
  wire  _EVAL_157;
  wire  _EVAL_207;
  wire  _EVAL_55;
  wire  _EVAL_113;
  wire  _EVAL_38;
  wire  _EVAL_180;
  wire  _EVAL_76;
  wire [9:0] _EVAL_135;
  wire  _EVAL_97;
  wire [7:0] _EVAL_223;
  wire [7:0] _EVAL_203;
  wire [8:0] _EVAL_87;
  wire [8:0] _EVAL_80;
  wire [9:0] _EVAL_111;
  wire [10:0] _EVAL_96;
  wire  _EVAL_50;
  wire [3:0] _EVAL_160;
  wire [3:0] _EVAL_216;
  wire  _EVAL_179;
  wire  _EVAL_145;
  wire  _EVAL_222;
  wire [5:0] _EVAL_109;
  wire  _EVAL_33;
  wire  _EVAL_69;
  wire  _EVAL_158;
  wire  _EVAL_143;
  wire  _EVAL_75;
  wire  _EVAL_108;
  wire  _EVAL_209;
  wire  _EVAL_32;
  wire  _EVAL_141;
  wire  _EVAL_176;
  wire  _EVAL_192;
  wire  _EVAL_64;
  wire  _EVAL_98;
  wire [23:0] _EVAL_184;
  wire [23:0] _EVAL_82;
  wire [25:0] _EVAL_166;
  wire [25:0] _EVAL_103;
  wire [29:0] _EVAL_58;
  wire [29:0] _EVAL_56;
  wire [29:0] _EVAL_49;
  wire [29:0] _EVAL_78;
  wire [29:0] _EVAL_214;
  wire [29:0] _EVAL_127;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_44;
  wire  _EVAL_123;
  wire  _EVAL_61;
  wire  _EVAL_189;
  wire  _EVAL_70;
  wire  _EVAL_150;
  wire [8:0] _EVAL_93;
  wire [9:0] _EVAL_91;
  wire [9:0] _EVAL_182;
  wire [9:0] _EVAL_41;
  wire  _EVAL_185;
  wire  _EVAL_104;
  wire  _EVAL_194;
  wire  _EVAL_62;
  wire  _EVAL_68;
  wire  _EVAL_52;
  wire [26:0] _EVAL_24;
  wire  _EVAL_77;
  wire  _EVAL_213;
  wire  _EVAL_28;
  wire [4:0] _EVAL_153;
  wire  _EVAL_79;
  wire  _EVAL_116;
  wire [4:0] _EVAL_183;
  wire  _EVAL_138;
  wire [4:0] _EVAL_74;
  wire [4:0] _EVAL_206;
  wire  _EVAL_125;
  wire  _EVAL_195;
  wire  _EVAL_73;
  wire  _EVAL_191;
  wire  _EVAL_22;
  wire  _EVAL_155;
  wire [4:0] _EVAL_193;
  wire [4:0] _EVAL_181;
  wire  _EVAL_196;
  wire [4:0] _EVAL_156;
  wire [4:0] _EVAL_67;
  wire  _EVAL_46;
  wire  _EVAL_212;
  wire [30:0] _EVAL_134;
  wire [30:0] _EVAL_201;
  wire  _EVAL_220;
  wire [22:0] _EVAL_178;
  wire  _EVAL_60;
  wire  _EVAL_136;
  wire  _EVAL_198;
  wire  _EVAL_162;
  wire  _EVAL_208;
  wire  _EVAL_197;
  wire  _EVAL_112;
  assign _EVAL_204 = {_EVAL_117, 1'h0};
  assign _EVAL_137 = _EVAL_224 <= 5'h1;
  assign _EVAL_133 = _EVAL_1[31:23];
  assign _EVAL_210 = {1'b0,$signed(_EVAL_133)};
  assign _EVAL_219 = _EVAL_210[0];
  assign _EVAL_169 = _EVAL_0 & _EVAL_219;
  assign _EVAL_152 = _EVAL_169 == 1'h0;
  assign _EVAL_88 = _EVAL_137 & _EVAL_152;
  assign _EVAL_36 = _EVAL_0 == 1'h0;
  assign _EVAL_217 = _EVAL_137 & _EVAL_36;
  assign _EVAL_30 = _EVAL_133[8:6];
  assign _EVAL_94 = _EVAL_30 == 3'h0;
  assign _EVAL_89 = _EVAL_94 == 1'h0;
  assign _EVAL_200 = _EVAL_1[22:0];
  assign _EVAL_102 = {1'h0,_EVAL_89,_EVAL_200};
  assign _EVAL_188 = {_EVAL_102, 1'h0};
  assign _EVAL_25 = _EVAL_88 ? _EVAL_188 : 26'h0;
  assign _EVAL_130 = {{1'd0}, _EVAL_25};
  assign _EVAL_84 = _EVAL_137 & _EVAL_169;
  assign _EVAL_21 = _EVAL_102[23:22];
  assign _EVAL_174 = _EVAL_21 - 2'h1;
  assign _EVAL_85 = _EVAL_102[21:0];
  assign _EVAL_190 = {_EVAL_85, 3'h0};
  assign _EVAL_99 = {_EVAL_174,_EVAL_190};
  assign _EVAL_126 = _EVAL_84 ? _EVAL_99 : 27'h0;
  assign _EVAL_31 = _EVAL_130 | _EVAL_126;
  assign _EVAL_27 = _EVAL_137 == 1'h0;
  assign _EVAL_51 = _EVAL_27 ? _EVAL_204 : 27'h0;
  assign _EVAL_131 = _EVAL_31 | _EVAL_51;
  assign _EVAL_118 = {1'b0,$signed(_EVAL_131)};
  assign _EVAL_29 = {{3{_EVAL_118[27]}},_EVAL_118};
  assign _EVAL_40 = _EVAL_15[31:23];
  assign _EVAL_48 = _EVAL_40[8:6];
  assign _EVAL_106 = _EVAL_48 == 3'h0;
  assign _EVAL_119 = _EVAL_106 == 1'h0;
  assign _EVAL_147 = _EVAL_15[22:0];
  assign _EVAL_164 = {1'h0,_EVAL_119,_EVAL_147};
  assign _EVAL_105 = {_EVAL_164, 1'h0};
  assign _EVAL_53 = _EVAL_217 ? _EVAL_105 : 26'h0;
  assign _EVAL_39 = _EVAL_219 == 1'h0;
  assign _EVAL_146 = _EVAL_0 & _EVAL_39;
  assign _EVAL_90 = _EVAL_137 & _EVAL_146;
  assign _EVAL_187 = _EVAL_90 ? 25'h1000000 : 25'h0;
  assign _EVAL_139 = {{1'd0}, _EVAL_187};
  assign _EVAL_167 = _EVAL_53 | _EVAL_139;
  assign _EVAL_45 = _EVAL_84 ? 26'h2800000 : 26'h0;
  assign _EVAL_124 = _EVAL_167 | _EVAL_45;
  assign _EVAL_171 = _EVAL_168 == 1'h0;
  assign _EVAL_35 = _EVAL_27 & _EVAL_171;
  assign _EVAL_43 = {1'h1,_EVAL_57};
  assign _EVAL_132 = {_EVAL_43, 1'h0};
  assign _EVAL_140 = _EVAL_35 ? _EVAL_132 : 25'h0;
  assign _EVAL_172 = {{1'd0}, _EVAL_140};
  assign _EVAL_144 = _EVAL_124 | _EVAL_172;
  assign _EVAL_34 = {{4'd0}, _EVAL_144};
  assign _EVAL_122 = _EVAL_27 & _EVAL_168;
  assign _EVAL_120 = {_EVAL_199, 1'h0};
  assign _EVAL_20 = {{3'd0}, _EVAL_120};
  assign _EVAL_37 = 32'h1 << _EVAL_224;
  assign _EVAL_63 = _EVAL_37[31:2];
  assign _EVAL_205 = _EVAL_20 | _EVAL_63;
  assign _EVAL_101 = _EVAL_122 ? _EVAL_205 : 30'h0;
  assign _EVAL_121 = _EVAL_34 | _EVAL_101;
  assign _EVAL_129 = {1'b0,$signed(_EVAL_121)};
  assign _EVAL_165 = $signed(_EVAL_29) - $signed(_EVAL_129);
  assign _EVAL_173 = $signed(_EVAL_165);
  assign _EVAL_71 = $signed(31'sh0) <= $signed(_EVAL_173);
  assign _EVAL_215 = {_EVAL_71, 25'h0};
  assign _EVAL_23 = _EVAL_217 ? _EVAL_215 : 26'h0;
  assign _EVAL_42 = _EVAL_137 & _EVAL_0;
  assign _EVAL_26 = _EVAL_42 ? 25'h1000000 : 25'h0;
  assign _EVAL_149 = {{1'd0}, _EVAL_26};
  assign _EVAL_65 = _EVAL_23 | _EVAL_149;
  assign _EVAL_100 = $unsigned(_EVAL_173);
  assign _EVAL_163 = _EVAL_133[8:7];
  assign _EVAL_186 = _EVAL_163 == 2'h3;
  assign _EVAL_95 = _EVAL_133[6];
  assign _EVAL_66 = _EVAL_95 == 1'h0;
  assign _EVAL_177 = _EVAL_186 & _EVAL_66;
  assign _EVAL_159 = _EVAL_40[8:7];
  assign _EVAL_47 = _EVAL_159 == 2'h3;
  assign _EVAL_72 = _EVAL_40[6];
  assign _EVAL_151 = _EVAL_72 == 1'h0;
  assign _EVAL_211 = _EVAL_47 & _EVAL_151;
  assign _EVAL_221 = _EVAL_177 & _EVAL_211;
  assign _EVAL_92 = _EVAL_219 ? 5'h18 : 5'h19;
  assign _EVAL_202 = _EVAL_0 ? _EVAL_92 : 5'h1a;
  assign _EVAL_157 = _EVAL_47 & _EVAL_72;
  assign _EVAL_207 = _EVAL_157 | _EVAL_211;
  assign _EVAL_55 = _EVAL_207 | _EVAL_106;
  assign _EVAL_113 = _EVAL_55 == 1'h0;
  assign _EVAL_38 = _EVAL_94 & _EVAL_106;
  assign _EVAL_180 = _EVAL_15[32];
  assign _EVAL_76 = _EVAL_177 == 1'h0;
  assign _EVAL_135 = {1'b0,$signed(_EVAL_40)};
  assign _EVAL_97 = _EVAL_135[8];
  assign _EVAL_223 = _EVAL_135[7:0];
  assign _EVAL_203 = ~ _EVAL_223;
  assign _EVAL_87 = {_EVAL_97,_EVAL_203};
  assign _EVAL_80 = $signed(_EVAL_87);
  assign _EVAL_111 = {{1{_EVAL_80[8]}},_EVAL_80};
  assign _EVAL_96 = $signed(_EVAL_210) + $signed(_EVAL_111);
  assign _EVAL_50 = $signed(11'sh1c0) <= $signed(_EVAL_96);
  assign _EVAL_160 = _EVAL_96[9:6];
  assign _EVAL_216 = _EVAL_50 ? 4'h6 : _EVAL_160;
  assign _EVAL_179 = _EVAL_102[22];
  assign _EVAL_145 = _EVAL_179 == 1'h0;
  assign _EVAL_222 = _EVAL_94 | _EVAL_211;
  assign _EVAL_109 = _EVAL_96[5:0];
  assign _EVAL_33 = _EVAL_137 & _EVAL_2;
  assign _EVAL_69 = _EVAL_186 & _EVAL_95;
  assign _EVAL_158 = _EVAL_69 | _EVAL_177;
  assign _EVAL_143 = _EVAL_158 | _EVAL_94;
  assign _EVAL_75 = _EVAL_143 == 1'h0;
  assign _EVAL_108 = _EVAL_1[32];
  assign _EVAL_209 = _EVAL_108 == 1'h0;
  assign _EVAL_32 = _EVAL_75 & _EVAL_209;
  assign _EVAL_141 = _EVAL_75 & _EVAL_113;
  assign _EVAL_176 = _EVAL_0 ? _EVAL_32 : _EVAL_141;
  assign _EVAL_192 = _EVAL_33 & _EVAL_176;
  assign _EVAL_64 = _EVAL_27 & _EVAL_71;
  assign _EVAL_98 = _EVAL_192 | _EVAL_64;
  assign _EVAL_184 = {_EVAL_71, 23'h0};
  assign _EVAL_82 = _EVAL_84 ? _EVAL_184 : 24'h0;
  assign _EVAL_166 = {{2'd0}, _EVAL_82};
  assign _EVAL_103 = _EVAL_65 | _EVAL_166;
  assign _EVAL_58 = {{4'd0}, _EVAL_103};
  assign _EVAL_56 = {{4'd0}, _EVAL_199};
  assign _EVAL_49 = _EVAL_56 | _EVAL_63;
  assign _EVAL_78 = _EVAL_27 ? _EVAL_49 : 30'h0;
  assign _EVAL_214 = _EVAL_58 | _EVAL_78;
  assign _EVAL_127 = _EVAL_98 ? _EVAL_214 : {{4'd0}, _EVAL_199};
  assign _EVAL_18 = _EVAL_176 == 1'h0;
  assign _EVAL_19 = _EVAL_36 & _EVAL_180;
  assign _EVAL_44 = _EVAL_108 ^ _EVAL_19;
  assign _EVAL_123 = _EVAL_69 & _EVAL_145;
  assign _EVAL_61 = _EVAL_164[22];
  assign _EVAL_189 = _EVAL_61 == 1'h0;
  assign _EVAL_70 = _EVAL_157 & _EVAL_189;
  assign _EVAL_150 = _EVAL_123 | _EVAL_70;
  assign _EVAL_93 = _EVAL_210[9:1];
  assign _EVAL_91 = $signed(_EVAL_93) + $signed(9'sh80);
  assign _EVAL_182 = {_EVAL_216,_EVAL_109};
  assign _EVAL_41 = $signed(_EVAL_182);
  assign _EVAL_185 = _EVAL_69 == 1'h0;
  assign _EVAL_104 = _EVAL_185 & _EVAL_76;
  assign _EVAL_194 = _EVAL_104 & _EVAL_106;
  assign _EVAL_62 = _EVAL_185 & _EVAL_89;
  assign _EVAL_68 = _EVAL_62 & _EVAL_108;
  assign _EVAL_52 = _EVAL_123 | _EVAL_68;
  assign _EVAL_24 = {{26'd0}, _EVAL_107};
  assign _EVAL_77 = _EVAL_38 | _EVAL_221;
  assign _EVAL_213 = _EVAL_150 | _EVAL_77;
  assign _EVAL_28 = _EVAL_213 | _EVAL_194;
  assign _EVAL_153 = _EVAL_224 - 5'h1;
  assign _EVAL_79 = _EVAL_69 | _EVAL_68;
  assign _EVAL_116 = _EVAL_224 == 5'h3;
  assign _EVAL_183 = _EVAL_192 ? _EVAL_202 : 5'h0;
  assign _EVAL_138 = _EVAL_33 & _EVAL_18;
  assign _EVAL_74 = {{4'd0}, _EVAL_138};
  assign _EVAL_206 = _EVAL_74 | _EVAL_183;
  assign _EVAL_125 = _EVAL_224 == 5'h0;
  assign _EVAL_195 = _EVAL_125 == 1'h0;
  assign _EVAL_73 = _EVAL_199[25];
  assign _EVAL_191 = _EVAL_116 & _EVAL_73;
  assign _EVAL_22 = _EVAL_191 == 1'h0;
  assign _EVAL_155 = _EVAL_195 & _EVAL_22;
  assign _EVAL_193 = _EVAL_155 ? _EVAL_153 : 5'h0;
  assign _EVAL_181 = _EVAL_206 | _EVAL_193;
  assign _EVAL_196 = _EVAL_195 & _EVAL_191;
  assign _EVAL_156 = {{4'd0}, _EVAL_196};
  assign _EVAL_67 = _EVAL_181 | _EVAL_156;
  assign _EVAL_46 = _EVAL_224 > 5'h2;
  assign _EVAL_212 = _EVAL_192 | _EVAL_46;
  assign _EVAL_134 = _EVAL_71 ? _EVAL_100 : {{4'd0}, _EVAL_131};
  assign _EVAL_201 = _EVAL_212 ? _EVAL_134 : {{5'd0}, _EVAL_117};
  assign _EVAL_220 = _EVAL_195 | _EVAL_2;
  assign _EVAL_178 = _EVAL_164[22:0];
  assign _EVAL_60 = _EVAL_192 & _EVAL_36;
  assign _EVAL_136 = _EVAL_86 == 1'h0;
  assign _EVAL_198 = _EVAL_177 | _EVAL_106;
  assign _EVAL_162 = _EVAL_69 | _EVAL_157;
  assign _EVAL_208 = _EVAL_162 | _EVAL_77;
  assign _EVAL_197 = _EVAL_224 == 5'h1;
  assign _EVAL_112 = $signed(_EVAL_173) != $signed(31'sh0);
  assign _EVAL_13 = _EVAL_81 & _EVAL_86;
  assign _EVAL_8 = _EVAL_197 & _EVAL_168;
  assign _EVAL_16 = _EVAL_83;
  assign _EVAL_10 = _EVAL_86;
  assign _EVAL_9 = _EVAL_120 | _EVAL_24;
  assign _EVAL_4 = _EVAL_59;
  assign _EVAL_14 = _EVAL_161;
  assign _EVAL_6 = _EVAL_110;
  assign _EVAL_3 = _EVAL_197 & _EVAL_171;
  assign _EVAL_11 = _EVAL_224 <= 5'h1;
  assign _EVAL = _EVAL_170;
  assign _EVAL_7 = _EVAL_81 & _EVAL_136;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_57 = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_59 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_81 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_83 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_86 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_107 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_110 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_117 = _RAND_7[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_161 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_168 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_170 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_199 = _RAND_11[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_224 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_12) begin
    if (_EVAL_60) begin
      _EVAL_57 <= _EVAL_178;
    end
    if (_EVAL_192) begin
      _EVAL_59 <= _EVAL_17;
    end
    if (_EVAL_33) begin
      if (_EVAL_0) begin
        _EVAL_81 <= _EVAL_52;
      end else begin
        _EVAL_81 <= _EVAL_28;
      end
    end
    if (_EVAL_192) begin
      if (_EVAL_0) begin
        _EVAL_83 <= _EVAL_91;
      end else begin
        _EVAL_83 <= _EVAL_41;
      end
    end
    if (_EVAL_33) begin
      if (_EVAL_0) begin
        _EVAL_86 <= _EVAL_79;
      end else begin
        _EVAL_86 <= _EVAL_208;
      end
    end
    if (_EVAL_98) begin
      _EVAL_107 <= _EVAL_112;
    end
    if (_EVAL_33) begin
      if (_EVAL_0) begin
        _EVAL_110 <= _EVAL_94;
      end else begin
        _EVAL_110 <= _EVAL_222;
      end
    end
    _EVAL_117 <= _EVAL_201[25:0];
    if (_EVAL_33) begin
      _EVAL_161 <= _EVAL_44;
    end
    if (_EVAL_33) begin
      _EVAL_168 <= _EVAL_0;
    end
    if (_EVAL_33) begin
      if (_EVAL_0) begin
        _EVAL_170 <= _EVAL_177;
      end else begin
        _EVAL_170 <= _EVAL_198;
      end
    end
    _EVAL_199 <= _EVAL_127[25:0];
    if (_EVAL_5) begin
      _EVAL_224 <= 5'h0;
    end else begin
      if (_EVAL_220) begin
        _EVAL_224 <= _EVAL_67;
      end
    end
  end
endmodule
