//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_217(
  output [1:0]  _EVAL,
  output        _EVAL_0,
  output [8:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output [1:0]  _EVAL_4,
  output        _EVAL_5,
  output [31:0] _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [2:0]  _EVAL_16,
  input  [8:0]  _EVAL_17,
  output        _EVAL_18,
  output [2:0]  _EVAL_19,
  output [3:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output        _EVAL_22,
  output [31:0] _EVAL_23,
  input  [1:0]  _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input  [31:0] _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  input  [3:0]  _EVAL_33
);
  wire  AsyncQueueSink__EVAL;
  wire  AsyncQueueSink__EVAL_0;
  wire  AsyncQueueSink__EVAL_1;
  wire [31:0] AsyncQueueSink__EVAL_2;
  wire  AsyncQueueSink__EVAL_3;
  wire  AsyncQueueSink__EVAL_4;
  wire [2:0] AsyncQueueSink__EVAL_5;
  wire [3:0] AsyncQueueSink__EVAL_6;
  wire [31:0] AsyncQueueSink__EVAL_7;
  wire [1:0] AsyncQueueSink__EVAL_8;
  wire [2:0] AsyncQueueSink__EVAL_9;
  wire  AsyncQueueSink__EVAL_10;
  wire  AsyncQueueSink__EVAL_11;
  wire  AsyncQueueSink__EVAL_12;
  wire [3:0] AsyncQueueSink__EVAL_13;
  wire [8:0] AsyncQueueSink__EVAL_14;
  wire [2:0] AsyncQueueSink__EVAL_15;
  wire  AsyncQueueSink__EVAL_16;
  wire [8:0] AsyncQueueSink__EVAL_17;
  wire  AsyncQueueSink__EVAL_18;
  wire  AsyncQueueSource__EVAL;
  wire  AsyncQueueSource__EVAL_0;
  wire [2:0] AsyncQueueSource__EVAL_1;
  wire [31:0] AsyncQueueSource__EVAL_2;
  wire [1:0] AsyncQueueSource__EVAL_3;
  wire [2:0] AsyncQueueSource__EVAL_4;
  wire  AsyncQueueSource__EVAL_5;
  wire  AsyncQueueSource__EVAL_6;
  wire  AsyncQueueSource__EVAL_7;
  wire  AsyncQueueSource__EVAL_8;
  wire [31:0] AsyncQueueSource__EVAL_9;
  wire  AsyncQueueSource__EVAL_10;
  wire  AsyncQueueSource__EVAL_11;
  wire [1:0] AsyncQueueSource__EVAL_12;
  wire  AsyncQueueSource__EVAL_13;
  wire  AsyncQueueSource__EVAL_14;
  SiFive__EVAL_215 AsyncQueueSink (
    ._EVAL(AsyncQueueSink__EVAL),
    ._EVAL_0(AsyncQueueSink__EVAL_0),
    ._EVAL_1(AsyncQueueSink__EVAL_1),
    ._EVAL_2(AsyncQueueSink__EVAL_2),
    ._EVAL_3(AsyncQueueSink__EVAL_3),
    ._EVAL_4(AsyncQueueSink__EVAL_4),
    ._EVAL_5(AsyncQueueSink__EVAL_5),
    ._EVAL_6(AsyncQueueSink__EVAL_6),
    ._EVAL_7(AsyncQueueSink__EVAL_7),
    ._EVAL_8(AsyncQueueSink__EVAL_8),
    ._EVAL_9(AsyncQueueSink__EVAL_9),
    ._EVAL_10(AsyncQueueSink__EVAL_10),
    ._EVAL_11(AsyncQueueSink__EVAL_11),
    ._EVAL_12(AsyncQueueSink__EVAL_12),
    ._EVAL_13(AsyncQueueSink__EVAL_13),
    ._EVAL_14(AsyncQueueSink__EVAL_14),
    ._EVAL_15(AsyncQueueSink__EVAL_15),
    ._EVAL_16(AsyncQueueSink__EVAL_16),
    ._EVAL_17(AsyncQueueSink__EVAL_17),
    ._EVAL_18(AsyncQueueSink__EVAL_18)
  );
  SiFive__EVAL_216 AsyncQueueSource (
    ._EVAL(AsyncQueueSource__EVAL),
    ._EVAL_0(AsyncQueueSource__EVAL_0),
    ._EVAL_1(AsyncQueueSource__EVAL_1),
    ._EVAL_2(AsyncQueueSource__EVAL_2),
    ._EVAL_3(AsyncQueueSource__EVAL_3),
    ._EVAL_4(AsyncQueueSource__EVAL_4),
    ._EVAL_5(AsyncQueueSource__EVAL_5),
    ._EVAL_6(AsyncQueueSource__EVAL_6),
    ._EVAL_7(AsyncQueueSource__EVAL_7),
    ._EVAL_8(AsyncQueueSource__EVAL_8),
    ._EVAL_9(AsyncQueueSource__EVAL_9),
    ._EVAL_10(AsyncQueueSource__EVAL_10),
    ._EVAL_11(AsyncQueueSource__EVAL_11),
    ._EVAL_12(AsyncQueueSource__EVAL_12),
    ._EVAL_13(AsyncQueueSource__EVAL_13),
    ._EVAL_14(AsyncQueueSource__EVAL_14)
  );
  assign AsyncQueueSink__EVAL_3 = _EVAL_2;
  assign AsyncQueueSource__EVAL_1 = _EVAL_15;
  assign AsyncQueueSource__EVAL_13 = _EVAL_9;
  assign AsyncQueueSink__EVAL_7 = _EVAL_29;
  assign _EVAL_5 = AsyncQueueSink__EVAL_11;
  assign _EVAL_4 = AsyncQueueSink__EVAL_8;
  assign _EVAL_25 = AsyncQueueSource__EVAL_10;
  assign AsyncQueueSink__EVAL = _EVAL_7;
  assign _EVAL = AsyncQueueSource__EVAL_12;
  assign _EVAL_1 = AsyncQueueSink__EVAL_14;
  assign _EVAL_0 = AsyncQueueSource__EVAL_0;
  assign _EVAL_22 = AsyncQueueSink__EVAL_12;
  assign _EVAL_32 = AsyncQueueSource__EVAL_11;
  assign _EVAL_19 = AsyncQueueSink__EVAL_15;
  assign AsyncQueueSink__EVAL_18 = _EVAL_12;
  assign _EVAL_20 = AsyncQueueSink__EVAL_13;
  assign AsyncQueueSink__EVAL_10 = _EVAL_3;
  assign _EVAL_23 = AsyncQueueSink__EVAL_2;
  assign _EVAL_16 = AsyncQueueSource__EVAL_4;
  assign AsyncQueueSource__EVAL_8 = _EVAL_13;
  assign _EVAL_31 = AsyncQueueSource__EVAL_7;
  assign AsyncQueueSource__EVAL_14 = _EVAL_26;
  assign _EVAL_18 = AsyncQueueSink__EVAL_16;
  assign _EVAL_6 = AsyncQueueSource__EVAL_9;
  assign AsyncQueueSource__EVAL = _EVAL_27;
  assign AsyncQueueSink__EVAL_4 = _EVAL_8;
  assign _EVAL_30 = AsyncQueueSink__EVAL_0;
  assign AsyncQueueSource__EVAL_3 = _EVAL_24;
  assign _EVAL_11 = AsyncQueueSink__EVAL_5;
  assign AsyncQueueSource__EVAL_5 = _EVAL_28;
  assign AsyncQueueSink__EVAL_9 = _EVAL_21;
  assign AsyncQueueSource__EVAL_2 = _EVAL_14;
  assign AsyncQueueSink__EVAL_6 = _EVAL_33;
  assign AsyncQueueSink__EVAL_17 = _EVAL_17;
  assign AsyncQueueSource__EVAL_6 = _EVAL_7;
  assign _EVAL_10 = AsyncQueueSink__EVAL_1;
endmodule
