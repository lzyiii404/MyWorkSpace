//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_187_assert(
  input  [2:0]  _EVAL,
  input  [11:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [25:0] _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [1:0]  _EVAL_17,
  input         _EVAL_18,
  input  [3:0]  _EVAL_19,
  input         _EVAL_33,
  input         _EVAL_196,
  input         _EVAL_195,
  input         _EVAL_92,
  input  [31:0] _EVAL_62,
  input  [7:0]  _EVAL_139,
  input         _EVAL_67,
  input  [7:0]  _EVAL_179,
  input         _EVAL_123,
  input  [7:0]  _EVAL_110,
  input         _EVAL_96,
  input  [7:0]  _EVAL_71,
  input         _EVAL_198,
  input         _EVAL_88,
  input         _EVAL_176,
  input         _EVAL_40,
  input         _EVAL_109,
  input         _EVAL_112,
  input         _EVAL_163,
  input         _EVAL_75,
  input         _EVAL_146,
  input         _EVAL_85,
  input         _EVAL_140,
  input         _EVAL_201,
  input         _EVAL_189,
  input         _EVAL_22,
  input  [13:0] _EVAL_24,
  input         _EVAL_29,
  input         _EVAL_194,
  input         _EVAL_121,
  input         _EVAL_104,
  input         _EVAL_135,
  input         _EVAL_157,
  input         _EVAL_74
);
  wire  TLMonitor__EVAL;
  wire [1:0] TLMonitor__EVAL_0;
  wire [3:0] TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire [11:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire [11:0] TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire [25:0] TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire [1:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire  _EVAL_181;
  wire  _EVAL_105;
  wire  _EVAL_39;
  wire  _EVAL_26;
  wire [30:0] _EVAL_36;
  wire  _EVAL_136;
  wire  _EVAL_44;
  wire  _EVAL_32;
  wire  _EVAL_175;
  wire  _EVAL_124;
  wire  _EVAL_58;
  wire  _EVAL_95;
  wire  _EVAL_97;
  wire  _EVAL_119;
  wire  _EVAL_186;
  wire  _EVAL_99;
  wire  _EVAL_80;
  wire  _EVAL_90;
  wire  _EVAL_154;
  wire  _EVAL_190;
  wire  _EVAL_102;
  wire  _EVAL_101;
  wire  _EVAL_191;
  wire  _EVAL_34;
  wire  _EVAL_199;
  wire  _EVAL_68;
  wire  _EVAL_63;
  wire  _EVAL_30;
  wire  _EVAL_23;
  wire  _EVAL_86;
  wire  _EVAL_77;
  wire  _EVAL_60;
  wire  _EVAL_125;
  wire  _EVAL_51;
  wire  _EVAL_70;
  wire  _EVAL_131;
  wire  _EVAL_115;
  wire  _EVAL_116;
  SiFive__EVAL_186_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  assign _EVAL_181 = _EVAL_33 & _EVAL_196;
  assign _EVAL_105 = _EVAL_181 & _EVAL_75;
  assign _EVAL_39 = _EVAL_181 & _EVAL_109;
  assign _EVAL_26 = _EVAL_181 & _EVAL_85;
  assign _EVAL_36 = _EVAL_62[31:1];
  assign _EVAL_136 = _EVAL_36 != 31'h0;
  assign _EVAL_44 = _EVAL_181 & _EVAL_195;
  assign _EVAL_32 = _EVAL_44 & _EVAL_92;
  assign _EVAL_175 = _EVAL_179 != 8'h0;
  assign _EVAL_124 = _EVAL_32 & _EVAL_175;
  assign _EVAL_58 = _EVAL_139 != 8'h0;
  assign _EVAL_95 = _EVAL_32 & _EVAL_58;
  assign _EVAL_97 = _EVAL_26 & _EVAL_112;
  assign _EVAL_119 = _EVAL_97 & _EVAL_58;
  assign _EVAL_186 = _EVAL_71 != 8'h0;
  assign _EVAL_99 = _EVAL_39 & _EVAL_112;
  assign _EVAL_80 = _EVAL_99 & _EVAL_186;
  assign _EVAL_90 = _EVAL_99 & _EVAL_58;
  assign _EVAL_154 = _EVAL_181 & _EVAL_88;
  assign _EVAL_190 = _EVAL_154 & _EVAL_92;
  assign _EVAL_102 = _EVAL_110 != 8'h0;
  assign _EVAL_101 = _EVAL_190 & _EVAL_102;
  assign _EVAL_191 = _EVAL_36 == 31'h7fffffff;
  assign _EVAL_34 = _EVAL_11 == 1'h0;
  assign _EVAL_199 = _EVAL_99 & _EVAL_175;
  assign _EVAL_68 = _EVAL_190 & _EVAL_186;
  assign _EVAL_63 = _EVAL_97 & _EVAL_102;
  assign _EVAL_30 = _EVAL_97 & _EVAL_175;
  assign _EVAL_23 = _EVAL_105 & _EVAL_92;
  assign _EVAL_86 = _EVAL_190 & _EVAL_58;
  assign _EVAL_77 = _EVAL_23 & _EVAL_135;
  assign _EVAL_60 = _EVAL_32 & _EVAL_186;
  assign _EVAL_125 = _EVAL_99 & _EVAL_102;
  assign _EVAL_51 = _EVAL_190 & _EVAL_175;
  assign _EVAL_70 = _EVAL_104 & _EVAL_191;
  assign _EVAL_131 = _EVAL_97 & _EVAL_186;
  assign _EVAL_115 = _EVAL_32 & _EVAL_102;
  assign _EVAL_116 = _EVAL_23 & _EVAL_136;
  assign TLMonitor__EVAL_11 = _EVAL;
  assign TLMonitor__EVAL_3 = _EVAL_16;
  assign TLMonitor__EVAL_13 = _EVAL_18;
  assign TLMonitor__EVAL_10 = _EVAL_15;
  assign TLMonitor__EVAL_2 = {{2'd0}, _EVAL_196};
  assign TLMonitor__EVAL_4 = _EVAL_24[13:2];
  assign TLMonitor__EVAL_6 = _EVAL_10;
  assign TLMonitor__EVAL_14 = _EVAL_3;
  assign TLMonitor__EVAL_8 = _EVAL_1;
  assign TLMonitor__EVAL_9 = _EVAL_2;
  assign TLMonitor__EVAL_12 = _EVAL_24[1:0];
  assign TLMonitor__EVAL_5 = _EVAL_11;
  assign TLMonitor__EVAL = _EVAL_3;
  assign TLMonitor__EVAL_7 = _EVAL_18;
  assign TLMonitor__EVAL_0 = _EVAL_17;
  assign TLMonitor__EVAL_1 = _EVAL_19;
  always @(posedge _EVAL_10) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a84d8f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fd17d52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d430dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e4e0946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed2cf2a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc70a10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cff64fa8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(457efe16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d4d3b4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35196506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fad4806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ae811ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99ffb4f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a9cfff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e366a758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aa7970e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef837cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55b9374)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc2e5035)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f628da97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9981b13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6655e6e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6bd2417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75035d07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55171fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3782bc8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1532b462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23d03a54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51583e47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6e8261)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9078fbcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a18bc4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d05e5692)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd73fd34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51513657)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d56cbf7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8edd1fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1665bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2165987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff3fe197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27a81a67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4010fd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a38033bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fd6e30f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fde38fac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf02c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6d3ac8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34619dd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d8c77f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9da3cd9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(612a7ca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472cd3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673b7792)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc445861)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e89c13ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e615b476)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96200104)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fe196f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7988edd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfd26e44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721c945d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a61fa49a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69cdd24a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64063857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4912e66b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c8caea4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f971138)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2464bf92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
