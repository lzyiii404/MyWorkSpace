//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_249(
  output        _EVAL,
  input         _EVAL_0,
  output [1:0]  _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  output [7:0]  _EVAL_4,
  output [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  output        _EVAL_8,
  input  [3:0]  _EVAL_9,
  output [31:0] _EVAL_10,
  output [24:0] _EVAL_11,
  output [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output [3:0]  _EVAL_17,
  input  [7:0]  _EVAL_18,
  input  [31:0] _EVAL_19,
  input         _EVAL_20,
  output [2:0]  _EVAL_21,
  input  [1:0]  _EVAL_22,
  output [31:0] _EVAL_23,
  output        _EVAL_24,
  input  [24:0] _EVAL_25,
  input  [2:0]  _EVAL_26,
  input         _EVAL_27,
  input  [12:0] _EVAL_28,
  output [2:0]  _EVAL_29,
  output [12:0] _EVAL_30,
  input  [2:0]  _EVAL_31,
  output        _EVAL_32
);
  wire  Repeater__EVAL;
  wire [2:0] Repeater__EVAL_0;
  wire [7:0] Repeater__EVAL_1;
  wire  Repeater__EVAL_2;
  wire [2:0] Repeater__EVAL_3;
  wire [2:0] Repeater__EVAL_4;
  wire  Repeater__EVAL_5;
  wire [24:0] Repeater__EVAL_6;
  wire [2:0] Repeater__EVAL_7;
  wire  Repeater__EVAL_8;
  wire  Repeater__EVAL_9;
  wire [3:0] Repeater__EVAL_10;
  wire  Repeater__EVAL_11;
  wire  Repeater__EVAL_12;
  wire [7:0] Repeater__EVAL_13;
  wire [3:0] Repeater__EVAL_14;
  wire [2:0] Repeater__EVAL_15;
  wire  Repeater__EVAL_16;
  wire  Repeater__EVAL_17;
  wire [24:0] Repeater__EVAL_18;
  wire [2:0] Repeater__EVAL_19;
  wire  Repeater__EVAL_20;
  reg [2:0] _EVAL_39;
  reg [31:0] _RAND_0;
  reg  _EVAL_67;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_73;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_94;
  reg [31:0] _RAND_3;
  reg  _EVAL_108;
  reg [31:0] _RAND_4;
  wire [12:0] _EVAL_99;
  wire [5:0] _EVAL_71;
  wire [5:0] _EVAL_54;
  wire [5:0] _EVAL_66;
  wire [3:0] _EVAL_84;
  wire [5:0] _EVAL_85;
  wire [4:0] _EVAL_92;
  wire [1:0] _EVAL_97;
  wire [1:0] _EVAL_79;
  wire [5:0] _EVAL_41;
  wire [5:0] _EVAL_57;
  wire [6:0] _EVAL_55;
  wire [6:0] _EVAL_72;
  wire  _EVAL_110;
  wire [3:0] _EVAL_51;
  wire [3:0] _EVAL_61;
  wire [3:0] _EVAL_69;
  wire [3:0] _EVAL_45;
  wire [3:0] _EVAL_107;
  wire  _EVAL_120;
  wire  _EVAL_74;
  wire  _EVAL_35;
  wire [8:0] _EVAL_122;
  wire [5:0] _EVAL_95;
  wire [5:0] _EVAL_44;
  wire [3:0] _EVAL_70;
  wire [2:0] _EVAL_87;
  wire  _EVAL_64;
  wire  _EVAL_77;
  wire [2:0] _EVAL_98;
  wire [8:0] _EVAL_65;
  wire [1:0] _EVAL_113;
  wire [1:0] _EVAL_93;
  wire [5:0] _EVAL_109;
  wire [5:0] _EVAL_53;
  wire [5:0] _EVAL_91;
  wire  _EVAL_49;
  wire  _EVAL_114;
  wire [3:0] _EVAL_48;
  wire  _EVAL_88;
  wire [6:0] _EVAL_76;
  wire [6:0] _EVAL_58;
  wire [6:0] _EVAL_52;
  wire [3:0] _EVAL_68;
  wire  _EVAL_111;
  wire  _EVAL_38;
  wire  _EVAL_90;
  wire  _EVAL_100;
  wire  _EVAL_115;
  wire  _EVAL_89;
  wire  _EVAL_81;
  wire [5:0] _EVAL_121;
  wire [24:0] _EVAL_75;
  wire  _EVAL_117;
  wire  _EVAL_82;
  wire  _EVAL_40;
  wire  _EVAL_33;
  wire [2:0] _EVAL_118;
  wire  _EVAL_103;
  wire  _EVAL_86;
  wire [3:0] _EVAL_112;
  wire [3:0] _EVAL_101;
  wire [3:0] _EVAL_123;
  wire [1:0] _EVAL_47;
  wire  _EVAL_62;
  wire [1:0] _EVAL_42;
  wire [1:0] _EVAL_96;
  wire  _EVAL_37;
  wire [2:0] _EVAL_56;
  wire  _EVAL_106;
  SiFive__EVAL_248 Repeater (
    ._EVAL(Repeater__EVAL),
    ._EVAL_0(Repeater__EVAL_0),
    ._EVAL_1(Repeater__EVAL_1),
    ._EVAL_2(Repeater__EVAL_2),
    ._EVAL_3(Repeater__EVAL_3),
    ._EVAL_4(Repeater__EVAL_4),
    ._EVAL_5(Repeater__EVAL_5),
    ._EVAL_6(Repeater__EVAL_6),
    ._EVAL_7(Repeater__EVAL_7),
    ._EVAL_8(Repeater__EVAL_8),
    ._EVAL_9(Repeater__EVAL_9),
    ._EVAL_10(Repeater__EVAL_10),
    ._EVAL_11(Repeater__EVAL_11),
    ._EVAL_12(Repeater__EVAL_12),
    ._EVAL_13(Repeater__EVAL_13),
    ._EVAL_14(Repeater__EVAL_14),
    ._EVAL_15(Repeater__EVAL_15),
    ._EVAL_16(Repeater__EVAL_16),
    ._EVAL_17(Repeater__EVAL_17),
    ._EVAL_18(Repeater__EVAL_18),
    ._EVAL_19(Repeater__EVAL_19),
    ._EVAL_20(Repeater__EVAL_20)
  );
  assign _EVAL_99 = 13'h3f << Repeater__EVAL_15;
  assign _EVAL_71 = _EVAL_99[5:0];
  assign _EVAL_54 = ~ _EVAL_71;
  assign _EVAL_66 = ~ _EVAL_54;
  assign _EVAL_84 = _EVAL_28[3:0];
  assign _EVAL_85 = {_EVAL_84, 2'h0};
  assign _EVAL_92 = 5'h3 << _EVAL_22;
  assign _EVAL_97 = _EVAL_92[1:0];
  assign _EVAL_79 = ~ _EVAL_97;
  assign _EVAL_41 = {{4'd0}, _EVAL_79};
  assign _EVAL_57 = _EVAL_85 | _EVAL_41;
  assign _EVAL_55 = {1'h0,_EVAL_57};
  assign _EVAL_72 = ~ _EVAL_55;
  assign _EVAL_110 = _EVAL_94 == 4'h0;
  assign _EVAL_51 = _EVAL_54[5:2];
  assign _EVAL_61 = _EVAL_94 - 4'h1;
  assign _EVAL_69 = _EVAL_110 ? _EVAL_51 : _EVAL_61;
  assign _EVAL_45 = ~ _EVAL_69;
  assign _EVAL_107 = ~ _EVAL_45;
  assign _EVAL_120 = _EVAL_107 != 4'h0;
  assign _EVAL_74 = _EVAL_110 ? _EVAL_108 : _EVAL_67;
  assign _EVAL_35 = _EVAL_74 == 1'h0;
  assign _EVAL_122 = {Repeater__EVAL_1,_EVAL_35};
  assign _EVAL_95 = {_EVAL_69, 2'h0};
  assign _EVAL_44 = _EVAL_95 | _EVAL_66;
  assign _EVAL_70 = 4'h1 << _EVAL_22;
  assign _EVAL_87 = _EVAL_70[2:0];
  assign _EVAL_64 = _EVAL_87[2:2];
  assign _EVAL_77 = Repeater__EVAL_15 > 3'h2;
  assign _EVAL_98 = _EVAL_77 ? 3'h2 : Repeater__EVAL_15;
  assign _EVAL_65 = 9'h3 << _EVAL_98;
  assign _EVAL_113 = _EVAL_65[1:0];
  assign _EVAL_93 = ~ _EVAL_113;
  assign _EVAL_109 = {{4'd0}, _EVAL_93};
  assign _EVAL_53 = _EVAL_44 | _EVAL_109;
  assign _EVAL_91 = _EVAL_53 | 6'h3;
  assign _EVAL_49 = _EVAL_13[0];
  assign _EVAL_114 = _EVAL_49 ? 1'h1 : _EVAL_64;
  assign _EVAL_48 = {{3'd0}, _EVAL_114};
  assign _EVAL_88 = _EVAL_49 == 1'h0;
  assign _EVAL_76 = {_EVAL_57, 1'h0};
  assign _EVAL_58 = _EVAL_76 | 7'h1;
  assign _EVAL_52 = _EVAL_58 & _EVAL_72;
  assign _EVAL_68 = _EVAL_52[3:0];
  assign _EVAL_111 = _EVAL_84 == 4'h0;
  assign _EVAL_38 = _EVAL_111 == 1'h0;
  assign _EVAL_90 = _EVAL_88 & _EVAL_38;
  assign _EVAL_100 = _EVAL_7 | _EVAL_90;
  assign _EVAL_115 = _EVAL_100 & _EVAL_20;
  assign _EVAL_89 = _EVAL_73 == 4'h0;
  assign _EVAL_81 = _EVAL_28[4];
  assign _EVAL_121 = ~ _EVAL_91;
  assign _EVAL_75 = {{19'd0}, _EVAL_121};
  assign _EVAL_117 = Repeater__EVAL_12;
  assign _EVAL_82 = Repeater__EVAL_0[2];
  assign _EVAL_40 = _EVAL_82 == 1'h0;
  assign _EVAL_33 = _EVAL_40 == 1'h0;
  assign _EVAL_118 = _EVAL_52[6:4];
  assign _EVAL_103 = _EVAL_118 != 3'h0;
  assign _EVAL_86 = _EVAL_16 & _EVAL_117;
  assign _EVAL_112 = {{1'd0}, _EVAL_118};
  assign _EVAL_101 = _EVAL_73 - _EVAL_48;
  assign _EVAL_123 = _EVAL_112 | _EVAL_68;
  assign _EVAL_47 = _EVAL_123[3:2];
  assign _EVAL_62 = _EVAL_47 != 2'h0;
  assign _EVAL_42 = _EVAL_123[1:0];
  assign _EVAL_96 = _EVAL_47 | _EVAL_42;
  assign _EVAL_37 = _EVAL_96[1];
  assign _EVAL_56 = {_EVAL_103,_EVAL_62,_EVAL_37};
  assign _EVAL_106 = _EVAL_90 == 1'h0;
  assign _EVAL_3 = _EVAL_20 & _EVAL_106;
  assign _EVAL_8 = _EVAL_7 | _EVAL_90;
  assign _EVAL_24 = Repeater__EVAL_5;
  assign _EVAL_12 = _EVAL_13;
  assign _EVAL_30 = {_EVAL_122,_EVAL_107};
  assign Repeater__EVAL_7 = _EVAL_6;
  assign _EVAL_21 = Repeater__EVAL_0;
  assign _EVAL_17 = Repeater__EVAL_17 ? 4'hf : _EVAL_9;
  assign Repeater__EVAL_11 = _EVAL_27;
  assign Repeater__EVAL_18 = _EVAL_25;
  assign _EVAL_1 = _EVAL_98[1:0];
  assign Repeater__EVAL_10 = _EVAL_9;
  assign _EVAL_5 = _EVAL_89 ? _EVAL_56 : _EVAL_39;
  assign Repeater__EVAL_13 = _EVAL_18;
  assign _EVAL_32 = Repeater__EVAL_2;
  assign _EVAL_29 = Repeater__EVAL_3;
  assign Repeater__EVAL = _EVAL_33 & _EVAL_120;
  assign Repeater__EVAL_20 = _EVAL_0;
  assign _EVAL_4 = _EVAL_28[12:5];
  assign Repeater__EVAL_16 = _EVAL_16;
  assign _EVAL_11 = Repeater__EVAL_6 | _EVAL_75;
  assign Repeater__EVAL_19 = _EVAL_26;
  assign Repeater__EVAL_9 = _EVAL_15;
  assign _EVAL_23 = _EVAL_14;
  assign _EVAL = Repeater__EVAL_12;
  assign _EVAL_10 = _EVAL_19;
  assign Repeater__EVAL_8 = _EVAL_2;
  assign Repeater__EVAL_4 = _EVAL_31;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_39 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_67 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_73 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_94 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_108 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_115) begin
      if (_EVAL_89) begin
        _EVAL_39 <= _EVAL_56;
      end
    end
    if (_EVAL_110) begin
      _EVAL_67 <= _EVAL_108;
    end
    if (_EVAL_15) begin
      _EVAL_73 <= 4'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_89) begin
          _EVAL_73 <= _EVAL_84;
        end else begin
          _EVAL_73 <= _EVAL_101;
        end
      end
    end
    if (_EVAL_15) begin
      _EVAL_94 <= 4'h0;
    end else begin
      if (_EVAL_86) begin
        _EVAL_94 <= _EVAL_107;
      end
    end
    if (_EVAL_15) begin
      _EVAL_108 <= 1'h0;
    end else begin
      if (_EVAL_115) begin
        if (_EVAL_89) begin
          _EVAL_108 <= _EVAL_81;
        end
      end
    end
  end
endmodule
