//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_30_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [6:0]  _EVAL_5,
  input         _EVAL_6,
  input  [6:0]  _EVAL_7,
  input  [30:0] _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [30:0] _EVAL_40;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_57;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_71;
  reg [31:0] _RAND_2;
  reg [6:0] _EVAL_78;
  reg [31:0] _RAND_3;
  reg [72:0] _EVAL_121;
  reg [95:0] _RAND_4;
  reg [2:0] _EVAL_140;
  reg [31:0] _RAND_5;
  reg  _EVAL_149;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_162;
  reg [31:0] _RAND_7;
  reg [31:0] _EVAL_169;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_175;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_190;
  reg [31:0] _RAND_10;
  reg [6:0] _EVAL_205;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_246;
  reg [31:0] _RAND_12;
  reg [3:0] _EVAL_252;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_292;
  reg [31:0] _RAND_14;
  wire  _EVAL_49;
  wire  _EVAL_148;
  wire  _EVAL_99;
  wire  _EVAL_296;
  wire  _EVAL_186;
  wire [3:0] _EVAL_68;
  wire  _EVAL_180;
  wire  _EVAL_112;
  wire  _EVAL_29;
  wire  _EVAL_136;
  wire  _EVAL_196;
  wire  _EVAL_215;
  wire  _EVAL_242;
  wire [127:0] _EVAL_18;
  wire [127:0] _EVAL_264;
  wire [72:0] _EVAL_43;
  wire  _EVAL_138;
  wire  _EVAL_234;
  wire  _EVAL_225;
  wire  _EVAL_187;
  wire  _EVAL_235;
  wire  _EVAL_36;
  wire  _EVAL_31;
  wire  _EVAL_275;
  wire  _EVAL_173;
  wire  _EVAL_84;
  wire [30:0] _EVAL_178;
  wire [31:0] _EVAL_207;
  wire [31:0] _EVAL_154;
  wire [31:0] _EVAL_201;
  wire  _EVAL_167;
  wire  _EVAL_109;
  wire  _EVAL_271;
  wire  _EVAL_293;
  wire  _EVAL_213;
  wire  _EVAL_193;
  wire [127:0] _EVAL_113;
  wire [127:0] _EVAL_142;
  wire [72:0] _EVAL_218;
  wire [3:0] _EVAL_303;
  wire  _EVAL_42;
  wire [72:0] _EVAL_279;
  wire  _EVAL_50;
  wire  _EVAL_69;
  wire [12:0] _EVAL_299;
  wire [5:0] _EVAL_41;
  wire [5:0] _EVAL_283;
  wire [30:0] _EVAL_300;
  wire  _EVAL_203;
  wire  _EVAL_222;
  wire  _EVAL_183;
  wire  _EVAL_230;
  wire  _EVAL_62;
  wire [1:0] _EVAL_120;
  wire [1:0] _EVAL_288;
  wire  _EVAL_184;
  wire  _EVAL_260;
  wire  _EVAL_72;
  wire  _EVAL_262;
  wire  _EVAL_133;
  wire  _EVAL_211;
  wire  _EVAL_268;
  wire  _EVAL_179;
  wire  _EVAL_23;
  wire  _EVAL_202;
  wire  _EVAL_259;
  wire  _EVAL_61;
  wire  _EVAL_47;
  wire  _EVAL_143;
  wire  _EVAL_44;
  wire  _EVAL_22;
  wire  _EVAL_130;
  wire  _EVAL_298;
  wire  _EVAL_155;
  wire  _EVAL_126;
  wire  _EVAL_282;
  wire [12:0] _EVAL_245;
  wire [5:0] _EVAL_297;
  wire [5:0] _EVAL_110;
  wire [3:0] _EVAL_129;
  wire  _EVAL_86;
  wire  _EVAL_94;
  wire  _EVAL_237;
  wire  _EVAL_77;
  wire  _EVAL_28;
  wire  _EVAL_81;
  wire  _EVAL_115;
  wire  _EVAL_21;
  wire  _EVAL_170;
  wire  _EVAL_147;
  wire  _EVAL_65;
  wire  _EVAL_165;
  wire  _EVAL_103;
  wire  _EVAL_152;
  wire [3:0] _EVAL_181;
  wire  _EVAL_192;
  wire  _EVAL_274;
  wire  _EVAL_161;
  wire  _EVAL_269;
  wire [2:0] _EVAL_265;
  wire  _EVAL_153;
  wire  _EVAL_64;
  wire  _EVAL_217;
  wire  _EVAL_88;
  wire  _EVAL_19;
  wire  _EVAL_104;
  wire  _EVAL_206;
  wire  _EVAL_189;
  wire  _EVAL_277;
  wire  _EVAL_34;
  wire [2:0] _EVAL_248;
  wire  _EVAL_106;
  wire  _EVAL_141;
  wire  _EVAL_281;
  wire  _EVAL_127;
  wire  _EVAL_53;
  wire [72:0] _EVAL_158;
  wire  _EVAL_157;
  wire  _EVAL_54;
  wire  _EVAL_107;
  wire  _EVAL_122;
  wire  _EVAL_76;
  wire  _EVAL_164;
  wire  _EVAL_80;
  wire  _EVAL_233;
  wire  _EVAL_240;
  wire  _EVAL_239;
  wire  _EVAL_156;
  wire [3:0] _EVAL_289;
  wire  _EVAL_291;
  wire  _EVAL_92;
  wire  _EVAL_219;
  wire [72:0] _EVAL_116;
  wire  _EVAL_75;
  wire  _EVAL_301;
  wire  _EVAL_123;
  wire  _EVAL_247;
  wire  _EVAL_254;
  wire  _EVAL_256;
  wire  _EVAL_290;
  wire  _EVAL_220;
  wire  _EVAL_236;
  wire  _EVAL_37;
  wire  _EVAL_46;
  wire  _EVAL_134;
  wire  _EVAL_124;
  wire [3:0] _EVAL_177;
  wire [3:0] _EVAL_232;
  wire [3:0] _EVAL_250;
  wire  _EVAL_89;
  wire  _EVAL_199;
  wire [3:0] _EVAL_228;
  wire  _EVAL_273;
  wire  _EVAL_114;
  wire  _EVAL_67;
  wire  _EVAL_60;
  wire  _EVAL_204;
  wire  _EVAL_258;
  wire  _EVAL_280;
  wire  _EVAL_135;
  wire  _EVAL_51;
  wire [30:0] _EVAL_223;
  wire  _EVAL_166;
  wire  _EVAL_185;
  wire  _EVAL_55;
  wire  _EVAL_209;
  wire  _EVAL_276;
  wire  _EVAL_214;
  wire  _EVAL_241;
  wire  _EVAL_272;
  wire  _EVAL_198;
  wire  _EVAL_63;
  wire  _EVAL_118;
  wire  _EVAL_168;
  wire  _EVAL_176;
  wire  _EVAL_238;
  wire  _EVAL_249;
  wire  _EVAL_79;
  wire [3:0] _EVAL_91;
  wire  _EVAL_263;
  wire [3:0] _EVAL_287;
  wire  _EVAL_111;
  wire  _EVAL_74;
  wire  _EVAL_231;
  wire  _EVAL_56;
  wire  _EVAL_119;
  wire  _EVAL_27;
  wire  _EVAL_159;
  wire  _EVAL_255;
  wire  _EVAL_128;
  wire  _EVAL_210;
  wire  _EVAL_208;
  wire  _EVAL_195;
  wire  _EVAL_24;
  wire  _EVAL_171;
  wire  _EVAL_216;
  wire  _EVAL_224;
  wire  _EVAL_96;
  wire  _EVAL_52;
  wire  _EVAL_286;
  wire  _EVAL_160;
  wire [31:0] _EVAL_58;
  wire  _EVAL_105;
  wire  _EVAL_95;
  wire  _EVAL_244;
  wire  _EVAL_25;
  wire  _EVAL_101;
  wire  _EVAL_243;
  wire  _EVAL_59;
  wire  _EVAL_137;
  wire [3:0] _EVAL_197;
  wire  _EVAL_188;
  wire  _EVAL_82;
  wire  _EVAL_270;
  wire  _EVAL_108;
  wire  _EVAL_20;
  wire [72:0] _EVAL_66;
  wire [72:0] _EVAL_100;
  wire  _EVAL_26;
  wire  _EVAL_221;
  wire  _EVAL_172;
  wire  _EVAL_257;
  wire  _EVAL_35;
  wire  _EVAL_295;
  wire  _EVAL_33;
  wire  _EVAL_32;
  wire  _EVAL_139;
  wire  _EVAL_212;
  wire  _EVAL_229;
  wire  _EVAL_251;
  wire  _EVAL_151;
  wire  _EVAL_132;
  wire  _EVAL_87;
  wire  _EVAL_278;
  wire  _EVAL_174;
  wire  _EVAL_117;
  wire  _EVAL_83;
  wire  _EVAL_30;
  wire  _EVAL_266;
  wire  _EVAL_182;
  wire  _EVAL_97;
  wire [72:0] _EVAL_93;
  wire  _EVAL_145;
  wire  _EVAL_48;
  wire  _EVAL_131;
  wire  _EVAL_85;
  wire  _EVAL_226;
  wire  _EVAL_253;
  wire  _EVAL_98;
  wire  _EVAL_90;
  wire  _EVAL_17;
  wire  _EVAL_102;
  wire  _EVAL_125;
  wire  _EVAL_227;
  wire  _EVAL_194;
  wire  _EVAL_70;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_49 = _EVAL_6 & _EVAL_1;
  assign _EVAL_148 = _EVAL_175 == 4'h0;
  assign _EVAL_99 = _EVAL_49 & _EVAL_148;
  assign _EVAL_296 = _EVAL_12 == 3'h5;
  assign _EVAL_186 = _EVAL_1 & _EVAL_296;
  assign _EVAL_68 = _EVAL_71 - 4'h1;
  assign _EVAL_180 = _EVAL_12 <= 3'h6;
  assign _EVAL_112 = _EVAL_180 | _EVAL_13;
  assign _EVAL_29 = _EVAL_292 == 4'h0;
  assign _EVAL_136 = _EVAL_49 & _EVAL_29;
  assign _EVAL_196 = _EVAL_12 == 3'h6;
  assign _EVAL_215 = _EVAL_196 == 1'h0;
  assign _EVAL_242 = _EVAL_136 & _EVAL_215;
  assign _EVAL_18 = 128'h1 << _EVAL_7;
  assign _EVAL_264 = _EVAL_242 ? _EVAL_18 : 128'h0;
  assign _EVAL_43 = _EVAL_264[72:0];
  assign _EVAL_138 = _EVAL == 1'h0;
  assign _EVAL_234 = _EVAL_138 | _EVAL_13;
  assign _EVAL_225 = _EVAL_234 == 1'h0;
  assign _EVAL_187 = _EVAL_9 == _EVAL_140;
  assign _EVAL_235 = _EVAL_187 | _EVAL_13;
  assign _EVAL_36 = _EVAL_8[1];
  assign _EVAL_31 = _EVAL_8[0];
  assign _EVAL_275 = _EVAL_31 == 1'h0;
  assign _EVAL_173 = _EVAL_36 & _EVAL_275;
  assign _EVAL_84 = _EVAL_9 <= 3'h6;
  assign _EVAL_178 = _EVAL_8 ^ 31'h40000000;
  assign _EVAL_207 = {1'b0,$signed(_EVAL_178)};
  assign _EVAL_154 = $signed(_EVAL_207) & $signed(-32'sh2000);
  assign _EVAL_201 = $signed(_EVAL_154);
  assign _EVAL_167 = $signed(_EVAL_201) == $signed(32'sh0);
  assign _EVAL_109 = _EVAL_84 & _EVAL_167;
  assign _EVAL_271 = _EVAL_109 | _EVAL_13;
  assign _EVAL_293 = _EVAL_15 & _EVAL_0;
  assign _EVAL_213 = _EVAL_71 == 4'h0;
  assign _EVAL_193 = _EVAL_293 & _EVAL_213;
  assign _EVAL_113 = 128'h1 << _EVAL_5;
  assign _EVAL_142 = _EVAL_193 ? _EVAL_113 : 128'h0;
  assign _EVAL_218 = _EVAL_142[72:0];
  assign _EVAL_303 = _EVAL_5[6:3];
  assign _EVAL_42 = _EVAL_303 == 4'h8;
  assign _EVAL_279 = _EVAL_121 >> _EVAL_5;
  assign _EVAL_50 = _EVAL_279[0];
  assign _EVAL_69 = _EVAL_50 == 1'h0;
  assign _EVAL_299 = 13'h3f << _EVAL_9;
  assign _EVAL_41 = _EVAL_299[5:0];
  assign _EVAL_283 = ~ _EVAL_41;
  assign _EVAL_300 = {{25'd0}, _EVAL_283};
  assign _EVAL_203 = _EVAL_252 == 4'h0;
  assign _EVAL_222 = _EVAL_293 & _EVAL_203;
  assign _EVAL_183 = _EVAL_10 == 3'h7;
  assign _EVAL_230 = _EVAL_9 >= 3'h2;
  assign _EVAL_62 = _EVAL_9[0];
  assign _EVAL_120 = 2'h1 << _EVAL_62;
  assign _EVAL_288 = _EVAL_120 | 2'h1;
  assign _EVAL_184 = _EVAL_288[1];
  assign _EVAL_260 = _EVAL_184 & _EVAL_36;
  assign _EVAL_72 = _EVAL_230 | _EVAL_260;
  assign _EVAL_262 = _EVAL_288[0];
  assign _EVAL_133 = _EVAL_36 & _EVAL_31;
  assign _EVAL_211 = _EVAL_262 & _EVAL_133;
  assign _EVAL_268 = _EVAL_72 | _EVAL_211;
  assign _EVAL_179 = _EVAL_218 != _EVAL_43;
  assign _EVAL_23 = _EVAL_218 != 73'h0;
  assign _EVAL_202 = _EVAL_23 == 1'h0;
  assign _EVAL_259 = _EVAL_179 | _EVAL_202;
  assign _EVAL_61 = _EVAL_259 | _EVAL_13;
  assign _EVAL_47 = _EVAL_10 == _EVAL_162;
  assign _EVAL_143 = _EVAL_47 | _EVAL_13;
  assign _EVAL_44 = _EVAL_7 == _EVAL_78;
  assign _EVAL_22 = _EVAL_12 == 3'h4;
  assign _EVAL_130 = _EVAL_1 & _EVAL_22;
  assign _EVAL_298 = _EVAL_10 == 3'h4;
  assign _EVAL_155 = _EVAL_0 & _EVAL_298;
  assign _EVAL_126 = _EVAL_2 >= 3'h2;
  assign _EVAL_282 = _EVAL_126 | _EVAL_13;
  assign _EVAL_245 = 13'h3f << _EVAL_2;
  assign _EVAL_297 = _EVAL_245[5:0];
  assign _EVAL_110 = ~ _EVAL_297;
  assign _EVAL_129 = _EVAL_110[5:2];
  assign _EVAL_86 = _EVAL_121 != 73'h0;
  assign _EVAL_94 = _EVAL_86 == 1'h0;
  assign _EVAL_237 = plusarg_reader_out == 32'h0;
  assign _EVAL_77 = _EVAL_94 | _EVAL_237;
  assign _EVAL_28 = _EVAL_169 < plusarg_reader_out;
  assign _EVAL_81 = _EVAL_77 | _EVAL_28;
  assign _EVAL_115 = _EVAL_81 | _EVAL_13;
  assign _EVAL_21 = _EVAL_12 == _EVAL_57;
  assign _EVAL_170 = _EVAL_21 | _EVAL_13;
  assign _EVAL_147 = _EVAL_10 == 3'h1;
  assign _EVAL_65 = _EVAL_0 & _EVAL_147;
  assign _EVAL_165 = _EVAL_10[2];
  assign _EVAL_103 = _EVAL_165 == 1'h0;
  assign _EVAL_152 = _EVAL_303 == 4'h0;
  assign _EVAL_181 = _EVAL_7[6:3];
  assign _EVAL_192 = _EVAL_181 == 4'h1;
  assign _EVAL_274 = _EVAL_5 == 7'h48;
  assign _EVAL_161 = _EVAL_5 == 7'h40;
  assign _EVAL_269 = _EVAL_274 | _EVAL_161;
  assign _EVAL_265 = _EVAL_5[2:0];
  assign _EVAL_153 = 3'h1 <= _EVAL_265;
  assign _EVAL_64 = _EVAL_42 & _EVAL_153;
  assign _EVAL_217 = _EVAL_269 | _EVAL_64;
  assign _EVAL_88 = _EVAL_5 == 7'h20;
  assign _EVAL_19 = _EVAL_217 | _EVAL_88;
  assign _EVAL_104 = _EVAL_19 | _EVAL_152;
  assign _EVAL_206 = _EVAL_7 == 7'h48;
  assign _EVAL_189 = _EVAL_7 == 7'h40;
  assign _EVAL_277 = _EVAL_206 | _EVAL_189;
  assign _EVAL_34 = _EVAL_181 == 4'h8;
  assign _EVAL_248 = _EVAL_7[2:0];
  assign _EVAL_106 = 3'h1 <= _EVAL_248;
  assign _EVAL_141 = _EVAL_34 & _EVAL_106;
  assign _EVAL_281 = _EVAL_277 | _EVAL_141;
  assign _EVAL_127 = _EVAL_7 == 7'h20;
  assign _EVAL_53 = _EVAL_281 | _EVAL_127;
  assign _EVAL_158 = ~ _EVAL_43;
  assign _EVAL_157 = _EVAL_3 == 3'h0;
  assign _EVAL_54 = _EVAL_181 == 4'h0;
  assign _EVAL_107 = _EVAL_53 | _EVAL_54;
  assign _EVAL_122 = _EVAL_107 | _EVAL_192;
  assign _EVAL_76 = _EVAL_181 == 4'h2;
  assign _EVAL_164 = _EVAL_122 | _EVAL_76;
  assign _EVAL_80 = _EVAL_181 == 4'h3;
  assign _EVAL_233 = _EVAL_164 | _EVAL_80;
  assign _EVAL_240 = _EVAL_233 | _EVAL_13;
  assign _EVAL_239 = _EVAL_240 == 1'h0;
  assign _EVAL_156 = _EVAL_12[0];
  assign _EVAL_289 = _EVAL_175 - 4'h1;
  assign _EVAL_291 = _EVAL_12 == 3'h2;
  assign _EVAL_92 = _EVAL_1 & _EVAL_291;
  assign _EVAL_219 = _EVAL_138 | _EVAL_16;
  assign _EVAL_116 = _EVAL_121 | _EVAL_218;
  assign _EVAL_75 = _EVAL_219 | _EVAL_13;
  assign _EVAL_301 = _EVAL_75 == 1'h0;
  assign _EVAL_123 = _EVAL_262 & _EVAL_173;
  assign _EVAL_247 = _EVAL_72 | _EVAL_123;
  assign _EVAL_254 = _EVAL_36 == 1'h0;
  assign _EVAL_256 = _EVAL_184 & _EVAL_254;
  assign _EVAL_290 = _EVAL_230 | _EVAL_256;
  assign _EVAL_220 = _EVAL_254 & _EVAL_31;
  assign _EVAL_236 = _EVAL_262 & _EVAL_220;
  assign _EVAL_37 = _EVAL_290 | _EVAL_236;
  assign _EVAL_46 = _EVAL_254 & _EVAL_275;
  assign _EVAL_134 = _EVAL_262 & _EVAL_46;
  assign _EVAL_124 = _EVAL_290 | _EVAL_134;
  assign _EVAL_177 = {_EVAL_268,_EVAL_247,_EVAL_37,_EVAL_124};
  assign _EVAL_232 = ~ _EVAL_177;
  assign _EVAL_250 = _EVAL_11 & _EVAL_232;
  assign _EVAL_89 = _EVAL_250 == 4'h0;
  assign _EVAL_199 = _EVAL_89 | _EVAL_13;
  assign _EVAL_228 = _EVAL_292 - 4'h1;
  assign _EVAL_273 = _EVAL_16 == 1'h0;
  assign _EVAL_114 = _EVAL_273 | _EVAL_13;
  assign _EVAL_67 = _EVAL_61 == 1'h0;
  assign _EVAL_60 = _EVAL_11 == _EVAL_177;
  assign _EVAL_204 = _EVAL_60 | _EVAL_13;
  assign _EVAL_258 = _EVAL_204 == 1'h0;
  assign _EVAL_280 = _EVAL_44 | _EVAL_13;
  assign _EVAL_135 = _EVAL_148 == 1'h0;
  assign _EVAL_51 = _EVAL_1 & _EVAL_135;
  assign _EVAL_223 = _EVAL_8 & _EVAL_300;
  assign _EVAL_166 = _EVAL_223 == 31'h0;
  assign _EVAL_185 = _EVAL_166 | _EVAL_13;
  assign _EVAL_55 = _EVAL_185 == 1'h0;
  assign _EVAL_209 = _EVAL_170 == 1'h0;
  assign _EVAL_276 = _EVAL_12 == 3'h1;
  assign _EVAL_214 = _EVAL_1 & _EVAL_276;
  assign _EVAL_241 = _EVAL_303 == 4'h1;
  assign _EVAL_272 = _EVAL_104 | _EVAL_241;
  assign _EVAL_198 = _EVAL_303 == 4'h2;
  assign _EVAL_63 = _EVAL_272 | _EVAL_198;
  assign _EVAL_118 = _EVAL_303 == 4'h3;
  assign _EVAL_168 = _EVAL_63 | _EVAL_118;
  assign _EVAL_176 = _EVAL_168 | _EVAL_13;
  assign _EVAL_238 = _EVAL_3 != 3'h0;
  assign _EVAL_249 = _EVAL_238 | _EVAL_13;
  assign _EVAL_79 = _EVAL_249 == 1'h0;
  assign _EVAL_91 = _EVAL_283[5:2];
  assign _EVAL_263 = _EVAL_10 == 3'h2;
  assign _EVAL_287 = ~ _EVAL_11;
  assign _EVAL_111 = _EVAL_287 == 4'h0;
  assign _EVAL_74 = 3'h6 == _EVAL_9;
  assign _EVAL_231 = _EVAL_161 ? _EVAL_74 : 1'h0;
  assign _EVAL_56 = _EVAL_231 | _EVAL_13;
  assign _EVAL_119 = _EVAL_56 == 1'h0;
  assign _EVAL_27 = _EVAL_203 == 1'h0;
  assign _EVAL_159 = _EVAL_115 == 1'h0;
  assign _EVAL_255 = _EVAL_293 | _EVAL_49;
  assign _EVAL_128 = _EVAL_10 == 3'h5;
  assign _EVAL_210 = _EVAL_0 & _EVAL_128;
  assign _EVAL_208 = _EVAL_111 | _EVAL_13;
  assign _EVAL_195 = _EVAL_208 == 1'h0;
  assign _EVAL_24 = _EVAL_280 == 1'h0;
  assign _EVAL_171 = _EVAL_282 == 1'h0;
  assign _EVAL_216 = _EVAL_3 == _EVAL_190;
  assign _EVAL_224 = _EVAL_216 | _EVAL_13;
  assign _EVAL_96 = _EVAL_2 == _EVAL_246;
  assign _EVAL_52 = _EVAL_96 | _EVAL_13;
  assign _EVAL_286 = _EVAL_52 == 1'h0;
  assign _EVAL_160 = _EVAL_157 | _EVAL_13;
  assign _EVAL_58 = _EVAL_169 + 32'h1;
  assign _EVAL_105 = _EVAL_3 <= 3'h2;
  assign _EVAL_95 = _EVAL_105 | _EVAL_13;
  assign _EVAL_244 = _EVAL_230 | _EVAL_13;
  assign _EVAL_25 = _EVAL_143 == 1'h0;
  assign _EVAL_101 = _EVAL_8 == _EVAL_40;
  assign _EVAL_243 = _EVAL_101 | _EVAL_13;
  assign _EVAL_59 = _EVAL_176 == 1'h0;
  assign _EVAL_137 = _EVAL == _EVAL_149;
  assign _EVAL_197 = _EVAL_252 - 4'h1;
  assign _EVAL_188 = _EVAL_14 == 1'h0;
  assign _EVAL_82 = _EVAL_188 | _EVAL_13;
  assign _EVAL_270 = _EVAL_82 == 1'h0;
  assign _EVAL_108 = _EVAL_160 == 1'h0;
  assign _EVAL_20 = _EVAL_5 == _EVAL_205;
  assign _EVAL_66 = _EVAL_218 | _EVAL_121;
  assign _EVAL_100 = _EVAL_66 >> _EVAL_7;
  assign _EVAL_26 = _EVAL_100[0];
  assign _EVAL_221 = _EVAL_26 | _EVAL_13;
  assign _EVAL_172 = _EVAL_221 == 1'h0;
  assign _EVAL_257 = _EVAL_10 == 3'h3;
  assign _EVAL_35 = _EVAL_0 & _EVAL_257;
  assign _EVAL_295 = _EVAL_271 == 1'h0;
  assign _EVAL_33 = _EVAL_12 == 3'h0;
  assign _EVAL_32 = _EVAL_1 & _EVAL_196;
  assign _EVAL_139 = _EVAL_95 == 1'h0;
  assign _EVAL_212 = _EVAL_69 | _EVAL_13;
  assign _EVAL_229 = _EVAL_212 == 1'h0;
  assign _EVAL_251 = _EVAL_3 <= 3'h3;
  assign _EVAL_151 = _EVAL_251 | _EVAL_13;
  assign _EVAL_132 = _EVAL_151 == 1'h0;
  assign _EVAL_87 = _EVAL_137 | _EVAL_13;
  assign _EVAL_278 = _EVAL_87 == 1'h0;
  assign _EVAL_174 = _EVAL_244 == 1'h0;
  assign _EVAL_117 = _EVAL_0 & _EVAL_183;
  assign _EVAL_83 = _EVAL_13 == 1'h0;
  assign _EVAL_30 = _EVAL_10 == 3'h0;
  assign _EVAL_266 = _EVAL_1 & _EVAL_33;
  assign _EVAL_182 = _EVAL_10 == 3'h6;
  assign _EVAL_97 = _EVAL_0 & _EVAL_182;
  assign _EVAL_93 = _EVAL_116 & _EVAL_158;
  assign _EVAL_145 = _EVAL_235 == 1'h0;
  assign _EVAL_48 = _EVAL_243 == 1'h0;
  assign _EVAL_131 = _EVAL_20 | _EVAL_13;
  assign _EVAL_85 = _EVAL_131 == 1'h0;
  assign _EVAL_226 = _EVAL_224 == 1'h0;
  assign _EVAL_253 = _EVAL_112 == 1'h0;
  assign _EVAL_98 = _EVAL_0 & _EVAL_27;
  assign _EVAL_90 = _EVAL_114 == 1'h0;
  assign _EVAL_17 = _EVAL_3 <= 3'h4;
  assign _EVAL_102 = _EVAL_17 | _EVAL_13;
  assign _EVAL_125 = _EVAL_0 & _EVAL_30;
  assign _EVAL_227 = _EVAL_0 & _EVAL_263;
  assign _EVAL_194 = _EVAL_199 == 1'h0;
  assign _EVAL_70 = _EVAL_102 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_40 = _RAND_0[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_57 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_71 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_78 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  _EVAL_121 = _RAND_4[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_140 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_149 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_162 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_169 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_175 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_190 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_205 = _RAND_11[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_246 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_252 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_292 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_222) begin
      _EVAL_40 <= _EVAL_8;
    end
    if (_EVAL_99) begin
      _EVAL_57 <= _EVAL_12;
    end
    if (_EVAL_13) begin
      _EVAL_71 <= 4'h0;
    end else begin
      if (_EVAL_293) begin
        if (_EVAL_213) begin
          if (_EVAL_103) begin
            _EVAL_71 <= _EVAL_91;
          end else begin
            _EVAL_71 <= 4'h0;
          end
        end else begin
          _EVAL_71 <= _EVAL_68;
        end
      end
    end
    if (_EVAL_99) begin
      _EVAL_78 <= _EVAL_7;
    end
    if (_EVAL_13) begin
      _EVAL_121 <= 73'h0;
    end else begin
      _EVAL_121 <= _EVAL_93;
    end
    if (_EVAL_222) begin
      _EVAL_140 <= _EVAL_9;
    end
    if (_EVAL_99) begin
      _EVAL_149 <= _EVAL;
    end
    if (_EVAL_222) begin
      _EVAL_162 <= _EVAL_10;
    end
    if (_EVAL_13) begin
      _EVAL_169 <= 32'h0;
    end else begin
      if (_EVAL_255) begin
        _EVAL_169 <= 32'h0;
      end else begin
        _EVAL_169 <= _EVAL_58;
      end
    end
    if (_EVAL_13) begin
      _EVAL_175 <= 4'h0;
    end else begin
      if (_EVAL_49) begin
        if (_EVAL_148) begin
          if (_EVAL_156) begin
            _EVAL_175 <= _EVAL_129;
          end else begin
            _EVAL_175 <= 4'h0;
          end
        end else begin
          _EVAL_175 <= _EVAL_289;
        end
      end
    end
    if (_EVAL_222) begin
      _EVAL_190 <= _EVAL_3;
    end
    if (_EVAL_222) begin
      _EVAL_205 <= _EVAL_5;
    end
    if (_EVAL_99) begin
      _EVAL_246 <= _EVAL_2;
    end
    if (_EVAL_13) begin
      _EVAL_252 <= 4'h0;
    end else begin
      if (_EVAL_293) begin
        if (_EVAL_203) begin
          if (_EVAL_103) begin
            _EVAL_252 <= _EVAL_91;
          end else begin
            _EVAL_252 <= 4'h0;
          end
        end else begin
          _EVAL_252 <= _EVAL_197;
        end
      end
    end
    if (_EVAL_13) begin
      _EVAL_292 <= 4'h0;
    end else begin
      if (_EVAL_49) begin
        if (_EVAL_29) begin
          if (_EVAL_156) begin
            _EVAL_292 <= _EVAL_129;
          end else begin
            _EVAL_292 <= 4'h0;
          end
        end else begin
          _EVAL_292 <= _EVAL_228;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a4f9179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd8beefc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f01144e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6934e7b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(852043e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16db40b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab104118)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(298429ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(305ff33b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b619d3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18aed00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e56d81f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33d13a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd9f8982)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f96225c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d66e03f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f3cccf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c52d786)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(764fe0df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38e775a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de0937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9401d31d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3db41353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(128cd404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7cbd3ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a74407f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(788dcbf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ada157b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f41dbbc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf7b4aea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4abb63a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80ed0412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ebd3e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c59fc98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f8e54cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79f15155)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d9e0d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cc751f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5973c421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75c6894a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6b4229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b62ac05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a9963f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c29ce2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65c12d87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc6f7efd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f69fe626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(382bd8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928433de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec7dc1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2e71f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d2f79c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a23dce3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(461d4869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6845e0d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a6d3b0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6486ad9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdb425f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3ee7b0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b607afc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4b13773)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b759a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7197070)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c7cbef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fadacc9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(984e3368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2caa6da2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0f1ad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(319f2bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c6d7dbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(712e6f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e9bb47c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc9b2a8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df5ce594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb7bdddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28f7b2d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1df0753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de4efa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a1110a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c64ea4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
