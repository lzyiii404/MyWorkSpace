//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_240(
  input         _EVAL,
  output [3:0]  _EVAL_0,
  input         _EVAL_1,
  input  [63:0] _EVAL_2,
  output [31:0] _EVAL_3,
  output [63:0] _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  output        _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [1:0]  _EVAL_13,
  output        _EVAL_14,
  output [2:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19
);
  assign _EVAL_0 = _EVAL_6;
  assign _EVAL_14 = _EVAL_17;
  assign _EVAL_15 = _EVAL_7;
  assign _EVAL_18 = _EVAL;
  assign _EVAL_3 = _EVAL_12;
  assign _EVAL_8 = _EVAL_5;
  assign _EVAL_4 = _EVAL_2;
  assign _EVAL_11 = _EVAL_9;
endmodule
