//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_291(
  output [32:0] _EVAL,
  input  [9:0]  _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  output [4:0]  _EVAL_4,
  input         _EVAL_5,
  input  [26:0] _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9
);
  wire [9:0] roundAnyRawFNToRecFN__EVAL;
  wire  roundAnyRawFNToRecFN__EVAL_0;
  wire [4:0] roundAnyRawFNToRecFN__EVAL_1;
  wire [32:0] roundAnyRawFNToRecFN__EVAL_2;
  wire  roundAnyRawFNToRecFN__EVAL_3;
  wire  roundAnyRawFNToRecFN__EVAL_4;
  wire  roundAnyRawFNToRecFN__EVAL_5;
  wire [26:0] roundAnyRawFNToRecFN__EVAL_6;
  wire [2:0] roundAnyRawFNToRecFN__EVAL_7;
  wire  roundAnyRawFNToRecFN__EVAL_8;
  wire  roundAnyRawFNToRecFN__EVAL_9;
  SiFive__EVAL_290 roundAnyRawFNToRecFN (
    ._EVAL(roundAnyRawFNToRecFN__EVAL),
    ._EVAL_0(roundAnyRawFNToRecFN__EVAL_0),
    ._EVAL_1(roundAnyRawFNToRecFN__EVAL_1),
    ._EVAL_2(roundAnyRawFNToRecFN__EVAL_2),
    ._EVAL_3(roundAnyRawFNToRecFN__EVAL_3),
    ._EVAL_4(roundAnyRawFNToRecFN__EVAL_4),
    ._EVAL_5(roundAnyRawFNToRecFN__EVAL_5),
    ._EVAL_6(roundAnyRawFNToRecFN__EVAL_6),
    ._EVAL_7(roundAnyRawFNToRecFN__EVAL_7),
    ._EVAL_8(roundAnyRawFNToRecFN__EVAL_8),
    ._EVAL_9(roundAnyRawFNToRecFN__EVAL_9)
  );
  assign _EVAL_4 = roundAnyRawFNToRecFN__EVAL_1;
  assign roundAnyRawFNToRecFN__EVAL = _EVAL_0;
  assign roundAnyRawFNToRecFN__EVAL_0 = _EVAL_1;
  assign roundAnyRawFNToRecFN__EVAL_3 = _EVAL_5;
  assign roundAnyRawFNToRecFN__EVAL_6 = _EVAL_6;
  assign roundAnyRawFNToRecFN__EVAL_9 = _EVAL_9;
  assign roundAnyRawFNToRecFN__EVAL_7 = _EVAL_2;
  assign roundAnyRawFNToRecFN__EVAL_4 = _EVAL_7;
  assign _EVAL = roundAnyRawFNToRecFN__EVAL_2;
  assign roundAnyRawFNToRecFN__EVAL_5 = _EVAL_8;
  assign roundAnyRawFNToRecFN__EVAL_8 = _EVAL_3;
endmodule
