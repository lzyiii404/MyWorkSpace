//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_152(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  output [6:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  output [6:0]  _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [31:0] _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [6:0]  _EVAL_13,
  output        _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [1:0]  _EVAL_18,
  output [1:0]  _EVAL_19,
  output        _EVAL_20,
  output [2:0]  _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [6:0]  _EVAL_24,
  output [3:0]  _EVAL_25,
  output [1:0]  _EVAL_26,
  output [2:0]  _EVAL_27,
  output        _EVAL_28,
  output [2:0]  _EVAL_29,
  output        _EVAL_30,
  input  [3:0]  _EVAL_31,
  output [1:0]  _EVAL_32,
  input  [2:0]  _EVAL_33,
  output        _EVAL_34,
  input  [24:0] _EVAL_35,
  output [6:0]  _EVAL_36,
  input         _EVAL_37,
  output [24:0] _EVAL_38,
  input         _EVAL_39,
  input  [6:0]  _EVAL_40,
  input         _EVAL_41,
  output [31:0] _EVAL_42,
  input         _EVAL_43,
  output [24:0] _EVAL_44,
  input  [31:0] _EVAL_45,
  input  [1:0]  _EVAL_46,
  input  [2:0]  _EVAL_47,
  output [2:0]  _EVAL_48,
  output        _EVAL_49,
  input  [1:0]  _EVAL_50,
  output [2:0]  _EVAL_51,
  output [2:0]  _EVAL_52,
  input         _EVAL_53,
  output [3:0]  _EVAL_54,
  output        _EVAL_55,
  input         _EVAL_56,
  input  [31:0] _EVAL_57,
  output [31:0] _EVAL_58,
  output [31:0] _EVAL_59,
  input         _EVAL_60
);
  wire  rsource__EVAL;
  wire  rsource__EVAL_0;
  wire [2:0] rsource__EVAL_1;
  wire  rsource__EVAL_2;
  wire [2:0] rsource__EVAL_3;
  wire [31:0] rsource__EVAL_4;
  wire  rsource__EVAL_5;
  wire [1:0] rsource__EVAL_6;
  wire  rsource__EVAL_7;
  wire [3:0] rsource__EVAL_8;
  wire  rsource__EVAL_9;
  wire [1:0] rsource__EVAL_10;
  wire [6:0] rsource__EVAL_11;
  wire [2:0] rsource__EVAL_12;
  wire  rsource__EVAL_13;
  wire  rsource__EVAL_14;
  wire  rsource__EVAL_15;
  wire [2:0] rsource__EVAL_16;
  wire  rsource__EVAL_17;
  wire [31:0] rsource__EVAL_18;
  wire [1:0] rsource__EVAL_19;
  wire [24:0] rsource__EVAL_20;
  wire [2:0] rsource__EVAL_21;
  wire  rsource__EVAL_22;
  wire [2:0] rsource__EVAL_23;
  wire  rsource__EVAL_24;
  wire [31:0] rsource__EVAL_25;
  wire [31:0] rsource__EVAL_26;
  wire  rsource__EVAL_27;
  wire [3:0] rsource__EVAL_28;
  wire [1:0] rsource__EVAL_29;
  wire  rsource__EVAL_30;
  wire [2:0] rsource__EVAL_31;
  wire [2:0] rsource__EVAL_32;
  wire  rsource__EVAL_33;
  wire [2:0] rsource__EVAL_34;
  wire [1:0] rsource__EVAL_35;
  wire [2:0] rsource__EVAL_36;
  wire [6:0] rsource__EVAL_37;
  wire [6:0] rsource__EVAL_38;
  wire [2:0] rsource__EVAL_39;
  wire [2:0] rsource__EVAL_40;
  wire [2:0] rsource__EVAL_41;
  wire  rsource__EVAL_42;
  wire [6:0] rsource__EVAL_43;
  wire [24:0] rsource__EVAL_44;
  wire [24:0] rsource__EVAL_45;
  wire  rsource__EVAL_46;
  wire  rsource__EVAL_47;
  wire [31:0] rsource__EVAL_48;
  wire [2:0] rsource__EVAL_49;
  wire  rsource__EVAL_50;
  wire [6:0] rsource__EVAL_51;
  wire [1:0] rsource__EVAL_52;
  wire  rsource__EVAL_53;
  wire [3:0] rsource__EVAL_54;
  wire  rsource__EVAL_55;
  wire [6:0] rsource__EVAL_56;
  wire [2:0] rsource__EVAL_57;
  wire [31:0] rsource__EVAL_58;
  wire [1:0] rsource__EVAL_59;
  wire  rsource__EVAL_60;
  wire [2:0] widget__EVAL;
  wire [2:0] widget__EVAL_0;
  wire [2:0] widget__EVAL_1;
  wire [31:0] widget__EVAL_2;
  wire  widget__EVAL_3;
  wire  widget__EVAL_4;
  wire  widget__EVAL_5;
  wire  widget__EVAL_6;
  wire  widget__EVAL_7;
  wire [31:0] widget__EVAL_8;
  wire [1:0] widget__EVAL_9;
  wire  widget__EVAL_10;
  wire  widget__EVAL_11;
  wire [1:0] widget__EVAL_12;
  wire [6:0] widget__EVAL_13;
  wire  widget__EVAL_14;
  wire  widget__EVAL_15;
  wire [2:0] widget__EVAL_16;
  wire [2:0] widget__EVAL_17;
  wire  widget__EVAL_18;
  wire  widget__EVAL_19;
  wire [3:0] widget__EVAL_20;
  wire [2:0] widget__EVAL_21;
  wire [31:0] widget__EVAL_22;
  wire [6:0] widget__EVAL_23;
  wire [3:0] widget__EVAL_24;
  wire  widget__EVAL_25;
  wire  widget__EVAL_26;
  wire  widget__EVAL_27;
  wire [2:0] widget__EVAL_28;
  wire [2:0] widget__EVAL_29;
  wire [24:0] widget__EVAL_30;
  wire  widget__EVAL_31;
  wire [31:0] widget__EVAL_32;
  wire  widget__EVAL_33;
  wire [2:0] widget__EVAL_34;
  wire [24:0] widget__EVAL_35;
  wire  widget__EVAL_36;
  wire  widget__EVAL_37;
  wire [6:0] widget__EVAL_38;
  wire [6:0] widget__EVAL_39;
  wire [2:0] widget__EVAL_40;
  wire  buffer__EVAL;
  wire [2:0] buffer__EVAL_0;
  wire [2:0] buffer__EVAL_1;
  wire [1:0] buffer__EVAL_2;
  wire [1:0] buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire [2:0] buffer__EVAL_5;
  wire [2:0] buffer__EVAL_6;
  wire [2:0] buffer__EVAL_7;
  wire [24:0] buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [2:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire [2:0] buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire [31:0] buffer__EVAL_14;
  wire [24:0] buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire [2:0] buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire [3:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire [6:0] buffer__EVAL_23;
  wire [2:0] buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire [6:0] buffer__EVAL_26;
  wire [6:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [2:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire [6:0] buffer__EVAL_32;
  wire [31:0] buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire  buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [31:0] buffer__EVAL_37;
  wire [31:0] buffer__EVAL_38;
  wire [3:0] buffer__EVAL_39;
  wire  buffer__EVAL_40;
  SiFive__EVAL_147 rsource (
    ._EVAL(rsource__EVAL),
    ._EVAL_0(rsource__EVAL_0),
    ._EVAL_1(rsource__EVAL_1),
    ._EVAL_2(rsource__EVAL_2),
    ._EVAL_3(rsource__EVAL_3),
    ._EVAL_4(rsource__EVAL_4),
    ._EVAL_5(rsource__EVAL_5),
    ._EVAL_6(rsource__EVAL_6),
    ._EVAL_7(rsource__EVAL_7),
    ._EVAL_8(rsource__EVAL_8),
    ._EVAL_9(rsource__EVAL_9),
    ._EVAL_10(rsource__EVAL_10),
    ._EVAL_11(rsource__EVAL_11),
    ._EVAL_12(rsource__EVAL_12),
    ._EVAL_13(rsource__EVAL_13),
    ._EVAL_14(rsource__EVAL_14),
    ._EVAL_15(rsource__EVAL_15),
    ._EVAL_16(rsource__EVAL_16),
    ._EVAL_17(rsource__EVAL_17),
    ._EVAL_18(rsource__EVAL_18),
    ._EVAL_19(rsource__EVAL_19),
    ._EVAL_20(rsource__EVAL_20),
    ._EVAL_21(rsource__EVAL_21),
    ._EVAL_22(rsource__EVAL_22),
    ._EVAL_23(rsource__EVAL_23),
    ._EVAL_24(rsource__EVAL_24),
    ._EVAL_25(rsource__EVAL_25),
    ._EVAL_26(rsource__EVAL_26),
    ._EVAL_27(rsource__EVAL_27),
    ._EVAL_28(rsource__EVAL_28),
    ._EVAL_29(rsource__EVAL_29),
    ._EVAL_30(rsource__EVAL_30),
    ._EVAL_31(rsource__EVAL_31),
    ._EVAL_32(rsource__EVAL_32),
    ._EVAL_33(rsource__EVAL_33),
    ._EVAL_34(rsource__EVAL_34),
    ._EVAL_35(rsource__EVAL_35),
    ._EVAL_36(rsource__EVAL_36),
    ._EVAL_37(rsource__EVAL_37),
    ._EVAL_38(rsource__EVAL_38),
    ._EVAL_39(rsource__EVAL_39),
    ._EVAL_40(rsource__EVAL_40),
    ._EVAL_41(rsource__EVAL_41),
    ._EVAL_42(rsource__EVAL_42),
    ._EVAL_43(rsource__EVAL_43),
    ._EVAL_44(rsource__EVAL_44),
    ._EVAL_45(rsource__EVAL_45),
    ._EVAL_46(rsource__EVAL_46),
    ._EVAL_47(rsource__EVAL_47),
    ._EVAL_48(rsource__EVAL_48),
    ._EVAL_49(rsource__EVAL_49),
    ._EVAL_50(rsource__EVAL_50),
    ._EVAL_51(rsource__EVAL_51),
    ._EVAL_52(rsource__EVAL_52),
    ._EVAL_53(rsource__EVAL_53),
    ._EVAL_54(rsource__EVAL_54),
    ._EVAL_55(rsource__EVAL_55),
    ._EVAL_56(rsource__EVAL_56),
    ._EVAL_57(rsource__EVAL_57),
    ._EVAL_58(rsource__EVAL_58),
    ._EVAL_59(rsource__EVAL_59),
    ._EVAL_60(rsource__EVAL_60)
  );
  SiFive__EVAL_149 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36),
    ._EVAL_37(widget__EVAL_37),
    ._EVAL_38(widget__EVAL_38),
    ._EVAL_39(widget__EVAL_39),
    ._EVAL_40(widget__EVAL_40)
  );
  SiFive__EVAL_151 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40)
  );
  assign buffer__EVAL_9 = _EVAL_39;
  assign widget__EVAL_0 = rsource__EVAL_16;
  assign rsource__EVAL = _EVAL_22;
  assign buffer__EVAL_24 = _EVAL_33;
  assign _EVAL_30 = buffer__EVAL_36;
  assign buffer__EVAL_11 = widget__EVAL_4;
  assign rsource__EVAL_34 = _EVAL_15;
  assign _EVAL_8 = rsource__EVAL_38;
  assign rsource__EVAL_53 = widget__EVAL_31;
  assign _EVAL_54 = rsource__EVAL_28;
  assign widget__EVAL_30 = buffer__EVAL_15;
  assign buffer__EVAL_39 = _EVAL_31;
  assign rsource__EVAL_25 = _EVAL_45;
  assign _EVAL_1 = buffer__EVAL_28;
  assign rsource__EVAL_59 = _EVAL_46;
  assign buffer__EVAL_8 = _EVAL_35;
  assign widget__EVAL_37 = rsource__EVAL_14;
  assign widget__EVAL_8 = rsource__EVAL_18;
  assign rsource__EVAL_6 = _EVAL_10;
  assign widget__EVAL_20 = buffer__EVAL_21;
  assign rsource__EVAL_47 = _EVAL_60;
  assign buffer__EVAL_29 = _EVAL_22;
  assign _EVAL_27 = rsource__EVAL_3;
  assign _EVAL_49 = buffer__EVAL_22;
  assign _EVAL_38 = rsource__EVAL_20;
  assign buffer__EVAL_2 = widget__EVAL_9;
  assign buffer__EVAL_31 = widget__EVAL_14;
  assign _EVAL_5 = buffer__EVAL_27;
  assign rsource__EVAL_17 = _EVAL_43;
  assign widget__EVAL_2 = buffer__EVAL_37;
  assign rsource__EVAL_10 = _EVAL_18;
  assign widget__EVAL_40 = buffer__EVAL_10;
  assign widget__EVAL_6 = buffer__EVAL_16;
  assign _EVAL_34 = rsource__EVAL_27;
  assign _EVAL_59 = buffer__EVAL_38;
  assign buffer__EVAL_33 = widget__EVAL_22;
  assign _EVAL_4 = buffer__EVAL_19;
  assign rsource__EVAL_37 = _EVAL_24;
  assign buffer__EVAL_13 = _EVAL_53;
  assign rsource__EVAL_13 = widget__EVAL_33;
  assign rsource__EVAL_4 = _EVAL_11;
  assign _EVAL_20 = rsource__EVAL_42;
  assign _EVAL_42 = rsource__EVAL_58;
  assign rsource__EVAL_21 = widget__EVAL_1;
  assign widget__EVAL_3 = _EVAL_56;
  assign widget__EVAL = rsource__EVAL_31;
  assign buffer__EVAL_40 = widget__EVAL_10;
  assign _EVAL_28 = rsource__EVAL_33;
  assign widget__EVAL_12 = rsource__EVAL_29;
  assign rsource__EVAL_8 = widget__EVAL_24;
  assign widget__EVAL_11 = buffer__EVAL_20;
  assign buffer__EVAL = _EVAL_41;
  assign rsource__EVAL_32 = widget__EVAL_16;
  assign _EVAL_51 = rsource__EVAL_36;
  assign rsource__EVAL_57 = _EVAL_12;
  assign _EVAL = rsource__EVAL_41;
  assign _EVAL_44 = rsource__EVAL_45;
  assign widget__EVAL_29 = buffer__EVAL_6;
  assign rsource__EVAL_43 = _EVAL_13;
  assign buffer__EVAL_32 = _EVAL_40;
  assign widget__EVAL_27 = _EVAL_22;
  assign widget__EVAL_19 = rsource__EVAL_7;
  assign rsource__EVAL_46 = _EVAL_17;
  assign _EVAL_23 = buffer__EVAL_4;
  assign rsource__EVAL_52 = _EVAL_50;
  assign rsource__EVAL_44 = widget__EVAL_35;
  assign widget__EVAL_26 = buffer__EVAL_18;
  assign buffer__EVAL_7 = widget__EVAL_21;
  assign buffer__EVAL_34 = widget__EVAL_18;
  assign _EVAL_48 = rsource__EVAL_39;
  assign rsource__EVAL_5 = _EVAL_6;
  assign _EVAL_19 = rsource__EVAL_35;
  assign rsource__EVAL_26 = widget__EVAL_32;
  assign _EVAL_21 = rsource__EVAL_49;
  assign widget__EVAL_38 = rsource__EVAL_56;
  assign _EVAL_36 = rsource__EVAL_51;
  assign widget__EVAL_36 = rsource__EVAL_55;
  assign buffer__EVAL_25 = _EVAL_56;
  assign rsource__EVAL_2 = _EVAL_9;
  assign rsource__EVAL_40 = _EVAL_2;
  assign rsource__EVAL_11 = widget__EVAL_13;
  assign rsource__EVAL_0 = _EVAL_37;
  assign _EVAL_58 = rsource__EVAL_48;
  assign rsource__EVAL_1 = _EVAL_3;
  assign widget__EVAL_17 = buffer__EVAL_0;
  assign _EVAL_25 = rsource__EVAL_54;
  assign _EVAL_55 = buffer__EVAL_17;
  assign buffer__EVAL_12 = _EVAL_47;
  assign buffer__EVAL_1 = _EVAL_7;
  assign _EVAL_26 = rsource__EVAL_19;
  assign buffer__EVAL_30 = widget__EVAL_34;
  assign buffer__EVAL_35 = widget__EVAL_15;
  assign rsource__EVAL_50 = _EVAL_16;
  assign buffer__EVAL_14 = _EVAL_57;
  assign widget__EVAL_5 = rsource__EVAL_22;
  assign _EVAL_32 = buffer__EVAL_3;
  assign widget__EVAL_7 = rsource__EVAL_9;
  assign widget__EVAL_23 = buffer__EVAL_23;
  assign _EVAL_29 = buffer__EVAL_5;
  assign _EVAL_14 = rsource__EVAL_15;
  assign rsource__EVAL_60 = widget__EVAL_25;
  assign buffer__EVAL_26 = widget__EVAL_39;
  assign rsource__EVAL_12 = widget__EVAL_28;
  assign rsource__EVAL_24 = _EVAL_56;
  assign _EVAL_52 = rsource__EVAL_23;
  assign rsource__EVAL_30 = _EVAL_0;
endmodule
