//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_264(
  input  [2:0]  _EVAL,
  output [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [7:0]  _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  output [31:0] _EVAL_5,
  input  [2:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output [3:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  output [1:0]  _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  output [31:0] _EVAL_18,
  output [2:0]  _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output [3:0]  _EVAL_25,
  output [1:0]  _EVAL_26,
  output        _EVAL_27,
  output [31:0] _EVAL_28,
  output [2:0]  _EVAL_29,
  output [63:0] _EVAL_30,
  output [2:0]  _EVAL_31,
  input  [3:0]  _EVAL_32,
  input  [63:0] _EVAL_33,
  output [2:0]  _EVAL_34,
  input  [63:0] _EVAL_35,
  output [3:0]  _EVAL_36,
  input  [63:0] _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  output [2:0]  _EVAL_40,
  input  [1:0]  _EVAL_41,
  output        _EVAL_42,
  output [2:0]  _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output        _EVAL_46,
  output [2:0]  _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  output        _EVAL_50,
  input  [2:0]  _EVAL_51,
  input  [3:0]  _EVAL_52,
  input         _EVAL_53,
  output        _EVAL_54,
  output        _EVAL_55,
  input  [31:0] _EVAL_56,
  input         _EVAL_57,
  input  [2:0]  _EVAL_58,
  output        _EVAL_59,
  input         _EVAL_60,
  input  [3:0]  _EVAL_61,
  output        _EVAL_62,
  output [63:0] _EVAL_63,
  input  [2:0]  _EVAL_64,
  output [63:0] _EVAL_65,
  input  [31:0] _EVAL_66,
  output        _EVAL_67,
  output [7:0]  _EVAL_68,
  input  [31:0] _EVAL_69,
  input  [2:0]  _EVAL_70,
  input  [2:0]  _EVAL_71,
  input         _EVAL_72
);
  assign _EVAL_43 = _EVAL_70;
  assign _EVAL_5 = _EVAL_69;
  assign _EVAL_24 = _EVAL_60;
  assign _EVAL_29 = _EVAL_58;
  assign _EVAL_63 = _EVAL_35;
  assign _EVAL_26 = _EVAL_41;
  assign _EVAL_27 = _EVAL_44;
  assign _EVAL_40 = _EVAL;
  assign _EVAL_30 = _EVAL_37;
  assign _EVAL_68 = _EVAL_2;
  assign _EVAL_21 = _EVAL_12;
  assign _EVAL_15 = _EVAL_11;
  assign _EVAL_23 = _EVAL_72;
  assign _EVAL_36 = _EVAL_61;
  assign _EVAL_62 = _EVAL_8;
  assign _EVAL_0 = _EVAL_71;
  assign _EVAL_65 = _EVAL_33;
  assign _EVAL_20 = _EVAL_14;
  assign _EVAL_47 = _EVAL_64;
  assign _EVAL_67 = _EVAL_57;
  assign _EVAL_46 = _EVAL_1;
  assign _EVAL_42 = _EVAL_53;
  assign _EVAL_50 = _EVAL_48;
  assign _EVAL_34 = _EVAL_51;
  assign _EVAL_55 = _EVAL_38;
  assign _EVAL_31 = _EVAL_13;
  assign _EVAL_16 = _EVAL_17;
  assign _EVAL_25 = _EVAL_52;
  assign _EVAL_10 = _EVAL_32;
  assign _EVAL_3 = _EVAL_22;
  assign _EVAL_54 = _EVAL_45;
  assign _EVAL_18 = _EVAL_56;
  assign _EVAL_28 = _EVAL_66;
  assign _EVAL_7 = _EVAL_9;
  assign _EVAL_19 = _EVAL_6;
  assign _EVAL_59 = _EVAL_4;
endmodule
