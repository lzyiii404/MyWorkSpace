//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_329(
  input         _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [10:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6
);
  reg  _EVAL_7;
  reg [31:0] _RAND_0;
  reg  _EVAL_13;
  reg [31:0] _RAND_1;
  reg  _EVAL_19;
  reg [31:0] _RAND_2;
  reg  _EVAL_24;
  reg [31:0] _RAND_3;
  reg  _EVAL_28;
  reg [31:0] _RAND_4;
  reg  _EVAL_29;
  reg [31:0] _RAND_5;
  reg  _EVAL_34;
  reg [31:0] _RAND_6;
  reg  _EVAL_37;
  reg [31:0] _RAND_7;
  reg  _EVAL_40;
  reg [31:0] _RAND_8;
  reg  _EVAL_42;
  reg [31:0] _RAND_9;
  reg  _EVAL_45;
  reg [31:0] _RAND_10;
  reg  _EVAL_52;
  reg [31:0] _RAND_11;
  reg  _EVAL_55;
  reg [31:0] _RAND_12;
  reg  _EVAL_57;
  reg [31:0] _RAND_13;
  reg  _EVAL_60;
  reg [31:0] _RAND_14;
  reg  _EVAL_67;
  reg [31:0] _RAND_15;
  reg  _EVAL_71;
  reg [31:0] _RAND_16;
  reg  _EVAL_73;
  reg [31:0] _RAND_17;
  reg  _EVAL_81;
  reg [31:0] _RAND_18;
  reg  _EVAL_84;
  reg [31:0] _RAND_19;
  reg  _EVAL_85;
  reg [31:0] _RAND_20;
  reg  _EVAL_88;
  reg [31:0] _RAND_21;
  reg  _EVAL_90;
  reg [31:0] _RAND_22;
  reg  _EVAL_91;
  reg [31:0] _RAND_23;
  reg  _EVAL_93;
  reg [31:0] _RAND_24;
  reg  _EVAL_95;
  reg [31:0] _RAND_25;
  reg  _EVAL_101;
  reg [31:0] _RAND_26;
  reg  _EVAL_102;
  reg [31:0] _RAND_27;
  reg  _EVAL_109;
  reg [31:0] _RAND_28;
  reg  _EVAL_110;
  reg [31:0] _RAND_29;
  reg  _EVAL_113;
  reg [31:0] _RAND_30;
  reg  _EVAL_114;
  reg [31:0] _RAND_31;
  wire [31:0] _EVAL_36;
  wire  _EVAL_14;
  wire  _EVAL_104;
  wire  _EVAL_22;
  wire  _EVAL_108;
  wire  _EVAL_100;
  wire  _EVAL_62;
  wire  _EVAL_69;
  wire  _EVAL_41;
  wire  _EVAL_77;
  wire  _EVAL_64;
  wire  _EVAL_53;
  wire  _EVAL_74;
  wire  _EVAL_12;
  wire  _EVAL_63;
  wire  _EVAL_103;
  wire  _EVAL_89;
  wire  _EVAL_16;
  wire  _EVAL_65;
  wire  _EVAL_92;
  wire  _EVAL_8;
  wire  _EVAL_32;
  wire  _EVAL_68;
  wire  _EVAL_33;
  wire  _EVAL_17;
  wire  _EVAL_30;
  wire  _EVAL_56;
  wire  _EVAL_35;
  wire  _EVAL_94;
  wire  _EVAL_20;
  wire  _EVAL_15;
  wire  _EVAL_39;
  wire  _EVAL_61;
  assign _EVAL_36 = {20'h20000,_EVAL_4,1'h1};
  assign _EVAL_14 = _EVAL_36[12];
  assign _EVAL_104 = _EVAL_36[11];
  assign _EVAL_22 = _EVAL_36[22];
  assign _EVAL_108 = _EVAL_36[14];
  assign _EVAL_100 = _EVAL_36[21];
  assign _EVAL_62 = _EVAL_36[26];
  assign _EVAL_69 = _EVAL_36[16];
  assign _EVAL_41 = _EVAL_36[0];
  assign _EVAL_77 = _EVAL_36[5];
  assign _EVAL_64 = _EVAL_36[3];
  assign _EVAL_53 = _EVAL_36[10];
  assign _EVAL_74 = _EVAL_36[8];
  assign _EVAL_12 = _EVAL_36[27];
  assign _EVAL_63 = _EVAL_36[2];
  assign _EVAL_103 = _EVAL_36[28];
  assign _EVAL_89 = _EVAL_36[7];
  assign _EVAL_16 = _EVAL_36[29];
  assign _EVAL_65 = _EVAL_36[19];
  assign _EVAL_92 = _EVAL_36[24];
  assign _EVAL_8 = _EVAL_36[20];
  assign _EVAL_32 = _EVAL_36[23];
  assign _EVAL_68 = _EVAL_36[9];
  assign _EVAL_33 = _EVAL_36[17];
  assign _EVAL_17 = _EVAL_36[25];
  assign _EVAL_30 = _EVAL_36[1];
  assign _EVAL_56 = _EVAL_36[31];
  assign _EVAL_35 = _EVAL_36[13];
  assign _EVAL_94 = _EVAL_36[4];
  assign _EVAL_20 = _EVAL_36[30];
  assign _EVAL_15 = _EVAL_36[15];
  assign _EVAL_39 = _EVAL_36[6];
  assign _EVAL_61 = _EVAL_36[18];
  assign _EVAL_0 = _EVAL_93;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_7 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_13 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_19 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_24 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_28 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_29 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_34 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_37 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_40 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_42 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_45 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_52 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_55 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_57 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_60 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_67 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_71 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_73 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_81 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_84 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_85 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_88 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_90 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_91 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_93 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_95 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_101 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_102 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_109 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_110 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_113 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_114 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_1) begin
    if (_EVAL_5) begin
      _EVAL_7 <= _EVAL_68;
    end else begin
      if (_EVAL_2) begin
        _EVAL_7 <= _EVAL_110;
      end
    end
    if (_EVAL_5) begin
      _EVAL_13 <= _EVAL_63;
    end else begin
      if (_EVAL_2) begin
        _EVAL_13 <= _EVAL_57;
      end
    end
    if (_EVAL_5) begin
      _EVAL_19 <= _EVAL_16;
    end else begin
      if (_EVAL_2) begin
        _EVAL_19 <= _EVAL_90;
      end
    end
    if (_EVAL_5) begin
      _EVAL_24 <= _EVAL_94;
    end else begin
      if (_EVAL_2) begin
        _EVAL_24 <= _EVAL_101;
      end
    end
    if (_EVAL_5) begin
      _EVAL_28 <= _EVAL_62;
    end else begin
      if (_EVAL_2) begin
        _EVAL_28 <= _EVAL_29;
      end
    end
    if (_EVAL_5) begin
      _EVAL_29 <= _EVAL_12;
    end else begin
      if (_EVAL_2) begin
        _EVAL_29 <= _EVAL_95;
      end
    end
    if (_EVAL_5) begin
      _EVAL_34 <= _EVAL_14;
    end else begin
      if (_EVAL_2) begin
        _EVAL_34 <= _EVAL_91;
      end
    end
    if (_EVAL_5) begin
      _EVAL_37 <= _EVAL_108;
    end else begin
      if (_EVAL_2) begin
        _EVAL_37 <= _EVAL_113;
      end
    end
    if (_EVAL_5) begin
      _EVAL_40 <= _EVAL_92;
    end else begin
      if (_EVAL_2) begin
        _EVAL_40 <= _EVAL_60;
      end
    end
    if (_EVAL_5) begin
      _EVAL_42 <= _EVAL_100;
    end else begin
      if (_EVAL_2) begin
        _EVAL_42 <= _EVAL_109;
      end
    end
    if (_EVAL_5) begin
      _EVAL_45 <= _EVAL_39;
    end else begin
      if (_EVAL_2) begin
        _EVAL_45 <= _EVAL_84;
      end
    end
    if (_EVAL_5) begin
      _EVAL_52 <= _EVAL_61;
    end else begin
      if (_EVAL_2) begin
        _EVAL_52 <= _EVAL_71;
      end
    end
    if (_EVAL_5) begin
      _EVAL_55 <= _EVAL_8;
    end else begin
      if (_EVAL_2) begin
        _EVAL_55 <= _EVAL_42;
      end
    end
    if (_EVAL_5) begin
      _EVAL_57 <= _EVAL_64;
    end else begin
      if (_EVAL_2) begin
        _EVAL_57 <= _EVAL_24;
      end
    end
    if (_EVAL_5) begin
      _EVAL_60 <= _EVAL_17;
    end else begin
      if (_EVAL_2) begin
        _EVAL_60 <= _EVAL_28;
      end
    end
    if (_EVAL_5) begin
      _EVAL_67 <= _EVAL_33;
    end else begin
      if (_EVAL_2) begin
        _EVAL_67 <= _EVAL_52;
      end
    end
    if (_EVAL_5) begin
      _EVAL_71 <= _EVAL_65;
    end else begin
      if (_EVAL_2) begin
        _EVAL_71 <= _EVAL_55;
      end
    end
    if (_EVAL_5) begin
      _EVAL_73 <= _EVAL_56;
    end else begin
      if (_EVAL_2) begin
        _EVAL_73 <= _EVAL_3;
      end
    end
    if (_EVAL_5) begin
      _EVAL_81 <= _EVAL_69;
    end else begin
      if (_EVAL_2) begin
        _EVAL_81 <= _EVAL_67;
      end
    end
    if (_EVAL_5) begin
      _EVAL_84 <= _EVAL_89;
    end else begin
      if (_EVAL_2) begin
        _EVAL_84 <= _EVAL_88;
      end
    end
    if (_EVAL_5) begin
      _EVAL_85 <= _EVAL_32;
    end else begin
      if (_EVAL_2) begin
        _EVAL_85 <= _EVAL_40;
      end
    end
    if (_EVAL_5) begin
      _EVAL_88 <= _EVAL_74;
    end else begin
      if (_EVAL_2) begin
        _EVAL_88 <= _EVAL_7;
      end
    end
    if (_EVAL_5) begin
      _EVAL_90 <= _EVAL_20;
    end else begin
      if (_EVAL_2) begin
        _EVAL_90 <= _EVAL_73;
      end
    end
    if (_EVAL_5) begin
      _EVAL_91 <= _EVAL_35;
    end else begin
      if (_EVAL_2) begin
        _EVAL_91 <= _EVAL_37;
      end
    end
    if (_EVAL_5) begin
      _EVAL_93 <= _EVAL_41;
    end else begin
      if (_EVAL_2) begin
        _EVAL_93 <= _EVAL_114;
      end
    end
    if (_EVAL_5) begin
      _EVAL_95 <= _EVAL_103;
    end else begin
      if (_EVAL_2) begin
        _EVAL_95 <= _EVAL_19;
      end
    end
    if (_EVAL_5) begin
      _EVAL_101 <= _EVAL_77;
    end else begin
      if (_EVAL_2) begin
        _EVAL_101 <= _EVAL_45;
      end
    end
    if (_EVAL_5) begin
      _EVAL_102 <= _EVAL_104;
    end else begin
      if (_EVAL_2) begin
        _EVAL_102 <= _EVAL_34;
      end
    end
    if (_EVAL_5) begin
      _EVAL_109 <= _EVAL_22;
    end else begin
      if (_EVAL_2) begin
        _EVAL_109 <= _EVAL_85;
      end
    end
    if (_EVAL_5) begin
      _EVAL_110 <= _EVAL_53;
    end else begin
      if (_EVAL_2) begin
        _EVAL_110 <= _EVAL_102;
      end
    end
    if (_EVAL_5) begin
      _EVAL_113 <= _EVAL_15;
    end else begin
      if (_EVAL_2) begin
        _EVAL_113 <= _EVAL_81;
      end
    end
    if (_EVAL_5) begin
      _EVAL_114 <= _EVAL_30;
    end else begin
      if (_EVAL_2) begin
        _EVAL_114 <= _EVAL_13;
      end
    end
  end
endmodule
