//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_81_assert(
  input  [5:0]  _EVAL,
  input         _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input  [5:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input  [31:0] _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_20;
  reg [31:0] _RAND_0;
  reg [5:0] _EVAL_22;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_30;
  reg [31:0] _RAND_2;
  reg  _EVAL_58;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_70;
  reg [31:0] _RAND_4;
  reg [5:0] _EVAL_82;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_105;
  reg [31:0] _RAND_6;
  reg [5:0] _EVAL_147;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_168;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_292;
  reg [31:0] _RAND_9;
  reg  _EVAL_304;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_306;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_314;
  reg [31:0] _RAND_12;
  reg [32:0] _EVAL_328;
  reg [63:0] _RAND_13;
  reg [5:0] _EVAL_347;
  reg [31:0] _RAND_14;
  reg [1:0] _EVAL_349;
  reg [31:0] _RAND_15;
  reg [5:0] _EVAL_363;
  reg [31:0] _RAND_16;
  wire  _EVAL_64;
  wire  _EVAL_124;
  wire  _EVAL_99;
  wire  _EVAL_223;
  wire  _EVAL_336;
  wire  _EVAL_84;
  wire  _EVAL_139;
  wire  _EVAL_212;
  wire  _EVAL_37;
  wire [31:0] _EVAL_264;
  wire [32:0] _EVAL_340;
  wire  _EVAL_106;
  wire  _EVAL_333;
  wire  _EVAL_40;
  wire [22:0] _EVAL_80;
  wire [7:0] _EVAL_32;
  wire [7:0] _EVAL_214;
  wire [5:0] _EVAL_252;
  wire [5:0] _EVAL_192;
  wire  _EVAL_361;
  wire  _EVAL_227;
  wire [1:0] _EVAL_182;
  wire [1:0] _EVAL_152;
  wire  _EVAL_158;
  wire  _EVAL_342;
  wire  _EVAL_153;
  wire  _EVAL_131;
  wire  _EVAL_109;
  wire  _EVAL_358;
  wire [2:0] _EVAL_102;
  wire  _EVAL_229;
  wire  _EVAL_324;
  wire  _EVAL_186;
  wire  _EVAL_52;
  wire  _EVAL_156;
  wire  _EVAL_85;
  wire  _EVAL_120;
  wire  _EVAL_261;
  wire  _EVAL_180;
  wire  _EVAL_195;
  wire  _EVAL_295;
  wire  _EVAL_81;
  wire  _EVAL_235;
  wire [32:0] _EVAL_239;
  wire [32:0] _EVAL_344;
  wire  _EVAL_123;
  wire  _EVAL_35;
  wire  _EVAL_268;
  wire  _EVAL_155;
  wire  _EVAL_283;
  wire  _EVAL_121;
  wire [31:0] _EVAL_50;
  wire [32:0] _EVAL_110;
  wire [32:0] _EVAL_219;
  wire [32:0] _EVAL_309;
  wire  _EVAL_202;
  wire  _EVAL_140;
  wire [63:0] _EVAL_28;
  wire  _EVAL_128;
  wire [22:0] _EVAL_220;
  wire [7:0] _EVAL_111;
  wire [7:0] _EVAL_162;
  wire [5:0] _EVAL_134;
  wire [31:0] _EVAL_93;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_273;
  wire [32:0] _EVAL_72;
  wire  _EVAL_126;
  wire  _EVAL_356;
  wire  _EVAL_245;
  wire [5:0] _EVAL_320;
  wire [31:0] _EVAL_298;
  wire [32:0] _EVAL_203;
  wire  _EVAL_281;
  wire  _EVAL_199;
  wire  _EVAL_250;
  wire  _EVAL_169;
  wire  _EVAL_200;
  wire  _EVAL_346;
  wire  _EVAL_94;
  wire  _EVAL_308;
  wire  _EVAL_209;
  wire  _EVAL_160;
  wire  _EVAL_62;
  wire  _EVAL_290;
  wire  _EVAL_142;
  wire  _EVAL_337;
  wire  _EVAL_318;
  wire  _EVAL_213;
  wire  _EVAL_132;
  wire [3:0] _EVAL_351;
  wire [3:0] _EVAL_315;
  wire [3:0] _EVAL_74;
  wire  _EVAL_232;
  wire  _EVAL_312;
  wire  _EVAL_260;
  wire [63:0] _EVAL_189;
  wire  _EVAL_159;
  wire [31:0] _EVAL_236;
  wire [32:0] _EVAL_77;
  wire [32:0] _EVAL_331;
  wire [32:0] _EVAL_263;
  wire  _EVAL_362;
  wire [31:0] _EVAL_329;
  wire [32:0] _EVAL_73;
  wire [32:0] _EVAL_248;
  wire [32:0] _EVAL_341;
  wire  _EVAL_231;
  wire  _EVAL_246;
  wire  _EVAL_364;
  wire  _EVAL_164;
  wire [32:0] _EVAL_143;
  wire [32:0] _EVAL_92;
  wire  _EVAL_319;
  wire  _EVAL_345;
  wire  _EVAL_230;
  wire  _EVAL_146;
  wire  _EVAL_301;
  wire  _EVAL_265;
  wire  _EVAL_357;
  wire  _EVAL_27;
  wire  _EVAL_338;
  wire  _EVAL_293;
  wire  _EVAL_233;
  wire  _EVAL_136;
  wire  _EVAL_208;
  wire  _EVAL_326;
  wire  _EVAL_332;
  wire  _EVAL_138;
  wire [32:0] _EVAL_45;
  wire [32:0] _EVAL_49;
  wire [32:0] _EVAL_278;
  wire  _EVAL_282;
  wire [31:0] _EVAL_95;
  wire [32:0] _EVAL_280;
  wire [32:0] _EVAL_47;
  wire  _EVAL_355;
  wire  _EVAL_23;
  wire  _EVAL_174;
  wire  _EVAL_104;
  wire  _EVAL_198;
  wire [63:0] _EVAL_48;
  wire [32:0] _EVAL_129;
  wire  _EVAL_55;
  wire  _EVAL_274;
  wire  _EVAL_135;
  wire  _EVAL_86;
  wire  _EVAL_352;
  wire [63:0] _EVAL_237;
  wire [32:0] _EVAL_191;
  wire  _EVAL_272;
  wire  _EVAL_316;
  wire  _EVAL_144;
  wire  _EVAL_218;
  wire  _EVAL_173;
  wire  _EVAL_38;
  wire  _EVAL_216;
  wire  _EVAL_127;
  wire  _EVAL_339;
  wire  _EVAL_217;
  wire  _EVAL_269;
  wire  _EVAL_90;
  wire  _EVAL_221;
  wire  _EVAL_194;
  wire [32:0] _EVAL_67;
  wire [32:0] _EVAL_175;
  wire [32:0] _EVAL_242;
  wire  _EVAL_42;
  wire  _EVAL_255;
  wire  _EVAL_310;
  wire  _EVAL_33;
  wire  _EVAL_228;
  wire  _EVAL_240;
  wire  _EVAL_226;
  wire [32:0] _EVAL_207;
  wire  _EVAL_97;
  wire  _EVAL_39;
  wire  _EVAL_353;
  wire  _EVAL_88;
  wire  _EVAL_154;
  wire  _EVAL_305;
  wire  _EVAL_63;
  wire  _EVAL_76;
  wire [32:0] _EVAL_57;
  wire  _EVAL_277;
  wire  _EVAL_150;
  wire [31:0] _EVAL_279;
  wire [32:0] _EVAL_36;
  wire [32:0] _EVAL_65;
  wire [32:0] _EVAL_322;
  wire  _EVAL_151;
  wire  _EVAL_299;
  wire  _EVAL_61;
  wire  _EVAL_19;
  wire [31:0] _EVAL_60;
  wire  _EVAL_53;
  wire [31:0] _EVAL_287;
  wire  _EVAL_204;
  wire  _EVAL_215;
  wire  _EVAL_112;
  wire  _EVAL_188;
  wire  _EVAL_161;
  wire [2:0] _EVAL_56;
  wire  _EVAL_270;
  wire  _EVAL_113;
  wire  _EVAL_26;
  wire  _EVAL_348;
  wire  _EVAL_354;
  wire  _EVAL_177;
  wire  _EVAL_107;
  wire  _EVAL_247;
  wire  _EVAL_87;
  wire  _EVAL_285;
  wire [5:0] _EVAL_176;
  wire  _EVAL_259;
  wire  _EVAL_78;
  wire  _EVAL_108;
  wire  _EVAL_313;
  wire  _EVAL_100;
  wire [32:0] _EVAL_271;
  wire [32:0] _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_311;
  wire  _EVAL_249;
  wire  _EVAL_251;
  wire  _EVAL_66;
  wire  _EVAL_266;
  wire  _EVAL_149;
  wire  _EVAL_238;
  wire  _EVAL_296;
  wire  _EVAL_288;
  wire  _EVAL_205;
  wire  _EVAL_335;
  wire  _EVAL_222;
  wire  _EVAL_257;
  wire [31:0] _EVAL_157;
  wire  _EVAL_130;
  wire  _EVAL_297;
  wire  _EVAL_114;
  wire  _EVAL_171;
  wire  _EVAL_234;
  wire  _EVAL_68;
  wire [5:0] _EVAL_183;
  wire  _EVAL_276;
  wire  _EVAL_34;
  wire  _EVAL_343;
  wire  _EVAL_225;
  wire  _EVAL_125;
  wire  _EVAL_211;
  wire  _EVAL_44;
  wire  _EVAL_286;
  wire  _EVAL_284;
  wire  _EVAL_46;
  wire [3:0] _EVAL_334;
  wire  _EVAL_166;
  wire  _EVAL_302;
  wire  _EVAL_167;
  wire  _EVAL_291;
  wire  _EVAL_165;
  wire  _EVAL_327;
  wire  _EVAL_256;
  wire  _EVAL_115;
  wire  _EVAL_323;
  wire  _EVAL_148;
  wire  _EVAL_119;
  wire  _EVAL_190;
  wire  _EVAL_184;
  wire  _EVAL_187;
  wire  _EVAL_197;
  wire  _EVAL_179;
  wire  _EVAL_141;
  wire  _EVAL_181;
  wire  _EVAL_71;
  wire  _EVAL_262;
  wire  _EVAL_206;
  wire  _EVAL_196;
  wire  _EVAL_31;
  wire  _EVAL_185;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_137;
  wire  _EVAL_317;
  wire  _EVAL_244;
  wire  _EVAL_258;
  wire  _EVAL_193;
  wire  _EVAL_122;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_41;
  wire  _EVAL_101;
  wire  _EVAL_178;
  wire  _EVAL_54;
  wire  _EVAL_29;
  wire  _EVAL_145;
  wire  _EVAL_98;
  wire  _EVAL_83;
  wire  _EVAL_91;
  wire  _EVAL_210;
  wire  _EVAL_303;
  wire  _EVAL_163;
  wire  _EVAL_254;
  wire  _EVAL_59;
  wire  _EVAL_75;
  wire  _EVAL_294;
  wire  _EVAL_103;
  wire  _EVAL_79;
  wire  _EVAL_201;
  wire  _EVAL_275;
  wire  _EVAL_224;
  wire  _EVAL_243;
  wire  _EVAL_21;
  wire  _EVAL_330;
  wire  _EVAL_51;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_64 = _EVAL_5 == 1'h0;
  assign _EVAL_124 = _EVAL_64 | _EVAL_12;
  assign _EVAL_99 = _EVAL_124 | _EVAL_15;
  assign _EVAL_223 = _EVAL_5 == _EVAL_58;
  assign _EVAL_336 = _EVAL_223 | _EVAL_15;
  assign _EVAL_84 = _EVAL_336 == 1'h0;
  assign _EVAL_139 = _EVAL_10 == 1'h0;
  assign _EVAL_212 = _EVAL_139 | _EVAL_15;
  assign _EVAL_37 = _EVAL_212 == 1'h0;
  assign _EVAL_264 = _EVAL_16 ^ 32'h1800000;
  assign _EVAL_340 = {1'b0,$signed(_EVAL_264)};
  assign _EVAL_106 = _EVAL_292 == 6'h0;
  assign _EVAL_333 = _EVAL_17[2];
  assign _EVAL_40 = _EVAL_333 == 1'h0;
  assign _EVAL_80 = 23'hff << _EVAL_11;
  assign _EVAL_32 = _EVAL_80[7:0];
  assign _EVAL_214 = ~ _EVAL_32;
  assign _EVAL_252 = _EVAL_214[7:2];
  assign _EVAL_192 = _EVAL_292 - 6'h1;
  assign _EVAL_361 = _EVAL_11 == _EVAL_30;
  assign _EVAL_227 = _EVAL_11[0];
  assign _EVAL_182 = 2'h1 << _EVAL_227;
  assign _EVAL_152 = _EVAL_182 | 2'h1;
  assign _EVAL_158 = _EVAL_152[1];
  assign _EVAL_342 = _EVAL_16[1];
  assign _EVAL_153 = _EVAL_342 == 1'h0;
  assign _EVAL_131 = _EVAL_158 & _EVAL_153;
  assign _EVAL_109 = _EVAL_11 >= 4'h2;
  assign _EVAL_358 = _EVAL_109 | _EVAL_131;
  assign _EVAL_102 = _EVAL[5:3];
  assign _EVAL_229 = _EVAL_102 == 3'h0;
  assign _EVAL_324 = _EVAL_17 == 3'h4;
  assign _EVAL_186 = _EVAL_3 & _EVAL_324;
  assign _EVAL_52 = _EVAL_328 != 33'h0;
  assign _EVAL_156 = _EVAL_52 == 1'h0;
  assign _EVAL_85 = plusarg_reader_out == 32'h0;
  assign _EVAL_120 = _EVAL_156 | _EVAL_85;
  assign _EVAL_261 = _EVAL_314 < plusarg_reader_out;
  assign _EVAL_180 = _EVAL_120 | _EVAL_261;
  assign _EVAL_195 = _EVAL_180 | _EVAL_15;
  assign _EVAL_295 = _EVAL_195 == 1'h0;
  assign _EVAL_81 = _EVAL_14 <= 3'h4;
  assign _EVAL_235 = _EVAL_81 | _EVAL_15;
  assign _EVAL_239 = $signed(_EVAL_340) & $signed(-33'sh8000);
  assign _EVAL_344 = $signed(_EVAL_239);
  assign _EVAL_123 = $signed(_EVAL_344) == $signed(33'sh0);
  assign _EVAL_35 = _EVAL_15 == 1'h0;
  assign _EVAL_268 = _EVAL_2 == 2'h0;
  assign _EVAL_155 = _EVAL_268 | _EVAL_15;
  assign _EVAL_283 = _EVAL_17 == 3'h2;
  assign _EVAL_121 = _EVAL_3 & _EVAL_283;
  assign _EVAL_50 = _EVAL_16 ^ 32'hc000000;
  assign _EVAL_110 = {1'b0,$signed(_EVAL_50)};
  assign _EVAL_219 = $signed(_EVAL_110) & $signed(-33'sh4000000);
  assign _EVAL_309 = $signed(_EVAL_219);
  assign _EVAL_202 = _EVAL == _EVAL_147;
  assign _EVAL_140 = _EVAL_202 | _EVAL_15;
  assign _EVAL_28 = 64'h1 << _EVAL_4;
  assign _EVAL_128 = _EVAL_7[0];
  assign _EVAL_220 = 23'hff << _EVAL_1;
  assign _EVAL_111 = _EVAL_220[7:0];
  assign _EVAL_162 = ~ _EVAL_111;
  assign _EVAL_134 = _EVAL_162[7:2];
  assign _EVAL_93 = _EVAL_16 ^ 32'h3000;
  assign _EVAL_172 = {1'b0,$signed(_EVAL_93)};
  assign _EVAL_273 = $signed(_EVAL_172) & $signed(-33'sh1000);
  assign _EVAL_72 = $signed(_EVAL_273);
  assign _EVAL_126 = $signed(_EVAL_72) == $signed(33'sh0);
  assign _EVAL_356 = _EVAL_13 & _EVAL_6;
  assign _EVAL_245 = _EVAL_82 == 6'h0;
  assign _EVAL_320 = _EVAL_82 - 6'h1;
  assign _EVAL_298 = _EVAL_16 ^ 32'h2000000;
  assign _EVAL_203 = {1'b0,$signed(_EVAL_298)};
  assign _EVAL_281 = _EVAL_158 & _EVAL_342;
  assign _EVAL_199 = _EVAL_109 | _EVAL_281;
  assign _EVAL_250 = _EVAL_152[0];
  assign _EVAL_169 = _EVAL_16[0];
  assign _EVAL_200 = _EVAL_342 & _EVAL_169;
  assign _EVAL_346 = _EVAL_250 & _EVAL_200;
  assign _EVAL_94 = _EVAL_199 | _EVAL_346;
  assign _EVAL_308 = _EVAL_169 == 1'h0;
  assign _EVAL_209 = _EVAL_342 & _EVAL_308;
  assign _EVAL_160 = _EVAL_250 & _EVAL_209;
  assign _EVAL_62 = _EVAL_199 | _EVAL_160;
  assign _EVAL_290 = _EVAL_153 & _EVAL_169;
  assign _EVAL_142 = _EVAL_250 & _EVAL_290;
  assign _EVAL_337 = _EVAL_358 | _EVAL_142;
  assign _EVAL_318 = _EVAL_153 & _EVAL_308;
  assign _EVAL_213 = _EVAL_250 & _EVAL_318;
  assign _EVAL_132 = _EVAL_358 | _EVAL_213;
  assign _EVAL_351 = {_EVAL_94,_EVAL_62,_EVAL_337,_EVAL_132};
  assign _EVAL_315 = ~ _EVAL_351;
  assign _EVAL_74 = _EVAL_9 & _EVAL_315;
  assign _EVAL_232 = _EVAL_74 == 4'h0;
  assign _EVAL_312 = _EVAL_232 | _EVAL_15;
  assign _EVAL_260 = _EVAL_312 == 1'h0;
  assign _EVAL_189 = 64'h1 << _EVAL;
  assign _EVAL_159 = _EVAL_7 == 3'h1;
  assign _EVAL_236 = _EVAL_16 ^ 32'h40000000;
  assign _EVAL_77 = {1'b0,$signed(_EVAL_236)};
  assign _EVAL_331 = $signed(_EVAL_77) & $signed(-33'sh2000);
  assign _EVAL_263 = $signed(_EVAL_331);
  assign _EVAL_362 = $signed(_EVAL_263) == $signed(33'sh0);
  assign _EVAL_329 = _EVAL_16 ^ 32'h80000000;
  assign _EVAL_73 = {1'b0,$signed(_EVAL_329)};
  assign _EVAL_248 = $signed(_EVAL_73) & $signed(-33'sh20000);
  assign _EVAL_341 = $signed(_EVAL_248);
  assign _EVAL_231 = $signed(_EVAL_341) == $signed(33'sh0);
  assign _EVAL_246 = _EVAL_362 | _EVAL_231;
  assign _EVAL_364 = $signed(_EVAL_309) == $signed(33'sh0);
  assign _EVAL_164 = _EVAL_246 | _EVAL_364;
  assign _EVAL_143 = $signed(_EVAL_203) & $signed(-33'sh10000);
  assign _EVAL_92 = $signed(_EVAL_143);
  assign _EVAL_319 = $signed(_EVAL_92) == $signed(33'sh0);
  assign _EVAL_345 = _EVAL_164 | _EVAL_319;
  assign _EVAL_230 = _EVAL_361 | _EVAL_15;
  assign _EVAL_146 = _EVAL_140 == 1'h0;
  assign _EVAL_301 = _EVAL == 6'h20;
  assign _EVAL_265 = _EVAL_301 | _EVAL_229;
  assign _EVAL_357 = _EVAL_102 == 3'h1;
  assign _EVAL_27 = _EVAL_265 | _EVAL_357;
  assign _EVAL_338 = _EVAL_102 == 3'h2;
  assign _EVAL_293 = _EVAL_27 | _EVAL_338;
  assign _EVAL_233 = _EVAL_11 <= 4'h8;
  assign _EVAL_136 = _EVAL_1 >= 4'h2;
  assign _EVAL_208 = _EVAL_17 == 3'h3;
  assign _EVAL_326 = _EVAL_3 & _EVAL_208;
  assign _EVAL_332 = _EVAL_8 & _EVAL_3;
  assign _EVAL_138 = _EVAL_4 == _EVAL_363;
  assign _EVAL_45 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_49 = $signed(_EVAL_45) & $signed(-33'sh5000);
  assign _EVAL_278 = $signed(_EVAL_49);
  assign _EVAL_282 = $signed(_EVAL_278) == $signed(33'sh0);
  assign _EVAL_95 = _EVAL_16 ^ 32'h1900000;
  assign _EVAL_280 = {1'b0,$signed(_EVAL_95)};
  assign _EVAL_47 = $signed(_EVAL_280) & $signed(-33'sh2000);
  assign _EVAL_355 = _EVAL_14 == 3'h0;
  assign _EVAL_23 = _EVAL_355 | _EVAL_15;
  assign _EVAL_174 = _EVAL_23 == 1'h0;
  assign _EVAL_104 = _EVAL_64 | _EVAL_15;
  assign _EVAL_198 = _EVAL_332 & _EVAL_106;
  assign _EVAL_48 = _EVAL_198 ? _EVAL_189 : 64'h0;
  assign _EVAL_129 = _EVAL_48[32:0];
  assign _EVAL_55 = _EVAL_22 == 6'h0;
  assign _EVAL_274 = _EVAL_356 & _EVAL_55;
  assign _EVAL_135 = _EVAL_7 == 3'h6;
  assign _EVAL_86 = _EVAL_135 == 1'h0;
  assign _EVAL_352 = _EVAL_274 & _EVAL_86;
  assign _EVAL_237 = _EVAL_352 ? _EVAL_28 : 64'h0;
  assign _EVAL_191 = _EVAL_237[32:0];
  assign _EVAL_272 = _EVAL_129 != _EVAL_191;
  assign _EVAL_316 = _EVAL_129 != 33'h0;
  assign _EVAL_144 = _EVAL_316 == 1'h0;
  assign _EVAL_218 = _EVAL_272 | _EVAL_144;
  assign _EVAL_173 = _EVAL_218 | _EVAL_15;
  assign _EVAL_38 = _EVAL_173 == 1'h0;
  assign _EVAL_216 = _EVAL_17 == _EVAL_105;
  assign _EVAL_127 = _EVAL_216 | _EVAL_15;
  assign _EVAL_339 = _EVAL_17 == 3'h6;
  assign _EVAL_217 = _EVAL_136 | _EVAL_15;
  assign _EVAL_269 = _EVAL_217 == 1'h0;
  assign _EVAL_90 = _EVAL_16 == _EVAL_70;
  assign _EVAL_221 = _EVAL_1 == _EVAL_168;
  assign _EVAL_194 = _EVAL_221 | _EVAL_15;
  assign _EVAL_67 = _EVAL_328 | _EVAL_129;
  assign _EVAL_175 = ~ _EVAL_191;
  assign _EVAL_242 = _EVAL_67 & _EVAL_175;
  assign _EVAL_42 = _EVAL_14 <= 3'h2;
  assign _EVAL_255 = _EVAL_42 | _EVAL_15;
  assign _EVAL_310 = _EVAL_9 == _EVAL_351;
  assign _EVAL_33 = _EVAL_310 | _EVAL_15;
  assign _EVAL_228 = _EVAL_0 == _EVAL_304;
  assign _EVAL_240 = _EVAL_228 | _EVAL_15;
  assign _EVAL_226 = _EVAL_356 & _EVAL_245;
  assign _EVAL_207 = _EVAL_328 >> _EVAL;
  assign _EVAL_97 = _EVAL_207[0];
  assign _EVAL_39 = _EVAL_97 == 1'h0;
  assign _EVAL_353 = _EVAL_6 & _EVAL_159;
  assign _EVAL_88 = _EVAL_11 <= 4'h2;
  assign _EVAL_154 = _EVAL_126 | _EVAL_364;
  assign _EVAL_305 = _EVAL_154 | _EVAL_319;
  assign _EVAL_63 = _EVAL_305 | _EVAL_282;
  assign _EVAL_76 = _EVAL_63 | _EVAL_123;
  assign _EVAL_57 = $signed(_EVAL_47);
  assign _EVAL_277 = $signed(_EVAL_57) == $signed(33'sh0);
  assign _EVAL_150 = _EVAL_76 | _EVAL_277;
  assign _EVAL_279 = _EVAL_16 ^ 32'h20000000;
  assign _EVAL_36 = {1'b0,$signed(_EVAL_279)};
  assign _EVAL_65 = $signed(_EVAL_36) & $signed(-33'sh2000);
  assign _EVAL_322 = $signed(_EVAL_65);
  assign _EVAL_151 = $signed(_EVAL_322) == $signed(33'sh0);
  assign _EVAL_299 = _EVAL_150 | _EVAL_151;
  assign _EVAL_61 = _EVAL_88 & _EVAL_299;
  assign _EVAL_19 = _EVAL_61 | _EVAL_15;
  assign _EVAL_60 = {{24'd0}, _EVAL_214};
  assign _EVAL_53 = _EVAL_17 == 3'h0;
  assign _EVAL_287 = _EVAL_314 + 32'h1;
  assign _EVAL_204 = _EVAL_2 <= 2'h2;
  assign _EVAL_215 = _EVAL_7 == 3'h5;
  assign _EVAL_112 = _EVAL_12 == 1'h0;
  assign _EVAL_188 = _EVAL_112 | _EVAL_15;
  assign _EVAL_161 = _EVAL_4 == 6'h20;
  assign _EVAL_56 = _EVAL_4[5:3];
  assign _EVAL_270 = _EVAL_56 == 3'h0;
  assign _EVAL_113 = _EVAL_161 | _EVAL_270;
  assign _EVAL_26 = _EVAL_56 == 3'h1;
  assign _EVAL_348 = _EVAL_113 | _EVAL_26;
  assign _EVAL_354 = _EVAL_56 == 3'h2;
  assign _EVAL_177 = _EVAL_348 | _EVAL_354;
  assign _EVAL_107 = _EVAL_233 & _EVAL_126;
  assign _EVAL_247 = _EVAL_107 | _EVAL_15;
  assign _EVAL_87 = _EVAL_247 == 1'h0;
  assign _EVAL_285 = _EVAL_347 == 6'h0;
  assign _EVAL_176 = _EVAL_347 - 6'h1;
  assign _EVAL_259 = _EVAL_56 == 3'h3;
  assign _EVAL_78 = _EVAL_177 | _EVAL_259;
  assign _EVAL_108 = _EVAL_78 | _EVAL_15;
  assign _EVAL_313 = _EVAL_108 == 1'h0;
  assign _EVAL_100 = _EVAL_245 == 1'h0;
  assign _EVAL_271 = _EVAL_129 | _EVAL_328;
  assign _EVAL_116 = _EVAL_271 >> _EVAL_4;
  assign _EVAL_118 = _EVAL_116[0];
  assign _EVAL_311 = _EVAL_39 | _EVAL_15;
  assign _EVAL_249 = _EVAL_311 == 1'h0;
  assign _EVAL_251 = _EVAL_7 == 3'h0;
  assign _EVAL_66 = _EVAL_7 <= 3'h6;
  assign _EVAL_266 = _EVAL_66 | _EVAL_15;
  assign _EVAL_149 = _EVAL_102 == 3'h3;
  assign _EVAL_238 = _EVAL_293 | _EVAL_149;
  assign _EVAL_296 = _EVAL_118 | _EVAL_15;
  assign _EVAL_288 = _EVAL_296 == 1'h0;
  assign _EVAL_205 = _EVAL_345 | _EVAL_282;
  assign _EVAL_335 = _EVAL_14 != 3'h0;
  assign _EVAL_222 = _EVAL_335 | _EVAL_15;
  assign _EVAL_257 = _EVAL_222 == 1'h0;
  assign _EVAL_157 = _EVAL_16 & _EVAL_60;
  assign _EVAL_130 = _EVAL_157 == 32'h0;
  assign _EVAL_297 = _EVAL_14 == _EVAL_306;
  assign _EVAL_114 = _EVAL_297 | _EVAL_15;
  assign _EVAL_171 = _EVAL_230 == 1'h0;
  assign _EVAL_234 = _EVAL_2 != 2'h2;
  assign _EVAL_68 = _EVAL_234 | _EVAL_15;
  assign _EVAL_183 = _EVAL_22 - 6'h1;
  assign _EVAL_276 = _EVAL_285 == 1'h0;
  assign _EVAL_34 = _EVAL_109 | _EVAL_15;
  assign _EVAL_343 = _EVAL_104 == 1'h0;
  assign _EVAL_225 = _EVAL_14 <= 3'h3;
  assign _EVAL_125 = _EVAL_225 | _EVAL_15;
  assign _EVAL_211 = _EVAL_204 | _EVAL_15;
  assign _EVAL_44 = _EVAL_235 == 1'h0;
  assign _EVAL_286 = _EVAL_205 | _EVAL_123;
  assign _EVAL_284 = _EVAL_286 | _EVAL_277;
  assign _EVAL_46 = _EVAL_284 | _EVAL_151;
  assign _EVAL_334 = ~ _EVAL_9;
  assign _EVAL_166 = _EVAL_334 == 4'h0;
  assign _EVAL_302 = _EVAL_166 | _EVAL_15;
  assign _EVAL_167 = _EVAL_302 == 1'h0;
  assign _EVAL_291 = _EVAL_155 == 1'h0;
  assign _EVAL_165 = _EVAL_7 == _EVAL_20;
  assign _EVAL_327 = _EVAL_165 | _EVAL_15;
  assign _EVAL_256 = _EVAL_332 & _EVAL_285;
  assign _EVAL_115 = _EVAL_17 == 3'h7;
  assign _EVAL_323 = _EVAL_3 & _EVAL_115;
  assign _EVAL_148 = _EVAL_90 | _EVAL_15;
  assign _EVAL_119 = _EVAL_148 == 1'h0;
  assign _EVAL_190 = _EVAL_6 & _EVAL_251;
  assign _EVAL_184 = _EVAL_255 == 1'h0;
  assign _EVAL_187 = _EVAL_127 == 1'h0;
  assign _EVAL_197 = _EVAL_114 == 1'h0;
  assign _EVAL_179 = _EVAL_99 == 1'h0;
  assign _EVAL_141 = _EVAL_7 == 3'h2;
  assign _EVAL_181 = _EVAL_17 == 3'h5;
  assign _EVAL_71 = _EVAL_6 & _EVAL_215;
  assign _EVAL_262 = _EVAL_7 == 3'h4;
  assign _EVAL_206 = _EVAL_6 & _EVAL_262;
  assign _EVAL_196 = _EVAL_11 <= 4'h6;
  assign _EVAL_31 = _EVAL_196 & _EVAL_231;
  assign _EVAL_185 = _EVAL_31 | _EVAL_15;
  assign _EVAL_24 = _EVAL_2 == _EVAL_349;
  assign _EVAL_25 = _EVAL_24 | _EVAL_15;
  assign _EVAL_137 = _EVAL_185 == 1'h0;
  assign _EVAL_317 = _EVAL_196 & _EVAL_46;
  assign _EVAL_244 = _EVAL_327 == 1'h0;
  assign _EVAL_258 = _EVAL_238 | _EVAL_15;
  assign _EVAL_193 = _EVAL_125 == 1'h0;
  assign _EVAL_122 = _EVAL_211 == 1'h0;
  assign _EVAL_359 = _EVAL_17 == 3'h1;
  assign _EVAL_360 = _EVAL_3 & _EVAL_359;
  assign _EVAL_41 = _EVAL_317 | _EVAL_107;
  assign _EVAL_101 = _EVAL_41 | _EVAL_15;
  assign _EVAL_178 = _EVAL_19 == 1'h0;
  assign _EVAL_54 = _EVAL_332 | _EVAL_356;
  assign _EVAL_29 = _EVAL_3 & _EVAL_339;
  assign _EVAL_145 = _EVAL_130 | _EVAL_15;
  assign _EVAL_98 = _EVAL_145 == 1'h0;
  assign _EVAL_83 = _EVAL_68 == 1'h0;
  assign _EVAL_91 = _EVAL_138 | _EVAL_15;
  assign _EVAL_210 = _EVAL_6 & _EVAL_135;
  assign _EVAL_303 = _EVAL_240 == 1'h0;
  assign _EVAL_163 = _EVAL_25 == 1'h0;
  assign _EVAL_254 = _EVAL_34 == 1'h0;
  assign _EVAL_59 = _EVAL_266 == 1'h0;
  assign _EVAL_75 = _EVAL_3 & _EVAL_53;
  assign _EVAL_294 = _EVAL_33 == 1'h0;
  assign _EVAL_103 = _EVAL_194 == 1'h0;
  assign _EVAL_79 = _EVAL_3 & _EVAL_181;
  assign _EVAL_201 = _EVAL_3 & _EVAL_276;
  assign _EVAL_275 = _EVAL_101 == 1'h0;
  assign _EVAL_224 = _EVAL_6 & _EVAL_141;
  assign _EVAL_243 = _EVAL_188 == 1'h0;
  assign _EVAL_21 = _EVAL_91 == 1'h0;
  assign _EVAL_330 = _EVAL_258 == 1'h0;
  assign _EVAL_51 = _EVAL_6 & _EVAL_100;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_22 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_30 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_58 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_70 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_82 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_105 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_147 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_168 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_292 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_304 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_306 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_314 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _EVAL_328 = _RAND_13[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_347 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_349 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_363 = _RAND_16[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_18) begin
    if (_EVAL_226) begin
      _EVAL_20 <= _EVAL_7;
    end
    if (_EVAL_15) begin
      _EVAL_22 <= 6'h0;
    end else begin
      if (_EVAL_356) begin
        if (_EVAL_55) begin
          if (_EVAL_128) begin
            _EVAL_22 <= _EVAL_134;
          end else begin
            _EVAL_22 <= 6'h0;
          end
        end else begin
          _EVAL_22 <= _EVAL_183;
        end
      end
    end
    if (_EVAL_256) begin
      _EVAL_30 <= _EVAL_11;
    end
    if (_EVAL_226) begin
      _EVAL_58 <= _EVAL_5;
    end
    if (_EVAL_256) begin
      _EVAL_70 <= _EVAL_16;
    end
    if (_EVAL_15) begin
      _EVAL_82 <= 6'h0;
    end else begin
      if (_EVAL_356) begin
        if (_EVAL_245) begin
          if (_EVAL_128) begin
            _EVAL_82 <= _EVAL_134;
          end else begin
            _EVAL_82 <= 6'h0;
          end
        end else begin
          _EVAL_82 <= _EVAL_320;
        end
      end
    end
    if (_EVAL_256) begin
      _EVAL_105 <= _EVAL_17;
    end
    if (_EVAL_256) begin
      _EVAL_147 <= _EVAL;
    end
    if (_EVAL_226) begin
      _EVAL_168 <= _EVAL_1;
    end
    if (_EVAL_15) begin
      _EVAL_292 <= 6'h0;
    end else begin
      if (_EVAL_332) begin
        if (_EVAL_106) begin
          if (_EVAL_40) begin
            _EVAL_292 <= _EVAL_252;
          end else begin
            _EVAL_292 <= 6'h0;
          end
        end else begin
          _EVAL_292 <= _EVAL_192;
        end
      end
    end
    if (_EVAL_226) begin
      _EVAL_304 <= _EVAL_0;
    end
    if (_EVAL_256) begin
      _EVAL_306 <= _EVAL_14;
    end
    if (_EVAL_15) begin
      _EVAL_314 <= 32'h0;
    end else begin
      if (_EVAL_54) begin
        _EVAL_314 <= 32'h0;
      end else begin
        _EVAL_314 <= _EVAL_287;
      end
    end
    if (_EVAL_15) begin
      _EVAL_328 <= 33'h0;
    end else begin
      _EVAL_328 <= _EVAL_242;
    end
    if (_EVAL_15) begin
      _EVAL_347 <= 6'h0;
    end else begin
      if (_EVAL_332) begin
        if (_EVAL_285) begin
          if (_EVAL_40) begin
            _EVAL_347 <= _EVAL_252;
          end else begin
            _EVAL_347 <= 6'h0;
          end
        end else begin
          _EVAL_347 <= _EVAL_176;
        end
      end
    end
    if (_EVAL_226) begin
      _EVAL_349 <= _EVAL_2;
    end
    if (_EVAL_226) begin
      _EVAL_363 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(deba35af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa37e639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(592d5321)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aa1cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1281c01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efd71a5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99fefbbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7546932c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(213f5c51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eff4b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(259765de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(578d37ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2788d1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b454771)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e74ef1dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b6fad07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_343) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bbe079c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(222282be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4930302c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29cc5e41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6de05f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20507d9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6c164a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a11943b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dc41ef1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be3f5c0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43dd6951)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9169cf9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c55f240)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25415047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33289358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1212fc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59a82dc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7a3b083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(526e8bfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13d9e082)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1aff926)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d61a42d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bfbd55d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ef83466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55a52060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec8fd1bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9520e399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9d8e780)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e403c574)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4892bb14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(405f75b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b316a10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1cb985)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9a8a9ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42228d6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(204a3ab6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_343) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9202acea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8525f103)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d322b9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89eb36d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78bb44f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6440e51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41a9310)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42ce6a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1da68d80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90bfcd45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb965243)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abe504eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83e086b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bd300a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5504ada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6433100)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1610e4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afef68fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d9e14d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54691b09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(899cd897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8139a25f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49349079)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a8b9d91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(962188e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4b881e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8bcc70d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59b4894f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c656a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9f986e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88a08f17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75e46542)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91880d65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(922367d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(630842d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7c286e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
