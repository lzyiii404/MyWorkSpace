//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_222(
  output [1:0]  _EVAL,
  input         _EVAL_0,
  output [2:0]  _EVAL_1,
  input  [11:0] _EVAL_2,
  input         _EVAL_3,
  input  [1:0]  _EVAL_4,
  input         _EVAL_5,
  input  [11:0] _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  output [1:0]  _EVAL_10,
  output [31:0] _EVAL_11,
  input         _EVAL_12,
  output [31:0] _EVAL_13,
  output [7:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [1:0]  _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output [31:0] _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  input  [7:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input         _EVAL_34,
  input  [6:0]  _EVAL_35,
  output        _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input  [3:0]  _EVAL_41,
  output [11:0] _EVAL_42,
  output        _EVAL_43
);
  wire  dmOuter__EVAL;
  wire  dmOuter__EVAL_0;
  wire  dmOuter__EVAL_1;
  wire  dmOuter__EVAL_2;
  wire  dmOuter__EVAL_3;
  wire [1:0] dmOuter__EVAL_4;
  wire [31:0] dmOuter__EVAL_5;
  wire [3:0] dmOuter__EVAL_6;
  wire  dmOuter__EVAL_7;
  wire  dmOuter__EVAL_8;
  wire  dmOuter__EVAL_9;
  wire  dmOuter__EVAL_10;
  wire  dmOuter__EVAL_11;
  wire [31:0] dmOuter__EVAL_12;
  wire [31:0] dmOuter__EVAL_13;
  wire [1:0] dmOuter__EVAL_14;
  wire  dmOuter__EVAL_15;
  wire  dmOuter__EVAL_16;
  wire  dmOuter__EVAL_17;
  wire  dmOuter__EVAL_18;
  wire  dmOuter__EVAL_19;
  wire  dmOuter__EVAL_20;
  wire  dmOuter__EVAL_21;
  wire  dmOuter__EVAL_22;
  wire [8:0] dmOuter__EVAL_23;
  wire  dmOuter__EVAL_24;
  wire [2:0] dmOuter__EVAL_25;
  wire  dmOuter__EVAL_26;
  wire [2:0] dmOuter__EVAL_27;
  wire  dmOuter__EVAL_28;
  wire [31:0] dmOuter__EVAL_29;
  wire  dmOuter__EVAL_30;
  wire  dmOuter__EVAL_31;
  wire [1:0] dmOuter__EVAL_32;
  wire  dmOuter__EVAL_33;
  wire  dmOuter__EVAL_34;
  wire  dmOuter__EVAL_35;
  wire  dmOuter__EVAL_36;
  wire  dmOuter__EVAL_37;
  wire [9:0] dmOuter__EVAL_38;
  wire  dmOuter__EVAL_39;
  wire  dmOuter__EVAL_40;
  wire [6:0] dmOuter__EVAL_41;
  wire  dmInner__EVAL;
  wire  dmInner__EVAL_0;
  wire [31:0] dmInner__EVAL_1;
  wire [2:0] dmInner__EVAL_2;
  wire  dmInner__EVAL_3;
  wire [1:0] dmInner__EVAL_4;
  wire  dmInner__EVAL_5;
  wire  dmInner__EVAL_6;
  wire  dmInner__EVAL_7;
  wire [31:0] dmInner__EVAL_8;
  wire [8:0] dmInner__EVAL_9;
  wire  dmInner__EVAL_10;
  wire [3:0] dmInner__EVAL_11;
  wire [3:0] dmInner__EVAL_12;
  wire  dmInner__EVAL_13;
  wire [1:0] dmInner__EVAL_14;
  wire [11:0] dmInner__EVAL_15;
  wire [1:0] dmInner__EVAL_16;
  wire  dmInner__EVAL_17;
  wire [2:0] dmInner__EVAL_18;
  wire  dmInner__EVAL_19;
  wire  dmInner__EVAL_20;
  wire  dmInner__EVAL_21;
  wire  dmInner__EVAL_22;
  wire [31:0] dmInner__EVAL_23;
  wire  dmInner__EVAL_24;
  wire  dmInner__EVAL_25;
  wire [2:0] dmInner__EVAL_26;
  wire [7:0] dmInner__EVAL_27;
  wire  dmInner__EVAL_28;
  wire  dmInner__EVAL_29;
  wire [11:0] dmInner__EVAL_30;
  wire  dmInner__EVAL_31;
  wire  dmInner__EVAL_32;
  wire [2:0] dmInner__EVAL_33;
  wire [31:0] dmInner__EVAL_34;
  wire  dmInner__EVAL_35;
  wire  dmInner__EVAL_36;
  wire  dmInner__EVAL_37;
  wire [11:0] dmInner__EVAL_38;
  wire  dmInner__EVAL_39;
  wire  dmInner__EVAL_40;
  wire  dmInner__EVAL_41;
  wire  dmInner__EVAL_42;
  wire  dmInner__EVAL_43;
  wire  dmInner__EVAL_44;
  wire  dmInner__EVAL_45;
  wire  dmInner__EVAL_46;
  wire [31:0] dmInner__EVAL_47;
  wire  dmInner__EVAL_48;
  wire [2:0] dmInner__EVAL_49;
  wire  dmInner__EVAL_50;
  wire [3:0] dmInner__EVAL_51;
  wire  dmInner__EVAL_52;
  wire [9:0] dmInner__EVAL_53;
  wire  dmInner__EVAL_54;
  wire  dmInner__EVAL_55;
  wire [2:0] dmInner__EVAL_56;
  wire [7:0] dmInner__EVAL_57;
  wire  dmInner__EVAL_58;
  wire  dmInner__EVAL_59;
  SiFive__EVAL_208 dmOuter (
    ._EVAL(dmOuter__EVAL),
    ._EVAL_0(dmOuter__EVAL_0),
    ._EVAL_1(dmOuter__EVAL_1),
    ._EVAL_2(dmOuter__EVAL_2),
    ._EVAL_3(dmOuter__EVAL_3),
    ._EVAL_4(dmOuter__EVAL_4),
    ._EVAL_5(dmOuter__EVAL_5),
    ._EVAL_6(dmOuter__EVAL_6),
    ._EVAL_7(dmOuter__EVAL_7),
    ._EVAL_8(dmOuter__EVAL_8),
    ._EVAL_9(dmOuter__EVAL_9),
    ._EVAL_10(dmOuter__EVAL_10),
    ._EVAL_11(dmOuter__EVAL_11),
    ._EVAL_12(dmOuter__EVAL_12),
    ._EVAL_13(dmOuter__EVAL_13),
    ._EVAL_14(dmOuter__EVAL_14),
    ._EVAL_15(dmOuter__EVAL_15),
    ._EVAL_16(dmOuter__EVAL_16),
    ._EVAL_17(dmOuter__EVAL_17),
    ._EVAL_18(dmOuter__EVAL_18),
    ._EVAL_19(dmOuter__EVAL_19),
    ._EVAL_20(dmOuter__EVAL_20),
    ._EVAL_21(dmOuter__EVAL_21),
    ._EVAL_22(dmOuter__EVAL_22),
    ._EVAL_23(dmOuter__EVAL_23),
    ._EVAL_24(dmOuter__EVAL_24),
    ._EVAL_25(dmOuter__EVAL_25),
    ._EVAL_26(dmOuter__EVAL_26),
    ._EVAL_27(dmOuter__EVAL_27),
    ._EVAL_28(dmOuter__EVAL_28),
    ._EVAL_29(dmOuter__EVAL_29),
    ._EVAL_30(dmOuter__EVAL_30),
    ._EVAL_31(dmOuter__EVAL_31),
    ._EVAL_32(dmOuter__EVAL_32),
    ._EVAL_33(dmOuter__EVAL_33),
    ._EVAL_34(dmOuter__EVAL_34),
    ._EVAL_35(dmOuter__EVAL_35),
    ._EVAL_36(dmOuter__EVAL_36),
    ._EVAL_37(dmOuter__EVAL_37),
    ._EVAL_38(dmOuter__EVAL_38),
    ._EVAL_39(dmOuter__EVAL_39),
    ._EVAL_40(dmOuter__EVAL_40),
    ._EVAL_41(dmOuter__EVAL_41)
  );
  SiFive__EVAL_221 dmInner (
    ._EVAL(dmInner__EVAL),
    ._EVAL_0(dmInner__EVAL_0),
    ._EVAL_1(dmInner__EVAL_1),
    ._EVAL_2(dmInner__EVAL_2),
    ._EVAL_3(dmInner__EVAL_3),
    ._EVAL_4(dmInner__EVAL_4),
    ._EVAL_5(dmInner__EVAL_5),
    ._EVAL_6(dmInner__EVAL_6),
    ._EVAL_7(dmInner__EVAL_7),
    ._EVAL_8(dmInner__EVAL_8),
    ._EVAL_9(dmInner__EVAL_9),
    ._EVAL_10(dmInner__EVAL_10),
    ._EVAL_11(dmInner__EVAL_11),
    ._EVAL_12(dmInner__EVAL_12),
    ._EVAL_13(dmInner__EVAL_13),
    ._EVAL_14(dmInner__EVAL_14),
    ._EVAL_15(dmInner__EVAL_15),
    ._EVAL_16(dmInner__EVAL_16),
    ._EVAL_17(dmInner__EVAL_17),
    ._EVAL_18(dmInner__EVAL_18),
    ._EVAL_19(dmInner__EVAL_19),
    ._EVAL_20(dmInner__EVAL_20),
    ._EVAL_21(dmInner__EVAL_21),
    ._EVAL_22(dmInner__EVAL_22),
    ._EVAL_23(dmInner__EVAL_23),
    ._EVAL_24(dmInner__EVAL_24),
    ._EVAL_25(dmInner__EVAL_25),
    ._EVAL_26(dmInner__EVAL_26),
    ._EVAL_27(dmInner__EVAL_27),
    ._EVAL_28(dmInner__EVAL_28),
    ._EVAL_29(dmInner__EVAL_29),
    ._EVAL_30(dmInner__EVAL_30),
    ._EVAL_31(dmInner__EVAL_31),
    ._EVAL_32(dmInner__EVAL_32),
    ._EVAL_33(dmInner__EVAL_33),
    ._EVAL_34(dmInner__EVAL_34),
    ._EVAL_35(dmInner__EVAL_35),
    ._EVAL_36(dmInner__EVAL_36),
    ._EVAL_37(dmInner__EVAL_37),
    ._EVAL_38(dmInner__EVAL_38),
    ._EVAL_39(dmInner__EVAL_39),
    ._EVAL_40(dmInner__EVAL_40),
    ._EVAL_41(dmInner__EVAL_41),
    ._EVAL_42(dmInner__EVAL_42),
    ._EVAL_43(dmInner__EVAL_43),
    ._EVAL_44(dmInner__EVAL_44),
    ._EVAL_45(dmInner__EVAL_45),
    ._EVAL_46(dmInner__EVAL_46),
    ._EVAL_47(dmInner__EVAL_47),
    ._EVAL_48(dmInner__EVAL_48),
    ._EVAL_49(dmInner__EVAL_49),
    ._EVAL_50(dmInner__EVAL_50),
    ._EVAL_51(dmInner__EVAL_51),
    ._EVAL_52(dmInner__EVAL_52),
    ._EVAL_53(dmInner__EVAL_53),
    ._EVAL_54(dmInner__EVAL_54),
    ._EVAL_55(dmInner__EVAL_55),
    ._EVAL_56(dmInner__EVAL_56),
    ._EVAL_57(dmInner__EVAL_57),
    ._EVAL_58(dmInner__EVAL_58),
    ._EVAL_59(dmInner__EVAL_59)
  );
  assign _EVAL_43 = dmOuter__EVAL_17;
  assign dmInner__EVAL_28 = dmOuter__EVAL_16;
  assign dmInner__EVAL_47 = _EVAL_27;
  assign _EVAL_30 = dmOuter__EVAL_0;
  assign dmInner__EVAL_18 = dmOuter__EVAL_25;
  assign _EVAL_23 = dmInner__EVAL_42;
  assign dmOuter__EVAL_10 = dmInner__EVAL_3;
  assign dmInner__EVAL_48 = dmOuter__EVAL_7;
  assign _EVAL_1 = dmInner__EVAL_2;
  assign dmInner__EVAL_26 = _EVAL_15;
  assign dmOuter__EVAL_35 = dmInner__EVAL_58;
  assign dmOuter__EVAL_12 = dmInner__EVAL_1;
  assign dmInner__EVAL_51 = dmOuter__EVAL_6;
  assign dmInner__EVAL_41 = dmOuter__EVAL_3;
  assign dmInner__EVAL_14 = _EVAL_18;
  assign dmInner__EVAL_55 = dmOuter__EVAL_8;
  assign dmOuter__EVAL_1 = _EVAL_40;
  assign dmOuter__EVAL_19 = dmInner__EVAL_32;
  assign dmInner__EVAL_8 = dmOuter__EVAL_13;
  assign dmInner__EVAL_35 = dmOuter__EVAL_34;
  assign _EVAL_36 = dmOuter__EVAL_40;
  assign _EVAL_14 = dmInner__EVAL_27;
  assign _EVAL_11 = dmInner__EVAL_34;
  assign _EVAL_29 = dmOuter__EVAL_33;
  assign dmInner__EVAL_40 = dmOuter__EVAL_26;
  assign dmInner__EVAL_7 = _EVAL_22;
  assign _EVAL_25 = dmInner__EVAL_23;
  assign dmInner__EVAL_0 = dmOuter__EVAL_21;
  assign dmOuter__EVAL_24 = dmInner__EVAL_52;
  assign _EVAL_13 = dmOuter__EVAL_5;
  assign _EVAL_42 = dmInner__EVAL_38;
  assign dmInner__EVAL_49 = _EVAL_17;
  assign dmOuter__EVAL_27 = dmInner__EVAL_56;
  assign dmInner__EVAL_31 = _EVAL_12;
  assign _EVAL_8 = dmOuter__EVAL_28;
  assign dmInner__EVAL_15 = _EVAL_6;
  assign dmOuter__EVAL_36 = _EVAL_39;
  assign dmInner__EVAL_54 = dmOuter__EVAL_22;
  assign dmOuter__EVAL_39 = dmInner__EVAL_19;
  assign _EVAL_16 = dmInner__EVAL_12;
  assign dmInner__EVAL_39 = _EVAL_19;
  assign dmInner__EVAL_9 = dmOuter__EVAL_23;
  assign dmOuter__EVAL_14 = dmInner__EVAL_4;
  assign dmOuter__EVAL_2 = _EVAL_9;
  assign dmInner__EVAL_30 = _EVAL_2;
  assign dmOuter__EVAL_31 = _EVAL_0;
  assign dmInner__EVAL_57 = _EVAL_32;
  assign _EVAL_10 = dmOuter__EVAL_32;
  assign dmOuter__EVAL_41 = _EVAL_35;
  assign dmOuter__EVAL_29 = _EVAL_33;
  assign dmOuter__EVAL_4 = _EVAL_4;
  assign dmInner__EVAL_5 = _EVAL_5;
  assign dmInner__EVAL_29 = dmOuter__EVAL_37;
  assign dmInner__EVAL_44 = _EVAL_38;
  assign dmOuter__EVAL_11 = dmInner__EVAL_6;
  assign dmInner__EVAL_11 = _EVAL_41;
  assign dmInner__EVAL_17 = _EVAL_20;
  assign dmOuter__EVAL = dmInner__EVAL_43;
  assign _EVAL_26 = dmInner__EVAL_33;
  assign dmInner__EVAL_45 = dmOuter__EVAL_9;
  assign dmInner__EVAL_24 = _EVAL_3;
  assign dmInner__EVAL_46 = _EVAL_31;
  assign dmInner__EVAL_22 = _EVAL_37;
  assign dmInner__EVAL_36 = dmOuter__EVAL_33;
  assign _EVAL_24 = dmInner__EVAL_20;
  assign _EVAL_28 = dmInner__EVAL_25;
  assign dmInner__EVAL_53 = dmOuter__EVAL_38;
  assign dmOuter__EVAL_15 = dmInner__EVAL;
  assign dmOuter__EVAL_20 = dmInner__EVAL_10;
  assign _EVAL_7 = dmInner__EVAL_59;
  assign dmInner__EVAL_37 = _EVAL_34;
  assign dmInner__EVAL_21 = dmOuter__EVAL_18;
  assign _EVAL = dmInner__EVAL_16;
  assign dmInner__EVAL_13 = _EVAL_21;
  assign dmInner__EVAL_50 = dmOuter__EVAL_30;
endmodule
