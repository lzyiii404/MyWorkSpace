//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_223_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [2:0]  _EVAL_10
);
  wire [31:0] plusarg_reader_out;
  reg [4:0] _EVAL_23;
  reg [31:0] _RAND_0;
  reg [4:0] _EVAL_28;
  reg [31:0] _RAND_1;
  reg  _EVAL_61;
  reg [31:0] _RAND_2;
  reg  _EVAL_63;
  reg [31:0] _RAND_3;
  reg [4:0] _EVAL_66;
  reg [31:0] _RAND_4;
  reg [1:0] _EVAL_112;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_139;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_143;
  reg [31:0] _RAND_7;
  reg [31:0] _EVAL_162;
  reg [31:0] _RAND_8;
  reg [4:0] _EVAL_188;
  reg [31:0] _RAND_9;
  reg  _EVAL_196;
  reg [31:0] _RAND_10;
  reg [31:0] _EVAL_198;
  reg [31:0] _RAND_11;
  wire [31:0] _EVAL_59;
  wire [32:0] _EVAL_171;
  wire [31:0] _EVAL_166;
  wire [32:0] _EVAL_35;
  wire [32:0] _EVAL_17;
  wire [32:0] _EVAL_175;
  wire  _EVAL_122;
  wire [31:0] _EVAL_103;
  wire [32:0] _EVAL_121;
  wire  _EVAL_70;
  wire  _EVAL_49;
  wire  _EVAL_68;
  wire [31:0] _EVAL_58;
  wire [32:0] _EVAL_79;
  wire [32:0] _EVAL_53;
  wire [32:0] _EVAL_20;
  wire  _EVAL_117;
  wire [31:0] _EVAL_47;
  wire [32:0] _EVAL_82;
  wire [32:0] _EVAL_144;
  wire [32:0] _EVAL_13;
  wire  _EVAL_132;
  wire  _EVAL_141;
  wire [31:0] _EVAL_111;
  wire [32:0] _EVAL_34;
  wire [32:0] _EVAL_179;
  wire [32:0] _EVAL_83;
  wire  _EVAL_50;
  wire  _EVAL_164;
  wire [32:0] _EVAL_44;
  wire [32:0] _EVAL_95;
  wire  _EVAL_18;
  wire  _EVAL_32;
  wire [32:0] _EVAL_98;
  wire [32:0] _EVAL_152;
  wire [32:0] _EVAL_38;
  wire  _EVAL_26;
  wire  _EVAL_89;
  wire  _EVAL_186;
  wire [31:0] _EVAL_120;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_97;
  wire [32:0] _EVAL_174;
  wire  _EVAL_45;
  wire  _EVAL_48;
  wire [32:0] _EVAL_24;
  wire [32:0] _EVAL_108;
  wire  _EVAL_12;
  wire  _EVAL_114;
  wire [31:0] _EVAL_87;
  wire [32:0] _EVAL_27;
  wire [32:0] _EVAL_194;
  wire [32:0] _EVAL_106;
  wire  _EVAL_40;
  wire  _EVAL_81;
  wire  _EVAL_41;
  wire  _EVAL_19;
  wire  _EVAL_29;
  wire  _EVAL_56;
  wire  _EVAL_39;
  wire  _EVAL_134;
  wire  _EVAL_16;
  wire [1:0] _EVAL_182;
  wire  _EVAL_192;
  wire  _EVAL_124;
  wire  _EVAL_133;
  wire  _EVAL_184;
  wire  _EVAL_52;
  wire  _EVAL_73;
  wire  _EVAL_193;
  wire  _EVAL_21;
  wire [1:0] _EVAL_60;
  wire  _EVAL_33;
  wire  _EVAL_105;
  wire  _EVAL_181;
  wire  _EVAL_37;
  wire  _EVAL_160;
  wire  _EVAL_36;
  wire [31:0] _EVAL_119;
  wire [4:0] _EVAL_90;
  wire  _EVAL_99;
  wire  _EVAL_189;
  wire  _EVAL_187;
  wire [22:0] _EVAL_85;
  wire [7:0] _EVAL_62;
  wire [7:0] _EVAL_135;
  wire [4:0] _EVAL_101;
  wire [4:0] _EVAL_110;
  wire  _EVAL_172;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_195;
  wire  _EVAL_167;
  wire  _EVAL_31;
  wire  _EVAL_127;
  wire  _EVAL_100;
  wire  _EVAL_177;
  wire  _EVAL_155;
  wire  _EVAL_185;
  wire  _EVAL_191;
  wire  _EVAL_128;
  wire  _EVAL_55;
  wire  _EVAL_51;
  wire [31:0] _EVAL_199;
  wire  _EVAL_137;
  wire  _EVAL_69;
  wire  _EVAL_150;
  wire [4:0] _EVAL_92;
  wire  _EVAL_151;
  wire  _EVAL_197;
  wire  _EVAL_94;
  wire  _EVAL_93;
  wire  _EVAL_42;
  wire  _EVAL_78;
  wire  _EVAL_75;
  wire  _EVAL_14;
  wire  _EVAL_30;
  wire  _EVAL_129;
  wire  _EVAL_65;
  wire  _EVAL_168;
  wire  _EVAL_67;
  wire  _EVAL_64;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_22;
  wire  _EVAL_57;
  wire  _EVAL_153;
  wire  _EVAL_107;
  wire  _EVAL_190;
  wire  _EVAL_46;
  wire  _EVAL_54;
  wire  _EVAL_159;
  wire  _EVAL_183;
  wire  _EVAL_102;
  wire [4:0] _EVAL_180;
  wire  _EVAL_178;
  wire  _EVAL_88;
  wire  _EVAL_142;
  wire  _EVAL_76;
  wire  _EVAL_118;
  wire  _EVAL_126;
  wire  _EVAL_96;
  wire  _EVAL_86;
  wire  _EVAL_136;
  wire  _EVAL_138;
  wire  _EVAL_163;
  wire  _EVAL_157;
  wire  _EVAL_109;
  wire  _EVAL_11;
  wire  _EVAL_123;
  wire  _EVAL_77;
  wire  _EVAL_84;
  wire  _EVAL_140;
  wire  _EVAL_15;
  wire  _EVAL_149;
  wire  _EVAL_131;
  wire  _EVAL_115;
  wire  _EVAL_165;
  wire  _EVAL_74;
  wire  _EVAL_104;
  wire  _EVAL_173;
  wire  _EVAL_147;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_59 = _EVAL_8 ^ 32'h20000000;
  assign _EVAL_171 = {1'b0,$signed(_EVAL_59)};
  assign _EVAL_166 = _EVAL_8 ^ 32'h1800000;
  assign _EVAL_35 = {1'b0,$signed(_EVAL_166)};
  assign _EVAL_17 = $signed(_EVAL_35) & $signed(-33'sh8000);
  assign _EVAL_175 = $signed(_EVAL_17);
  assign _EVAL_122 = $signed(_EVAL_175) == $signed(33'sh0);
  assign _EVAL_103 = _EVAL_8 ^ 32'h2000000;
  assign _EVAL_121 = {1'b0,$signed(_EVAL_103)};
  assign _EVAL_70 = _EVAL_7 <= 2'h2;
  assign _EVAL_49 = _EVAL_70 | _EVAL_2;
  assign _EVAL_68 = _EVAL_49 == 1'h0;
  assign _EVAL_58 = _EVAL_8 ^ 32'h40000000;
  assign _EVAL_79 = {1'b0,$signed(_EVAL_58)};
  assign _EVAL_53 = $signed(_EVAL_79) & $signed(-33'sh2000);
  assign _EVAL_20 = $signed(_EVAL_53);
  assign _EVAL_117 = $signed(_EVAL_20) == $signed(33'sh0);
  assign _EVAL_47 = _EVAL_8 ^ 32'h80000000;
  assign _EVAL_82 = {1'b0,$signed(_EVAL_47)};
  assign _EVAL_144 = $signed(_EVAL_82) & $signed(-33'sh20000);
  assign _EVAL_13 = $signed(_EVAL_144);
  assign _EVAL_132 = $signed(_EVAL_13) == $signed(33'sh0);
  assign _EVAL_141 = _EVAL_117 | _EVAL_132;
  assign _EVAL_111 = _EVAL_8 ^ 32'hc000000;
  assign _EVAL_34 = {1'b0,$signed(_EVAL_111)};
  assign _EVAL_179 = $signed(_EVAL_34) & $signed(-33'sh4000000);
  assign _EVAL_83 = $signed(_EVAL_179);
  assign _EVAL_50 = $signed(_EVAL_83) == $signed(33'sh0);
  assign _EVAL_164 = _EVAL_141 | _EVAL_50;
  assign _EVAL_44 = $signed(_EVAL_121) & $signed(-33'sh10000);
  assign _EVAL_95 = $signed(_EVAL_44);
  assign _EVAL_18 = $signed(_EVAL_95) == $signed(33'sh0);
  assign _EVAL_32 = _EVAL_164 | _EVAL_18;
  assign _EVAL_98 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_152 = $signed(_EVAL_98) & $signed(-33'sh5000);
  assign _EVAL_38 = $signed(_EVAL_152);
  assign _EVAL_26 = $signed(_EVAL_38) == $signed(33'sh0);
  assign _EVAL_89 = _EVAL_32 | _EVAL_26;
  assign _EVAL_186 = _EVAL_89 | _EVAL_122;
  assign _EVAL_120 = _EVAL_8 ^ 32'h1900000;
  assign _EVAL_130 = {1'b0,$signed(_EVAL_120)};
  assign _EVAL_97 = $signed(_EVAL_130) & $signed(-33'sh2000);
  assign _EVAL_174 = $signed(_EVAL_97);
  assign _EVAL_45 = $signed(_EVAL_174) == $signed(33'sh0);
  assign _EVAL_48 = _EVAL_186 | _EVAL_45;
  assign _EVAL_24 = $signed(_EVAL_171) & $signed(-33'sh2000);
  assign _EVAL_108 = $signed(_EVAL_24);
  assign _EVAL_12 = $signed(_EVAL_108) == $signed(33'sh0);
  assign _EVAL_114 = _EVAL_48 | _EVAL_12;
  assign _EVAL_87 = _EVAL_8 ^ 32'h3000;
  assign _EVAL_27 = {1'b0,$signed(_EVAL_87)};
  assign _EVAL_194 = $signed(_EVAL_27) & $signed(-33'sh1000);
  assign _EVAL_106 = $signed(_EVAL_194);
  assign _EVAL_40 = $signed(_EVAL_106) == $signed(33'sh0);
  assign _EVAL_81 = _EVAL_114 | _EVAL_40;
  assign _EVAL_41 = _EVAL_81 | _EVAL_2;
  assign _EVAL_19 = _EVAL_41 == 1'h0;
  assign _EVAL_29 = _EVAL_188 == 5'h0;
  assign _EVAL_56 = _EVAL_5 & _EVAL_29;
  assign _EVAL_39 = _EVAL_10 == 3'h6;
  assign _EVAL_134 = _EVAL_39 == 1'h0;
  assign _EVAL_16 = _EVAL_56 & _EVAL_134;
  assign _EVAL_182 = _EVAL_16 ? 2'h1 : 2'h0;
  assign _EVAL_192 = _EVAL_23 == 5'h0;
  assign _EVAL_124 = _EVAL_192 == 1'h0;
  assign _EVAL_133 = _EVAL_7 == 2'h0;
  assign _EVAL_184 = _EVAL_133 | _EVAL_2;
  assign _EVAL_52 = _EVAL_184 == 1'h0;
  assign _EVAL_73 = _EVAL_6 & _EVAL_4;
  assign _EVAL_193 = _EVAL_66 == 5'h0;
  assign _EVAL_21 = _EVAL_73 & _EVAL_193;
  assign _EVAL_60 = _EVAL_21 ? 2'h1 : 2'h0;
  assign _EVAL_33 = _EVAL_60[0];
  assign _EVAL_105 = _EVAL_10[0];
  assign _EVAL_181 = _EVAL_63 == 1'h0;
  assign _EVAL_37 = _EVAL_10 == _EVAL_139;
  assign _EVAL_160 = _EVAL_73 & _EVAL_192;
  assign _EVAL_36 = _EVAL_73 | _EVAL_5;
  assign _EVAL_119 = _EVAL_162 + 32'h1;
  assign _EVAL_90 = _EVAL_23 - 5'h1;
  assign _EVAL_99 = plusarg_reader_out == 32'h0;
  assign _EVAL_189 = _EVAL_181 | _EVAL_99;
  assign _EVAL_187 = _EVAL_28 == 5'h0;
  assign _EVAL_85 = 23'hff << _EVAL_9;
  assign _EVAL_62 = _EVAL_85[7:0];
  assign _EVAL_135 = ~ _EVAL_62;
  assign _EVAL_101 = _EVAL_135[7:3];
  assign _EVAL_110 = _EVAL_28 - 5'h1;
  assign _EVAL_172 = _EVAL_162 < plusarg_reader_out;
  assign _EVAL_145 = _EVAL_189 | _EVAL_172;
  assign _EVAL_146 = _EVAL_8 == _EVAL_198;
  assign _EVAL_195 = _EVAL_146 | _EVAL_2;
  assign _EVAL_167 = _EVAL_195 == 1'h0;
  assign _EVAL_31 = _EVAL_5 & _EVAL_39;
  assign _EVAL_127 = _EVAL_10 == 3'h2;
  assign _EVAL_100 = _EVAL_37 | _EVAL_2;
  assign _EVAL_177 = _EVAL_0 == _EVAL_61;
  assign _EVAL_155 = _EVAL_177 | _EVAL_2;
  assign _EVAL_185 = _EVAL == _EVAL_196;
  assign _EVAL_191 = _EVAL_185 | _EVAL_2;
  assign _EVAL_128 = _EVAL == 1'h0;
  assign _EVAL_55 = _EVAL_128 | _EVAL_1;
  assign _EVAL_51 = _EVAL_10 <= 3'h6;
  assign _EVAL_199 = _EVAL_8 & 32'h3f;
  assign _EVAL_137 = _EVAL_199 == 32'h0;
  assign _EVAL_69 = _EVAL_10 == 3'h4;
  assign _EVAL_150 = _EVAL_182[0];
  assign _EVAL_92 = _EVAL_66 - 5'h1;
  assign _EVAL_151 = ~ _EVAL_150;
  assign _EVAL_197 = _EVAL_187 == 1'h0;
  assign _EVAL_94 = _EVAL_5 & _EVAL_197;
  assign _EVAL_93 = _EVAL_10 == 3'h0;
  assign _EVAL_42 = _EVAL_5 & _EVAL_93;
  assign _EVAL_78 = _EVAL_7 == _EVAL_112;
  assign _EVAL_75 = _EVAL_5 & _EVAL_127;
  assign _EVAL_14 = _EVAL_9 >= 4'h3;
  assign _EVAL_30 = _EVAL_14 | _EVAL_2;
  assign _EVAL_129 = _EVAL_33 | _EVAL_63;
  assign _EVAL_65 = _EVAL_129 | _EVAL_2;
  assign _EVAL_168 = _EVAL_65 == 1'h0;
  assign _EVAL_67 = _EVAL_33 != _EVAL_150;
  assign _EVAL_64 = _EVAL_33 == 1'h0;
  assign _EVAL_71 = _EVAL_67 | _EVAL_64;
  assign _EVAL_72 = _EVAL_71 | _EVAL_2;
  assign _EVAL_22 = _EVAL_72 == 1'h0;
  assign _EVAL_57 = _EVAL_51 | _EVAL_2;
  assign _EVAL_153 = _EVAL_57 == 1'h0;
  assign _EVAL_107 = _EVAL_10 == 3'h1;
  assign _EVAL_190 = _EVAL_10 == 3'h5;
  assign _EVAL_46 = _EVAL_1 == 1'h0;
  assign _EVAL_54 = _EVAL_128 | _EVAL_2;
  assign _EVAL_159 = _EVAL_55 | _EVAL_2;
  assign _EVAL_183 = _EVAL_159 == 1'h0;
  assign _EVAL_102 = _EVAL_63 | _EVAL_33;
  assign _EVAL_180 = _EVAL_188 - 5'h1;
  assign _EVAL_178 = _EVAL_4 & _EVAL_124;
  assign _EVAL_88 = _EVAL_137 | _EVAL_2;
  assign _EVAL_142 = _EVAL_88 == 1'h0;
  assign _EVAL_76 = _EVAL_7 != 2'h2;
  assign _EVAL_118 = _EVAL_5 & _EVAL_107;
  assign _EVAL_126 = _EVAL_46 | _EVAL_2;
  assign _EVAL_96 = _EVAL_126 == 1'h0;
  assign _EVAL_86 = _EVAL_5 & _EVAL_187;
  assign _EVAL_136 = _EVAL_5 & _EVAL_190;
  assign _EVAL_138 = _EVAL_155 == 1'h0;
  assign _EVAL_163 = _EVAL_30 == 1'h0;
  assign _EVAL_157 = _EVAL_54 == 1'h0;
  assign _EVAL_109 = _EVAL_76 | _EVAL_2;
  assign _EVAL_11 = _EVAL_9 == _EVAL_143;
  assign _EVAL_123 = _EVAL_11 | _EVAL_2;
  assign _EVAL_77 = _EVAL_123 == 1'h0;
  assign _EVAL_84 = _EVAL_109 == 1'h0;
  assign _EVAL_140 = _EVAL_145 | _EVAL_2;
  assign _EVAL_15 = _EVAL_140 == 1'h0;
  assign _EVAL_149 = _EVAL_100 == 1'h0;
  assign _EVAL_131 = _EVAL_191 == 1'h0;
  assign _EVAL_115 = _EVAL_181 | _EVAL_2;
  assign _EVAL_165 = _EVAL_78 | _EVAL_2;
  assign _EVAL_74 = _EVAL_5 & _EVAL_69;
  assign _EVAL_104 = _EVAL_102 & _EVAL_151;
  assign _EVAL_173 = _EVAL_115 == 1'h0;
  assign _EVAL_147 = _EVAL_165 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_28 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_61 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_63 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_66 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_112 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_139 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_143 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_162 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_188 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_196 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_198 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_2) begin
      _EVAL_23 <= 5'h0;
    end else begin
      if (_EVAL_73) begin
        if (_EVAL_192) begin
          _EVAL_23 <= 5'h0;
        end else begin
          _EVAL_23 <= _EVAL_90;
        end
      end
    end
    if (_EVAL_2) begin
      _EVAL_28 <= 5'h0;
    end else begin
      if (_EVAL_5) begin
        if (_EVAL_187) begin
          if (_EVAL_105) begin
            _EVAL_28 <= _EVAL_101;
          end else begin
            _EVAL_28 <= 5'h0;
          end
        end else begin
          _EVAL_28 <= _EVAL_110;
        end
      end
    end
    if (_EVAL_86) begin
      _EVAL_61 <= _EVAL_0;
    end
    if (_EVAL_2) begin
      _EVAL_63 <= 1'h0;
    end else begin
      _EVAL_63 <= _EVAL_104;
    end
    if (_EVAL_2) begin
      _EVAL_66 <= 5'h0;
    end else begin
      if (_EVAL_73) begin
        if (_EVAL_193) begin
          _EVAL_66 <= 5'h0;
        end else begin
          _EVAL_66 <= _EVAL_92;
        end
      end
    end
    if (_EVAL_86) begin
      _EVAL_112 <= _EVAL_7;
    end
    if (_EVAL_86) begin
      _EVAL_139 <= _EVAL_10;
    end
    if (_EVAL_86) begin
      _EVAL_143 <= _EVAL_9;
    end
    if (_EVAL_2) begin
      _EVAL_162 <= 32'h0;
    end else begin
      if (_EVAL_36) begin
        _EVAL_162 <= 32'h0;
      end else begin
        _EVAL_162 <= _EVAL_119;
      end
    end
    if (_EVAL_2) begin
      _EVAL_188 <= 5'h0;
    end else begin
      if (_EVAL_5) begin
        if (_EVAL_29) begin
          if (_EVAL_105) begin
            _EVAL_188 <= _EVAL_101;
          end else begin
            _EVAL_188 <= 5'h0;
          end
        end else begin
          _EVAL_188 <= _EVAL_180;
        end
      end
    end
    if (_EVAL_86) begin
      _EVAL_196 <= _EVAL;
    end
    if (_EVAL_160) begin
      _EVAL_198 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cdcfd4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e50e4ac7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4fe31b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7073e7eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(906dc4c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba0d0aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2c2b330)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f6feb84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3613a503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f79f9ae6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c1db80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a45e3b9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5887ef22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d62c994a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f482be3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c26ab32d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816565ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e2ed64b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29788c9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b97fa2d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b55ace6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(465b8e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e249754)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41c5d24b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9f657a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46850ad7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ba3477f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecd92db4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da675380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7072c383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3de39e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
