//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_188_assert(
  input        _EVAL,
  input  [1:0] _EVAL_0,
  input        _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input  [2:0] _EVAL_4,
  input        _EVAL_5,
  input  [8:0] _EVAL_6,
  input        _EVAL_7,
  input  [3:0] _EVAL_8,
  input  [1:0] _EVAL_9,
  input        _EVAL_10,
  input  [2:0] _EVAL_11,
  input        _EVAL_12,
  input        _EVAL_13
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_15;
  reg [31:0] _RAND_0;
  reg  _EVAL_17;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_22;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_26;
  reg [31:0] _RAND_3;
  reg  _EVAL_31;
  reg [31:0] _RAND_4;
  reg  _EVAL_50;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_97;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_109;
  reg [31:0] _RAND_7;
  reg  _EVAL_110;
  reg [31:0] _RAND_8;
  reg [1:0] _EVAL_118;
  reg [31:0] _RAND_9;
  reg  _EVAL_145;
  reg [31:0] _RAND_10;
  reg [8:0] _EVAL_147;
  reg [31:0] _RAND_11;
  reg  _EVAL_155;
  reg [31:0] _RAND_12;
  wire  _EVAL_76;
  wire  _EVAL_170;
  wire  _EVAL_74;
  wire  _EVAL_77;
  wire  _EVAL_116;
  wire  _EVAL_104;
  wire  _EVAL_98;
  wire  _EVAL_100;
  wire  _EVAL_33;
  wire  _EVAL_71;
  wire  _EVAL_49;
  wire [1:0] _EVAL_88;
  wire  _EVAL_60;
  wire  _EVAL_157;
  wire  _EVAL_53;
  wire  _EVAL_126;
  wire  _EVAL_121;
  wire  _EVAL_103;
  wire  _EVAL_108;
  wire  _EVAL_161;
  wire [1:0] _EVAL_81;
  wire  _EVAL_43;
  wire  _EVAL_99;
  wire  _EVAL_89;
  wire [3:0] _EVAL_149;
  wire  _EVAL_144;
  wire  _EVAL_163;
  wire  _EVAL_70;
  wire [8:0] _EVAL_141;
  wire  _EVAL_58;
  wire  _EVAL_32;
  wire  _EVAL_164;
  wire  _EVAL_21;
  wire  _EVAL_111;
  wire  _EVAL_24;
  wire  _EVAL_134;
  wire  _EVAL_36;
  wire  _EVAL_127;
  wire  _EVAL_23;
  wire  _EVAL_72;
  wire  _EVAL_51;
  wire  _EVAL_171;
  wire [9:0] _EVAL_38;
  wire  _EVAL_25;
  wire [9:0] _EVAL_64;
  wire [9:0] _EVAL_45;
  wire  _EVAL_82;
  wire  _EVAL_150;
  wire  _EVAL_29;
  wire  _EVAL_140;
  wire  _EVAL_80;
  wire  _EVAL_27;
  wire  _EVAL_158;
  wire  _EVAL_57;
  wire  _EVAL_79;
  wire [31:0] _EVAL_59;
  wire  _EVAL_151;
  wire  _EVAL_135;
  wire  _EVAL_34;
  wire  _EVAL_172;
  wire  _EVAL_18;
  wire  _EVAL_146;
  wire  _EVAL_148;
  wire  _EVAL_19;
  wire  _EVAL_55;
  wire  _EVAL_166;
  wire  _EVAL_132;
  wire  _EVAL_159;
  wire  _EVAL_67;
  wire  _EVAL_133;
  wire  _EVAL_125;
  wire  _EVAL_56;
  wire  _EVAL_115;
  wire  _EVAL_69;
  wire  _EVAL_68;
  wire  _EVAL_83;
  wire  _EVAL_105;
  wire  _EVAL_42;
  wire  _EVAL_46;
  wire  _EVAL_40;
  wire  _EVAL_66;
  wire  _EVAL_47;
  wire  _EVAL_61;
  wire  _EVAL_131;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_107;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_124;
  wire  _EVAL_52;
  wire  _EVAL_63;
  wire  _EVAL_54;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_165;
  wire  _EVAL_44;
  wire  _EVAL_35;
  wire  _EVAL_102;
  wire  _EVAL_41;
  wire  _EVAL_14;
  wire  _EVAL_37;
  wire  _EVAL_73;
  wire  _EVAL_87;
  wire  _EVAL_48;
  wire  _EVAL_122;
  wire  _EVAL_113;
  wire  _EVAL_95;
  wire  _EVAL_106;
  wire  _EVAL_28;
  wire  _EVAL_94;
  wire  _EVAL_75;
  wire  _EVAL_39;
  wire  _EVAL_78;
  wire  _EVAL_117;
  wire  _EVAL_112;
  wire  _EVAL_156;
  wire  _EVAL_169;
  wire  _EVAL_168;
  wire  _EVAL_91;
  wire  _EVAL_160;
  wire  _EVAL_65;
  wire  _EVAL_96;
  wire  _EVAL_92;
  wire  _EVAL_120;
  wire  _EVAL_62;
  wire  _EVAL_130;
  wire  _EVAL_128;
  wire  _EVAL_90;
  wire  _EVAL_152;
  wire  _EVAL_30;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_76 = _EVAL == 1'h0;
  assign _EVAL_170 = _EVAL_76 | _EVAL_1;
  assign _EVAL_74 = _EVAL_170 == 1'h0;
  assign _EVAL_77 = _EVAL_12 & _EVAL_5;
  assign _EVAL_116 = _EVAL_15 == 1'h0;
  assign _EVAL_104 = _EVAL_77 & _EVAL_116;
  assign _EVAL_98 = _EVAL_155 - 1'h1;
  assign _EVAL_100 = _EVAL_4 <= 3'h6;
  assign _EVAL_33 = _EVAL_100 | _EVAL_1;
  assign _EVAL_71 = _EVAL_31 == 1'h0;
  assign _EVAL_49 = _EVAL_77 & _EVAL_71;
  assign _EVAL_88 = _EVAL_49 ? 2'h1 : 2'h0;
  assign _EVAL_60 = _EVAL_88[0];
  assign _EVAL_157 = _EVAL_50 | _EVAL_60;
  assign _EVAL_53 = _EVAL_2 & _EVAL_7;
  assign _EVAL_126 = _EVAL_145 == 1'h0;
  assign _EVAL_121 = _EVAL_53 & _EVAL_126;
  assign _EVAL_103 = _EVAL_4 == 3'h6;
  assign _EVAL_108 = _EVAL_103 == 1'h0;
  assign _EVAL_161 = _EVAL_121 & _EVAL_108;
  assign _EVAL_81 = _EVAL_161 ? 2'h1 : 2'h0;
  assign _EVAL_43 = _EVAL_81[0];
  assign _EVAL_99 = ~ _EVAL_43;
  assign _EVAL_89 = _EVAL_157 & _EVAL_99;
  assign _EVAL_149 = ~ _EVAL_8;
  assign _EVAL_144 = _EVAL_149 == 4'h0;
  assign _EVAL_163 = _EVAL_144 | _EVAL_1;
  assign _EVAL_70 = _EVAL_163 == 1'h0;
  assign _EVAL_141 = _EVAL_6 & 9'h3;
  assign _EVAL_58 = _EVAL_9 != 2'h2;
  assign _EVAL_32 = _EVAL_7 & _EVAL_103;
  assign _EVAL_164 = _EVAL_9 == 2'h0;
  assign _EVAL_21 = _EVAL_164 | _EVAL_1;
  assign _EVAL_111 = _EVAL_60 | _EVAL_50;
  assign _EVAL_24 = _EVAL_11 == 3'h5;
  assign _EVAL_134 = _EVAL_145 - 1'h1;
  assign _EVAL_36 = _EVAL_155 == 1'h0;
  assign _EVAL_127 = _EVAL_36 == 1'h0;
  assign _EVAL_23 = _EVAL_7 & _EVAL_127;
  assign _EVAL_72 = _EVAL_6 == _EVAL_147;
  assign _EVAL_51 = _EVAL_72 | _EVAL_1;
  assign _EVAL_171 = _EVAL_1 == 1'h0;
  assign _EVAL_38 = {1'b0,$signed(_EVAL_6)};
  assign _EVAL_25 = _EVAL_4 == _EVAL_22;
  assign _EVAL_64 = $signed(_EVAL_38) & $signed(-10'sh200);
  assign _EVAL_45 = $signed(_EVAL_64);
  assign _EVAL_82 = $signed(_EVAL_45) == $signed(10'sh0);
  assign _EVAL_150 = _EVAL_82 | _EVAL_1;
  assign _EVAL_29 = _EVAL_150 == 1'h0;
  assign _EVAL_140 = _EVAL_8 == 4'hf;
  assign _EVAL_80 = _EVAL_9 == _EVAL_26;
  assign _EVAL_27 = _EVAL_80 | _EVAL_1;
  assign _EVAL_158 = _EVAL_11 == _EVAL_97;
  assign _EVAL_57 = _EVAL_158 | _EVAL_1;
  assign _EVAL_79 = _EVAL_57 == 1'h0;
  assign _EVAL_59 = _EVAL_109 + 32'h1;
  assign _EVAL_151 = _EVAL_4 == 3'h2;
  assign _EVAL_135 = _EVAL_7 & _EVAL_151;
  assign _EVAL_34 = _EVAL_31 - 1'h1;
  assign _EVAL_172 = _EVAL_9 <= 2'h2;
  assign _EVAL_18 = _EVAL_172 | _EVAL_1;
  assign _EVAL_146 = _EVAL_18 == 1'h0;
  assign _EVAL_148 = _EVAL_116 == 1'h0;
  assign _EVAL_19 = _EVAL_5 & _EVAL_148;
  assign _EVAL_55 = _EVAL_27 == 1'h0;
  assign _EVAL_166 = _EVAL_58 | _EVAL_1;
  assign _EVAL_132 = _EVAL_166 == 1'h0;
  assign _EVAL_159 = _EVAL_76 | _EVAL_3;
  assign _EVAL_67 = _EVAL_159 | _EVAL_1;
  assign _EVAL_133 = _EVAL_67 == 1'h0;
  assign _EVAL_125 = _EVAL_50 == 1'h0;
  assign _EVAL_56 = _EVAL_125 | _EVAL_1;
  assign _EVAL_115 = _EVAL_56 == 1'h0;
  assign _EVAL_69 = _EVAL_4 == 3'h0;
  assign _EVAL_68 = _EVAL_7 & _EVAL_69;
  assign _EVAL_83 = _EVAL_111 | _EVAL_1;
  assign _EVAL_105 = _EVAL_140 | _EVAL_1;
  assign _EVAL_42 = _EVAL_13 == _EVAL_110;
  assign _EVAL_46 = _EVAL_42 | _EVAL_1;
  assign _EVAL_40 = _EVAL_46 == 1'h0;
  assign _EVAL_66 = _EVAL_25 | _EVAL_1;
  assign _EVAL_47 = _EVAL_66 == 1'h0;
  assign _EVAL_61 = _EVAL_5 & _EVAL_24;
  assign _EVAL_131 = _EVAL_11 == 3'h6;
  assign _EVAL_138 = _EVAL_4 == 3'h1;
  assign _EVAL_139 = _EVAL_0 == _EVAL_118;
  assign _EVAL_107 = _EVAL_139 | _EVAL_1;
  assign _EVAL_84 = _EVAL_107 == 1'h0;
  assign _EVAL_85 = _EVAL_4 == 3'h4;
  assign _EVAL_86 = _EVAL_11 == 3'h0;
  assign _EVAL_124 = _EVAL_5 & _EVAL_86;
  assign _EVAL_52 = _EVAL_11 == 3'h7;
  assign _EVAL_63 = _EVAL_5 & _EVAL_52;
  assign _EVAL_54 = _EVAL_53 & _EVAL_36;
  assign _EVAL_153 = _EVAL_83 == 1'h0;
  assign _EVAL_154 = _EVAL_11 == 3'h4;
  assign _EVAL_165 = _EVAL_5 & _EVAL_154;
  assign _EVAL_44 = plusarg_reader_out == 32'h0;
  assign _EVAL_35 = _EVAL_125 | _EVAL_44;
  assign _EVAL_102 = _EVAL_109 < plusarg_reader_out;
  assign _EVAL_41 = _EVAL_35 | _EVAL_102;
  assign _EVAL_14 = _EVAL_41 | _EVAL_1;
  assign _EVAL_37 = _EVAL_3 == 1'h0;
  assign _EVAL_73 = _EVAL_37 | _EVAL_1;
  assign _EVAL_87 = _EVAL_73 == 1'h0;
  assign _EVAL_48 = _EVAL == _EVAL_17;
  assign _EVAL_122 = _EVAL_48 | _EVAL_1;
  assign _EVAL_113 = _EVAL_51 == 1'h0;
  assign _EVAL_95 = _EVAL_21 == 1'h0;
  assign _EVAL_106 = _EVAL_11 == 3'h2;
  assign _EVAL_28 = _EVAL_5 & _EVAL_106;
  assign _EVAL_94 = _EVAL_141 == 9'h0;
  assign _EVAL_75 = _EVAL_4 == 3'h5;
  assign _EVAL_39 = _EVAL_11 == 3'h1;
  assign _EVAL_78 = _EVAL_15 - 1'h1;
  assign _EVAL_117 = _EVAL_5 & _EVAL_131;
  assign _EVAL_112 = _EVAL_77 | _EVAL_53;
  assign _EVAL_156 = _EVAL_7 & _EVAL_138;
  assign _EVAL_169 = _EVAL_7 & _EVAL_85;
  assign _EVAL_168 = _EVAL_122 == 1'h0;
  assign _EVAL_91 = _EVAL_0 >= 2'h2;
  assign _EVAL_160 = _EVAL_91 | _EVAL_1;
  assign _EVAL_65 = _EVAL_160 == 1'h0;
  assign _EVAL_96 = _EVAL_33 == 1'h0;
  assign _EVAL_92 = _EVAL_5 & _EVAL_39;
  assign _EVAL_120 = _EVAL_105 == 1'h0;
  assign _EVAL_62 = _EVAL_11 == 3'h3;
  assign _EVAL_130 = _EVAL_5 & _EVAL_62;
  assign _EVAL_128 = _EVAL_14 == 1'h0;
  assign _EVAL_90 = _EVAL_94 | _EVAL_1;
  assign _EVAL_152 = _EVAL_7 & _EVAL_75;
  assign _EVAL_30 = _EVAL_90 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_17 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_22 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_26 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_50 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_97 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_109 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_110 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_118 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_145 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_147 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_155 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_10) begin
    if (_EVAL_1) begin
      _EVAL_15 <= 1'h0;
    end else begin
      if (_EVAL_77) begin
        if (_EVAL_116) begin
          _EVAL_15 <= 1'h0;
        end else begin
          _EVAL_15 <= _EVAL_78;
        end
      end
    end
    if (_EVAL_54) begin
      _EVAL_17 <= _EVAL;
    end
    if (_EVAL_54) begin
      _EVAL_22 <= _EVAL_4;
    end
    if (_EVAL_54) begin
      _EVAL_26 <= _EVAL_9;
    end
    if (_EVAL_1) begin
      _EVAL_31 <= 1'h0;
    end else begin
      if (_EVAL_77) begin
        if (_EVAL_71) begin
          _EVAL_31 <= 1'h0;
        end else begin
          _EVAL_31 <= _EVAL_34;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_50 <= 1'h0;
    end else begin
      _EVAL_50 <= _EVAL_89;
    end
    if (_EVAL_104) begin
      _EVAL_97 <= _EVAL_11;
    end
    if (_EVAL_1) begin
      _EVAL_109 <= 32'h0;
    end else begin
      if (_EVAL_112) begin
        _EVAL_109 <= 32'h0;
      end else begin
        _EVAL_109 <= _EVAL_59;
      end
    end
    if (_EVAL_54) begin
      _EVAL_110 <= _EVAL_13;
    end
    if (_EVAL_54) begin
      _EVAL_118 <= _EVAL_0;
    end
    if (_EVAL_1) begin
      _EVAL_145 <= 1'h0;
    end else begin
      if (_EVAL_53) begin
        if (_EVAL_126) begin
          _EVAL_145 <= 1'h0;
        end else begin
          _EVAL_145 <= _EVAL_134;
        end
      end
    end
    if (_EVAL_104) begin
      _EVAL_147 <= _EVAL_6;
    end
    if (_EVAL_1) begin
      _EVAL_155 <= 1'h0;
    end else begin
      if (_EVAL_53) begin
        if (_EVAL_36) begin
          _EVAL_155 <= 1'h0;
        end else begin
          _EVAL_155 <= _EVAL_98;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22454922)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(475e1b88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30567319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49efc219)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51c60b41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d42e0e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d148629f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a994b26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1380d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ccd65d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b36aa0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(535489e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2b947dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(766117a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd0ca711)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(145f7aea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e8341af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d00735)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a108a0c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2e8359b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd30f76a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9eda2e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84e258fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0bdf165)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb55cd58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac6ba691)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e783499c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab262b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(878f95d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15110901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84b29069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2ab1bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a189a10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(759503f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff7f7f58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b970e1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b30b6a45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed0e83f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69038b1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(780daca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1eaae19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c981d62d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23ab40f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de03659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(250b6d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5e0b8ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b75ccb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45e6341f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22f0326c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66705792)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbdffccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98b35050)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa9686f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66cd0d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a94a0185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e122a93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ebe8462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d14d8464)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67f9d9a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cfa3340)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ba8f6af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e97e6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
