//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_159_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [6:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [6:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [29:0] _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_26;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_53;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_60;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_75;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_94;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_96;
  reg [31:0] _RAND_5;
  reg [29:0] _EVAL_101;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_112;
  reg [31:0] _RAND_7;
  reg [6:0] _EVAL_116;
  reg [31:0] _RAND_8;
  reg  _EVAL_147;
  reg [31:0] _RAND_9;
  reg [31:0] _EVAL_159;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_163;
  reg [31:0] _RAND_11;
  reg [6:0] _EVAL_168;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_261;
  reg [31:0] _RAND_13;
  reg [72:0] _EVAL_295;
  reg [95:0] _RAND_14;
  wire  _EVAL_285;
  wire  _EVAL_174;
  wire  _EVAL_258;
  wire  _EVAL_134;
  wire [1:0] _EVAL_148;
  wire [1:0] _EVAL_142;
  wire  _EVAL_92;
  wire  _EVAL_291;
  wire  _EVAL_47;
  wire  _EVAL_160;
  wire  _EVAL_32;
  wire  _EVAL_263;
  wire  _EVAL_266;
  wire  _EVAL_193;
  wire  _EVAL_69;
  wire  _EVAL_108;
  wire  _EVAL_278;
  wire  _EVAL_74;
  wire  _EVAL_244;
  wire  _EVAL_103;
  wire  _EVAL_282;
  wire  _EVAL_98;
  wire  _EVAL_149;
  wire  _EVAL_83;
  wire  _EVAL_138;
  wire  _EVAL_250;
  wire  _EVAL_186;
  wire  _EVAL_238;
  wire  _EVAL_245;
  wire  _EVAL_162;
  wire  _EVAL_280;
  wire  _EVAL_216;
  wire  _EVAL_218;
  wire  _EVAL_80;
  wire  _EVAL_50;
  wire  _EVAL_264;
  wire  _EVAL_156;
  wire  _EVAL_68;
  wire  _EVAL_145;
  wire  _EVAL_279;
  wire  _EVAL_166;
  wire  _EVAL_213;
  wire  _EVAL_120;
  wire [3:0] _EVAL_234;
  wire  _EVAL_196;
  wire  _EVAL_136;
  wire  _EVAL_58;
  wire  _EVAL_27;
  wire  _EVAL_281;
  wire  _EVAL_204;
  wire  _EVAL_104;
  wire  _EVAL_229;
  wire  _EVAL_184;
  wire  _EVAL_65;
  wire  _EVAL_203;
  wire [127:0] _EVAL_144;
  wire [127:0] _EVAL_257;
  wire [72:0] _EVAL_81;
  wire [72:0] _EVAL_301;
  wire  _EVAL_33;
  wire  _EVAL_167;
  wire  _EVAL_151;
  wire [127:0] _EVAL_165;
  wire [127:0] _EVAL_241;
  wire [72:0] _EVAL_208;
  wire [72:0] _EVAL_293;
  wire [72:0] _EVAL_220;
  wire  _EVAL_265;
  wire  _EVAL_130;
  wire [29:0] _EVAL_290;
  wire [30:0] _EVAL_84;
  wire [30:0] _EVAL_70;
  wire [30:0] _EVAL_109;
  wire  _EVAL_243;
  wire [3:0] _EVAL_198;
  wire  _EVAL_106;
  wire  _EVAL_18;
  wire  _EVAL_253;
  wire [12:0] _EVAL_199;
  wire [5:0] _EVAL_276;
  wire [5:0] _EVAL_226;
  wire [3:0] _EVAL_77;
  wire  _EVAL_248;
  wire [3:0] _EVAL_128;
  wire [3:0] _EVAL_217;
  wire  _EVAL_158;
  wire  _EVAL_71;
  wire  _EVAL_105;
  wire  _EVAL_172;
  wire  _EVAL_209;
  wire  _EVAL_121;
  wire  _EVAL_197;
  wire  _EVAL_122;
  wire  _EVAL_54;
  wire  _EVAL_17;
  wire  _EVAL_179;
  wire [2:0] _EVAL_230;
  wire  _EVAL_55;
  wire  _EVAL_195;
  wire  _EVAL_61;
  wire  _EVAL_274;
  wire  _EVAL_46;
  wire  _EVAL_177;
  wire  _EVAL_155;
  wire  _EVAL_249;
  wire  _EVAL_247;
  wire  _EVAL_189;
  wire  _EVAL_173;
  wire  _EVAL_185;
  wire  _EVAL_119;
  wire  _EVAL_237;
  wire  _EVAL_303;
  wire [3:0] _EVAL_111;
  wire [3:0] _EVAL_153;
  wire  _EVAL_262;
  wire  _EVAL_251;
  wire  _EVAL_182;
  wire  _EVAL_117;
  wire  _EVAL_200;
  wire  _EVAL_43;
  wire  _EVAL_202;
  wire  _EVAL_49;
  wire  _EVAL_20;
  wire  _EVAL_272;
  wire  _EVAL_52;
  wire  _EVAL_224;
  wire  _EVAL_223;
  wire  _EVAL_59;
  wire  _EVAL_79;
  wire  _EVAL_87;
  wire  _EVAL_154;
  wire [31:0] _EVAL_273;
  wire  _EVAL_164;
  wire  _EVAL_275;
  wire  _EVAL_294;
  wire  _EVAL_161;
  wire [3:0] _EVAL_125;
  wire  _EVAL_236;
  wire [2:0] _EVAL_35;
  wire  _EVAL_45;
  wire  _EVAL_110;
  wire  _EVAL_57;
  wire  _EVAL_206;
  wire  _EVAL_221;
  wire  _EVAL_132;
  wire  _EVAL_211;
  wire  _EVAL_194;
  wire  _EVAL_242;
  wire  _EVAL_268;
  wire  _EVAL_288;
  wire  _EVAL_91;
  wire  _EVAL_231;
  wire  _EVAL_292;
  wire  _EVAL_300;
  wire  _EVAL_42;
  wire  _EVAL_175;
  wire  _EVAL_40;
  wire  _EVAL_180;
  wire [3:0] _EVAL_270;
  wire  _EVAL_118;
  wire [12:0] _EVAL_170;
  wire [5:0] _EVAL_95;
  wire [5:0] _EVAL_107;
  wire [3:0] _EVAL_259;
  wire  _EVAL_48;
  wire  _EVAL_232;
  wire  _EVAL_219;
  wire  _EVAL_254;
  wire  _EVAL_24;
  wire [3:0] _EVAL_124;
  wire [29:0] _EVAL_214;
  wire [72:0] _EVAL_135;
  wire  _EVAL_192;
  wire  _EVAL_85;
  wire  _EVAL_140;
  wire  _EVAL_212;
  wire  _EVAL_289;
  wire  _EVAL_62;
  wire  _EVAL_28;
  wire  _EVAL_99;
  wire  _EVAL_246;
  wire  _EVAL_56;
  wire  _EVAL_127;
  wire  _EVAL_255;
  wire  _EVAL_283;
  wire  _EVAL_21;
  wire  _EVAL_64;
  wire  _EVAL_210;
  wire  _EVAL_114;
  wire  _EVAL_25;
  wire  _EVAL_123;
  wire  _EVAL_67;
  wire  _EVAL_181;
  wire  _EVAL_183;
  wire  _EVAL_228;
  wire  _EVAL_171;
  wire  _EVAL_73;
  wire  _EVAL_201;
  wire  _EVAL_222;
  wire  _EVAL_34;
  wire  _EVAL_30;
  wire  _EVAL_299;
  wire  _EVAL_29;
  wire  _EVAL_240;
  wire  _EVAL_302;
  wire  _EVAL_252;
  wire  _EVAL_137;
  wire  _EVAL_89;
  wire [3:0] _EVAL_37;
  wire  _EVAL_41;
  wire  _EVAL_100;
  wire  _EVAL_139;
  wire  _EVAL_267;
  wire  _EVAL_178;
  wire  _EVAL_19;
  wire  _EVAL_115;
  wire  _EVAL_39;
  wire  _EVAL_287;
  wire  _EVAL_22;
  wire  _EVAL_169;
  wire  _EVAL_76;
  wire [29:0] _EVAL_235;
  wire  _EVAL_97;
  wire  _EVAL_126;
  wire  _EVAL_215;
  wire  _EVAL_143;
  wire [72:0] _EVAL_298;
  wire [72:0] _EVAL_82;
  wire  _EVAL_188;
  wire  _EVAL_78;
  wire  _EVAL_271;
  wire  _EVAL_191;
  wire  _EVAL_205;
  wire  _EVAL_131;
  wire  _EVAL_260;
  wire  _EVAL_157;
  wire  _EVAL_225;
  wire  _EVAL_297;
  wire  _EVAL_90;
  wire  _EVAL_129;
  wire  _EVAL_88;
  wire  _EVAL_187;
  wire  _EVAL_152;
  wire  _EVAL_146;
  wire  _EVAL_284;
  wire  _EVAL_66;
  wire  _EVAL_93;
  wire  _EVAL_141;
  wire  _EVAL_239;
  wire  _EVAL_207;
  wire  _EVAL_286;
  wire  _EVAL_113;
  wire  _EVAL_190;
  wire  _EVAL_296;
  wire  _EVAL_38;
  wire  _EVAL_51;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_285 = _EVAL_295 != 73'h0;
  assign _EVAL_174 = _EVAL_13 <= 3'h4;
  assign _EVAL_258 = _EVAL_1 >= 3'h2;
  assign _EVAL_134 = _EVAL_1[0];
  assign _EVAL_148 = 2'h1 << _EVAL_134;
  assign _EVAL_142 = _EVAL_148 | 2'h1;
  assign _EVAL_92 = _EVAL_142[1];
  assign _EVAL_291 = _EVAL_11[1];
  assign _EVAL_47 = _EVAL_291 == 1'h0;
  assign _EVAL_160 = _EVAL_92 & _EVAL_47;
  assign _EVAL_32 = _EVAL_258 | _EVAL_160;
  assign _EVAL_263 = _EVAL_142[0];
  assign _EVAL_266 = _EVAL_11[0];
  assign _EVAL_193 = _EVAL_266 == 1'h0;
  assign _EVAL_69 = _EVAL_47 & _EVAL_193;
  assign _EVAL_108 = _EVAL_263 & _EVAL_69;
  assign _EVAL_278 = _EVAL_32 | _EVAL_108;
  assign _EVAL_74 = _EVAL_13 <= 3'h3;
  assign _EVAL_244 = _EVAL_74 | _EVAL_6;
  assign _EVAL_103 = _EVAL_0 == _EVAL_147;
  assign _EVAL_282 = _EVAL_75 == 4'h0;
  assign _EVAL_98 = _EVAL_282 == 1'h0;
  assign _EVAL_149 = _EVAL_285 == 1'h0;
  assign _EVAL_83 = plusarg_reader_out == 32'h0;
  assign _EVAL_138 = _EVAL_149 | _EVAL_83;
  assign _EVAL_250 = _EVAL_159 < plusarg_reader_out;
  assign _EVAL_186 = _EVAL_138 | _EVAL_250;
  assign _EVAL_238 = _EVAL_186 | _EVAL_6;
  assign _EVAL_245 = _EVAL_238 == 1'h0;
  assign _EVAL_162 = _EVAL_0 == 1'h0;
  assign _EVAL_280 = _EVAL_162 | _EVAL_6;
  assign _EVAL_216 = _EVAL_280 == 1'h0;
  assign _EVAL_218 = _EVAL_92 & _EVAL_291;
  assign _EVAL_80 = _EVAL_258 | _EVAL_218;
  assign _EVAL_50 = _EVAL_291 & _EVAL_266;
  assign _EVAL_264 = _EVAL_263 & _EVAL_50;
  assign _EVAL_156 = _EVAL_80 | _EVAL_264;
  assign _EVAL_68 = _EVAL_291 & _EVAL_193;
  assign _EVAL_145 = _EVAL_263 & _EVAL_68;
  assign _EVAL_279 = _EVAL_80 | _EVAL_145;
  assign _EVAL_166 = _EVAL_47 & _EVAL_266;
  assign _EVAL_213 = _EVAL_263 & _EVAL_166;
  assign _EVAL_120 = _EVAL_32 | _EVAL_213;
  assign _EVAL_234 = {_EVAL_156,_EVAL_279,_EVAL_120,_EVAL_278};
  assign _EVAL_196 = _EVAL_8 == _EVAL_234;
  assign _EVAL_136 = _EVAL_196 | _EVAL_6;
  assign _EVAL_58 = _EVAL_136 == 1'h0;
  assign _EVAL_27 = _EVAL_7 & _EVAL_16;
  assign _EVAL_281 = _EVAL_112 == 4'h0;
  assign _EVAL_204 = _EVAL_27 & _EVAL_281;
  assign _EVAL_104 = _EVAL_10 == 3'h1;
  assign _EVAL_229 = _EVAL & _EVAL_104;
  assign _EVAL_184 = _EVAL_12 & _EVAL;
  assign _EVAL_65 = _EVAL_163 == 4'h0;
  assign _EVAL_203 = _EVAL_184 & _EVAL_65;
  assign _EVAL_144 = 128'h1 << _EVAL_4;
  assign _EVAL_257 = _EVAL_203 ? _EVAL_144 : 128'h0;
  assign _EVAL_81 = _EVAL_257[72:0];
  assign _EVAL_301 = _EVAL_295 | _EVAL_81;
  assign _EVAL_33 = _EVAL_14 == 3'h6;
  assign _EVAL_167 = _EVAL_33 == 1'h0;
  assign _EVAL_151 = _EVAL_204 & _EVAL_167;
  assign _EVAL_165 = 128'h1 << _EVAL_9;
  assign _EVAL_241 = _EVAL_151 ? _EVAL_165 : 128'h0;
  assign _EVAL_208 = _EVAL_241[72:0];
  assign _EVAL_293 = ~ _EVAL_208;
  assign _EVAL_220 = _EVAL_301 & _EVAL_293;
  assign _EVAL_265 = _EVAL_14 == 3'h5;
  assign _EVAL_130 = _EVAL_16 & _EVAL_265;
  assign _EVAL_290 = _EVAL_11 ^ 30'h20000000;
  assign _EVAL_84 = {1'b0,$signed(_EVAL_290)};
  assign _EVAL_70 = $signed(_EVAL_84) & $signed(-31'sh2000);
  assign _EVAL_109 = $signed(_EVAL_70);
  assign _EVAL_243 = $signed(_EVAL_109) == $signed(31'sh0);
  assign _EVAL_198 = _EVAL_9[6:3];
  assign _EVAL_106 = _EVAL_198 == 4'h2;
  assign _EVAL_18 = _EVAL_10[2];
  assign _EVAL_253 = _EVAL_18 == 1'h0;
  assign _EVAL_199 = 13'h3f << _EVAL_1;
  assign _EVAL_276 = _EVAL_199[5:0];
  assign _EVAL_226 = ~ _EVAL_276;
  assign _EVAL_77 = _EVAL_226[5:2];
  assign _EVAL_248 = _EVAL_9 == _EVAL_116;
  assign _EVAL_128 = ~ _EVAL_234;
  assign _EVAL_217 = _EVAL_8 & _EVAL_128;
  assign _EVAL_158 = _EVAL_217 == 4'h0;
  assign _EVAL_71 = _EVAL_158 | _EVAL_6;
  assign _EVAL_105 = _EVAL_71 == 1'h0;
  assign _EVAL_172 = _EVAL_2 == _EVAL_26;
  assign _EVAL_209 = _EVAL_14 <= 3'h6;
  assign _EVAL_121 = _EVAL_209 | _EVAL_6;
  assign _EVAL_197 = _EVAL_121 == 1'h0;
  assign _EVAL_122 = _EVAL_9 == 7'h48;
  assign _EVAL_54 = _EVAL_9 == 7'h40;
  assign _EVAL_17 = _EVAL_122 | _EVAL_54;
  assign _EVAL_179 = _EVAL_198 == 4'h8;
  assign _EVAL_230 = _EVAL_9[2:0];
  assign _EVAL_55 = 3'h1 <= _EVAL_230;
  assign _EVAL_195 = _EVAL_179 & _EVAL_55;
  assign _EVAL_61 = _EVAL_17 | _EVAL_195;
  assign _EVAL_274 = _EVAL_9 == 7'h20;
  assign _EVAL_46 = _EVAL_61 | _EVAL_274;
  assign _EVAL_177 = _EVAL_198 == 4'h0;
  assign _EVAL_155 = _EVAL_46 | _EVAL_177;
  assign _EVAL_249 = _EVAL_198 == 4'h1;
  assign _EVAL_247 = _EVAL_155 | _EVAL_249;
  assign _EVAL_189 = _EVAL_15 == 1'h0;
  assign _EVAL_173 = _EVAL_189 | _EVAL_6;
  assign _EVAL_185 = _EVAL_173 == 1'h0;
  assign _EVAL_119 = _EVAL_2 >= 3'h2;
  assign _EVAL_237 = _EVAL_119 | _EVAL_6;
  assign _EVAL_303 = _EVAL_237 == 1'h0;
  assign _EVAL_111 = _EVAL_60 - 4'h1;
  assign _EVAL_153 = ~ _EVAL_8;
  assign _EVAL_262 = _EVAL_153 == 4'h0;
  assign _EVAL_251 = _EVAL_103 | _EVAL_6;
  assign _EVAL_182 = _EVAL_251 == 1'h0;
  assign _EVAL_117 = _EVAL_4 == 7'h40;
  assign _EVAL_200 = 3'h6 == _EVAL_1;
  assign _EVAL_43 = _EVAL_117 ? _EVAL_200 : 1'h0;
  assign _EVAL_202 = _EVAL_43 | _EVAL_6;
  assign _EVAL_49 = _EVAL_247 | _EVAL_106;
  assign _EVAL_20 = _EVAL_198 == 4'h3;
  assign _EVAL_272 = _EVAL_49 | _EVAL_20;
  assign _EVAL_52 = _EVAL_10 == 3'h0;
  assign _EVAL_224 = _EVAL & _EVAL_52;
  assign _EVAL_223 = _EVAL_14[0];
  assign _EVAL_59 = _EVAL_14 == _EVAL_96;
  assign _EVAL_79 = _EVAL_10 == 3'h5;
  assign _EVAL_87 = _EVAL & _EVAL_79;
  assign _EVAL_154 = _EVAL_184 | _EVAL_27;
  assign _EVAL_273 = _EVAL_159 + 32'h1;
  assign _EVAL_164 = _EVAL_10 == _EVAL_261;
  assign _EVAL_275 = _EVAL_164 | _EVAL_6;
  assign _EVAL_294 = _EVAL_4 == 7'h48;
  assign _EVAL_161 = _EVAL_294 | _EVAL_117;
  assign _EVAL_125 = _EVAL_4[6:3];
  assign _EVAL_236 = _EVAL_125 == 4'h8;
  assign _EVAL_35 = _EVAL_4[2:0];
  assign _EVAL_45 = 3'h1 <= _EVAL_35;
  assign _EVAL_110 = _EVAL_236 & _EVAL_45;
  assign _EVAL_57 = _EVAL_161 | _EVAL_110;
  assign _EVAL_206 = _EVAL_4 == 7'h20;
  assign _EVAL_221 = _EVAL_57 | _EVAL_206;
  assign _EVAL_132 = _EVAL_125 == 4'h0;
  assign _EVAL_211 = _EVAL_221 | _EVAL_132;
  assign _EVAL_194 = _EVAL_125 == 4'h1;
  assign _EVAL_242 = _EVAL_211 | _EVAL_194;
  assign _EVAL_268 = _EVAL_125 == 4'h2;
  assign _EVAL_288 = _EVAL_242 | _EVAL_268;
  assign _EVAL_91 = _EVAL_125 == 4'h3;
  assign _EVAL_231 = _EVAL_288 | _EVAL_91;
  assign _EVAL_292 = _EVAL_1 == _EVAL_53;
  assign _EVAL_300 = _EVAL_292 | _EVAL_6;
  assign _EVAL_42 = _EVAL_300 == 1'h0;
  assign _EVAL_175 = _EVAL_13 == _EVAL_94;
  assign _EVAL_40 = _EVAL_175 | _EVAL_6;
  assign _EVAL_180 = _EVAL_40 == 1'h0;
  assign _EVAL_270 = _EVAL_75 - 4'h1;
  assign _EVAL_118 = _EVAL_60 == 4'h0;
  assign _EVAL_170 = 13'h3f << _EVAL_2;
  assign _EVAL_95 = _EVAL_170[5:0];
  assign _EVAL_107 = ~ _EVAL_95;
  assign _EVAL_259 = _EVAL_107[5:2];
  assign _EVAL_48 = _EVAL_1 <= 3'h6;
  assign _EVAL_232 = _EVAL_48 & _EVAL_243;
  assign _EVAL_219 = _EVAL_232 | _EVAL_6;
  assign _EVAL_254 = _EVAL_219 == 1'h0;
  assign _EVAL_24 = _EVAL_272 | _EVAL_6;
  assign _EVAL_124 = _EVAL_163 - 4'h1;
  assign _EVAL_214 = {{24'd0}, _EVAL_226};
  assign _EVAL_135 = _EVAL_295 >> _EVAL_4;
  assign _EVAL_192 = _EVAL_3 == 1'h0;
  assign _EVAL_85 = _EVAL_192 | _EVAL_6;
  assign _EVAL_140 = _EVAL_135[0];
  assign _EVAL_212 = _EVAL_262 | _EVAL_6;
  assign _EVAL_289 = _EVAL_162 | _EVAL_3;
  assign _EVAL_62 = _EVAL_289 | _EVAL_6;
  assign _EVAL_28 = _EVAL_62 == 1'h0;
  assign _EVAL_99 = _EVAL_140 == 1'h0;
  assign _EVAL_246 = _EVAL_99 | _EVAL_6;
  assign _EVAL_56 = _EVAL_13 <= 3'h2;
  assign _EVAL_127 = _EVAL_56 | _EVAL_6;
  assign _EVAL_255 = _EVAL_127 == 1'h0;
  assign _EVAL_283 = _EVAL_172 | _EVAL_6;
  assign _EVAL_21 = _EVAL_81 != _EVAL_208;
  assign _EVAL_64 = _EVAL_81 != 73'h0;
  assign _EVAL_210 = _EVAL_64 == 1'h0;
  assign _EVAL_114 = _EVAL_21 | _EVAL_210;
  assign _EVAL_25 = _EVAL_13 != 3'h0;
  assign _EVAL_123 = _EVAL_25 | _EVAL_6;
  assign _EVAL_67 = _EVAL_11 == _EVAL_101;
  assign _EVAL_181 = _EVAL_67 | _EVAL_6;
  assign _EVAL_183 = _EVAL_231 | _EVAL_6;
  assign _EVAL_228 = _EVAL_183 == 1'h0;
  assign _EVAL_171 = _EVAL_184 & _EVAL_282;
  assign _EVAL_73 = _EVAL_246 == 1'h0;
  assign _EVAL_201 = _EVAL_248 | _EVAL_6;
  assign _EVAL_222 = _EVAL_201 == 1'h0;
  assign _EVAL_34 = _EVAL_244 == 1'h0;
  assign _EVAL_30 = _EVAL_14 == 3'h4;
  assign _EVAL_299 = _EVAL_16 & _EVAL_30;
  assign _EVAL_29 = _EVAL_59 | _EVAL_6;
  assign _EVAL_240 = _EVAL_29 == 1'h0;
  assign _EVAL_302 = _EVAL_6 == 1'h0;
  assign _EVAL_252 = _EVAL_275 == 1'h0;
  assign _EVAL_137 = _EVAL_10 == 3'h2;
  assign _EVAL_89 = _EVAL & _EVAL_137;
  assign _EVAL_37 = _EVAL_112 - 4'h1;
  assign _EVAL_41 = _EVAL_4 == _EVAL_168;
  assign _EVAL_100 = _EVAL & _EVAL_98;
  assign _EVAL_139 = _EVAL_283 == 1'h0;
  assign _EVAL_267 = _EVAL_10 == 3'h6;
  assign _EVAL_178 = _EVAL_14 == 3'h1;
  assign _EVAL_19 = _EVAL_10 == 3'h3;
  assign _EVAL_115 = _EVAL_258 | _EVAL_6;
  assign _EVAL_39 = _EVAL_115 == 1'h0;
  assign _EVAL_287 = _EVAL_114 | _EVAL_6;
  assign _EVAL_22 = _EVAL_287 == 1'h0;
  assign _EVAL_169 = _EVAL_41 | _EVAL_6;
  assign _EVAL_76 = _EVAL_10 == 3'h7;
  assign _EVAL_235 = _EVAL_11 & _EVAL_214;
  assign _EVAL_97 = _EVAL_235 == 30'h0;
  assign _EVAL_126 = _EVAL_97 | _EVAL_6;
  assign _EVAL_215 = _EVAL_202 == 1'h0;
  assign _EVAL_143 = _EVAL_212 == 1'h0;
  assign _EVAL_298 = _EVAL_81 | _EVAL_295;
  assign _EVAL_82 = _EVAL_298 >> _EVAL_9;
  assign _EVAL_188 = _EVAL_82[0];
  assign _EVAL_78 = _EVAL_169 == 1'h0;
  assign _EVAL_271 = _EVAL_126 == 1'h0;
  assign _EVAL_191 = _EVAL_14 == 3'h0;
  assign _EVAL_205 = _EVAL & _EVAL_267;
  assign _EVAL_131 = _EVAL_174 | _EVAL_6;
  assign _EVAL_260 = _EVAL_10 == 3'h4;
  assign _EVAL_157 = _EVAL & _EVAL_260;
  assign _EVAL_225 = _EVAL_14 == 3'h2;
  assign _EVAL_297 = _EVAL_16 & _EVAL_225;
  assign _EVAL_90 = _EVAL_16 & _EVAL_191;
  assign _EVAL_129 = _EVAL_85 == 1'h0;
  assign _EVAL_88 = _EVAL_131 == 1'h0;
  assign _EVAL_187 = _EVAL_118 == 1'h0;
  assign _EVAL_152 = _EVAL_16 & _EVAL_33;
  assign _EVAL_146 = _EVAL_123 == 1'h0;
  assign _EVAL_284 = _EVAL_13 == 3'h0;
  assign _EVAL_66 = _EVAL_284 | _EVAL_6;
  assign _EVAL_93 = _EVAL_16 & _EVAL_178;
  assign _EVAL_141 = _EVAL_188 | _EVAL_6;
  assign _EVAL_239 = _EVAL_141 == 1'h0;
  assign _EVAL_207 = _EVAL_27 & _EVAL_118;
  assign _EVAL_286 = _EVAL & _EVAL_76;
  assign _EVAL_113 = _EVAL_181 == 1'h0;
  assign _EVAL_190 = _EVAL_24 == 1'h0;
  assign _EVAL_296 = _EVAL_66 == 1'h0;
  assign _EVAL_38 = _EVAL & _EVAL_19;
  assign _EVAL_51 = _EVAL_16 & _EVAL_187;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_53 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_60 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_75 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_94 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_96 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_101 = _RAND_6[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_112 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_116 = _RAND_8[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_147 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_159 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_163 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_168 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_261 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {3{`RANDOM}};
  _EVAL_295 = _RAND_14[72:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_5) begin
    if (_EVAL_207) begin
      _EVAL_26 <= _EVAL_2;
    end
    if (_EVAL_171) begin
      _EVAL_53 <= _EVAL_1;
    end
    if (_EVAL_6) begin
      _EVAL_60 <= 4'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_118) begin
          if (_EVAL_223) begin
            _EVAL_60 <= _EVAL_259;
          end else begin
            _EVAL_60 <= 4'h0;
          end
        end else begin
          _EVAL_60 <= _EVAL_111;
        end
      end
    end
    if (_EVAL_6) begin
      _EVAL_75 <= 4'h0;
    end else begin
      if (_EVAL_184) begin
        if (_EVAL_282) begin
          if (_EVAL_253) begin
            _EVAL_75 <= _EVAL_77;
          end else begin
            _EVAL_75 <= 4'h0;
          end
        end else begin
          _EVAL_75 <= _EVAL_270;
        end
      end
    end
    if (_EVAL_171) begin
      _EVAL_94 <= _EVAL_13;
    end
    if (_EVAL_207) begin
      _EVAL_96 <= _EVAL_14;
    end
    if (_EVAL_171) begin
      _EVAL_101 <= _EVAL_11;
    end
    if (_EVAL_6) begin
      _EVAL_112 <= 4'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_281) begin
          if (_EVAL_223) begin
            _EVAL_112 <= _EVAL_259;
          end else begin
            _EVAL_112 <= 4'h0;
          end
        end else begin
          _EVAL_112 <= _EVAL_37;
        end
      end
    end
    if (_EVAL_207) begin
      _EVAL_116 <= _EVAL_9;
    end
    if (_EVAL_207) begin
      _EVAL_147 <= _EVAL_0;
    end
    if (_EVAL_6) begin
      _EVAL_159 <= 32'h0;
    end else begin
      if (_EVAL_154) begin
        _EVAL_159 <= 32'h0;
      end else begin
        _EVAL_159 <= _EVAL_273;
      end
    end
    if (_EVAL_6) begin
      _EVAL_163 <= 4'h0;
    end else begin
      if (_EVAL_184) begin
        if (_EVAL_65) begin
          if (_EVAL_253) begin
            _EVAL_163 <= _EVAL_77;
          end else begin
            _EVAL_163 <= 4'h0;
          end
        end else begin
          _EVAL_163 <= _EVAL_124;
        end
      end
    end
    if (_EVAL_171) begin
      _EVAL_168 <= _EVAL_4;
    end
    if (_EVAL_171) begin
      _EVAL_261 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_295 <= 73'h0;
    end else begin
      _EVAL_295 <= _EVAL_220;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a49d58d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1ca035c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2be3696)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da0df18a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c984872)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74a443cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e85e3bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73cba4b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b948d4f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a37a3f53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b908e00b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53b0b0c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d60b01d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f31f29cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83a77fc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0f9d7ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71760da1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db657f3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb81df06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51147d37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0c7013e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e329abf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d25dbf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96020b89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24670b47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c4260d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3fef5ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14aacde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a2a396c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6997956f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bddacaa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36211997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36739b68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f7dd11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(988f12cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34e06f35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb9106c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5146df60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b6e7827)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3510cd5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b41a9cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30a3a270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cc19e32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7740d27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c673c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a499825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2988185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(420a2c6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78d04c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3305d58d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1869541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6e8b82f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b879ba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c16ea186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c54adf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddbb480c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18c54783)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(544c950f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb2de4aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29d54bdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1569b24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2be88b74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8c69adb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b5bb1d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebfefc10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c254a658)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b544420a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da98189d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3756e266)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(345b0e09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cf5b90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(266f2e84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8f2106c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71d7014b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb90b53e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a587d44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(393e8044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77487cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb96e96b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbe2c0f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
