//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_287(
  input  [29:0] _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  output [1:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output [31:0] _EVAL_6,
  input  [29:0] _EVAL_7,
  input         _EVAL_8,
  output [1:0]  _EVAL_9,
  output [29:0] _EVAL_10,
  output        _EVAL_11,
  output [31:0] _EVAL_12,
  input  [29:0] _EVAL_13,
  output [1:0]  _EVAL_14,
  output [31:0] _EVAL_15,
  input         _EVAL_16,
  output [29:0] _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input  [31:0] _EVAL_21,
  output [31:0] _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output [1:0]  _EVAL_25,
  output [31:0] _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [31:0] _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  output [1:0]  _EVAL_31,
  output        _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input  [29:0] _EVAL_35,
  output        _EVAL_36,
  input         _EVAL_37,
  input  [1:0]  _EVAL_38,
  output        _EVAL_39,
  output        _EVAL_40,
  output [29:0] _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  output        _EVAL_45,
  output        _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  input  [1:0]  _EVAL_49,
  output [29:0] _EVAL_50,
  output        _EVAL_51,
  input         _EVAL_52,
  output [1:0]  _EVAL_53,
  output        _EVAL_54,
  output [29:0] _EVAL_55,
  input  [1:0]  _EVAL_56,
  output        _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  output        _EVAL_60,
  output        _EVAL_61,
  output [1:0]  _EVAL_62,
  output [1:0]  _EVAL_63,
  input         _EVAL_64,
  output [1:0]  _EVAL_65,
  output        _EVAL_66,
  input         _EVAL_67,
  output        _EVAL_68,
  input  [31:0] _EVAL_69,
  input         _EVAL_70,
  output [1:0]  _EVAL_71,
  input         _EVAL_72,
  input         _EVAL_73,
  output [29:0] _EVAL_74,
  output        _EVAL_75,
  output        _EVAL_76,
  input         _EVAL_77,
  output [31:0] _EVAL_78,
  output [1:0]  _EVAL_79,
  output        _EVAL_80,
  input         _EVAL_81,
  output [31:0] _EVAL_82,
  input         _EVAL_83,
  input  [29:0] _EVAL_84,
  output        _EVAL_85,
  output        _EVAL_86,
  output        _EVAL_87,
  output [1:0]  _EVAL_88,
  output [29:0] _EVAL_89,
  output [1:0]  _EVAL_90,
  output        _EVAL_91,
  output        _EVAL_92,
  output        _EVAL_93,
  output [31:0] _EVAL_94,
  output        _EVAL_95,
  input  [31:0] _EVAL_96,
  output        _EVAL_97,
  input  [29:0] _EVAL_98,
  input  [1:0]  _EVAL_99,
  output        _EVAL_100,
  input         _EVAL_101,
  output [29:0] _EVAL_102,
  output [1:0]  _EVAL_103,
  output [31:0] _EVAL_104,
  input         _EVAL_105,
  output [31:0] _EVAL_106,
  output [1:0]  _EVAL_107,
  output [31:0] _EVAL_108,
  input         _EVAL_109,
  output        _EVAL_110,
  output        _EVAL_111,
  input  [29:0] _EVAL_112,
  output        _EVAL_113,
  input         _EVAL_114,
  input         _EVAL_115,
  output        _EVAL_116,
  output [31:0] _EVAL_117,
  output        _EVAL_118,
  input  [1:0]  _EVAL_119,
  output        _EVAL_120,
  input         _EVAL_121,
  output [29:0] _EVAL_122,
  output        _EVAL_123,
  output        _EVAL_124,
  input  [1:0]  _EVAL_125,
  output        _EVAL_126,
  output        _EVAL_127,
  output        _EVAL_128,
  output [31:0] _EVAL_129,
  output [29:0] _EVAL_130,
  output        _EVAL_131,
  input  [1:0]  _EVAL_132,
  input  [31:0] _EVAL_133,
  output        _EVAL_134,
  output        _EVAL_135,
  output [29:0] _EVAL_136,
  output        _EVAL_137,
  output        _EVAL_138,
  output        _EVAL_139,
  output        _EVAL_140,
  input  [31:0] _EVAL_141,
  input         _EVAL_142,
  output        _EVAL_143,
  input         _EVAL_144,
  output [31:0] _EVAL_145,
  output        _EVAL_146,
  input         _EVAL_147,
  input  [1:0]  _EVAL_148,
  output        _EVAL_149,
  output [29:0] _EVAL_150,
  output [1:0]  _EVAL_151,
  output [1:0]  _EVAL_152,
  output        _EVAL_153,
  output [31:0] _EVAL_154,
  output [31:0] _EVAL_155,
  input  [29:0] _EVAL_156,
  output [1:0]  _EVAL_157,
  output        _EVAL_158,
  input  [31:0] _EVAL_159,
  output [29:0] _EVAL_160,
  input  [1:0]  _EVAL_161,
  input         _EVAL_162,
  output        _EVAL_163,
  output        _EVAL_164,
  input  [1:0]  _EVAL_165,
  output        _EVAL_166,
  output        _EVAL_167,
  output [31:0] _EVAL_168,
  input  [31:0] _EVAL_169,
  output        _EVAL_170,
  output [29:0] _EVAL_171,
  output        _EVAL_172,
  output [29:0] _EVAL_173,
  output        _EVAL_174,
  output [29:0] _EVAL_175,
  output        _EVAL_176,
  input         _EVAL_177,
  input         _EVAL_178,
  input         _EVAL_179
);
  wire  arb__EVAL;
  wire  arb__EVAL_0;
  wire  arb__EVAL_1;
  wire [2:0] packageanon1__EVAL;
  wire [2:0] packageanon1__EVAL_0;
  reg [2:0] _EVAL_185;
  reg [31:0] _RAND_0;
  wire  _EVAL_189;
  wire  _EVAL_182;
  wire  _EVAL_188;
  wire  _EVAL_187;
  wire [2:0] _EVAL_181;
  wire [2:0] _EVAL_184;
  wire [2:0] _EVAL_186;
  wire [2:0] _EVAL_183;
  wire  _EVAL_180;
  SiFive__EVAL_285 arb (
    ._EVAL(arb__EVAL),
    ._EVAL_0(arb__EVAL_0),
    ._EVAL_1(arb__EVAL_1)
  );
  SiFive__EVAL_286 packageanon1 (
    ._EVAL(packageanon1__EVAL),
    ._EVAL_0(packageanon1__EVAL_0)
  );
  assign _EVAL_189 = 3'h4 == _EVAL_185;
  assign _EVAL_182 = 3'h2 == _EVAL_185;
  assign _EVAL_188 = 3'h1 == _EVAL_185;
  assign _EVAL_187 = 3'h7 == _EVAL_185;
  assign _EVAL_181 = _EVAL_187 ? 3'h0 : _EVAL_185;
  assign _EVAL_184 = _EVAL_189 ? 3'h5 : _EVAL_181;
  assign _EVAL_186 = _EVAL_182 ? 3'h4 : _EVAL_184;
  assign _EVAL_183 = _EVAL_188 ? 3'h1 : _EVAL_186;
  assign _EVAL_180 = 3'h0 == _EVAL_185;
  assign _EVAL_23 = _EVAL_179;
  assign _EVAL_61 = _EVAL_67;
  assign _EVAL_130 = _EVAL_13;
  assign _EVAL_158 = _EVAL_178;
  assign _EVAL_12 = _EVAL_21;
  assign _EVAL_152 = _EVAL_132;
  assign _EVAL_65 = _EVAL_119;
  assign _EVAL_155 = _EVAL_141;
  assign _EVAL_3 = _EVAL_165;
  assign _EVAL_140 = _EVAL_142;
  assign _EVAL_68 = _EVAL_77;
  assign _EVAL_108 = _EVAL_69;
  assign _EVAL_127 = _EVAL_0;
  assign _EVAL_24 = _EVAL_33;
  assign _EVAL_60 = _EVAL_67;
  assign _EVAL_146 = _EVAL_72;
  assign _EVAL_166 = _EVAL_177;
  assign _EVAL_46 = _EVAL_121;
  assign _EVAL_120 = _EVAL_4;
  assign _EVAL_71 = _EVAL_119;
  assign _EVAL_145 = _EVAL_28;
  assign _EVAL_110 = _EVAL_59;
  assign _EVAL_163 = _EVAL_72;
  assign _EVAL_39 = _EVAL_64;
  assign _EVAL_93 = _EVAL_70;
  assign _EVAL_160 = _EVAL_7;
  assign _EVAL_48 = _EVAL_8;
  assign _EVAL_129 = _EVAL_27;
  assign _EVAL_131 = _EVAL_52;
  assign _EVAL_9 = _EVAL_49;
  assign _EVAL_143 = _EVAL_83;
  assign _EVAL_44 = _EVAL_121;
  assign _EVAL_135 = _EVAL_105;
  assign _EVAL_170 = _EVAL_147;
  assign _EVAL_89 = _EVAL_35;
  assign _EVAL_55 = _EVAL;
  assign _EVAL_168 = _EVAL_28;
  assign _EVAL_25 = _EVAL_99;
  assign _EVAL_14 = _EVAL_49;
  assign _EVAL_51 = _EVAL_59;
  assign _EVAL_126 = _EVAL_34;
  assign _EVAL_47 = _EVAL_77;
  assign _EVAL_103 = _EVAL_148;
  assign _EVAL_153 = _EVAL_58;
  assign _EVAL_100 = _EVAL_5;
  assign _EVAL_134 = _EVAL_5;
  assign _EVAL_82 = _EVAL_133;
  assign _EVAL_173 = _EVAL_112;
  assign _EVAL_6 = _EVAL_159;
  assign _EVAL_171 = _EVAL_35;
  assign _EVAL_85 = _EVAL_70;
  assign _EVAL_88 = _EVAL_38;
  assign _EVAL_32 = _EVAL_115;
  assign _EVAL_111 = _EVAL_20;
  assign _EVAL_42 = _EVAL_144;
  assign _EVAL_136 = _EVAL_112;
  assign _EVAL_167 = _EVAL_16;
  assign _EVAL_19 = _EVAL_16;
  assign _EVAL_31 = _EVAL_56;
  assign _EVAL_50 = _EVAL_98;
  assign _EVAL_139 = _EVAL_20;
  assign _EVAL_74 = _EVAL_7;
  assign _EVAL_91 = arb__EVAL_1;
  assign arb__EVAL_0 = _EVAL_185 == 3'h0;
  assign _EVAL_15 = _EVAL_96;
  assign _EVAL_10 = _EVAL_156;
  assign _EVAL_154 = _EVAL_96;
  assign _EVAL_117 = _EVAL_133;
  assign _EVAL_116 = _EVAL_114;
  assign _EVAL_63 = _EVAL_38;
  assign _EVAL_90 = _EVAL_148;
  assign _EVAL_174 = _EVAL_142;
  assign _EVAL_150 = _EVAL_156;
  assign _EVAL_113 = _EVAL_64;
  assign _EVAL_175 = _EVAL_98;
  assign _EVAL_102 = _EVAL_84;
  assign _EVAL_92 = _EVAL_0;
  assign packageanon1__EVAL_0 = _EVAL_180 ? _EVAL_185 : _EVAL_183;
  assign _EVAL_157 = _EVAL_165;
  assign _EVAL_164 = _EVAL_34;
  assign _EVAL_17 = _EVAL;
  assign _EVAL_87 = _EVAL_37;
  assign _EVAL_40 = _EVAL_109;
  assign _EVAL_122 = _EVAL_13;
  assign _EVAL_118 = _EVAL_43;
  assign _EVAL_97 = _EVAL_8;
  assign _EVAL_149 = _EVAL_105;
  assign _EVAL_62 = _EVAL_125;
  assign _EVAL_107 = _EVAL_161;
  assign _EVAL_106 = _EVAL_69;
  assign _EVAL_22 = _EVAL_169;
  assign _EVAL_80 = _EVAL_4;
  assign _EVAL_137 = _EVAL_52;
  assign _EVAL_36 = _EVAL_81;
  assign _EVAL_53 = _EVAL_125;
  assign _EVAL_138 = _EVAL_162;
  assign _EVAL_54 = _EVAL_162;
  assign _EVAL_95 = _EVAL_144;
  assign _EVAL_26 = _EVAL_159;
  assign _EVAL_30 = _EVAL_114;
  assign _EVAL_66 = _EVAL_58;
  assign _EVAL_86 = _EVAL_73;
  assign _EVAL_123 = _EVAL_115;
  assign _EVAL_41 = _EVAL_84;
  assign _EVAL_11 = _EVAL_81;
  assign _EVAL_104 = _EVAL_141;
  assign _EVAL_176 = _EVAL_178;
  assign _EVAL_94 = _EVAL_27;
  assign _EVAL_128 = _EVAL_179;
  assign _EVAL_76 = _EVAL_109;
  assign _EVAL_124 = _EVAL_33;
  assign _EVAL_79 = _EVAL_99;
  assign _EVAL_45 = _EVAL_83;
  assign _EVAL_172 = _EVAL_147;
  assign _EVAL_78 = _EVAL_169;
  assign _EVAL_18 = arb__EVAL;
  assign _EVAL_29 = _EVAL_177;
  assign _EVAL_57 = _EVAL_43;
  assign _EVAL_1 = _EVAL_37;
  assign _EVAL_75 = _EVAL_73;
  assign _EVAL_151 = _EVAL_132;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_185 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_2) begin
    if (_EVAL_101) begin
      _EVAL_185 <= 3'h0;
    end else begin
      _EVAL_185 <= packageanon1__EVAL;
    end
  end
endmodule
