//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_252_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [31:0] _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  input         _EVAL_20,
  input  [2:0]  _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [2:0]  _EVAL_25,
  input  [31:0] _EVAL_26,
  input  [1:0]  _EVAL_27,
  input  [7:0]  _EVAL_28,
  input  [3:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [31:0] _EVAL_33
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_74;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_80;
  reg [31:0] _RAND_1;
  reg [1:0] _EVAL_90;
  reg [31:0] _RAND_2;
  reg [4:0] _EVAL_111;
  reg [31:0] _RAND_3;
  reg [31:0] _EVAL_159;
  reg [31:0] _RAND_4;
  reg [4:0] _EVAL_164;
  reg [31:0] _RAND_5;
  reg [4:0] _EVAL_174;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_180;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_201;
  reg [31:0] _RAND_8;
  reg [4:0] _EVAL_243;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_253;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_277;
  reg [31:0] _RAND_11;
  reg [4:0] _EVAL_296;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_356;
  reg [31:0] _RAND_13;
  reg [1:0] _EVAL_390;
  reg [31:0] _RAND_14;
  reg [4:0] _EVAL_406;
  reg [31:0] _RAND_15;
  reg  _EVAL_437;
  reg [31:0] _RAND_16;
  reg [31:0] _EVAL_446;
  reg [31:0] _RAND_17;
  reg  _EVAL_456;
  reg [31:0] _RAND_18;
  reg [2:0] _EVAL_478;
  reg [31:0] _RAND_19;
  reg [31:0] _EVAL_492;
  reg [31:0] _RAND_20;
  reg [3:0] _EVAL_500;
  reg [31:0] _RAND_21;
  reg [31:0] _EVAL_551;
  reg [31:0] _RAND_22;
  reg [2:0] _EVAL_552;
  reg [31:0] _RAND_23;
  reg [4:0] _EVAL_557;
  reg [31:0] _RAND_24;
  reg [7:0] _EVAL_566;
  reg [31:0] _RAND_25;
  reg [1:0] _EVAL_567;
  reg [31:0] _RAND_26;
  reg [2:0] _EVAL_644;
  reg [31:0] _RAND_27;
  wire  _EVAL_317;
  wire  _EVAL_423;
  wire  _EVAL_403;
  wire [31:0] _EVAL_285;
  wire [32:0] _EVAL_618;
  wire [32:0] _EVAL_355;
  wire [32:0] _EVAL_324;
  wire  _EVAL_626;
  wire  _EVAL_625;
  wire  _EVAL_522;
  wire [22:0] _EVAL_431;
  wire [7:0] _EVAL_602;
  wire [7:0] _EVAL_586;
  wire [31:0] _EVAL_509;
  wire [31:0] _EVAL_571;
  wire [32:0] _EVAL_128;
  wire [32:0] _EVAL_614;
  wire [32:0] _EVAL_224;
  wire  _EVAL_234;
  wire [31:0] _EVAL_595;
  wire  _EVAL_358;
  wire [1:0] _EVAL_579;
  wire [3:0] _EVAL_177;
  wire [2:0] _EVAL_176;
  wire [2:0] _EVAL_455;
  wire  _EVAL_261;
  wire  _EVAL_382;
  wire  _EVAL_611;
  wire [31:0] _EVAL_638;
  wire [32:0] _EVAL_501;
  wire [32:0] _EVAL_134;
  wire [32:0] _EVAL_83;
  wire  _EVAL_152;
  wire [31:0] _EVAL_172;
  wire [32:0] _EVAL_233;
  wire [32:0] _EVAL_142;
  wire [22:0] _EVAL_475;
  wire [7:0] _EVAL_599;
  wire [7:0] _EVAL_291;
  wire [31:0] _EVAL_604;
  wire [31:0] _EVAL_531;
  wire  _EVAL_636;
  wire  _EVAL_131;
  wire  _EVAL_310;
  wire  _EVAL_60;
  wire  _EVAL_52;
  wire  _EVAL_512;
  wire  _EVAL_284;
  wire  _EVAL_578;
  wire  _EVAL_589;
  wire  _EVAL_487;
  wire [1:0] _EVAL_556;
  wire [1:0] _EVAL_535;
  wire [1:0] _EVAL_210;
  wire [1:0] _EVAL_235;
  wire  _EVAL_102;
  wire  _EVAL_425;
  wire  _EVAL_649;
  wire  _EVAL_273;
  wire  _EVAL_464;
  wire  _EVAL_191;
  wire  _EVAL_86;
  wire  _EVAL_384;
  wire  _EVAL_219;
  wire  _EVAL_267;
  wire [32:0] _EVAL_247;
  wire [32:0] _EVAL_352;
  wire [32:0] _EVAL_278;
  wire [31:0] _EVAL_603;
  wire [32:0] _EVAL_213;
  wire [32:0] _EVAL_183;
  wire [32:0] _EVAL_438;
  wire  _EVAL_440;
  wire  _EVAL_443;
  wire  _EVAL_133;
  wire  _EVAL_272;
  wire [31:0] _EVAL_282;
  wire [32:0] _EVAL_195;
  wire [32:0] _EVAL_650;
  wire [32:0] _EVAL_511;
  wire  _EVAL_519;
  wire [31:0] _EVAL_612;
  wire [32:0] _EVAL_517;
  wire [32:0] _EVAL_262;
  wire [32:0] _EVAL_76;
  wire  _EVAL_196;
  wire  _EVAL_157;
  wire  _EVAL_570;
  wire  _EVAL_258;
  wire  _EVAL_392;
  wire  _EVAL_114;
  wire  _EVAL_184;
  wire  _EVAL_375;
  wire  _EVAL_583;
  wire  _EVAL_479;
  wire  _EVAL_146;
  wire  _EVAL_504;
  wire  _EVAL_387;
  wire  _EVAL_232;
  wire  _EVAL_394;
  wire  _EVAL_476;
  wire  _EVAL_226;
  wire  _EVAL_365;
  wire  _EVAL_628;
  wire  _EVAL_484;
  wire [31:0] _EVAL_275;
  wire [32:0] _EVAL_572;
  wire [32:0] _EVAL_155;
  wire [32:0] _EVAL_140;
  wire [7:0] _EVAL_533;
  wire [31:0] _EVAL_75;
  wire [32:0] _EVAL_354;
  wire [32:0] _EVAL_491;
  wire [32:0] _EVAL_477;
  wire [1:0] _EVAL_441;
  wire  _EVAL_153;
  wire  _EVAL_71;
  wire  _EVAL_574;
  wire  _EVAL_208;
  wire [32:0] _EVAL_444;
  wire [32:0] _EVAL_601;
  wire [32:0] _EVAL_245;
  wire  _EVAL_434;
  wire [31:0] _EVAL_345;
  wire [32:0] _EVAL_320;
  wire [32:0] _EVAL_591;
  wire [32:0] _EVAL_199;
  wire  _EVAL_150;
  wire  _EVAL_359;
  wire [31:0] _EVAL_106;
  wire [32:0] _EVAL_417;
  wire [32:0] _EVAL_268;
  wire [32:0] _EVAL_427;
  wire  _EVAL_182;
  wire  _EVAL_369;
  wire [31:0] _EVAL_353;
  wire [32:0] _EVAL_53;
  wire [32:0] _EVAL_383;
  wire [32:0] _EVAL_115;
  wire  _EVAL_46;
  wire  _EVAL_577;
  wire  _EVAL_581;
  wire  _EVAL_373;
  wire [31:0] _EVAL_316;
  wire [32:0] _EVAL_116;
  wire [32:0] _EVAL_460;
  wire [32:0] _EVAL_85;
  wire  _EVAL_540;
  wire  _EVAL_147;
  wire [31:0] _EVAL_592;
  wire [32:0] _EVAL_113;
  wire [32:0] _EVAL_607;
  wire [32:0] _EVAL_309;
  wire  _EVAL_294;
  wire  _EVAL_388;
  wire [31:0] _EVAL_158;
  wire [32:0] _EVAL_209;
  wire [32:0] _EVAL_483;
  wire [32:0] _EVAL_279;
  wire  _EVAL_582;
  wire  _EVAL_429;
  wire  _EVAL_276;
  wire  _EVAL_585;
  wire  _EVAL_205;
  wire  _EVAL_162;
  wire  _EVAL_445;
  wire  _EVAL_206;
  wire  _EVAL_154;
  wire  _EVAL_421;
  wire  _EVAL_178;
  wire  _EVAL_536;
  wire  _EVAL_346;
  wire  _EVAL_218;
  wire  _EVAL_584;
  wire [31:0] _EVAL_493;
  wire [32:0] _EVAL_494;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_610;
  wire  _EVAL_143;
  wire  _EVAL_41;
  wire [31:0] _EVAL_343;
  wire [32:0] _EVAL_188;
  wire [32:0] _EVAL_553;
  wire [32:0] _EVAL_596;
  wire  _EVAL_404;
  wire  _EVAL_170;
  wire  _EVAL_313;
  wire  _EVAL_331;
  wire  _EVAL_333;
  wire [31:0] _EVAL_399;
  wire [32:0] _EVAL_528;
  wire [32:0] _EVAL_319;
  wire [32:0] _EVAL_575;
  wire  _EVAL_211;
  wire  _EVAL_499;
  wire  _EVAL_393;
  wire  _EVAL_400;
  wire [31:0] _EVAL_190;
  wire [32:0] _EVAL_600;
  wire [32:0] _EVAL_468;
  wire [32:0] _EVAL_486;
  wire  _EVAL_503;
  wire  _EVAL_56;
  wire [31:0] _EVAL_264;
  wire [32:0] _EVAL_237;
  wire [32:0] _EVAL_148;
  wire [32:0] _EVAL_192;
  wire  _EVAL_633;
  wire  _EVAL_651;
  wire [31:0] _EVAL_368;
  wire [32:0] _EVAL_588;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_89;
  wire  _EVAL_70;
  wire  _EVAL_629;
  wire  _EVAL_250;
  wire  _EVAL_79;
  wire  _EVAL_415;
  wire [4:0] _EVAL_168;
  wire [4:0] _EVAL_545;
  wire  _EVAL_424;
  wire  _EVAL_334;
  wire [32:0] _EVAL_520;
  wire  _EVAL_458;
  wire [31:0] _EVAL_380;
  wire [32:0] _EVAL_121;
  wire [32:0] _EVAL_321;
  wire [32:0] _EVAL_179;
  wire  _EVAL_40;
  wire  _EVAL_127;
  wire [31:0] _EVAL_318;
  wire [32:0] _EVAL_221;
  wire [32:0] _EVAL_336;
  wire [32:0] _EVAL_330;
  wire  _EVAL_305;
  wire  _EVAL_559;
  wire [31:0] _EVAL_467;
  wire [32:0] _EVAL_81;
  wire [32:0] _EVAL_169;
  wire [32:0] _EVAL_546;
  wire  _EVAL_255;
  wire  _EVAL_271;
  wire  _EVAL_547;
  wire  _EVAL_544;
  wire [32:0] _EVAL_481;
  wire [32:0] _EVAL_634;
  wire [32:0] _EVAL_510;
  wire  _EVAL_529;
  wire  _EVAL_292;
  wire  _EVAL_107;
  wire [31:0] _EVAL_307;
  wire [32:0] _EVAL_560;
  wire [32:0] _EVAL_428;
  wire [32:0] _EVAL_489;
  wire  _EVAL_43;
  wire  _EVAL_236;
  wire  _EVAL_418;
  wire  _EVAL_653;
  wire [31:0] _EVAL_370;
  wire [32:0] _EVAL_357;
  wire [32:0] _EVAL_42;
  wire [32:0] _EVAL_68;
  wire  _EVAL_91;
  wire  _EVAL_624;
  wire  _EVAL_364;
  wire  _EVAL_442;
  wire  _EVAL_381;
  wire  _EVAL_516;
  wire  _EVAL_340;
  wire  _EVAL_93;
  wire  _EVAL_525;
  wire  _EVAL_621;
  wire  _EVAL_300;
  wire  _EVAL_97;
  wire [22:0] _EVAL_351;
  wire [7:0] _EVAL_376;
  wire [7:0] _EVAL_457;
  wire [4:0] _EVAL_61;
  wire [4:0] _EVAL_401;
  wire  _EVAL_362;
  wire  _EVAL_590;
  wire  _EVAL_502;
  wire [7:0] _EVAL_101;
  wire  _EVAL_216;
  wire  _EVAL_405;
  wire  _EVAL_136;
  wire  _EVAL_57;
  wire  _EVAL_378;
  wire  _EVAL_266;
  wire  _EVAL_120;
  wire  _EVAL_96;
  wire  _EVAL_341;
  wire  _EVAL_123;
  wire  _EVAL_514;
  wire  _EVAL_426;
  wire  _EVAL_198;
  wire  _EVAL_637;
  wire  _EVAL_422;
  wire  _EVAL_145;
  wire  _EVAL_549;
  wire  _EVAL_608;
  wire  _EVAL_366;
  wire  _EVAL_204;
  wire [31:0] _EVAL_409;
  wire  _EVAL_265;
  wire  _EVAL_543;
  wire  _EVAL_248;
  wire  _EVAL_200;
  wire  _EVAL_451;
  wire  _EVAL_413;
  wire  _EVAL_328;
  wire  _EVAL_58;
  wire  _EVAL_173;
  wire  _EVAL_646;
  wire  _EVAL_408;
  wire  _EVAL_249;
  wire  _EVAL_523;
  wire [4:0] _EVAL_623;
  wire  _EVAL_436;
  wire  _EVAL_214;
  wire  _EVAL_447;
  wire  _EVAL_227;
  wire  _EVAL_78;
  wire  _EVAL_297;
  wire  _EVAL_295;
  wire  _EVAL_87;
  wire  _EVAL_642;
  wire  _EVAL_54;
  wire  _EVAL_532;
  wire  _EVAL_555;
  wire  _EVAL_342;
  wire  _EVAL_160;
  wire  _EVAL_45;
  wire  _EVAL_565;
  wire  _EVAL_548;
  wire [1:0] _EVAL_312;
  wire  _EVAL_505;
  wire  _EVAL_315;
  wire  _EVAL_507;
  wire  _EVAL_374;
  wire  _EVAL_361;
  wire  _EVAL_161;
  wire  _EVAL_474;
  wire  _EVAL_407;
  wire  _EVAL_117;
  wire  _EVAL_251;
  wire  _EVAL_62;
  wire  _EVAL_640;
  wire  _EVAL_537;
  wire  _EVAL_303;
  wire  _EVAL_149;
  wire  _EVAL_402;
  wire  _EVAL_482;
  wire  _EVAL_371;
  wire  _EVAL_135;
  wire  _EVAL_461;
  wire  _EVAL_124;
  wire  _EVAL_449;
  wire  _EVAL_508;
  wire  _EVAL_605;
  wire  _EVAL_433;
  wire  _EVAL_524;
  wire  _EVAL_470;
  wire [7:0] _EVAL_410;
  wire [7:0] _EVAL_187;
  wire  _EVAL_84;
  wire  _EVAL_207;
  wire  _EVAL_241;
  wire  _EVAL_263;
  wire  _EVAL_229;
  wire  _EVAL_647;
  wire  _EVAL_452;
  wire  _EVAL_125;
  wire  _EVAL_239;
  wire  _EVAL_432;
  wire  _EVAL_66;
  wire  _EVAL_521;
  wire  _EVAL_412;
  wire  _EVAL_166;
  wire  _EVAL_64;
  wire  _EVAL_118;
  wire  _EVAL_306;
  wire  _EVAL_573;
  wire [7:0] _EVAL_82;
  wire [7:0] _EVAL_337;
  wire [7:0] _EVAL_367;
  wire [7:0] _EVAL_550;
  wire  _EVAL_513;
  wire  _EVAL_472;
  wire  _EVAL_526;
  wire  _EVAL_126;
  wire  _EVAL_119;
  wire  _EVAL_506;
  wire  _EVAL_238;
  wire  _EVAL_181;
  wire  _EVAL_349;
  wire [7:0] _EVAL_109;
  wire [7:0] _EVAL_288;
  wire  _EVAL_420;
  wire  _EVAL_220;
  wire  _EVAL_454;
  wire  _EVAL_73;
  wire [1:0] _EVAL_648;
  wire [1:0] _EVAL_338;
  wire [1:0] _EVAL_391;
  wire [1:0] _EVAL_652;
  wire  _EVAL_99;
  wire  _EVAL_274;
  wire [4:0] _EVAL_465;
  wire  _EVAL_230;
  wire  _EVAL_260;
  wire  _EVAL_643;
  wire  _EVAL_348;
  wire  _EVAL_463;
  wire [4:0] _EVAL_459;
  wire  _EVAL_534;
  wire  _EVAL_498;
  wire  _EVAL_372;
  wire [4:0] _EVAL_593;
  wire  _EVAL_252;
  wire  _EVAL_223;
  wire  _EVAL_63;
  wire  _EVAL_194;
  wire  _EVAL_576;
  wire  _EVAL_50;
  wire  _EVAL_598;
  wire  _EVAL_298;
  wire  _EVAL_217;
  wire [7:0] _EVAL_613;
  wire [7:0] _EVAL_301;
  wire [7:0] _EVAL_473;
  wire  _EVAL_137;
  wire  _EVAL_606;
  wire  _EVAL_645;
  wire  _EVAL_554;
  wire  _EVAL_397;
  wire  _EVAL_385;
  wire  _EVAL_497;
  wire  _EVAL_563;
  wire  _EVAL_488;
  wire  _EVAL_419;
  wire  _EVAL_396;
  wire  _EVAL_171;
  wire  _EVAL_228;
  wire  _EVAL_49;
  wire  _EVAL_395;
  wire  _EVAL_344;
  wire  _EVAL_203;
  wire  _EVAL_414;
  wire  _EVAL_72;
  wire  _EVAL_495;
  wire  _EVAL_332;
  wire [7:0] _EVAL_322;
  wire  _EVAL_65;
  wire  _EVAL_35;
  wire  _EVAL_518;
  wire  _EVAL_244;
  wire  _EVAL_530;
  wire  _EVAL_110;
  wire  _EVAL_108;
  wire  _EVAL_311;
  wire  _EVAL_287;
  wire  _EVAL_202;
  wire  _EVAL_269;
  wire  _EVAL_293;
  wire [4:0] _EVAL_335;
  wire  _EVAL_471;
  wire  _EVAL_558;
  wire  _EVAL_639;
  wire  _EVAL_100;
  wire  _EVAL_541;
  wire  _EVAL_222;
  wire  _EVAL_37;
  wire  _EVAL_44;
  wire [4:0] _EVAL_416;
  wire  _EVAL_435;
  wire  _EVAL_430;
  wire  _EVAL_641;
  wire  _EVAL_36;
  wire  _EVAL_151;
  wire  _EVAL_485;
  wire  _EVAL_254;
  wire  _EVAL_167;
  wire  _EVAL_122;
  wire  _EVAL_242;
  wire  _EVAL_615;
  wire  _EVAL_619;
  wire  _EVAL_308;
  wire  _EVAL_620;
  wire  _EVAL_363;
  wire  _EVAL_92;
  wire  _EVAL_186;
  wire  _EVAL_246;
  wire  _EVAL_389;
  wire  _EVAL_386;
  wire [31:0] _EVAL_339;
  wire  _EVAL_597;
  wire  _EVAL_286;
  wire  _EVAL_462;
  wire  _EVAL_347;
  wire  _EVAL_377;
  wire  _EVAL_329;
  wire  _EVAL_314;
  wire  _EVAL_569;
  wire  _EVAL_48;
  wire  _EVAL_156;
  wire  _EVAL_594;
  wire  _EVAL_627;
  wire  _EVAL_59;
  wire  _EVAL_231;
  wire  _EVAL_496;
  wire  _EVAL_67;
  wire  _EVAL_34;
  wire  _EVAL_225;
  wire  _EVAL_259;
  wire  _EVAL_95;
  wire  _EVAL_129;
  wire  _EVAL_580;
  wire  _EVAL_175;
  wire  _EVAL_466;
  wire  _EVAL_281;
  wire  _EVAL_561;
  wire  _EVAL_302;
  wire  _EVAL_144;
  wire  _EVAL_379;
  wire  _EVAL_212;
  wire  _EVAL_88;
  wire  _EVAL_448;
  wire  _EVAL_568;
  wire  _EVAL_39;
  wire  _EVAL_360;
  wire  _EVAL_631;
  wire  _EVAL_289;
  wire  _EVAL_564;
  wire  _EVAL_630;
  wire  _EVAL_240;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_139;
  wire  _EVAL_350;
  wire  _EVAL_617;
  wire  _EVAL_165;
  wire  _EVAL_280;
  wire  _EVAL_163;
  wire  _EVAL_98;
  wire  _EVAL_327;
  wire  _EVAL_635;
  wire  _EVAL_632;
  wire  _EVAL_304;
  wire  _EVAL_323;
  wire  _EVAL_103;
  wire  _EVAL_450;
  wire  _EVAL_469;
  wire  _EVAL_132;
  wire  _EVAL_283;
  wire  _EVAL_527;
  wire  _EVAL_38;
  wire  _EVAL_515;
  wire  _EVAL_215;
  wire  _EVAL_138;
  wire  _EVAL_299;
  wire  _EVAL_256;
  wire  _EVAL_562;
  wire  _EVAL_189;
  wire  _EVAL_587;
  wire  _EVAL_622;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_317 = _EVAL_13 == 2'h0;
  assign _EVAL_423 = _EVAL_317 | _EVAL_22;
  assign _EVAL_403 = plusarg_reader_out == 32'h0;
  assign _EVAL_285 = _EVAL_33 ^ 32'h2000000;
  assign _EVAL_618 = {1'b0,$signed(_EVAL_285)};
  assign _EVAL_355 = $signed(_EVAL_618) & $signed(-33'sh10000);
  assign _EVAL_324 = $signed(_EVAL_355);
  assign _EVAL_626 = _EVAL_15 == _EVAL_500;
  assign _EVAL_625 = _EVAL_626 | _EVAL_22;
  assign _EVAL_522 = _EVAL_18 == 3'h0;
  assign _EVAL_431 = 23'hff << _EVAL_15;
  assign _EVAL_602 = _EVAL_431[7:0];
  assign _EVAL_586 = ~ _EVAL_602;
  assign _EVAL_509 = {{24'd0}, _EVAL_586};
  assign _EVAL_571 = _EVAL_26 ^ 32'h80000000;
  assign _EVAL_128 = {1'b0,$signed(_EVAL_571)};
  assign _EVAL_614 = $signed(_EVAL_128) & $signed(-33'sh20000);
  assign _EVAL_224 = $signed(_EVAL_614);
  assign _EVAL_234 = $signed(_EVAL_224) == $signed(33'sh0);
  assign _EVAL_595 = _EVAL_3 & _EVAL_509;
  assign _EVAL_358 = _EVAL_595 == 32'h0;
  assign _EVAL_579 = _EVAL_29[1:0];
  assign _EVAL_177 = 4'h1 << _EVAL_579;
  assign _EVAL_176 = _EVAL_177[2:0];
  assign _EVAL_455 = _EVAL_176 | 3'h1;
  assign _EVAL_261 = _EVAL_455[1];
  assign _EVAL_382 = _EVAL_566 != 8'h0;
  assign _EVAL_611 = _EVAL_382 == 1'h0;
  assign _EVAL_638 = _EVAL_33 ^ 32'h1800000;
  assign _EVAL_501 = {1'b0,$signed(_EVAL_638)};
  assign _EVAL_134 = $signed(_EVAL_501) & $signed(-33'sh8000);
  assign _EVAL_83 = $signed(_EVAL_134);
  assign _EVAL_152 = $signed(_EVAL_83) == $signed(33'sh0);
  assign _EVAL_172 = _EVAL_33 ^ 32'h1900000;
  assign _EVAL_233 = {1'b0,$signed(_EVAL_172)};
  assign _EVAL_142 = $signed(_EVAL_233) & $signed(-33'sh2000);
  assign _EVAL_475 = 23'hff << _EVAL_29;
  assign _EVAL_599 = _EVAL_475[7:0];
  assign _EVAL_291 = ~ _EVAL_599;
  assign _EVAL_604 = {{24'd0}, _EVAL_291};
  assign _EVAL_531 = _EVAL_33 & _EVAL_604;
  assign _EVAL_636 = _EVAL_10 == 3'h4;
  assign _EVAL_131 = _EVAL_24 & _EVAL_636;
  assign _EVAL_310 = _EVAL_30 & _EVAL_1;
  assign _EVAL_60 = _EVAL_296 == 5'h0;
  assign _EVAL_52 = _EVAL_310 & _EVAL_60;
  assign _EVAL_512 = _EVAL_25[2];
  assign _EVAL_284 = _EVAL_25[1];
  assign _EVAL_578 = _EVAL_284 == 1'h0;
  assign _EVAL_589 = _EVAL_512 & _EVAL_578;
  assign _EVAL_487 = _EVAL_52 & _EVAL_589;
  assign _EVAL_556 = 2'h1 << _EVAL_6;
  assign _EVAL_535 = _EVAL_487 ? _EVAL_556 : 2'h0;
  assign _EVAL_210 = _EVAL_535 | _EVAL_90;
  assign _EVAL_235 = _EVAL_210 >> _EVAL_11;
  assign _EVAL_102 = _EVAL_235[0];
  assign _EVAL_425 = _EVAL_102 | _EVAL_22;
  assign _EVAL_649 = _EVAL_425 == 1'h0;
  assign _EVAL_273 = _EVAL_13 <= 2'h2;
  assign _EVAL_464 = _EVAL_9 & _EVAL_24;
  assign _EVAL_191 = _EVAL_557 == 5'h0;
  assign _EVAL_86 = _EVAL_464 & _EVAL_191;
  assign _EVAL_384 = _EVAL_26 == _EVAL_159;
  assign _EVAL_219 = _EVAL_33[1];
  assign _EVAL_267 = _EVAL_219 == 1'h0;
  assign _EVAL_247 = {1'b0,$signed(_EVAL_26)};
  assign _EVAL_352 = $signed(_EVAL_247) & $signed(-33'sh1000);
  assign _EVAL_278 = $signed(_EVAL_352);
  assign _EVAL_603 = _EVAL_3 ^ 32'h3000;
  assign _EVAL_213 = {1'b0,$signed(_EVAL_603)};
  assign _EVAL_183 = $signed(_EVAL_213) & $signed(-33'sh1000);
  assign _EVAL_438 = $signed(_EVAL_183);
  assign _EVAL_440 = $signed(_EVAL_438) == $signed(33'sh0);
  assign _EVAL_443 = _EVAL_12 == 3'h2;
  assign _EVAL_133 = _EVAL_31 & _EVAL_443;
  assign _EVAL_272 = 3'h1 <= _EVAL_21;
  assign _EVAL_282 = _EVAL_26 ^ 32'h1900000;
  assign _EVAL_195 = {1'b0,$signed(_EVAL_282)};
  assign _EVAL_650 = $signed(_EVAL_195) & $signed(-33'sh2000);
  assign _EVAL_511 = $signed(_EVAL_650);
  assign _EVAL_519 = $signed(_EVAL_511) == $signed(33'sh0);
  assign _EVAL_612 = _EVAL_26 ^ 32'h40000000;
  assign _EVAL_517 = {1'b0,$signed(_EVAL_612)};
  assign _EVAL_262 = $signed(_EVAL_517) & $signed(-33'sh2000);
  assign _EVAL_76 = $signed(_EVAL_262);
  assign _EVAL_196 = $signed(_EVAL_76) == $signed(33'sh0);
  assign _EVAL_157 = _EVAL_519 | _EVAL_196;
  assign _EVAL_570 = _EVAL_21 == 3'h0;
  assign _EVAL_258 = _EVAL_570 | _EVAL_272;
  assign _EVAL_392 = _EVAL_455[0];
  assign _EVAL_114 = _EVAL_33[2];
  assign _EVAL_184 = _EVAL_114 == 1'h0;
  assign _EVAL_375 = _EVAL_184 & _EVAL_267;
  assign _EVAL_583 = _EVAL_33[0];
  assign _EVAL_479 = _EVAL_583 == 1'h0;
  assign _EVAL_146 = _EVAL_375 & _EVAL_479;
  assign _EVAL_504 = _EVAL_392 & _EVAL_146;
  assign _EVAL_387 = _EVAL_29 == _EVAL_180;
  assign _EVAL_232 = _EVAL_21 == _EVAL_80;
  assign _EVAL_394 = _EVAL_232 | _EVAL_22;
  assign _EVAL_476 = _EVAL_394 == 1'h0;
  assign _EVAL_226 = 4'h6 == _EVAL_15;
  assign _EVAL_365 = _EVAL_19 == _EVAL_277;
  assign _EVAL_628 = _EVAL_365 | _EVAL_22;
  assign _EVAL_484 = _EVAL_628 == 1'h0;
  assign _EVAL_275 = _EVAL_3 ^ 32'hc000000;
  assign _EVAL_572 = {1'b0,$signed(_EVAL_275)};
  assign _EVAL_155 = $signed(_EVAL_572) & $signed(-33'sh4000000);
  assign _EVAL_140 = $signed(_EVAL_155);
  assign _EVAL_533 = ~ _EVAL_28;
  assign _EVAL_75 = _EVAL_3 ^ 32'h1900000;
  assign _EVAL_354 = {1'b0,$signed(_EVAL_75)};
  assign _EVAL_491 = $signed(_EVAL_354) & $signed(-33'sh2000);
  assign _EVAL_477 = $signed(_EVAL_491);
  assign _EVAL_441 = _EVAL_90 >> _EVAL_6;
  assign _EVAL_153 = _EVAL_441[0];
  assign _EVAL_71 = _EVAL_153 == 1'h0;
  assign _EVAL_574 = _EVAL_71 | _EVAL_22;
  assign _EVAL_208 = _EVAL_574 == 1'h0;
  assign _EVAL_444 = {1'b0,$signed(_EVAL_3)};
  assign _EVAL_601 = $signed(_EVAL_444) & $signed(-33'sh1000);
  assign _EVAL_245 = $signed(_EVAL_601);
  assign _EVAL_434 = _EVAL_157 | _EVAL_234;
  assign _EVAL_345 = _EVAL_26 ^ 32'h3000;
  assign _EVAL_320 = {1'b0,$signed(_EVAL_345)};
  assign _EVAL_591 = $signed(_EVAL_320) & $signed(-33'sh1000);
  assign _EVAL_199 = $signed(_EVAL_591);
  assign _EVAL_150 = $signed(_EVAL_199) == $signed(33'sh0);
  assign _EVAL_359 = _EVAL_434 | _EVAL_150;
  assign _EVAL_106 = _EVAL_26 ^ 32'hc000000;
  assign _EVAL_417 = {1'b0,$signed(_EVAL_106)};
  assign _EVAL_268 = $signed(_EVAL_417) & $signed(-33'sh4000000);
  assign _EVAL_427 = $signed(_EVAL_268);
  assign _EVAL_182 = $signed(_EVAL_427) == $signed(33'sh0);
  assign _EVAL_369 = _EVAL_359 | _EVAL_182;
  assign _EVAL_353 = _EVAL_26 ^ 32'h2000000;
  assign _EVAL_53 = {1'b0,$signed(_EVAL_353)};
  assign _EVAL_383 = $signed(_EVAL_53) & $signed(-33'sh10000);
  assign _EVAL_115 = $signed(_EVAL_383);
  assign _EVAL_46 = $signed(_EVAL_115) == $signed(33'sh0);
  assign _EVAL_577 = _EVAL_369 | _EVAL_46;
  assign _EVAL_581 = $signed(_EVAL_278) == $signed(33'sh0);
  assign _EVAL_373 = _EVAL_577 | _EVAL_581;
  assign _EVAL_316 = _EVAL_26 ^ 32'h1800000;
  assign _EVAL_116 = {1'b0,$signed(_EVAL_316)};
  assign _EVAL_460 = $signed(_EVAL_116) & $signed(-33'sh8000);
  assign _EVAL_85 = $signed(_EVAL_460);
  assign _EVAL_540 = $signed(_EVAL_85) == $signed(33'sh0);
  assign _EVAL_147 = _EVAL_373 | _EVAL_540;
  assign _EVAL_592 = _EVAL_26 ^ 32'h4000;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_592)};
  assign _EVAL_607 = $signed(_EVAL_113) & $signed(-33'sh1000);
  assign _EVAL_309 = $signed(_EVAL_607);
  assign _EVAL_294 = $signed(_EVAL_309) == $signed(33'sh0);
  assign _EVAL_388 = _EVAL_147 | _EVAL_294;
  assign _EVAL_158 = _EVAL_26 ^ 32'h20000000;
  assign _EVAL_209 = {1'b0,$signed(_EVAL_158)};
  assign _EVAL_483 = $signed(_EVAL_209) & $signed(-33'sh2000);
  assign _EVAL_279 = $signed(_EVAL_483);
  assign _EVAL_582 = $signed(_EVAL_279) == $signed(33'sh0);
  assign _EVAL_429 = _EVAL_388 | _EVAL_582;
  assign _EVAL_276 = _EVAL_429 | _EVAL_22;
  assign _EVAL_585 = _EVAL_14 >= 4'h3;
  assign _EVAL_205 = _EVAL_29 >= 4'h3;
  assign _EVAL_162 = _EVAL_455[2];
  assign _EVAL_445 = _EVAL_162 & _EVAL_114;
  assign _EVAL_206 = _EVAL_205 | _EVAL_445;
  assign _EVAL_154 = _EVAL_114 & _EVAL_267;
  assign _EVAL_421 = _EVAL_261 & _EVAL_154;
  assign _EVAL_178 = _EVAL_206 | _EVAL_421;
  assign _EVAL_536 = _EVAL_25 <= 3'h6;
  assign _EVAL_346 = _EVAL_536 | _EVAL_22;
  assign _EVAL_218 = _EVAL_346 == 1'h0;
  assign _EVAL_584 = $signed(_EVAL_477) == $signed(33'sh0);
  assign _EVAL_493 = _EVAL_3 ^ 32'h40000000;
  assign _EVAL_494 = {1'b0,$signed(_EVAL_493)};
  assign _EVAL_104 = $signed(_EVAL_494) & $signed(-33'sh2000);
  assign _EVAL_610 = $signed(_EVAL_104);
  assign _EVAL_143 = $signed(_EVAL_610) == $signed(33'sh0);
  assign _EVAL_41 = _EVAL_584 | _EVAL_143;
  assign _EVAL_343 = _EVAL_3 ^ 32'h80000000;
  assign _EVAL_188 = {1'b0,$signed(_EVAL_343)};
  assign _EVAL_553 = $signed(_EVAL_188) & $signed(-33'sh20000);
  assign _EVAL_596 = $signed(_EVAL_553);
  assign _EVAL_404 = $signed(_EVAL_596) == $signed(33'sh0);
  assign _EVAL_170 = _EVAL_41 | _EVAL_404;
  assign _EVAL_313 = _EVAL_170 | _EVAL_440;
  assign _EVAL_331 = $signed(_EVAL_140) == $signed(33'sh0);
  assign _EVAL_333 = _EVAL_313 | _EVAL_331;
  assign _EVAL_399 = _EVAL_3 ^ 32'h2000000;
  assign _EVAL_528 = {1'b0,$signed(_EVAL_399)};
  assign _EVAL_319 = $signed(_EVAL_528) & $signed(-33'sh10000);
  assign _EVAL_575 = $signed(_EVAL_319);
  assign _EVAL_211 = $signed(_EVAL_575) == $signed(33'sh0);
  assign _EVAL_499 = _EVAL_333 | _EVAL_211;
  assign _EVAL_393 = $signed(_EVAL_245) == $signed(33'sh0);
  assign _EVAL_400 = _EVAL_499 | _EVAL_393;
  assign _EVAL_190 = _EVAL_3 ^ 32'h1800000;
  assign _EVAL_600 = {1'b0,$signed(_EVAL_190)};
  assign _EVAL_468 = $signed(_EVAL_600) & $signed(-33'sh8000);
  assign _EVAL_486 = $signed(_EVAL_468);
  assign _EVAL_503 = $signed(_EVAL_486) == $signed(33'sh0);
  assign _EVAL_56 = _EVAL_400 | _EVAL_503;
  assign _EVAL_264 = _EVAL_3 ^ 32'h4000;
  assign _EVAL_237 = {1'b0,$signed(_EVAL_264)};
  assign _EVAL_148 = $signed(_EVAL_237) & $signed(-33'sh1000);
  assign _EVAL_192 = $signed(_EVAL_148);
  assign _EVAL_633 = $signed(_EVAL_192) == $signed(33'sh0);
  assign _EVAL_651 = _EVAL_56 | _EVAL_633;
  assign _EVAL_368 = _EVAL_3 ^ 32'h20000000;
  assign _EVAL_588 = {1'b0,$signed(_EVAL_368)};
  assign _EVAL_130 = $signed(_EVAL_588) & $signed(-33'sh2000);
  assign _EVAL_89 = $signed(_EVAL_130);
  assign _EVAL_70 = $signed(_EVAL_89) == $signed(33'sh0);
  assign _EVAL_629 = _EVAL_651 | _EVAL_70;
  assign _EVAL_250 = _EVAL_243 == 5'h0;
  assign _EVAL_79 = _EVAL_10[2];
  assign _EVAL_415 = _EVAL_79 == 1'h0;
  assign _EVAL_168 = _EVAL_291[7:3];
  assign _EVAL_545 = _EVAL_243 - 5'h1;
  assign _EVAL_424 = _EVAL_27 <= 2'h2;
  assign _EVAL_334 = _EVAL_29 <= 4'h6;
  assign _EVAL_520 = $signed(_EVAL_142);
  assign _EVAL_458 = $signed(_EVAL_520) == $signed(33'sh0);
  assign _EVAL_380 = _EVAL_33 ^ 32'h40000000;
  assign _EVAL_121 = {1'b0,$signed(_EVAL_380)};
  assign _EVAL_321 = $signed(_EVAL_121) & $signed(-33'sh2000);
  assign _EVAL_179 = $signed(_EVAL_321);
  assign _EVAL_40 = $signed(_EVAL_179) == $signed(33'sh0);
  assign _EVAL_127 = _EVAL_458 | _EVAL_40;
  assign _EVAL_318 = _EVAL_33 ^ 32'h80000000;
  assign _EVAL_221 = {1'b0,$signed(_EVAL_318)};
  assign _EVAL_336 = $signed(_EVAL_221) & $signed(-33'sh20000);
  assign _EVAL_330 = $signed(_EVAL_336);
  assign _EVAL_305 = $signed(_EVAL_330) == $signed(33'sh0);
  assign _EVAL_559 = _EVAL_127 | _EVAL_305;
  assign _EVAL_467 = _EVAL_33 ^ 32'hc000000;
  assign _EVAL_81 = {1'b0,$signed(_EVAL_467)};
  assign _EVAL_169 = $signed(_EVAL_81) & $signed(-33'sh4000000);
  assign _EVAL_546 = $signed(_EVAL_169);
  assign _EVAL_255 = $signed(_EVAL_546) == $signed(33'sh0);
  assign _EVAL_271 = _EVAL_559 | _EVAL_255;
  assign _EVAL_547 = $signed(_EVAL_324) == $signed(33'sh0);
  assign _EVAL_544 = _EVAL_271 | _EVAL_547;
  assign _EVAL_481 = {1'b0,$signed(_EVAL_33)};
  assign _EVAL_634 = $signed(_EVAL_481) & $signed(-33'sh5000);
  assign _EVAL_510 = $signed(_EVAL_634);
  assign _EVAL_529 = $signed(_EVAL_510) == $signed(33'sh0);
  assign _EVAL_292 = _EVAL_544 | _EVAL_529;
  assign _EVAL_107 = _EVAL_292 | _EVAL_152;
  assign _EVAL_307 = _EVAL_33 ^ 32'h20000000;
  assign _EVAL_560 = {1'b0,$signed(_EVAL_307)};
  assign _EVAL_428 = $signed(_EVAL_560) & $signed(-33'sh2000);
  assign _EVAL_489 = $signed(_EVAL_428);
  assign _EVAL_43 = $signed(_EVAL_489) == $signed(33'sh0);
  assign _EVAL_236 = _EVAL_107 | _EVAL_43;
  assign _EVAL_418 = _EVAL_334 & _EVAL_236;
  assign _EVAL_653 = _EVAL_29 <= 4'h8;
  assign _EVAL_370 = _EVAL_33 ^ 32'h3000;
  assign _EVAL_357 = {1'b0,$signed(_EVAL_370)};
  assign _EVAL_42 = $signed(_EVAL_357) & $signed(-33'sh1000);
  assign _EVAL_68 = $signed(_EVAL_42);
  assign _EVAL_91 = $signed(_EVAL_68) == $signed(33'sh0);
  assign _EVAL_624 = _EVAL_653 & _EVAL_91;
  assign _EVAL_364 = _EVAL_418 | _EVAL_624;
  assign _EVAL_442 = _EVAL_10 == 3'h7;
  assign _EVAL_381 = 4'h6 == _EVAL_29;
  assign _EVAL_516 = _EVAL_570 ? _EVAL_381 : 1'h0;
  assign _EVAL_340 = _EVAL_516 | _EVAL_22;
  assign _EVAL_93 = _EVAL_174 == 5'h0;
  assign _EVAL_525 = _EVAL_93 == 1'h0;
  assign _EVAL_621 = _EVAL_1 & _EVAL_525;
  assign _EVAL_300 = _EVAL_23 == 1'h0;
  assign _EVAL_97 = _EVAL_25[0];
  assign _EVAL_351 = 23'hff << _EVAL_14;
  assign _EVAL_376 = _EVAL_351[7:0];
  assign _EVAL_457 = ~ _EVAL_376;
  assign _EVAL_61 = _EVAL_457[7:3];
  assign _EVAL_401 = _EVAL_296 - 5'h1;
  assign _EVAL_362 = _EVAL_358 | _EVAL_22;
  assign _EVAL_590 = _EVAL_7 == 1'h0;
  assign _EVAL_502 = _EVAL_590 | _EVAL_22;
  assign _EVAL_101 = _EVAL_566 >> _EVAL_21;
  assign _EVAL_216 = _EVAL_101[0];
  assign _EVAL_405 = _EVAL_216 == 1'h0;
  assign _EVAL_136 = _EVAL_405 | _EVAL_22;
  assign _EVAL_57 = _EVAL_136 == 1'h0;
  assign _EVAL_378 = _EVAL_154 & _EVAL_583;
  assign _EVAL_266 = _EVAL_392 & _EVAL_378;
  assign _EVAL_120 = _EVAL_12 == 3'h7;
  assign _EVAL_96 = _EVAL_387 | _EVAL_22;
  assign _EVAL_341 = _EVAL_96 == 1'h0;
  assign _EVAL_123 = 3'h1 <= _EVAL_19;
  assign _EVAL_514 = _EVAL_164 == 5'h0;
  assign _EVAL_426 = _EVAL_611 | _EVAL_403;
  assign _EVAL_198 = _EVAL_590 | _EVAL_2;
  assign _EVAL_637 = _EVAL_7 == _EVAL_456;
  assign _EVAL_422 = _EVAL_637 | _EVAL_22;
  assign _EVAL_145 = _EVAL_422 == 1'h0;
  assign _EVAL_549 = _EVAL_13 != 2'h2;
  assign _EVAL_608 = _EVAL_19 == 3'h0;
  assign _EVAL_366 = _EVAL_608 | _EVAL_123;
  assign _EVAL_204 = _EVAL_32 == _EVAL_552;
  assign _EVAL_409 = _EVAL_26 & 32'h3f;
  assign _EVAL_265 = _EVAL_409 == 32'h0;
  assign _EVAL_543 = _EVAL_29 <= 4'h2;
  assign _EVAL_248 = _EVAL_10 == 3'h2;
  assign _EVAL_200 = _EVAL_458 | _EVAL_91;
  assign _EVAL_451 = _EVAL_200 | _EVAL_255;
  assign _EVAL_413 = _EVAL_451 | _EVAL_547;
  assign _EVAL_328 = _EVAL_413 | _EVAL_529;
  assign _EVAL_58 = _EVAL_328 | _EVAL_152;
  assign _EVAL_173 = _EVAL_58 | _EVAL_43;
  assign _EVAL_646 = _EVAL_543 & _EVAL_173;
  assign _EVAL_408 = _EVAL_646 | _EVAL_22;
  assign _EVAL_249 = _EVAL_408 == 1'h0;
  assign _EVAL_523 = _EVAL_178 | _EVAL_266;
  assign _EVAL_623 = _EVAL_164 - 5'h1;
  assign _EVAL_436 = _EVAL_0 <= 3'h2;
  assign _EVAL_214 = _EVAL_436 | _EVAL_22;
  assign _EVAL_447 = _EVAL_214 == 1'h0;
  assign _EVAL_227 = _EVAL_608 ? _EVAL_226 : 1'h0;
  assign _EVAL_78 = _EVAL_227 | _EVAL_22;
  assign _EVAL_297 = _EVAL_78 == 1'h0;
  assign _EVAL_295 = _EVAL_10 == 3'h5;
  assign _EVAL_87 = _EVAL_629 | _EVAL_22;
  assign _EVAL_642 = _EVAL_87 == 1'h0;
  assign _EVAL_54 = _EVAL_16 & _EVAL_20;
  assign _EVAL_532 = _EVAL_364 | _EVAL_22;
  assign _EVAL_555 = _EVAL_154 & _EVAL_479;
  assign _EVAL_342 = _EVAL_392 & _EVAL_555;
  assign _EVAL_160 = _EVAL_178 | _EVAL_342;
  assign _EVAL_45 = _EVAL_12 == 3'h0;
  assign _EVAL_565 = _EVAL_31 & _EVAL_45;
  assign _EVAL_548 = _EVAL_366 | _EVAL_22;
  assign _EVAL_312 = _EVAL_90 | _EVAL_535;
  assign _EVAL_505 = _EVAL_362 == 1'h0;
  assign _EVAL_315 = _EVAL_114 & _EVAL_219;
  assign _EVAL_507 = _EVAL_261 & _EVAL_315;
  assign _EVAL_374 = _EVAL_206 | _EVAL_507;
  assign _EVAL_361 = _EVAL_315 & _EVAL_583;
  assign _EVAL_161 = _EVAL_392 & _EVAL_361;
  assign _EVAL_474 = _EVAL_374 | _EVAL_161;
  assign _EVAL_407 = _EVAL_315 & _EVAL_479;
  assign _EVAL_117 = _EVAL_392 & _EVAL_407;
  assign _EVAL_251 = _EVAL_374 | _EVAL_117;
  assign _EVAL_62 = _EVAL_162 & _EVAL_184;
  assign _EVAL_640 = _EVAL_205 | _EVAL_62;
  assign _EVAL_537 = _EVAL_184 & _EVAL_219;
  assign _EVAL_303 = _EVAL_261 & _EVAL_537;
  assign _EVAL_149 = _EVAL_640 | _EVAL_303;
  assign _EVAL_402 = _EVAL_537 & _EVAL_583;
  assign _EVAL_482 = _EVAL_392 & _EVAL_402;
  assign _EVAL_371 = _EVAL_149 | _EVAL_482;
  assign _EVAL_135 = _EVAL_537 & _EVAL_479;
  assign _EVAL_461 = _EVAL_392 & _EVAL_135;
  assign _EVAL_124 = _EVAL_149 | _EVAL_461;
  assign _EVAL_449 = _EVAL_261 & _EVAL_375;
  assign _EVAL_508 = _EVAL_640 | _EVAL_449;
  assign _EVAL_605 = _EVAL_375 & _EVAL_583;
  assign _EVAL_433 = _EVAL_392 & _EVAL_605;
  assign _EVAL_524 = _EVAL_508 | _EVAL_433;
  assign _EVAL_470 = _EVAL_508 | _EVAL_504;
  assign _EVAL_410 = {_EVAL_474,_EVAL_251,_EVAL_523,_EVAL_160,_EVAL_371,_EVAL_124,_EVAL_524,_EVAL_470};
  assign _EVAL_187 = ~ _EVAL_410;
  assign _EVAL_84 = _EVAL_6 == _EVAL_437;
  assign _EVAL_207 = _EVAL_84 | _EVAL_22;
  assign _EVAL_241 = _EVAL_207 == 1'h0;
  assign _EVAL_263 = _EVAL_25 == 3'h2;
  assign _EVAL_229 = _EVAL_624 | _EVAL_22;
  assign _EVAL_647 = _EVAL_549 | _EVAL_22;
  assign _EVAL_452 = _EVAL_111 == 5'h0;
  assign _EVAL_125 = _EVAL_452 == 1'h0;
  assign _EVAL_239 = _EVAL_18 == _EVAL_478;
  assign _EVAL_432 = _EVAL_334 & _EVAL_305;
  assign _EVAL_66 = _EVAL_432 | _EVAL_22;
  assign _EVAL_521 = _EVAL_66 == 1'h0;
  assign _EVAL_412 = _EVAL_15 >= 4'h3;
  assign _EVAL_166 = _EVAL_205 | _EVAL_22;
  assign _EVAL_64 = _EVAL_8 & _EVAL;
  assign _EVAL_118 = _EVAL_10 == _EVAL_644;
  assign _EVAL_306 = _EVAL_118 | _EVAL_22;
  assign _EVAL_573 = _EVAL & _EVAL_125;
  assign _EVAL_82 = 8'h1 << _EVAL_21;
  assign _EVAL_337 = _EVAL_86 ? _EVAL_82 : 8'h0;
  assign _EVAL_367 = _EVAL_337 | _EVAL_566;
  assign _EVAL_550 = _EVAL_367 >> _EVAL_32;
  assign _EVAL_513 = _EVAL_550[0];
  assign _EVAL_472 = _EVAL_2 == 1'h0;
  assign _EVAL_526 = _EVAL_472 | _EVAL_22;
  assign _EVAL_126 = _EVAL_24 & _EVAL_295;
  assign _EVAL_119 = 3'h1 <= _EVAL_32;
  assign _EVAL_506 = _EVAL_310 & _EVAL_514;
  assign _EVAL_238 = _EVAL_25 == 3'h6;
  assign _EVAL_181 = _EVAL_238 == 1'h0;
  assign _EVAL_349 = _EVAL_506 & _EVAL_181;
  assign _EVAL_109 = 8'h1 << _EVAL_32;
  assign _EVAL_288 = _EVAL_349 ? _EVAL_109 : 8'h0;
  assign _EVAL_420 = _EVAL_337 != _EVAL_288;
  assign _EVAL_220 = _EVAL_15 <= 4'h6;
  assign _EVAL_454 = _EVAL_220 & _EVAL_404;
  assign _EVAL_73 = _EVAL_548 == 1'h0;
  assign _EVAL_648 = 2'h1 << _EVAL_11;
  assign _EVAL_338 = _EVAL_54 ? _EVAL_648 : 2'h0;
  assign _EVAL_391 = ~ _EVAL_338;
  assign _EVAL_652 = _EVAL_312 & _EVAL_391;
  assign _EVAL_99 = _EVAL_533 == 8'h0;
  assign _EVAL_274 = _EVAL_99 | _EVAL_22;
  assign _EVAL_465 = _EVAL_111 - 5'h1;
  assign _EVAL_230 = _EVAL_10 == 3'h0;
  assign _EVAL_260 = _EVAL_10 == 3'h6;
  assign _EVAL_643 = _EVAL_24 & _EVAL_260;
  assign _EVAL_348 = _EVAL_28 == _EVAL_410;
  assign _EVAL_463 = _EVAL_348 | _EVAL_22;
  assign _EVAL_459 = _EVAL_174 - 5'h1;
  assign _EVAL_534 = _EVAL_25 == 3'h5;
  assign _EVAL_498 = _EVAL_33 == _EVAL_446;
  assign _EVAL_372 = _EVAL_498 | _EVAL_22;
  assign _EVAL_593 = _EVAL_557 - 5'h1;
  assign _EVAL_252 = _EVAL_306 == 1'h0;
  assign _EVAL_223 = _EVAL_340 == 1'h0;
  assign _EVAL_63 = _EVAL_14 == _EVAL_253;
  assign _EVAL_194 = _EVAL_63 | _EVAL_22;
  assign _EVAL_576 = _EVAL_300 | _EVAL_22;
  assign _EVAL_50 = _EVAL_576 == 1'h0;
  assign _EVAL_598 = _EVAL_32 == 3'h0;
  assign _EVAL_298 = _EVAL_25 == 3'h0;
  assign _EVAL_217 = _EVAL_239 | _EVAL_22;
  assign _EVAL_613 = _EVAL_566 | _EVAL_337;
  assign _EVAL_301 = ~ _EVAL_288;
  assign _EVAL_473 = _EVAL_613 & _EVAL_301;
  assign _EVAL_137 = _EVAL_502 == 1'h0;
  assign _EVAL_606 = _EVAL_10 == 3'h1;
  assign _EVAL_645 = _EVAL_24 & _EVAL_606;
  assign _EVAL_554 = _EVAL_27 == _EVAL_390;
  assign _EVAL_397 = _EVAL_554 | _EVAL_22;
  assign _EVAL_385 = _EVAL_273 | _EVAL_22;
  assign _EVAL_497 = _EVAL_385 == 1'h0;
  assign _EVAL_563 = _EVAL_424 | _EVAL_22;
  assign _EVAL_488 = _EVAL_12 == 3'h6;
  assign _EVAL_419 = _EVAL_250 == 1'h0;
  assign _EVAL_396 = _EVAL_24 & _EVAL_419;
  assign _EVAL_171 = _EVAL_531 == 32'h0;
  assign _EVAL_228 = _EVAL_171 | _EVAL_22;
  assign _EVAL_49 = _EVAL_406 == 5'h0;
  assign _EVAL_395 = _EVAL_49 == 1'h0;
  assign _EVAL_344 = _EVAL_31 & _EVAL_395;
  assign _EVAL_203 = _EVAL_513 | _EVAL_22;
  assign _EVAL_414 = _EVAL_337 != 8'h0;
  assign _EVAL_72 = _EVAL_414 == 1'h0;
  assign _EVAL_495 = _EVAL_420 | _EVAL_72;
  assign _EVAL_332 = _EVAL_495 | _EVAL_22;
  assign _EVAL_322 = _EVAL_28 & _EVAL_187;
  assign _EVAL_65 = _EVAL_322 == 8'h0;
  assign _EVAL_35 = _EVAL_229 == 1'h0;
  assign _EVAL_518 = _EVAL_25 == _EVAL_74;
  assign _EVAL_244 = _EVAL_518 | _EVAL_22;
  assign _EVAL_530 = _EVAL_244 == 1'h0;
  assign _EVAL_110 = _EVAL_198 | _EVAL_22;
  assign _EVAL_108 = _EVAL_110 == 1'h0;
  assign _EVAL_311 = _EVAL_0 <= 3'h5;
  assign _EVAL_287 = _EVAL_412 | _EVAL_22;
  assign _EVAL_202 = _EVAL_287 == 1'h0;
  assign _EVAL_269 = _EVAL_17 == 1'h0;
  assign _EVAL_293 = _EVAL_647 == 1'h0;
  assign _EVAL_335 = _EVAL_406 - 5'h1;
  assign _EVAL_471 = _EVAL_0 == _EVAL_201;
  assign _EVAL_558 = _EVAL_471 | _EVAL_22;
  assign _EVAL_639 = _EVAL_12 == 3'h1;
  assign _EVAL_100 = _EVAL_31 & _EVAL_639;
  assign _EVAL_541 = _EVAL_18 != 3'h0;
  assign _EVAL_222 = _EVAL_541 | _EVAL_22;
  assign _EVAL_37 = _EVAL_18 <= 3'h3;
  assign _EVAL_44 = _EVAL_12[0];
  assign _EVAL_416 = _EVAL_586[7:3];
  assign _EVAL_435 = _EVAL_258 | _EVAL_22;
  assign _EVAL_430 = _EVAL_384 | _EVAL_22;
  assign _EVAL_641 = _EVAL_430 == 1'h0;
  assign _EVAL_36 = _EVAL_24 & _EVAL_248;
  assign _EVAL_151 = _EVAL_5 & _EVAL_31;
  assign _EVAL_485 = _EVAL_463 == 1'h0;
  assign _EVAL_254 = _EVAL_492 < plusarg_reader_out;
  assign _EVAL_167 = _EVAL_426 | _EVAL_254;
  assign _EVAL_122 = _EVAL_532 == 1'h0;
  assign _EVAL_242 = _EVAL_18 <= 3'h4;
  assign _EVAL_615 = _EVAL_526 == 1'h0;
  assign _EVAL_619 = _EVAL_12 == 3'h4;
  assign _EVAL_308 = _EVAL_31 & _EVAL_619;
  assign _EVAL_620 = _EVAL_24 & _EVAL_442;
  assign _EVAL_363 = _EVAL_585 | _EVAL_22;
  assign _EVAL_92 = _EVAL_217 == 1'h0;
  assign _EVAL_186 = _EVAL_454 | _EVAL_22;
  assign _EVAL_246 = _EVAL_186 == 1'h0;
  assign _EVAL_389 = _EVAL_558 == 1'h0;
  assign _EVAL_386 = _EVAL_464 | _EVAL_310;
  assign _EVAL_339 = _EVAL_492 + 32'h1;
  assign _EVAL_597 = _EVAL_37 | _EVAL_22;
  assign _EVAL_286 = _EVAL_65 | _EVAL_22;
  assign _EVAL_462 = _EVAL_1 & _EVAL_534;
  assign _EVAL_347 = _EVAL_0 == 3'h0;
  assign _EVAL_377 = _EVAL_347 | _EVAL_22;
  assign _EVAL_329 = _EVAL_151 & _EVAL_49;
  assign _EVAL_314 = _EVAL_3 == _EVAL_551;
  assign _EVAL_569 = _EVAL_242 | _EVAL_22;
  assign _EVAL_48 = _EVAL_311 | _EVAL_22;
  assign _EVAL_156 = _EVAL_18 <= 3'h2;
  assign _EVAL_594 = _EVAL_156 | _EVAL_22;
  assign _EVAL_627 = _EVAL_594 == 1'h0;
  assign _EVAL_59 = _EVAL_25 == 3'h4;
  assign _EVAL_231 = _EVAL_522 | _EVAL_22;
  assign _EVAL_496 = _EVAL_598 | _EVAL_119;
  assign _EVAL_67 = _EVAL_496 | _EVAL_22;
  assign _EVAL_34 = _EVAL_269 | _EVAL_22;
  assign _EVAL_225 = _EVAL_597 == 1'h0;
  assign _EVAL_259 = _EVAL_274 == 1'h0;
  assign _EVAL_95 = _EVAL_423 == 1'h0;
  assign _EVAL_129 = _EVAL_276 == 1'h0;
  assign _EVAL_580 = _EVAL_363 == 1'h0;
  assign _EVAL_175 = _EVAL_1 & _EVAL_263;
  assign _EVAL_466 = _EVAL_48 == 1'h0;
  assign _EVAL_281 = _EVAL_310 & _EVAL_93;
  assign _EVAL_561 = _EVAL_13 == _EVAL_567;
  assign _EVAL_302 = _EVAL_12 == _EVAL_356;
  assign _EVAL_144 = _EVAL_302 | _EVAL_22;
  assign _EVAL_379 = _EVAL_464 & _EVAL_250;
  assign _EVAL_212 = _EVAL_561 | _EVAL_22;
  assign _EVAL_88 = _EVAL_212 == 1'h0;
  assign _EVAL_448 = _EVAL_31 & _EVAL_488;
  assign _EVAL_568 = _EVAL_563 == 1'h0;
  assign _EVAL_39 = _EVAL_265 | _EVAL_22;
  assign _EVAL_360 = _EVAL_39 == 1'h0;
  assign _EVAL_631 = _EVAL_25 == 3'h1;
  assign _EVAL_289 = _EVAL_1 & _EVAL_631;
  assign _EVAL_564 = _EVAL_144 == 1'h0;
  assign _EVAL_630 = _EVAL_397 == 1'h0;
  assign _EVAL_240 = _EVAL_1 & _EVAL_298;
  assign _EVAL_325 = _EVAL_204 | _EVAL_22;
  assign _EVAL_326 = _EVAL_325 == 1'h0;
  assign _EVAL_139 = _EVAL_228 == 1'h0;
  assign _EVAL_350 = _EVAL_31 & _EVAL_120;
  assign _EVAL_617 = _EVAL_1 & _EVAL_238;
  assign _EVAL_165 = _EVAL_569 == 1'h0;
  assign _EVAL_280 = _EVAL_167 | _EVAL_22;
  assign _EVAL_163 = _EVAL_280 == 1'h0;
  assign _EVAL_98 = _EVAL_1 & _EVAL_59;
  assign _EVAL_327 = _EVAL_34 == 1'h0;
  assign _EVAL_635 = _EVAL_332 == 1'h0;
  assign _EVAL_632 = _EVAL_24 & _EVAL_230;
  assign _EVAL_304 = _EVAL_231 == 1'h0;
  assign _EVAL_323 = _EVAL_314 | _EVAL_22;
  assign _EVAL_103 = _EVAL_323 == 1'h0;
  assign _EVAL_450 = _EVAL_372 == 1'h0;
  assign _EVAL_469 = _EVAL_10 == 3'h3;
  assign _EVAL_132 = _EVAL_67 == 1'h0;
  assign _EVAL_283 = _EVAL_203 == 1'h0;
  assign _EVAL_527 = _EVAL_625 == 1'h0;
  assign _EVAL_38 = _EVAL_12 == 3'h5;
  assign _EVAL_515 = _EVAL_31 & _EVAL_38;
  assign _EVAL_215 = _EVAL_286 == 1'h0;
  assign _EVAL_138 = _EVAL_222 == 1'h0;
  assign _EVAL_299 = _EVAL_166 == 1'h0;
  assign _EVAL_256 = _EVAL_435 == 1'h0;
  assign _EVAL_562 = _EVAL_24 & _EVAL_469;
  assign _EVAL_189 = _EVAL_64 & _EVAL_452;
  assign _EVAL_587 = _EVAL_377 == 1'h0;
  assign _EVAL_622 = _EVAL_194 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_74 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_80 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_90 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_111 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_159 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_164 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_174 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_180 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_201 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_243 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_253 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_277 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_296 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_356 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_390 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_406 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_437 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_446 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_456 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_478 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_492 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_500 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_551 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_552 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_557 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_566 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_567 = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_644 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_281) begin
      _EVAL_74 <= _EVAL_25;
    end
    if (_EVAL_379) begin
      _EVAL_80 <= _EVAL_21;
    end
    if (_EVAL_22) begin
      _EVAL_90 <= 2'h0;
    end else begin
      _EVAL_90 <= _EVAL_652;
    end
    if (_EVAL_22) begin
      _EVAL_111 <= 5'h0;
    end else begin
      if (_EVAL_64) begin
        if (_EVAL_452) begin
          _EVAL_111 <= 5'h0;
        end else begin
          _EVAL_111 <= _EVAL_465;
        end
      end
    end
    if (_EVAL_189) begin
      _EVAL_159 <= _EVAL_26;
    end
    if (_EVAL_22) begin
      _EVAL_164 <= 5'h0;
    end else begin
      if (_EVAL_310) begin
        if (_EVAL_514) begin
          if (_EVAL_97) begin
            _EVAL_164 <= _EVAL_61;
          end else begin
            _EVAL_164 <= 5'h0;
          end
        end else begin
          _EVAL_164 <= _EVAL_623;
        end
      end
    end
    if (_EVAL_22) begin
      _EVAL_174 <= 5'h0;
    end else begin
      if (_EVAL_310) begin
        if (_EVAL_93) begin
          if (_EVAL_97) begin
            _EVAL_174 <= _EVAL_61;
          end else begin
            _EVAL_174 <= 5'h0;
          end
        end else begin
          _EVAL_174 <= _EVAL_459;
        end
      end
    end
    if (_EVAL_379) begin
      _EVAL_180 <= _EVAL_29;
    end
    if (_EVAL_329) begin
      _EVAL_201 <= _EVAL_0;
    end
    if (_EVAL_22) begin
      _EVAL_243 <= 5'h0;
    end else begin
      if (_EVAL_464) begin
        if (_EVAL_250) begin
          if (_EVAL_415) begin
            _EVAL_243 <= _EVAL_168;
          end else begin
            _EVAL_243 <= 5'h0;
          end
        end else begin
          _EVAL_243 <= _EVAL_545;
        end
      end
    end
    if (_EVAL_281) begin
      _EVAL_253 <= _EVAL_14;
    end
    if (_EVAL_329) begin
      _EVAL_277 <= _EVAL_19;
    end
    if (_EVAL_22) begin
      _EVAL_296 <= 5'h0;
    end else begin
      if (_EVAL_310) begin
        if (_EVAL_60) begin
          if (_EVAL_97) begin
            _EVAL_296 <= _EVAL_61;
          end else begin
            _EVAL_296 <= 5'h0;
          end
        end else begin
          _EVAL_296 <= _EVAL_401;
        end
      end
    end
    if (_EVAL_329) begin
      _EVAL_356 <= _EVAL_12;
    end
    if (_EVAL_189) begin
      _EVAL_390 <= _EVAL_27;
    end
    if (_EVAL_22) begin
      _EVAL_406 <= 5'h0;
    end else begin
      if (_EVAL_151) begin
        if (_EVAL_49) begin
          if (_EVAL_44) begin
            _EVAL_406 <= _EVAL_416;
          end else begin
            _EVAL_406 <= 5'h0;
          end
        end else begin
          _EVAL_406 <= _EVAL_335;
        end
      end
    end
    if (_EVAL_281) begin
      _EVAL_437 <= _EVAL_6;
    end
    if (_EVAL_379) begin
      _EVAL_446 <= _EVAL_33;
    end
    if (_EVAL_281) begin
      _EVAL_456 <= _EVAL_7;
    end
    if (_EVAL_379) begin
      _EVAL_478 <= _EVAL_18;
    end
    if (_EVAL_22) begin
      _EVAL_492 <= 32'h0;
    end else begin
      if (_EVAL_386) begin
        _EVAL_492 <= 32'h0;
      end else begin
        _EVAL_492 <= _EVAL_339;
      end
    end
    if (_EVAL_329) begin
      _EVAL_500 <= _EVAL_15;
    end
    if (_EVAL_329) begin
      _EVAL_551 <= _EVAL_3;
    end
    if (_EVAL_281) begin
      _EVAL_552 <= _EVAL_32;
    end
    if (_EVAL_22) begin
      _EVAL_557 <= 5'h0;
    end else begin
      if (_EVAL_464) begin
        if (_EVAL_191) begin
          if (_EVAL_415) begin
            _EVAL_557 <= _EVAL_168;
          end else begin
            _EVAL_557 <= 5'h0;
          end
        end else begin
          _EVAL_557 <= _EVAL_593;
        end
      end
    end
    if (_EVAL_22) begin
      _EVAL_566 <= 8'h0;
    end else begin
      _EVAL_566 <= _EVAL_473;
    end
    if (_EVAL_281) begin
      _EVAL_567 <= _EVAL_13;
    end
    if (_EVAL_379) begin
      _EVAL_644 <= _EVAL_10;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d017517)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_497) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_630) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe61af5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cffb273)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_615) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_447) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae04e9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_630) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_615) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30691ca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e69098e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_466) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91e0c8ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2782f1c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f69a9ab1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a013b91d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_622) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dafd9e10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_521) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_521) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c528cf83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(823a6d6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b02c80a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a983ba8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecdab1a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e6a907d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_447) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab7c578e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b84aed4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcc29f2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(645da0f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_641) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e2eabb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfd14b4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc284e12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71bd8955)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_622) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_641) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8df1124d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_587) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8bd04d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84fd20ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c7c6eab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c1c228)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_450) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a58d5300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_587) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_615) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7b1b2ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e219aa61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_627) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c64ae498)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_635) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da2f4c2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7532678b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecb6cad8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_487 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc59bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_487 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f016d8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_649) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3010a7f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2953b19f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37e7e4d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_521) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f32202db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed59eaca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8fd5acd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_627) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380413a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f0a3c14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0603f7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_349 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_466) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(566caa74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_476) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_587) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38f5a261)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_580) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e92d26e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20c54025)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8bda9c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_497) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_627) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ccfcb60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3a2fa9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_530) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b411fa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de15b8ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(429f00ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d36751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1053c399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22255405)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee89fac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_527) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a09276)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11652404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab8bd231)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_450) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e35578fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8513397e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_635) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2052f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a03c2650)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff67a4dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(852a6132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b68677e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_389) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ba9f0b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(594c7403)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_476) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de3b787b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_627) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b82b34a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6400bcbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f289a5c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb0a5c66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f474571a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_527) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2b46703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48dce570)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816fffd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_447) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4d3274b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff063702)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a369a9d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_530) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da2207ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d07a441)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_568) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d7606d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_505) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8faf5748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caab3d31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf24ca05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_505) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_568) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_649) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12440d4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(317c2867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_389) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_521) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e011c662)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_349 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a14a0950)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f83619d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_615) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee740fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a7136f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_580) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab8586f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf6ef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1515d304)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_447) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_615) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b78eaf26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_466) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bee98561)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_587) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(663dfa05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dedc093)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d74e7e3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(481fc4e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_564) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5590195f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_617 & _EVAL_615) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c3dc008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb4e8d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcd3b06c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61b983ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa2207ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_615) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d45e1bb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8837af0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_587) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0c6cf7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8541bf76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(debb83f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_485) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc57296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4cb9db2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45b344e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(398982cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed5d78eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_484) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0f4818f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_564) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9066652)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_484) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_587) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_466) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68e75052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3b9ae96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_497) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f009e110)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(369033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_615) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a2db40a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f8f954e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c83b6350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_497) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9954469)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_580) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad5c41df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93949318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8346338d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1da963f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
