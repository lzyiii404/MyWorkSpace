//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_94(
  output [2:0]  _EVAL,
  output [3:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  output        _EVAL_2,
  input  [4:0]  _EVAL_3,
  input  [4:0]  _EVAL_4,
  input  [3:0]  _EVAL_5,
  output        _EVAL_6,
  input  [3:0]  _EVAL_7,
  output        _EVAL_8,
  output [7:0]  _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  input  [1:0]  _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input  [7:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output [3:0]  _EVAL_20,
  input  [63:0] _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [63:0] _EVAL_24,
  input         _EVAL_25,
  output [1:0]  _EVAL_26,
  input  [4:0]  _EVAL_27,
  output        _EVAL_28,
  input  [31:0] _EVAL_29,
  input  [3:0]  _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [4:0]  _EVAL_33,
  output [1:0]  _EVAL_34,
  input         _EVAL_35,
  input  [1:0]  _EVAL_36,
  input         _EVAL_37,
  output [4:0]  _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  output [1:0]  _EVAL_41,
  output [2:0]  _EVAL_42,
  output        _EVAL_43,
  input         _EVAL_44,
  output [31:0] _EVAL_45,
  output        _EVAL_46,
  input  [7:0]  _EVAL_47,
  input  [3:0]  _EVAL_48,
  input  [3:0]  _EVAL_49,
  input  [2:0]  _EVAL_50,
  output [3:0]  _EVAL_51,
  output [31:0] _EVAL_52,
  input         _EVAL_53,
  output [7:0]  _EVAL_54,
  input  [3:0]  _EVAL_55,
  output [3:0]  _EVAL_56,
  output [7:0]  _EVAL_57,
  input  [1:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  output [2:0]  _EVAL_60,
  input         _EVAL_61,
  input  [4:0]  _EVAL_62,
  input  [7:0]  _EVAL_63,
  output [3:0]  _EVAL_64,
  input  [3:0]  _EVAL_65,
  output        _EVAL_66,
  output [3:0]  _EVAL_67,
  input         _EVAL_68,
  input         _EVAL_69,
  input  [2:0]  _EVAL_70,
  input         _EVAL_71,
  output [4:0]  _EVAL_72,
  input         _EVAL_73,
  output        _EVAL_74,
  output [1:0]  _EVAL_75,
  output [4:0]  _EVAL_76,
  output [63:0] _EVAL_77,
  input  [2:0]  _EVAL_78,
  output [3:0]  _EVAL_79,
  output [63:0] _EVAL_80,
  output        _EVAL_81,
  output [2:0]  _EVAL_82,
  input  [31:0] _EVAL_83,
  input         _EVAL_84
);
  wire [1:0] Queue__EVAL;
  wire  Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire [63:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire [63:0] Queue__EVAL_6;
  wire [4:0] Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire [3:0] Queue__EVAL_9;
  wire [1:0] Queue__EVAL_10;
  wire [4:0] Queue__EVAL_11;
  wire  Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire [3:0] Queue__EVAL_14;
  wire [1:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire [63:0] Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire [63:0] Queue_1__EVAL_6;
  wire [4:0] Queue_1__EVAL_7;
  wire  Queue_1__EVAL_8;
  wire [3:0] Queue_1__EVAL_9;
  wire [1:0] Queue_1__EVAL_10;
  wire [4:0] Queue_1__EVAL_11;
  wire  Queue_1__EVAL_12;
  wire  Queue_1__EVAL_13;
  wire [3:0] Queue_1__EVAL_14;
  reg  _EVAL_178;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_206;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_207;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_267;
  reg [31:0] _RAND_3;
  wire [15:0] _EVAL_90;
  wire  _EVAL_126;
  wire  _EVAL_114;
  wire  _EVAL_234;
  wire  _EVAL_202;
  wire  _EVAL_190;
  wire  _EVAL_225;
  wire  _EVAL_138;
  wire  _EVAL_96;
  wire  _EVAL_276;
  wire  _EVAL_209;
  wire  _EVAL_139;
  wire  _EVAL_112;
  wire  _EVAL_156;
  wire  _EVAL_167;
  wire  _EVAL_172;
  wire  _EVAL_142;
  wire  _EVAL_247;
  wire  _EVAL_132;
  wire  _EVAL_195;
  wire  _EVAL_271;
  wire  _EVAL_194;
  wire [3:0] _EVAL_128;
  wire [3:0] _EVAL_237;
  wire [15:0] _EVAL_157;
  wire  _EVAL_175;
  wire  _EVAL_208;
  wire  _EVAL_151;
  wire  _EVAL_113;
  wire  _EVAL_189;
  wire  _EVAL_124;
  wire  _EVAL_213;
  wire  _EVAL_201;
  wire  _EVAL_143;
  wire  _EVAL_259;
  wire  _EVAL_199;
  wire  _EVAL_99;
  wire  _EVAL_163;
  wire  _EVAL_192;
  wire  _EVAL_130;
  wire  _EVAL_118;
  wire  _EVAL_171;
  wire  _EVAL_253;
  wire  _EVAL_212;
  wire  _EVAL_125;
  wire  _EVAL_219;
  wire  _EVAL_226;
  wire  _EVAL_216;
  wire  _EVAL_229;
  wire [3:0] _EVAL_197;
  wire [3:0] _EVAL_165;
  wire  _EVAL_144;
  wire  _EVAL_266;
  wire  _EVAL_155;
  wire [3:0] _EVAL_230;
  wire [3:0] _EVAL_205;
  wire  _EVAL_141;
  wire [3:0] _EVAL_94;
  wire [3:0] _EVAL_240;
  wire  _EVAL_258;
  wire [15:0] _EVAL_115;
  wire [16:0] _EVAL_136;
  wire [16:0] _EVAL_273;
  wire [15:0] _EVAL_117;
  wire [15:0] _EVAL_152;
  wire [17:0] _EVAL_173;
  wire [15:0] _EVAL_243;
  wire [15:0] _EVAL_135;
  wire [19:0] _EVAL_262;
  wire [15:0] _EVAL_121;
  wire [15:0] _EVAL_214;
  wire [23:0] _EVAL_210;
  wire [15:0] _EVAL_134;
  wire [15:0] _EVAL_277;
  wire [16:0] _EVAL_133;
  wire [16:0] _EVAL_275;
  wire [16:0] _EVAL_223;
  wire  _EVAL_248;
  wire [15:0] _EVAL_261;
  wire [15:0] _EVAL_217;
  wire [15:0] _EVAL_269;
  wire [7:0] _EVAL_227;
  wire  _EVAL_88;
  wire [1:0] _EVAL_109;
  wire [1:0] _EVAL_154;
  wire [1:0] _EVAL_218;
  wire [1:0] _EVAL_250;
  wire [1:0] _EVAL_119;
  wire [1:0] _EVAL_252;
  wire [1:0] _EVAL_127;
  wire [1:0] _EVAL_245;
  wire [1:0] _EVAL_89;
  wire [1:0] _EVAL_95;
  wire [1:0] _EVAL_107;
  wire [1:0] _EVAL_149;
  wire  _EVAL_272;
  wire  _EVAL_224;
  wire  _EVAL_196;
  wire [63:0] _EVAL_102;
  wire [4:0] _EVAL_198;
  wire [4:0] _EVAL_184;
  wire [4:0] _EVAL_233;
  wire [4:0] _EVAL_93;
  wire [4:0] _EVAL_129;
  wire [4:0] _EVAL_92;
  wire [4:0] _EVAL_249;
  wire [4:0] _EVAL_241;
  wire [7:0] _EVAL_185;
  wire [7:0] _EVAL_161;
  wire [3:0] _EVAL_203;
  wire [3:0] _EVAL_103;
  wire [3:0] _EVAL_191;
  wire [1:0] _EVAL_257;
  wire  _EVAL_86;
  wire [3:0] _EVAL_87;
  wire [3:0] _EVAL_215;
  wire [3:0] _EVAL_222;
  wire [3:0] _EVAL_123;
  wire [3:0] _EVAL_187;
  wire [3:0] _EVAL_186;
  wire [3:0] _EVAL_146;
  wire [3:0] _EVAL_255;
  wire [3:0] _EVAL_182;
  wire [3:0] _EVAL_251;
  wire [3:0] _EVAL_211;
  wire [3:0] _EVAL_204;
  wire [3:0] _EVAL_158;
  wire [3:0] _EVAL_111;
  wire [3:0] _EVAL_244;
  wire [63:0] _EVAL_181;
  wire [63:0] _EVAL_236;
  wire [63:0] _EVAL_263;
  wire [63:0] _EVAL_174;
  wire [63:0] _EVAL_168;
  wire [63:0] _EVAL_176;
  wire [63:0] _EVAL_104;
  wire [63:0] _EVAL_228;
  wire [63:0] _EVAL_160;
  wire [63:0] _EVAL_238;
  wire [63:0] _EVAL_122;
  wire [63:0] _EVAL_268;
  wire [63:0] _EVAL_169;
  wire [63:0] _EVAL_162;
  wire [63:0] _EVAL_105;
  wire  _EVAL_179;
  wire [3:0] _EVAL_180;
  wire [1:0] _EVAL_170;
  wire [1:0] _EVAL_264;
  wire [1:0] _EVAL_183;
  wire [1:0] _EVAL_231;
  wire  _EVAL_260;
  wire [4:0] _EVAL_110;
  wire [4:0] _EVAL_145;
  wire [4:0] _EVAL_137;
  wire [1:0] _EVAL_166;
  wire [1:0] _EVAL_188;
  wire  _EVAL_120;
  wire [4:0] _EVAL_246;
  wire [4:0] _EVAL_91;
  wire [4:0] _EVAL_147;
  wire [4:0] _EVAL_164;
  wire [4:0] _EVAL_85;
  wire [4:0] _EVAL_153;
  wire [4:0] _EVAL_256;
  SiFive__EVAL_93 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14)
  );
  SiFive__EVAL_93 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14)
  );
  assign _EVAL_90 = 16'h1 << _EVAL_5;
  assign _EVAL_126 = _EVAL_90[0];
  assign _EVAL_114 = Queue_1__EVAL_2;
  assign _EVAL_234 = Queue__EVAL_2;
  assign _EVAL_202 = 4'h1 == _EVAL_5 ? _EVAL_114 : _EVAL_234;
  assign _EVAL_190 = 4'h2 == _EVAL_5 ? 1'h0 : _EVAL_202;
  assign _EVAL_225 = 4'h3 == _EVAL_5 ? 1'h0 : _EVAL_190;
  assign _EVAL_138 = 4'h4 == _EVAL_5 ? 1'h0 : _EVAL_225;
  assign _EVAL_96 = 4'h5 == _EVAL_5 ? 1'h0 : _EVAL_138;
  assign _EVAL_276 = 4'h6 == _EVAL_5 ? 1'h0 : _EVAL_96;
  assign _EVAL_209 = 4'h7 == _EVAL_5 ? 1'h0 : _EVAL_276;
  assign _EVAL_139 = 4'h8 == _EVAL_5 ? 1'h0 : _EVAL_209;
  assign _EVAL_112 = 4'h9 == _EVAL_5 ? 1'h0 : _EVAL_139;
  assign _EVAL_156 = 4'ha == _EVAL_5 ? 1'h0 : _EVAL_112;
  assign _EVAL_167 = 4'hb == _EVAL_5 ? 1'h0 : _EVAL_156;
  assign _EVAL_172 = 4'hc == _EVAL_5 ? 1'h0 : _EVAL_167;
  assign _EVAL_142 = 4'hd == _EVAL_5 ? 1'h0 : _EVAL_172;
  assign _EVAL_247 = 4'he == _EVAL_5 ? 1'h0 : _EVAL_142;
  assign _EVAL_132 = 4'hf == _EVAL_5 ? 1'h0 : _EVAL_247;
  assign _EVAL_195 = _EVAL_132 & _EVAL_22;
  assign _EVAL_271 = _EVAL_126 & _EVAL_195;
  assign _EVAL_194 = _EVAL_271 & _EVAL_53;
  assign _EVAL_128 = {{3'd0}, _EVAL_194};
  assign _EVAL_237 = _EVAL_267 + _EVAL_128;
  assign _EVAL_157 = 16'h1 << _EVAL_207;
  assign _EVAL_175 = _EVAL_157[0];
  assign _EVAL_208 = _EVAL_44 & _EVAL_178;
  assign _EVAL_151 = _EVAL_175 & _EVAL_208;
  assign _EVAL_113 = Queue_1__EVAL_13;
  assign _EVAL_189 = Queue__EVAL_13;
  assign _EVAL_124 = 4'h1 == _EVAL_207 ? _EVAL_113 : _EVAL_189;
  assign _EVAL_213 = 4'h2 == _EVAL_207 ? 1'h0 : _EVAL_124;
  assign _EVAL_201 = 4'h3 == _EVAL_207 ? 1'h0 : _EVAL_213;
  assign _EVAL_143 = 4'h4 == _EVAL_207 ? 1'h0 : _EVAL_201;
  assign _EVAL_259 = 4'h5 == _EVAL_207 ? 1'h0 : _EVAL_143;
  assign _EVAL_199 = 4'h6 == _EVAL_207 ? 1'h0 : _EVAL_259;
  assign _EVAL_99 = 4'h7 == _EVAL_207 ? 1'h0 : _EVAL_199;
  assign _EVAL_163 = 4'h8 == _EVAL_207 ? 1'h0 : _EVAL_99;
  assign _EVAL_192 = 4'h9 == _EVAL_207 ? 1'h0 : _EVAL_163;
  assign _EVAL_130 = 4'ha == _EVAL_207 ? 1'h0 : _EVAL_192;
  assign _EVAL_118 = 4'hb == _EVAL_207 ? 1'h0 : _EVAL_130;
  assign _EVAL_171 = 4'hc == _EVAL_207 ? 1'h0 : _EVAL_118;
  assign _EVAL_253 = 4'hd == _EVAL_207 ? 1'h0 : _EVAL_171;
  assign _EVAL_212 = 4'he == _EVAL_207 ? 1'h0 : _EVAL_253;
  assign _EVAL_125 = 4'hf == _EVAL_207 ? 1'h0 : _EVAL_212;
  assign _EVAL_219 = _EVAL_151 & _EVAL_125;
  assign _EVAL_226 = _EVAL_90[1];
  assign _EVAL_216 = _EVAL_226 & _EVAL_195;
  assign _EVAL_229 = _EVAL_216 & _EVAL_53;
  assign _EVAL_197 = {{3'd0}, _EVAL_229};
  assign _EVAL_165 = _EVAL_206 + _EVAL_197;
  assign _EVAL_144 = _EVAL_157[1];
  assign _EVAL_266 = _EVAL_144 & _EVAL_208;
  assign _EVAL_155 = _EVAL_266 & _EVAL_125;
  assign _EVAL_230 = {{3'd0}, _EVAL_155};
  assign _EVAL_205 = _EVAL_165 - _EVAL_230;
  assign _EVAL_141 = _EVAL_205 != 4'h0;
  assign _EVAL_94 = {{3'd0}, _EVAL_219};
  assign _EVAL_240 = _EVAL_237 - _EVAL_94;
  assign _EVAL_258 = _EVAL_240 != 4'h0;
  assign _EVAL_115 = {8'h0,4'h0,2'h0,_EVAL_141,_EVAL_258};
  assign _EVAL_136 = {{1'd0}, _EVAL_115};
  assign _EVAL_273 = {_EVAL_115, 1'h0};
  assign _EVAL_117 = _EVAL_273[15:0];
  assign _EVAL_152 = _EVAL_115 | _EVAL_117;
  assign _EVAL_173 = {_EVAL_152, 2'h0};
  assign _EVAL_243 = _EVAL_173[15:0];
  assign _EVAL_135 = _EVAL_152 | _EVAL_243;
  assign _EVAL_262 = {_EVAL_135, 4'h0};
  assign _EVAL_121 = _EVAL_262[15:0];
  assign _EVAL_214 = _EVAL_135 | _EVAL_121;
  assign _EVAL_210 = {_EVAL_214, 8'h0};
  assign _EVAL_134 = _EVAL_210[15:0];
  assign _EVAL_277 = _EVAL_214 | _EVAL_134;
  assign _EVAL_133 = {_EVAL_277, 1'h0};
  assign _EVAL_275 = ~ _EVAL_133;
  assign _EVAL_223 = _EVAL_136 & _EVAL_275;
  assign _EVAL_248 = _EVAL_223[16];
  assign _EVAL_261 = {{15'd0}, _EVAL_248};
  assign _EVAL_217 = _EVAL_223[15:0];
  assign _EVAL_269 = _EVAL_261 | _EVAL_217;
  assign _EVAL_227 = _EVAL_269[15:8];
  assign _EVAL_88 = _EVAL_227 != 8'h0;
  assign _EVAL_109 = Queue_1__EVAL_10;
  assign _EVAL_154 = Queue__EVAL_10;
  assign _EVAL_218 = 4'h1 == _EVAL_207 ? _EVAL_109 : _EVAL_154;
  assign _EVAL_250 = 4'h2 == _EVAL_207 ? 2'h0 : _EVAL_218;
  assign _EVAL_119 = 4'h3 == _EVAL_207 ? 2'h0 : _EVAL_250;
  assign _EVAL_252 = 4'h4 == _EVAL_207 ? 2'h0 : _EVAL_119;
  assign _EVAL_127 = 4'h5 == _EVAL_207 ? 2'h0 : _EVAL_252;
  assign _EVAL_245 = 4'h6 == _EVAL_207 ? 2'h0 : _EVAL_127;
  assign _EVAL_89 = 4'h7 == _EVAL_207 ? 2'h0 : _EVAL_245;
  assign _EVAL_95 = 4'h8 == _EVAL_207 ? 2'h0 : _EVAL_89;
  assign _EVAL_107 = 4'h9 == _EVAL_207 ? 2'h0 : _EVAL_95;
  assign _EVAL_149 = 4'ha == _EVAL_207 ? 2'h0 : _EVAL_107;
  assign _EVAL_272 = _EVAL_178 == 1'h0;
  assign _EVAL_224 = _EVAL_208 & _EVAL_125;
  assign _EVAL_196 = _EVAL_272 | _EVAL_224;
  assign _EVAL_102 = Queue__EVAL_6;
  assign _EVAL_198 = Queue_1__EVAL_7;
  assign _EVAL_184 = Queue__EVAL_7;
  assign _EVAL_233 = 4'h1 == _EVAL_207 ? _EVAL_198 : _EVAL_184;
  assign _EVAL_93 = 4'h2 == _EVAL_207 ? 5'h0 : _EVAL_233;
  assign _EVAL_129 = 4'h3 == _EVAL_207 ? 5'h0 : _EVAL_93;
  assign _EVAL_92 = 4'h4 == _EVAL_207 ? 5'h0 : _EVAL_129;
  assign _EVAL_249 = 4'h5 == _EVAL_207 ? 5'h0 : _EVAL_92;
  assign _EVAL_241 = 4'h6 == _EVAL_207 ? 5'h0 : _EVAL_249;
  assign _EVAL_185 = _EVAL_269[7:0];
  assign _EVAL_161 = _EVAL_227 | _EVAL_185;
  assign _EVAL_203 = _EVAL_161[7:4];
  assign _EVAL_103 = _EVAL_161[3:0];
  assign _EVAL_191 = _EVAL_203 | _EVAL_103;
  assign _EVAL_257 = _EVAL_191[3:2];
  assign _EVAL_86 = _EVAL_257 != 2'h0;
  assign _EVAL_87 = Queue_1__EVAL_14;
  assign _EVAL_215 = Queue__EVAL_14;
  assign _EVAL_222 = 4'h1 == _EVAL_207 ? _EVAL_87 : _EVAL_215;
  assign _EVAL_123 = 4'h2 == _EVAL_207 ? 4'h0 : _EVAL_222;
  assign _EVAL_187 = 4'h3 == _EVAL_207 ? 4'h0 : _EVAL_123;
  assign _EVAL_186 = 4'h4 == _EVAL_207 ? 4'h0 : _EVAL_187;
  assign _EVAL_146 = 4'h5 == _EVAL_207 ? 4'h0 : _EVAL_186;
  assign _EVAL_255 = 4'h6 == _EVAL_207 ? 4'h0 : _EVAL_146;
  assign _EVAL_182 = 4'h7 == _EVAL_207 ? 4'h0 : _EVAL_255;
  assign _EVAL_251 = 4'h8 == _EVAL_207 ? 4'h0 : _EVAL_182;
  assign _EVAL_211 = 4'h9 == _EVAL_207 ? 4'h0 : _EVAL_251;
  assign _EVAL_204 = 4'ha == _EVAL_207 ? 4'h0 : _EVAL_211;
  assign _EVAL_158 = 4'hb == _EVAL_207 ? 4'h0 : _EVAL_204;
  assign _EVAL_111 = 4'hc == _EVAL_207 ? 4'h0 : _EVAL_158;
  assign _EVAL_244 = 4'hd == _EVAL_207 ? 4'h0 : _EVAL_111;
  assign _EVAL_181 = Queue_1__EVAL_6;
  assign _EVAL_236 = 4'h1 == _EVAL_207 ? _EVAL_181 : _EVAL_102;
  assign _EVAL_263 = 4'h2 == _EVAL_207 ? 64'h0 : _EVAL_236;
  assign _EVAL_174 = 4'h3 == _EVAL_207 ? 64'h0 : _EVAL_263;
  assign _EVAL_168 = 4'h4 == _EVAL_207 ? 64'h0 : _EVAL_174;
  assign _EVAL_176 = 4'h5 == _EVAL_207 ? 64'h0 : _EVAL_168;
  assign _EVAL_104 = 4'h6 == _EVAL_207 ? 64'h0 : _EVAL_176;
  assign _EVAL_228 = 4'h7 == _EVAL_207 ? 64'h0 : _EVAL_104;
  assign _EVAL_160 = 4'h8 == _EVAL_207 ? 64'h0 : _EVAL_228;
  assign _EVAL_238 = 4'h9 == _EVAL_207 ? 64'h0 : _EVAL_160;
  assign _EVAL_122 = 4'ha == _EVAL_207 ? 64'h0 : _EVAL_238;
  assign _EVAL_268 = 4'hb == _EVAL_207 ? 64'h0 : _EVAL_122;
  assign _EVAL_169 = 4'hc == _EVAL_207 ? 64'h0 : _EVAL_268;
  assign _EVAL_162 = 4'hd == _EVAL_207 ? 64'h0 : _EVAL_169;
  assign _EVAL_105 = 4'he == _EVAL_207 ? 64'h0 : _EVAL_162;
  assign _EVAL_179 = _EVAL_115 != 16'h0;
  assign _EVAL_180 = 4'he == _EVAL_207 ? 4'h0 : _EVAL_244;
  assign _EVAL_170 = 4'hb == _EVAL_207 ? 2'h0 : _EVAL_149;
  assign _EVAL_264 = 4'hc == _EVAL_207 ? 2'h0 : _EVAL_170;
  assign _EVAL_183 = 4'hd == _EVAL_207 ? 2'h0 : _EVAL_264;
  assign _EVAL_231 = 4'he == _EVAL_207 ? 2'h0 : _EVAL_183;
  assign _EVAL_260 = _EVAL_203 != 4'h0;
  assign _EVAL_110 = 4'h7 == _EVAL_207 ? 5'h0 : _EVAL_241;
  assign _EVAL_145 = 4'h8 == _EVAL_207 ? 5'h0 : _EVAL_110;
  assign _EVAL_137 = 4'h9 == _EVAL_207 ? 5'h0 : _EVAL_145;
  assign _EVAL_166 = _EVAL_191[1:0];
  assign _EVAL_188 = _EVAL_257 | _EVAL_166;
  assign _EVAL_120 = _EVAL_188[1];
  assign _EVAL_246 = {_EVAL_248,_EVAL_88,_EVAL_260,_EVAL_86,_EVAL_120};
  assign _EVAL_91 = _EVAL_196 ? _EVAL_246 : {{1'd0}, _EVAL_207};
  assign _EVAL_147 = 4'ha == _EVAL_207 ? 5'h0 : _EVAL_137;
  assign _EVAL_164 = 4'hb == _EVAL_207 ? 5'h0 : _EVAL_147;
  assign _EVAL_85 = 4'hc == _EVAL_207 ? 5'h0 : _EVAL_164;
  assign _EVAL_153 = 4'hd == _EVAL_207 ? 5'h0 : _EVAL_85;
  assign _EVAL_256 = 4'he == _EVAL_207 ? 5'h0 : _EVAL_153;
  assign _EVAL_6 = _EVAL_68;
  assign _EVAL_43 = _EVAL_31;
  assign _EVAL_34 = _EVAL_1;
  assign Queue_1__EVAL_3 = _EVAL_24;
  assign _EVAL_51 = _EVAL_7;
  assign Queue_1__EVAL_12 = _EVAL_226 & _EVAL_22;
  assign _EVAL_0 = _EVAL_48;
  assign _EVAL_66 = _EVAL_35;
  assign _EVAL_45 = _EVAL_83;
  assign _EVAL_8 = _EVAL_84;
  assign _EVAL_19 = _EVAL_178;
  assign _EVAL_23 = _EVAL_25;
  assign _EVAL_33 = 4'hf == _EVAL_207 ? 5'h0 : _EVAL_256;
  assign Queue_1__EVAL_0 = _EVAL_53;
  assign _EVAL = _EVAL_17;
  assign _EVAL_82 = _EVAL_70;
  assign Queue_1__EVAL_1 = _EVAL_144 & _EVAL_208;
  assign Queue__EVAL_8 = _EVAL_71;
  assign _EVAL_79 = _EVAL_30;
  assign Queue_1__EVAL = _EVAL_12;
  assign _EVAL_42 = _EVAL_78;
  assign _EVAL_13 = _EVAL_40;
  assign _EVAL_64 = _EVAL_49;
  assign _EVAL_56 = 4'hf == _EVAL_207 ? 4'h0 : _EVAL_180;
  assign Queue_1__EVAL_4 = _EVAL_32;
  assign Queue_1__EVAL_9 = _EVAL_5;
  assign Queue_1__EVAL_11 = _EVAL_62;
  assign _EVAL_57 = _EVAL_47;
  assign _EVAL_74 = 4'hf == _EVAL_207 ? 1'h0 : _EVAL_212;
  assign _EVAL_72 = _EVAL_4;
  assign Queue__EVAL_12 = _EVAL_126 & _EVAL_22;
  assign Queue__EVAL_1 = _EVAL_175 & _EVAL_208;
  assign Queue__EVAL_9 = _EVAL_5;
  assign Queue__EVAL = _EVAL_12;
  assign _EVAL_9 = _EVAL_15;
  assign _EVAL_52 = _EVAL_29;
  assign _EVAL_10 = _EVAL_69;
  assign _EVAL_76 = _EVAL_27;
  assign _EVAL_60 = _EVAL_50;
  assign _EVAL_46 = _EVAL_73;
  assign Queue__EVAL_0 = _EVAL_53;
  assign _EVAL_59 = _EVAL_55;
  assign _EVAL_26 = _EVAL_58;
  assign _EVAL_80 = 4'hf == _EVAL_207 ? 64'h0 : _EVAL_105;
  assign Queue__EVAL_4 = _EVAL_32;
  assign _EVAL_54 = _EVAL_63;
  assign _EVAL_75 = _EVAL_36;
  assign _EVAL_38 = _EVAL_3;
  assign _EVAL_28 = _EVAL_37;
  assign _EVAL_39 = 4'hf == _EVAL_5 ? 1'h0 : _EVAL_247;
  assign _EVAL_11 = _EVAL_61;
  assign Queue_1__EVAL_8 = _EVAL_71;
  assign _EVAL_77 = _EVAL_21;
  assign _EVAL_20 = _EVAL_65;
  assign _EVAL_2 = _EVAL_18;
  assign _EVAL_81 = _EVAL_14;
  assign Queue__EVAL_3 = _EVAL_24;
  assign _EVAL_67 = _EVAL_16;
  assign _EVAL_41 = 4'hf == _EVAL_207 ? 2'h0 : _EVAL_231;
  assign Queue__EVAL_11 = _EVAL_62;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_178 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_206 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_207 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_267 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_32) begin
    if (_EVAL_71) begin
      _EVAL_178 <= 1'h0;
    end else begin
      if (_EVAL_196) begin
        _EVAL_178 <= _EVAL_179;
      end
    end
    if (_EVAL_71) begin
      _EVAL_206 <= 4'h0;
    end else begin
      _EVAL_206 <= _EVAL_205;
    end
    _EVAL_207 <= _EVAL_91[3:0];
    if (_EVAL_71) begin
      _EVAL_267 <= 4'h0;
    end else begin
      _EVAL_267 <= _EVAL_240;
    end
  end
endmodule
