//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_307_assert(
  input        _EVAL_24,
  input        _EVAL_36,
  input        _EVAL_60,
  input        _EVAL_63,
  input        _EVAL_95,
  input        _EVAL_123,
  input        _EVAL_156,
  input        _EVAL_174,
  input        _EVAL_246,
  input        _EVAL_1647,
  input        _EVAL_2506,
  input        _EVAL_3448,
  input        _EVAL_4721,
  input        _EVAL_890,
  input        _EVAL_4820,
  input        _EVAL_1162,
  input        _EVAL_4072,
  input        _EVAL_854,
  input        _EVAL_3672,
  input        _EVAL_5329,
  input        _EVAL_4150,
  input        _EVAL_4474,
  input        _EVAL_4139,
  input        _EVAL_5120,
  input        _EVAL_781,
  input  [2:0] _EVAL_4776,
  input        _EVAL_1246,
  input        _EVAL_2004,
  input        _EVAL_4405,
  input        _EVAL_2963,
  input        _EVAL_3812,
  input  [2:0] _EVAL_3579,
  input        _EVAL_995,
  input        _EVAL_3496,
  input        _EVAL_1691,
  input        _EVAL_686,
  input        _EVAL_646,
  input        _EVAL_2557,
  input        _EVAL_4223,
  input        _EVAL_2402,
  input        _EVAL_1118,
  input        _EVAL_4435,
  input        _EVAL_3592,
  input        _EVAL_3009,
  input        _EVAL_4225,
  input        _EVAL_4788,
  input        _EVAL_2001,
  input        _EVAL_3873,
  input        _EVAL_4671,
  input        _EVAL_1840,
  input        _EVAL_4189,
  input        _EVAL_4125,
  input        _EVAL_2541,
  input        _EVAL_2604,
  input        _EVAL_4149,
  input        _EVAL_4704,
  input        _EVAL_4296,
  input        _EVAL_1852,
  input        _EVAL_5272,
  input        _EVAL_4543,
  input        _EVAL_1034,
  input        _EVAL_1163,
  input        _EVAL_3821,
  input        _EVAL_5276,
  input        _EVAL_1732,
  input        bullet_clock_gate_out
);
  reg  _EVAL_289;
  reg [31:0] _RAND_0;
  reg  _EVAL_295;
  reg [31:0] _RAND_1;
  reg  _EVAL_542;
  reg [31:0] _RAND_2;
  reg  _EVAL_580;
  reg [31:0] _RAND_3;
  reg  _EVAL_763;
  reg [31:0] _RAND_4;
  reg  _EVAL_778;
  reg [31:0] _RAND_5;
  reg  _EVAL_844;
  reg [31:0] _RAND_6;
  reg  _EVAL_877;
  reg [31:0] _RAND_7;
  reg  _EVAL_898;
  reg [31:0] _RAND_8;
  reg  _EVAL_1219;
  reg [31:0] _RAND_9;
  reg  _EVAL_1516;
  reg [31:0] _RAND_10;
  reg  _EVAL_1532;
  reg [31:0] _RAND_11;
  reg  _EVAL_1541;
  reg [31:0] _RAND_12;
  reg  _EVAL_1544;
  reg [31:0] _RAND_13;
  reg  _EVAL_1783;
  reg [31:0] _RAND_14;
  reg  _EVAL_1785;
  reg [31:0] _RAND_15;
  reg  _EVAL_1984;
  reg [31:0] _RAND_16;
  reg  _EVAL_2014;
  reg [31:0] _RAND_17;
  reg  _EVAL_2113;
  reg [31:0] _RAND_18;
  reg  _EVAL_2241;
  reg [31:0] _RAND_19;
  reg  _EVAL_2290;
  reg [31:0] _RAND_20;
  reg  _EVAL_2315;
  reg [31:0] _RAND_21;
  reg  _EVAL_2360;
  reg [31:0] _RAND_22;
  reg  _EVAL_2490;
  reg [31:0] _RAND_23;
  reg  _EVAL_2648;
  reg [31:0] _RAND_24;
  reg  _EVAL_2692;
  reg [31:0] _RAND_25;
  reg  _EVAL_2793;
  reg [31:0] _RAND_26;
  reg  _EVAL_2960;
  reg [31:0] _RAND_27;
  reg  _EVAL_3099;
  reg [31:0] _RAND_28;
  reg  _EVAL_3146;
  reg [31:0] _RAND_29;
  reg  _EVAL_3314;
  reg [31:0] _RAND_30;
  reg  _EVAL_3424;
  reg [31:0] _RAND_31;
  reg  _EVAL_3454;
  reg [31:0] _RAND_32;
  reg  _EVAL_3505;
  reg [31:0] _RAND_33;
  reg  _EVAL_3652;
  reg [31:0] _RAND_34;
  reg  _EVAL_3667;
  reg [31:0] _RAND_35;
  reg  _EVAL_3999;
  reg [31:0] _RAND_36;
  reg  _EVAL_4181;
  reg [31:0] _RAND_37;
  reg  _EVAL_4364;
  reg [31:0] _RAND_38;
  reg  _EVAL_4419;
  reg [31:0] _RAND_39;
  reg  _EVAL_4566;
  reg [31:0] _RAND_40;
  reg  _EVAL_4609;
  reg [31:0] _RAND_41;
  reg  _EVAL_4655;
  reg [31:0] _RAND_42;
  reg  _EVAL_4674;
  reg [31:0] _RAND_43;
  reg  _EVAL_4817;
  reg [31:0] _RAND_44;
  reg  _EVAL_4822;
  reg [31:0] _RAND_45;
  reg  _EVAL_4899;
  reg [31:0] _RAND_46;
  reg  _EVAL_5140;
  reg [31:0] _RAND_47;
  reg  _EVAL_5166;
  reg [31:0] _RAND_48;
  wire [2:0] _EVAL_4904;
  wire [1:0] _EVAL_2501;
  wire [1:0] _EVAL_1035;
  wire [7:0] _EVAL_4113;
  wire [7:0] _EVAL_4891;
  wire [17:0] _EVAL_1172;
  wire [17:0] _EVAL_4558;
  wire [10:0] _EVAL_374;
  wire [10:0] _EVAL_1638;
  wire [2:0] _EVAL_3363;
  wire [3:0] _EVAL_4466;
  wire  _EVAL_4984;
  wire  _EVAL_2680;
  wire  _EVAL_2527;
  wire  _EVAL_3239;
  wire  _EVAL_2502;
  wire [11:0] _EVAL_3062;
  wire  _EVAL_3660;
  wire  _EVAL_3678;
  wire [2:0] _EVAL_914;
  wire  _EVAL_3976;
  wire  _EVAL_2441;
  wire  _EVAL_1256;
  wire [1:0] _EVAL_1719;
  wire [1:0] _EVAL_5301;
  wire [4:0] _EVAL_1611;
  wire [4:0] _EVAL_2328;
  wire [10:0] _EVAL_3627;
  wire [4:0] _EVAL_5159;
  wire [14:0] _EVAL_3668;
  wire [7:0] _EVAL_2518;
  wire [1:0] _EVAL_4087;
  wire [1:0] _EVAL_304;
  wire [3:0] _EVAL_3774;
  wire  _EVAL_3586;
  wire [15:0] _EVAL_2361;
  wire [15:0] _EVAL_355;
  wire [5:0] _EVAL_3203;
  wire [5:0] _EVAL_4976;
  wire  _EVAL_4989;
  wire  _EVAL_1276;
  wire  _EVAL_4289;
  wire  _EVAL_645;
  wire  _EVAL_3766;
  wire [10:0] _EVAL_1606;
  wire [10:0] _EVAL_2505;
  wire [4:0] _EVAL_1626;
  wire  _EVAL_2016;
  wire  _EVAL_5058;
  wire  _EVAL_3140;
  wire [3:0] _EVAL_2856;
  wire [3:0] _EVAL_4833;
  wire [16:0] _EVAL_787;
  wire [16:0] _EVAL_608;
  wire [8:0] _EVAL_2786;
  wire [8:0] _EVAL_3315;
  wire  _EVAL_1537;
  wire [9:0] _EVAL_752;
  wire [9:0] _EVAL_4110;
  wire  _EVAL_5392;
  wire  _EVAL_3114;
  wire [5:0] _EVAL_446;
  wire [5:0] _EVAL_1147;
  wire  _EVAL_3087;
  wire  _EVAL_865;
  wire [12:0] _EVAL_1337;
  wire  _EVAL_5079;
  wire  _EVAL_3802;
  wire  _EVAL_3556;
  wire  _EVAL_3516;
  wire  _EVAL_5247;
  wire [4:0] _EVAL_2688;
  wire  _EVAL_1596;
  wire [4:0] _EVAL_1878;
  wire [10:0] _EVAL_3005;
  wire [12:0] _EVAL_2476;
  wire  _EVAL_5325;
  wire [4:0] _EVAL_1409;
  wire [5:0] _EVAL_2018;
  wire [5:0] _EVAL_913;
  wire  _EVAL_1053;
  wire [2:0] _EVAL_5256;
  wire [2:0] _EVAL_3634;
  wire [8:0] _EVAL_2513;
  wire [8:0] _EVAL_2966;
  wire [9:0] _EVAL_1850;
  wire [3:0] _EVAL_3636;
  wire  _EVAL_1164;
  wire  _EVAL_376;
  wire  _EVAL_3718;
  wire [8:0] _EVAL_5044;
  wire [8:0] _EVAL_3436;
  wire  _EVAL_5314;
  wire [1:0] _EVAL_312;
  wire [6:0] _EVAL_4695;
  wire [6:0] _EVAL_3772;
  wire [9:0] _EVAL_485;
  wire  _EVAL_287;
  wire [1:0] _EVAL_2222;
  wire [10:0] _EVAL_3887;
  wire  _EVAL_4799;
  wire [7:0] _EVAL_2678;
  wire [3:0] _EVAL_1681;
  wire [3:0] _EVAL_3441;
  wire  _EVAL_4185;
  wire  _EVAL_4720;
  wire  _EVAL_2811;
  wire  _EVAL_1342;
  wire [6:0] _EVAL_3968;
  wire [6:0] _EVAL_3352;
  wire  _EVAL_5165;
  wire  _EVAL_652;
  wire  _EVAL_3767;
  wire  _EVAL_4054;
  wire  _EVAL_1590;
  wire [10:0] _EVAL_2968;
  wire [11:0] _EVAL_1811;
  wire  _EVAL_4876;
  wire [7:0] _EVAL_2651;
  wire [7:0] _EVAL_1351;
  wire  _EVAL_488;
  wire  _EVAL_2261;
  wire  _EVAL_3590;
  wire [9:0] _EVAL_2209;
  wire  _EVAL_3838;
  wire [14:0] _EVAL_2285;
  wire  _EVAL_3451;
  wire [13:0] _EVAL_3687;
  wire [13:0] _EVAL_4711;
  wire  _EVAL_5307;
  wire [9:0] _EVAL_1884;
  wire [4:0] _EVAL_5212;
  wire [3:0] _EVAL_1077;
  assign _EVAL_4904 = {_EVAL_4072, 2'h0};
  assign _EVAL_2501 = {_EVAL_246, 1'h0};
  assign _EVAL_1035 = 2'h2 & _EVAL_2501;
  assign _EVAL_4113 = {_EVAL_5120, 7'h0};
  assign _EVAL_4891 = 8'h80 & _EVAL_4113;
  assign _EVAL_1172 = {_EVAL_1246, 17'h0};
  assign _EVAL_4558 = 18'h20000 & _EVAL_1172;
  assign _EVAL_374 = {_EVAL_3812, 10'h0};
  assign _EVAL_1638 = 11'h400 & _EVAL_374;
  assign _EVAL_3363 = {{2'd0}, _EVAL_1647};
  assign _EVAL_4466 = _EVAL_3579 + _EVAL_3363;
  assign _EVAL_4984 = _EVAL_4466 <= 4'h2;
  assign _EVAL_2680 = _EVAL_4984 | _EVAL_63;
  assign _EVAL_2527 = _EVAL_2680 == 1'h0;
  assign _EVAL_3239 = _EVAL_995 | _EVAL_4139;
  assign _EVAL_2502 = _EVAL_3239 == 1'h0;
  assign _EVAL_3062 = {_EVAL_3496, 11'h0};
  assign _EVAL_3660 = _EVAL_890 & _EVAL_2290;
  assign _EVAL_3678 = _EVAL_890 & _EVAL_2648;
  assign _EVAL_914 = 3'h4 & _EVAL_4904;
  assign _EVAL_3976 = _EVAL_4721 & _EVAL_3652;
  assign _EVAL_2441 = _EVAL_3009 & _EVAL_3672;
  assign _EVAL_1256 = _EVAL_890 & _EVAL_1541;
  assign _EVAL_1719 = {_EVAL_3592, 1'h0};
  assign _EVAL_5301 = {_EVAL_2001, 1'h0};
  assign _EVAL_1611 = {_EVAL_854, 4'h0};
  assign _EVAL_2328 = 5'h10 & _EVAL_1611;
  assign _EVAL_3627 = {_EVAL_4189, 10'h0};
  assign _EVAL_5159 = {_EVAL_2604, 4'h0};
  assign _EVAL_3668 = {_EVAL_646, 14'h0};
  assign _EVAL_2518 = {_EVAL_4149, 7'h0};
  assign _EVAL_4087 = {_EVAL_2402, 1'h0};
  assign _EVAL_304 = 2'h2 & _EVAL_4087;
  assign _EVAL_3774 = {_EVAL_1840, 3'h0};
  assign _EVAL_3586 = _EVAL_4721 & _EVAL_3505;
  assign _EVAL_2361 = {_EVAL_686, 15'h0};
  assign _EVAL_355 = 16'h8000 & _EVAL_2361;
  assign _EVAL_3203 = {_EVAL_1852, 5'h0};
  assign _EVAL_4976 = 6'h20 & _EVAL_3203;
  assign _EVAL_4989 = _EVAL_5272 == 1'h0;
  assign _EVAL_1276 = _EVAL_4989 | _EVAL_4543;
  assign _EVAL_4289 = _EVAL_1276 | _EVAL_63;
  assign _EVAL_645 = _EVAL_4721 & _EVAL_4566;
  assign _EVAL_3766 = _EVAL_2502 | _EVAL_4474;
  assign _EVAL_1606 = {_EVAL_4125, 10'h0};
  assign _EVAL_2505 = 11'h400 & _EVAL_1606;
  assign _EVAL_1626 = {_EVAL_24, 4'h0};
  assign _EVAL_2016 = _EVAL_3821 == 1'h0;
  assign _EVAL_5058 = _EVAL_2016 | _EVAL_5276;
  assign _EVAL_3140 = _EVAL_5058 | _EVAL_63;
  assign _EVAL_2856 = {_EVAL_95, 3'h0};
  assign _EVAL_4833 = 4'h8 & _EVAL_2856;
  assign _EVAL_787 = {_EVAL_1691, 16'h0};
  assign _EVAL_608 = 17'h10000 & _EVAL_787;
  assign _EVAL_2786 = {_EVAL_4435, 8'h0};
  assign _EVAL_3315 = 9'h100 & _EVAL_2786;
  assign _EVAL_1537 = _EVAL_890 & _EVAL_4817;
  assign _EVAL_752 = {_EVAL_1163, 9'h0};
  assign _EVAL_4110 = 10'h200 & _EVAL_752;
  assign _EVAL_5392 = _EVAL_890 & _EVAL_3314;
  assign _EVAL_3114 = _EVAL_4721 & _EVAL_2793;
  assign _EVAL_446 = {_EVAL_4223, 5'h0};
  assign _EVAL_1147 = 6'h20 & _EVAL_446;
  assign _EVAL_3087 = _EVAL_3766 | _EVAL_63;
  assign _EVAL_865 = _EVAL_3087 == 1'h0;
  assign _EVAL_1337 = {_EVAL_1162, 12'h0};
  assign _EVAL_5079 = _EVAL_890 & _EVAL_1532;
  assign _EVAL_3802 = _EVAL_4820 == 1'h0;
  assign _EVAL_3556 = _EVAL_3448 | _EVAL_1732;
  assign _EVAL_3516 = _EVAL_3802 | _EVAL_3556;
  assign _EVAL_5247 = _EVAL_3516 | _EVAL_63;
  assign _EVAL_2688 = {_EVAL_4671, 4'h0};
  assign _EVAL_1596 = _EVAL_4721 & _EVAL_2315;
  assign _EVAL_1878 = 5'h10 & _EVAL_5159;
  assign _EVAL_3005 = 11'h400 & _EVAL_3627;
  assign _EVAL_2476 = 13'h1000 & _EVAL_1337;
  assign _EVAL_5325 = _EVAL_2506 & _EVAL_4704;
  assign _EVAL_1409 = 5'h10 & _EVAL_1626;
  assign _EVAL_2018 = {_EVAL_3873, 5'h0};
  assign _EVAL_913 = 6'h20 & _EVAL_2018;
  assign _EVAL_1053 = _EVAL_4721 & _EVAL_3667;
  assign _EVAL_5256 = {_EVAL_174, 2'h0};
  assign _EVAL_3634 = 3'h4 & _EVAL_5256;
  assign _EVAL_2513 = {_EVAL_4405, 8'h0};
  assign _EVAL_2966 = 9'h100 & _EVAL_2513;
  assign _EVAL_1850 = {_EVAL_2541, 9'h0};
  assign _EVAL_3636 = _EVAL_4776 + _EVAL_3363;
  assign _EVAL_1164 = _EVAL_3636 <= 4'h2;
  assign _EVAL_376 = _EVAL_1164 | _EVAL_63;
  assign _EVAL_3718 = _EVAL_376 == 1'h0;
  assign _EVAL_5044 = {_EVAL_4225, 8'h0};
  assign _EVAL_3436 = 9'h100 & _EVAL_5044;
  assign _EVAL_5314 = _EVAL_2441 == 1'h0;
  assign _EVAL_312 = 2'h2 & _EVAL_1719;
  assign _EVAL_4695 = {_EVAL_5329, 6'h0};
  assign _EVAL_3772 = 7'h40 & _EVAL_4695;
  assign _EVAL_485 = 10'h200 & _EVAL_1850;
  assign _EVAL_287 = _EVAL_4721 & _EVAL_5166;
  assign _EVAL_2222 = 2'h2 & _EVAL_5301;
  assign _EVAL_3887 = {_EVAL_781, 10'h0};
  assign _EVAL_4799 = _EVAL_890 & _EVAL_580;
  assign _EVAL_2678 = 8'h80 & _EVAL_2518;
  assign _EVAL_1681 = {_EVAL_156, 3'h0};
  assign _EVAL_3441 = 4'h8 & _EVAL_1681;
  assign _EVAL_4185 = _EVAL_4289 == 1'h0;
  assign _EVAL_4720 = _EVAL_890 & _EVAL_1783;
  assign _EVAL_2811 = _EVAL_5314 | _EVAL_63;
  assign _EVAL_1342 = _EVAL_2811 == 1'h0;
  assign _EVAL_3968 = {_EVAL_1034, 6'h0};
  assign _EVAL_3352 = 7'h40 & _EVAL_3968;
  assign _EVAL_5165 = _EVAL_5325 == 1'h0;
  assign _EVAL_652 = _EVAL_5165 | _EVAL_63;
  assign _EVAL_3767 = _EVAL_3140 == 1'h0;
  assign _EVAL_4054 = _EVAL_4721 & _EVAL_2490;
  assign _EVAL_1590 = _EVAL_890 & _EVAL_4822;
  assign _EVAL_2968 = 11'h400 & _EVAL_3887;
  assign _EVAL_1811 = 12'h800 & _EVAL_3062;
  assign _EVAL_4876 = _EVAL_652 == 1'h0;
  assign _EVAL_2651 = {_EVAL_2004, 7'h0};
  assign _EVAL_1351 = 8'h80 & _EVAL_2651;
  assign _EVAL_488 = _EVAL_890 & _EVAL_1516;
  assign _EVAL_2261 = _EVAL_63 == 1'h0;
  assign _EVAL_3590 = _EVAL_4721 & _EVAL_1785;
  assign _EVAL_2209 = {_EVAL_4150, 9'h0};
  assign _EVAL_3838 = _EVAL_890 & _EVAL_4674;
  assign _EVAL_2285 = 15'h4000 & _EVAL_3668;
  assign _EVAL_3451 = _EVAL_5247 == 1'h0;
  assign _EVAL_3687 = {_EVAL_2557, 13'h0};
  assign _EVAL_4711 = 14'h2000 & _EVAL_3687;
  assign _EVAL_5307 = _EVAL_890 & _EVAL_2014;
  assign _EVAL_1884 = 10'h200 & _EVAL_2209;
  assign _EVAL_5212 = 5'h10 & _EVAL_2688;
  assign _EVAL_1077 = 4'h8 & _EVAL_3774;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_289 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_295 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_542 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_580 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_763 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_778 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_844 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_877 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_898 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_1219 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_1516 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_1532 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_1541 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_1544 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_1783 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_1785 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_1984 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_2014 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_2113 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_2241 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_2290 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_2315 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_2360 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_2490 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_2648 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_2692 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_2793 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_2960 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_3099 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_3146 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_3314 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_3424 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_3454 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_3505 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_3652 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_3667 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_3999 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_4181 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_4364 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_4419 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_4566 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_4609 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_4655 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_4674 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_4817 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_4822 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_4899 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_5140 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_5166 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge bullet_clock_gate_out) begin
    _EVAL_289 <= _EVAL_4110 != 10'h0;
    _EVAL_295 <= _EVAL_2222 != 2'h0;
    _EVAL_542 <= _EVAL_4833 != 4'h0;
    _EVAL_580 <= _EVAL_2285 != 15'h0;
    _EVAL_763 <= _EVAL_304 != 2'h0;
    _EVAL_778 <= _EVAL_1638 != 11'h0;
    _EVAL_844 <= _EVAL_1409 != 5'h0;
    _EVAL_877 <= _EVAL_1351 != 8'h0;
    _EVAL_898 <= _EVAL_3441 != 4'h0;
    _EVAL_1219 <= _EVAL_1878 != 5'h0;
    _EVAL_1516 <= _EVAL_2966 != 9'h0;
    _EVAL_1532 <= _EVAL_2968 != 11'h0;
    _EVAL_1541 <= _EVAL_355 != 16'h0;
    _EVAL_1544 <= _EVAL_3634 != 3'h0;
    _EVAL_1783 <= _EVAL_1884 != 10'h0;
    _EVAL_1785 <= _EVAL_2505 != 11'h0;
    _EVAL_1984 <= _EVAL_36;
    _EVAL_2014 <= _EVAL_1147 != 6'h0;
    _EVAL_2113 <= _EVAL_3441 != 4'h0;
    _EVAL_2241 <= _EVAL_3436 != 9'h0;
    _EVAL_2290 <= _EVAL_608 != 17'h0;
    _EVAL_2315 <= _EVAL_914 != 3'h0;
    _EVAL_2360 <= _EVAL_3634 != 3'h0;
    _EVAL_2490 <= _EVAL_1077 != 4'h0;
    _EVAL_2648 <= _EVAL_4558 != 18'h0;
    _EVAL_2692 <= _EVAL_2963 & _EVAL_1118;
    _EVAL_2793 <= _EVAL_312 != 2'h0;
    _EVAL_2960 <= _EVAL_36;
    _EVAL_3099 <= _EVAL_4976 != 6'h0;
    _EVAL_3146 <= _EVAL_4833 != 4'h0;
    _EVAL_3314 <= _EVAL_4891 != 8'h0;
    _EVAL_3424 <= _EVAL_3315 != 9'h0;
    _EVAL_3454 <= _EVAL_1409 != 5'h0;
    _EVAL_3505 <= _EVAL_2476 != 13'h0;
    _EVAL_3652 <= _EVAL_5212 != 5'h0;
    _EVAL_3667 <= _EVAL_1811 != 12'h0;
    _EVAL_3999 <= _EVAL_3005 != 11'h0;
    _EVAL_4181 <= _EVAL_3352 != 7'h0;
    _EVAL_4364 <= _EVAL_2678 != 8'h0;
    _EVAL_4419 <= _EVAL_4788 & _EVAL_4296;
    _EVAL_4566 <= _EVAL_913 != 6'h0;
    _EVAL_4609 <= _EVAL_3352 != 7'h0;
    _EVAL_4655 <= _EVAL_4976 != 6'h0;
    _EVAL_4674 <= _EVAL_4711 != 14'h0;
    _EVAL_4817 <= _EVAL_2328 != 5'h0;
    _EVAL_4822 <= _EVAL_3772 != 7'h0;
    _EVAL_4899 <= _EVAL_1035 != 2'h0;
    _EVAL_5140 <= _EVAL_1035 != 2'h0;
    _EVAL_5166 <= _EVAL_485 != 10'h0;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4054 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1fb4482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2527) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5392 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb685a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2692 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff19b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4899 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93b71033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5307 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(197905c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3451) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2960 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e69b87d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_763 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d5b70e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4364 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8382174d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3451) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd5aef2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1544 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1b6662a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_898 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dcbf071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1537 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c734ac48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3114 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c699316)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3767) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1647 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53d47da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3999 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daffcba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3590 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(537ee5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bd5f96c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3424 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef528e66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d5b70e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4799 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cc4951a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2360 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1b6662a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4720 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10857e91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4181 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a243b90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3718) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5a8a247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1256 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62bbe377)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1984 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e69b87d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3678 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec6fd407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2527) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5a8a247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3099 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4af3784)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3838 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18df66e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac6f5d54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3146 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f355195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1053 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82a80c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_877 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8382174d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2113 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dcbf071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f355195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4609 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a243b90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4876) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44500821)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_865) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28be6844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_778 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daffcba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1219 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0a15140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3767) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bd5f96c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1590 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a0821e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9193043b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3454 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ea25701)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3976 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c734ac48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_865) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2241 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef528e66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4655 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4af3784)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4876) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2efaad1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5079 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(537ee5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(197905c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44500821)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c75b07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3586 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2122785e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3660 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(372e1772)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1596 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a01b668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_844 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ea25701)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3718) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4419 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff19b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10857e91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5140 & _EVAL_2261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93b71033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
