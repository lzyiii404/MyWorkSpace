//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_100_assert(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [7:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_26;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_39;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_52;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_56;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_65;
  reg [31:0] _RAND_4;
  reg  _EVAL_82;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_133;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_134;
  reg [31:0] _RAND_7;
  reg  _EVAL_137;
  reg [31:0] _RAND_8;
  reg [1:0] _EVAL_154;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_162;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_170;
  reg [31:0] _RAND_11;
  reg [31:0] _EVAL_185;
  reg [31:0] _RAND_12;
  reg  _EVAL_248;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_269;
  reg [31:0] _RAND_14;
  wire  _EVAL_254;
  wire  _EVAL_276;
  wire  _EVAL_221;
  wire [1:0] _EVAL_128;
  wire  _EVAL_22;
  wire  _EVAL_106;
  wire  _EVAL_224;
  wire  _EVAL_96;
  wire [1:0] _EVAL_47;
  wire [3:0] _EVAL_207;
  wire [2:0] _EVAL_84;
  wire [2:0] _EVAL_21;
  wire  _EVAL_220;
  wire  _EVAL_211;
  wire  _EVAL_118;
  wire  _EVAL_37;
  wire  _EVAL_274;
  wire  _EVAL_174;
  wire  _EVAL_193;
  wire  _EVAL_237;
  wire  _EVAL_251;
  wire  _EVAL_127;
  wire  _EVAL_230;
  wire  _EVAL_271;
  wire  _EVAL_245;
  wire  _EVAL_204;
  wire  _EVAL_100;
  wire  _EVAL_192;
  wire  _EVAL_242;
  wire  _EVAL_142;
  wire  _EVAL_167;
  wire  _EVAL_30;
  wire  _EVAL_250;
  wire  _EVAL_114;
  wire  _EVAL_119;
  wire  _EVAL_189;
  wire  _EVAL_120;
  wire  _EVAL_234;
  wire  _EVAL_93;
  wire  _EVAL_163;
  wire  _EVAL_268;
  wire  _EVAL_223;
  wire  _EVAL_90;
  wire  _EVAL_178;
  wire  _EVAL_91;
  wire  _EVAL_176;
  wire  _EVAL_227;
  wire  _EVAL_99;
  wire  _EVAL_101;
  wire  _EVAL_74;
  wire  _EVAL_66;
  wire  _EVAL_214;
  wire  _EVAL_156;
  wire  _EVAL_67;
  wire  _EVAL_173;
  wire  _EVAL_249;
  wire  _EVAL_41;
  wire  _EVAL_35;
  wire  _EVAL_168;
  wire  _EVAL_64;
  wire  _EVAL_136;
  wire [7:0] _EVAL_217;
  wire  _EVAL_46;
  wire  _EVAL_171;
  wire  _EVAL_213;
  wire  _EVAL_81;
  wire  _EVAL_144;
  wire  _EVAL_195;
  wire [1:0] _EVAL_257;
  wire [1:0] _EVAL_72;
  wire  _EVAL_228;
  wire  _EVAL_265;
  wire  _EVAL_277;
  wire  _EVAL_86;
  wire  _EVAL_20;
  wire  _EVAL_205;
  wire [1:0] _EVAL_222;
  wire [1:0] _EVAL_50;
  wire  _EVAL_78;
  wire [12:0] _EVAL_104;
  wire [5:0] _EVAL_203;
  wire  _EVAL_43;
  wire  _EVAL_243;
  wire [1:0] _EVAL_209;
  wire [1:0] _EVAL_25;
  wire  _EVAL_105;
  wire  _EVAL_151;
  wire  _EVAL_182;
  wire  _EVAL_129;
  wire  _EVAL_139;
  wire  _EVAL_191;
  wire  _EVAL_34;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_272;
  wire  _EVAL_115;
  wire  _EVAL_113;
  wire  _EVAL_190;
  wire  _EVAL_273;
  wire  _EVAL_94;
  wire [7:0] _EVAL_282;
  wire [7:0] _EVAL_117;
  wire  _EVAL_164;
  wire  _EVAL_17;
  wire  _EVAL_280;
  wire  _EVAL_38;
  wire  _EVAL_215;
  wire  _EVAL_212;
  wire [31:0] _EVAL_264;
  wire [32:0] _EVAL_161;
  wire [32:0] _EVAL_218;
  wire [32:0] _EVAL_68;
  wire  _EVAL_145;
  wire  _EVAL_77;
  wire  _EVAL_53;
  wire [7:0] _EVAL_80;
  wire  _EVAL_231;
  wire  _EVAL_179;
  wire  _EVAL_97;
  wire  _EVAL_103;
  wire  _EVAL_98;
  wire  _EVAL_19;
  wire  _EVAL_180;
  wire  _EVAL_76;
  wire  _EVAL_123;
  wire  _EVAL_186;
  wire  _EVAL_69;
  wire  _EVAL_126;
  wire [12:0] _EVAL_92;
  wire [5:0] _EVAL_88;
  wire [5:0] _EVAL_229;
  wire [2:0] _EVAL_208;
  wire [2:0] _EVAL_225;
  wire  _EVAL_149;
  wire  _EVAL_157;
  wire  _EVAL_262;
  wire [31:0] _EVAL_122;
  wire [31:0] _EVAL_18;
  wire  _EVAL_42;
  wire  _EVAL_159;
  wire  _EVAL_226;
  wire  _EVAL_219;
  wire  _EVAL_244;
  wire  _EVAL_263;
  wire  _EVAL_172;
  wire  _EVAL_70;
  wire [31:0] _EVAL_131;
  wire  _EVAL_89;
  wire  _EVAL_200;
  wire  _EVAL_110;
  wire  _EVAL_141;
  wire  _EVAL_51;
  wire  _EVAL_201;
  wire  _EVAL_239;
  wire  _EVAL_188;
  wire  _EVAL_169;
  wire  _EVAL_36;
  wire  _EVAL_246;
  wire  _EVAL_198;
  wire  _EVAL_177;
  wire  _EVAL_54;
  wire  _EVAL_102;
  wire  _EVAL_132;
  wire  _EVAL_233;
  wire  _EVAL_252;
  wire  _EVAL_75;
  wire  _EVAL_116;
  wire  _EVAL_121;
  wire  _EVAL_235;
  wire  _EVAL_194;
  wire  _EVAL_73;
  wire  _EVAL_140;
  wire  _EVAL_147;
  wire  _EVAL_241;
  wire  _EVAL_183;
  wire [1:0] _EVAL_267;
  wire  _EVAL_87;
  wire  _EVAL_279;
  wire  _EVAL_278;
  wire  _EVAL_253;
  wire  _EVAL_256;
  wire  _EVAL_146;
  wire  _EVAL_27;
  wire  _EVAL_232;
  wire  _EVAL_150;
  wire  _EVAL_32;
  wire  _EVAL_48;
  wire  _EVAL_109;
  wire  _EVAL_28;
  wire  _EVAL_59;
  wire  _EVAL_24;
  wire [2:0] _EVAL_71;
  wire  _EVAL_238;
  wire  _EVAL_112;
  wire  _EVAL_152;
  wire  _EVAL_187;
  wire  _EVAL_196;
  wire  _EVAL_261;
  wire  _EVAL_199;
  wire  _EVAL_281;
  wire  _EVAL_57;
  wire  _EVAL_85;
  wire  _EVAL_247;
  wire  _EVAL_255;
  wire  _EVAL_40;
  wire  _EVAL_143;
  wire  _EVAL_33;
  wire  _EVAL_49;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_181;
  wire [1:0] _EVAL_108;
  wire  _EVAL_23;
  wire  _EVAL_83;
  wire  _EVAL_197;
  wire  _EVAL_165;
  wire  _EVAL_184;
  wire [1:0] _EVAL_58;
  wire [5:0] _EVAL_155;
  wire  _EVAL_124;
  wire  _EVAL_29;
  wire  _EVAL_130;
  wire  _EVAL_260;
  wire [2:0] _EVAL_63;
  wire [2:0] _EVAL_111;
  wire  _EVAL_270;
  wire  _EVAL_259;
  wire  _EVAL_236;
  wire  _EVAL_283;
  wire  _EVAL_206;
  wire  _EVAL_266;
  wire  _EVAL_138;
  wire  _EVAL_148;
  wire [2:0] _EVAL_175;
  wire  _EVAL_31;
  wire  _EVAL_79;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_254 = _EVAL_3 == _EVAL_52;
  assign _EVAL_276 = _EVAL_254 | _EVAL_0;
  assign _EVAL_221 = _EVAL_276 == 1'h0;
  assign _EVAL_128 = _EVAL_154 >> _EVAL_16;
  assign _EVAL_22 = _EVAL_128[0];
  assign _EVAL_106 = _EVAL_2 >= 3'h3;
  assign _EVAL_224 = _EVAL_106 | _EVAL_0;
  assign _EVAL_96 = _EVAL_224 == 1'h0;
  assign _EVAL_47 = _EVAL_2[1:0];
  assign _EVAL_207 = 4'h1 << _EVAL_47;
  assign _EVAL_84 = _EVAL_207[2:0];
  assign _EVAL_21 = _EVAL_84 | 3'h1;
  assign _EVAL_220 = _EVAL_21[1];
  assign _EVAL_211 = _EVAL[2];
  assign _EVAL_118 = _EVAL_211 == 1'h0;
  assign _EVAL_37 = _EVAL[1];
  assign _EVAL_274 = _EVAL_37 == 1'h0;
  assign _EVAL_174 = _EVAL_118 & _EVAL_274;
  assign _EVAL_193 = _EVAL_220 & _EVAL_174;
  assign _EVAL_237 = _EVAL_21[2];
  assign _EVAL_251 = _EVAL_237 & _EVAL_211;
  assign _EVAL_127 = _EVAL_106 | _EVAL_251;
  assign _EVAL_230 = _EVAL_211 & _EVAL_37;
  assign _EVAL_271 = _EVAL_220 & _EVAL_230;
  assign _EVAL_245 = _EVAL_127 | _EVAL_271;
  assign _EVAL_204 = _EVAL_21[0];
  assign _EVAL_100 = _EVAL[0];
  assign _EVAL_192 = _EVAL_230 & _EVAL_100;
  assign _EVAL_242 = _EVAL_204 & _EVAL_192;
  assign _EVAL_142 = _EVAL_245 | _EVAL_242;
  assign _EVAL_167 = _EVAL_100 == 1'h0;
  assign _EVAL_30 = _EVAL_230 & _EVAL_167;
  assign _EVAL_250 = _EVAL_204 & _EVAL_30;
  assign _EVAL_114 = _EVAL_245 | _EVAL_250;
  assign _EVAL_119 = _EVAL_211 & _EVAL_274;
  assign _EVAL_189 = _EVAL_220 & _EVAL_119;
  assign _EVAL_120 = _EVAL_127 | _EVAL_189;
  assign _EVAL_234 = _EVAL_119 & _EVAL_100;
  assign _EVAL_93 = _EVAL_204 & _EVAL_234;
  assign _EVAL_163 = _EVAL_120 | _EVAL_93;
  assign _EVAL_268 = _EVAL_119 & _EVAL_167;
  assign _EVAL_223 = _EVAL_204 & _EVAL_268;
  assign _EVAL_90 = _EVAL_120 | _EVAL_223;
  assign _EVAL_178 = _EVAL_237 & _EVAL_118;
  assign _EVAL_91 = _EVAL_106 | _EVAL_178;
  assign _EVAL_176 = _EVAL_118 & _EVAL_37;
  assign _EVAL_227 = _EVAL_220 & _EVAL_176;
  assign _EVAL_99 = _EVAL_91 | _EVAL_227;
  assign _EVAL_101 = _EVAL_176 & _EVAL_100;
  assign _EVAL_74 = _EVAL_204 & _EVAL_101;
  assign _EVAL_66 = _EVAL_99 | _EVAL_74;
  assign _EVAL_214 = _EVAL_176 & _EVAL_167;
  assign _EVAL_156 = _EVAL_204 & _EVAL_214;
  assign _EVAL_67 = _EVAL_99 | _EVAL_156;
  assign _EVAL_173 = _EVAL_91 | _EVAL_193;
  assign _EVAL_249 = _EVAL_174 & _EVAL_100;
  assign _EVAL_41 = _EVAL_204 & _EVAL_249;
  assign _EVAL_35 = _EVAL_173 | _EVAL_41;
  assign _EVAL_168 = _EVAL_174 & _EVAL_167;
  assign _EVAL_64 = _EVAL_204 & _EVAL_168;
  assign _EVAL_136 = _EVAL_173 | _EVAL_64;
  assign _EVAL_217 = {_EVAL_142,_EVAL_114,_EVAL_163,_EVAL_90,_EVAL_66,_EVAL_67,_EVAL_35,_EVAL_136};
  assign _EVAL_46 = _EVAL_15 <= 3'h2;
  assign _EVAL_171 = _EVAL_46 | _EVAL_0;
  assign _EVAL_213 = _EVAL_171 == 1'h0;
  assign _EVAL_81 = _EVAL_14 & _EVAL_8;
  assign _EVAL_144 = _EVAL_39 == 3'h0;
  assign _EVAL_195 = _EVAL_81 & _EVAL_144;
  assign _EVAL_257 = 2'h1 << _EVAL_16;
  assign _EVAL_72 = _EVAL_195 ? _EVAL_257 : 2'h0;
  assign _EVAL_228 = _EVAL_7 & _EVAL_12;
  assign _EVAL_265 = _EVAL_65 == 3'h0;
  assign _EVAL_277 = _EVAL_228 & _EVAL_265;
  assign _EVAL_86 = _EVAL_3 == 3'h6;
  assign _EVAL_20 = _EVAL_86 == 1'h0;
  assign _EVAL_205 = _EVAL_277 & _EVAL_20;
  assign _EVAL_222 = 2'h1 << _EVAL_5;
  assign _EVAL_50 = _EVAL_205 ? _EVAL_222 : 2'h0;
  assign _EVAL_78 = _EVAL_72 != _EVAL_50;
  assign _EVAL_104 = 13'h3f << _EVAL_9;
  assign _EVAL_203 = _EVAL_104[5:0];
  assign _EVAL_43 = _EVAL_1 == 1'h0;
  assign _EVAL_243 = _EVAL_43 | _EVAL_4;
  assign _EVAL_209 = _EVAL_72 | _EVAL_154;
  assign _EVAL_25 = _EVAL_209 >> _EVAL_5;
  assign _EVAL_105 = _EVAL_25[0];
  assign _EVAL_151 = _EVAL_105 | _EVAL_0;
  assign _EVAL_182 = _EVAL_151 == 1'h0;
  assign _EVAL_129 = _EVAL_1 == _EVAL_82;
  assign _EVAL_139 = _EVAL_129 | _EVAL_0;
  assign _EVAL_191 = _EVAL_139 == 1'h0;
  assign _EVAL_34 = _EVAL_15 <= 3'h4;
  assign _EVAL_60 = _EVAL_34 | _EVAL_0;
  assign _EVAL_62 = _EVAL_81 | _EVAL_228;
  assign _EVAL_272 = _EVAL_3 == 3'h0;
  assign _EVAL_115 = _EVAL_5 == _EVAL_137;
  assign _EVAL_113 = _EVAL_26 == 3'h0;
  assign _EVAL_190 = _EVAL_6 == 3'h1;
  assign _EVAL_273 = _EVAL_43 | _EVAL_0;
  assign _EVAL_94 = _EVAL_273 == 1'h0;
  assign _EVAL_282 = ~ _EVAL_217;
  assign _EVAL_117 = _EVAL_10 & _EVAL_282;
  assign _EVAL_164 = _EVAL_115 | _EVAL_0;
  assign _EVAL_17 = _EVAL_164 == 1'h0;
  assign _EVAL_280 = _EVAL_72 != 2'h0;
  assign _EVAL_38 = _EVAL_280 == 1'h0;
  assign _EVAL_215 = _EVAL_78 | _EVAL_38;
  assign _EVAL_212 = _EVAL_2 <= 3'h6;
  assign _EVAL_264 = _EVAL ^ 32'h80000000;
  assign _EVAL_161 = {1'b0,$signed(_EVAL_264)};
  assign _EVAL_218 = $signed(_EVAL_161) & $signed(-33'sh20000);
  assign _EVAL_68 = $signed(_EVAL_218);
  assign _EVAL_145 = $signed(_EVAL_68) == $signed(33'sh0);
  assign _EVAL_77 = _EVAL_212 & _EVAL_145;
  assign _EVAL_53 = _EVAL_9 == _EVAL_56;
  assign _EVAL_80 = ~ _EVAL_10;
  assign _EVAL_231 = _EVAL_80 == 8'h0;
  assign _EVAL_179 = _EVAL_231 | _EVAL_0;
  assign _EVAL_97 = _EVAL_179 == 1'h0;
  assign _EVAL_103 = _EVAL_6 == 3'h4;
  assign _EVAL_98 = _EVAL_228 & _EVAL_113;
  assign _EVAL_19 = _EVAL_6 == _EVAL_269;
  assign _EVAL_180 = _EVAL_19 | _EVAL_0;
  assign _EVAL_76 = _EVAL_215 | _EVAL_0;
  assign _EVAL_123 = _EVAL_76 == 1'h0;
  assign _EVAL_186 = _EVAL_2 == _EVAL_170;
  assign _EVAL_69 = _EVAL_6[2];
  assign _EVAL_126 = _EVAL_69 == 1'h0;
  assign _EVAL_92 = 13'h3f << _EVAL_2;
  assign _EVAL_88 = _EVAL_92[5:0];
  assign _EVAL_229 = ~ _EVAL_88;
  assign _EVAL_208 = _EVAL_229[5:3];
  assign _EVAL_225 = _EVAL_39 - 3'h1;
  assign _EVAL_149 = _EVAL_6 == 3'h3;
  assign _EVAL_157 = _EVAL_10 == _EVAL_217;
  assign _EVAL_262 = _EVAL_157 | _EVAL_0;
  assign _EVAL_122 = {{26'd0}, _EVAL_229};
  assign _EVAL_18 = _EVAL & _EVAL_122;
  assign _EVAL_42 = _EVAL_18 == 32'h0;
  assign _EVAL_159 = _EVAL_42 | _EVAL_0;
  assign _EVAL_226 = _EVAL_159 == 1'h0;
  assign _EVAL_219 = _EVAL_22 == 1'h0;
  assign _EVAL_244 = _EVAL_219 | _EVAL_0;
  assign _EVAL_263 = _EVAL_15 == _EVAL_133;
  assign _EVAL_172 = _EVAL_263 | _EVAL_0;
  assign _EVAL_70 = _EVAL_172 == 1'h0;
  assign _EVAL_131 = _EVAL_185 + 32'h1;
  assign _EVAL_89 = _EVAL == _EVAL_134;
  assign _EVAL_200 = _EVAL_162 == 3'h0;
  assign _EVAL_110 = _EVAL_81 & _EVAL_200;
  assign _EVAL_141 = _EVAL_15 <= 3'h3;
  assign _EVAL_51 = _EVAL_141 | _EVAL_0;
  assign _EVAL_201 = _EVAL_15 != 3'h0;
  assign _EVAL_239 = _EVAL_201 | _EVAL_0;
  assign _EVAL_188 = _EVAL_53 | _EVAL_0;
  assign _EVAL_169 = _EVAL_188 == 1'h0;
  assign _EVAL_36 = _EVAL_113 == 1'h0;
  assign _EVAL_246 = _EVAL_12 & _EVAL_36;
  assign _EVAL_198 = _EVAL_15 == 3'h0;
  assign _EVAL_177 = _EVAL_244 == 1'h0;
  assign _EVAL_54 = _EVAL_16 == _EVAL_248;
  assign _EVAL_102 = _EVAL_54 | _EVAL_0;
  assign _EVAL_132 = _EVAL_102 == 1'h0;
  assign _EVAL_233 = _EVAL_3 == 3'h5;
  assign _EVAL_252 = _EVAL_12 & _EVAL_233;
  assign _EVAL_75 = _EVAL_12 & _EVAL_272;
  assign _EVAL_116 = _EVAL_243 | _EVAL_0;
  assign _EVAL_121 = _EVAL_3 == 3'h4;
  assign _EVAL_235 = _EVAL_154 != 2'h0;
  assign _EVAL_194 = _EVAL_235 == 1'h0;
  assign _EVAL_73 = _EVAL_77 | _EVAL_0;
  assign _EVAL_140 = _EVAL_3[0];
  assign _EVAL_147 = _EVAL_117 == 8'h0;
  assign _EVAL_241 = _EVAL_200 == 1'h0;
  assign _EVAL_183 = _EVAL_8 & _EVAL_241;
  assign _EVAL_267 = _EVAL_154 | _EVAL_72;
  assign _EVAL_87 = _EVAL_0 == 1'h0;
  assign _EVAL_279 = _EVAL_89 | _EVAL_0;
  assign _EVAL_278 = _EVAL_279 == 1'h0;
  assign _EVAL_253 = plusarg_reader_out == 32'h0;
  assign _EVAL_256 = _EVAL_194 | _EVAL_253;
  assign _EVAL_146 = _EVAL_6 == 3'h0;
  assign _EVAL_27 = _EVAL_6 == 3'h5;
  assign _EVAL_232 = _EVAL_8 & _EVAL_27;
  assign _EVAL_150 = _EVAL_185 < plusarg_reader_out;
  assign _EVAL_32 = _EVAL_256 | _EVAL_150;
  assign _EVAL_48 = _EVAL_32 | _EVAL_0;
  assign _EVAL_109 = _EVAL_48 == 1'h0;
  assign _EVAL_28 = _EVAL_3 == 3'h2;
  assign _EVAL_59 = _EVAL_12 & _EVAL_86;
  assign _EVAL_24 = _EVAL_239 == 1'h0;
  assign _EVAL_71 = _EVAL_162 - 3'h1;
  assign _EVAL_238 = _EVAL_4 == 1'h0;
  assign _EVAL_112 = _EVAL_238 | _EVAL_0;
  assign _EVAL_152 = _EVAL_112 == 1'h0;
  assign _EVAL_187 = _EVAL_8 & _EVAL_103;
  assign _EVAL_196 = _EVAL_186 | _EVAL_0;
  assign _EVAL_261 = _EVAL_196 == 1'h0;
  assign _EVAL_199 = _EVAL_147 | _EVAL_0;
  assign _EVAL_281 = _EVAL_116 == 1'h0;
  assign _EVAL_57 = _EVAL_180 == 1'h0;
  assign _EVAL_85 = _EVAL_262 == 1'h0;
  assign _EVAL_247 = _EVAL_8 & _EVAL_190;
  assign _EVAL_255 = _EVAL_6 == 3'h7;
  assign _EVAL_40 = _EVAL_8 & _EVAL_255;
  assign _EVAL_143 = _EVAL_3 == 3'h1;
  assign _EVAL_33 = _EVAL_12 & _EVAL_143;
  assign _EVAL_49 = _EVAL_11 == 1'h0;
  assign _EVAL_44 = _EVAL_49 | _EVAL_0;
  assign _EVAL_45 = _EVAL_44 == 1'h0;
  assign _EVAL_181 = _EVAL_198 | _EVAL_0;
  assign _EVAL_108 = ~ _EVAL_50;
  assign _EVAL_23 = _EVAL_6 == 3'h2;
  assign _EVAL_83 = _EVAL_3 <= 3'h6;
  assign _EVAL_197 = _EVAL_83 | _EVAL_0;
  assign _EVAL_165 = _EVAL_197 == 1'h0;
  assign _EVAL_184 = _EVAL_181 == 1'h0;
  assign _EVAL_58 = _EVAL_267 & _EVAL_108;
  assign _EVAL_155 = ~ _EVAL_203;
  assign _EVAL_124 = _EVAL_12 & _EVAL_28;
  assign _EVAL_29 = _EVAL_9 >= 3'h3;
  assign _EVAL_130 = _EVAL_29 | _EVAL_0;
  assign _EVAL_260 = _EVAL_130 == 1'h0;
  assign _EVAL_63 = _EVAL_26 - 3'h1;
  assign _EVAL_111 = _EVAL_155[5:3];
  assign _EVAL_270 = _EVAL_8 & _EVAL_23;
  assign _EVAL_259 = _EVAL_199 == 1'h0;
  assign _EVAL_236 = _EVAL_8 & _EVAL_146;
  assign _EVAL_283 = _EVAL_51 == 1'h0;
  assign _EVAL_206 = _EVAL_6 == 3'h6;
  assign _EVAL_266 = _EVAL_8 & _EVAL_206;
  assign _EVAL_138 = _EVAL_73 == 1'h0;
  assign _EVAL_148 = _EVAL_8 & _EVAL_149;
  assign _EVAL_175 = _EVAL_65 - 3'h1;
  assign _EVAL_31 = _EVAL_12 & _EVAL_121;
  assign _EVAL_79 = _EVAL_60 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_39 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_52 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_56 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_65 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_82 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_133 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_134 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_137 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_154 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_162 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_170 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_185 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_248 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_269 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_13) begin
    if (_EVAL_0) begin
      _EVAL_26 <= 3'h0;
    end else begin
      if (_EVAL_228) begin
        if (_EVAL_113) begin
          if (_EVAL_140) begin
            _EVAL_26 <= _EVAL_111;
          end else begin
            _EVAL_26 <= 3'h0;
          end
        end else begin
          _EVAL_26 <= _EVAL_63;
        end
      end
    end
    if (_EVAL_0) begin
      _EVAL_39 <= 3'h0;
    end else begin
      if (_EVAL_81) begin
        if (_EVAL_144) begin
          if (_EVAL_126) begin
            _EVAL_39 <= _EVAL_208;
          end else begin
            _EVAL_39 <= 3'h0;
          end
        end else begin
          _EVAL_39 <= _EVAL_225;
        end
      end
    end
    if (_EVAL_98) begin
      _EVAL_52 <= _EVAL_3;
    end
    if (_EVAL_98) begin
      _EVAL_56 <= _EVAL_9;
    end
    if (_EVAL_0) begin
      _EVAL_65 <= 3'h0;
    end else begin
      if (_EVAL_228) begin
        if (_EVAL_265) begin
          if (_EVAL_140) begin
            _EVAL_65 <= _EVAL_111;
          end else begin
            _EVAL_65 <= 3'h0;
          end
        end else begin
          _EVAL_65 <= _EVAL_175;
        end
      end
    end
    if (_EVAL_98) begin
      _EVAL_82 <= _EVAL_1;
    end
    if (_EVAL_110) begin
      _EVAL_133 <= _EVAL_15;
    end
    if (_EVAL_110) begin
      _EVAL_134 <= _EVAL;
    end
    if (_EVAL_98) begin
      _EVAL_137 <= _EVAL_5;
    end
    if (_EVAL_0) begin
      _EVAL_154 <= 2'h0;
    end else begin
      _EVAL_154 <= _EVAL_58;
    end
    if (_EVAL_0) begin
      _EVAL_162 <= 3'h0;
    end else begin
      if (_EVAL_81) begin
        if (_EVAL_200) begin
          if (_EVAL_126) begin
            _EVAL_162 <= _EVAL_208;
          end else begin
            _EVAL_162 <= 3'h0;
          end
        end else begin
          _EVAL_162 <= _EVAL_71;
        end
      end
    end
    if (_EVAL_110) begin
      _EVAL_170 <= _EVAL_2;
    end
    if (_EVAL_0) begin
      _EVAL_185 <= 32'h0;
    end else begin
      if (_EVAL_62) begin
        _EVAL_185 <= 32'h0;
      end else begin
        _EVAL_185 <= _EVAL_131;
      end
    end
    if (_EVAL_110) begin
      _EVAL_248 <= _EVAL_16;
    end
    if (_EVAL_110) begin
      _EVAL_269 <= _EVAL_6;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad211e21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2020b61d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(217b1fda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc06e1be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d53c907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8960a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e333ca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a07141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52ce0e85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(755d09e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3a62b4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4a6b978)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97a3b6c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35765e19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b34d98a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80497d1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ae3ab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c88e0a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac777df8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(887c2edb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c5c7c0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49e9866b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(501810a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3b1a522)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38606243)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4ccf5c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dc4adfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85b2a0eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ce00edc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30440a8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78777c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9467a6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(741cb012)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffc12f5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93348f8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4fcf3eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(210af7fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a93377)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c43f77f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52bb05f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd19096a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(372c914)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(415f456e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82e28c1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2daf7a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(502aa5f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fef1cf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8e75e94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fce969b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8370af5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d85ea0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf57aed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4617a778)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6efab23d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee4869b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceda3794)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59a89033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86dc7dcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(681ed0fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3137070c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d437b720)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60f8c90d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c55538a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(285e18ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bffbbfaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f4f6164)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
