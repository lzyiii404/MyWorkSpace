//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_251(
  output        _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input  [24:0] _EVAL_2,
  input  [2:0]  _EVAL_3,
  output [31:0] _EVAL_4,
  output [31:0] _EVAL_5,
  output [2:0]  _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [7:0]  _EVAL_10,
  output [2:0]  _EVAL_11,
  output [3:0]  _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  output [7:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18,
  input  [31:0] _EVAL_19,
  input  [7:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  input  [2:0]  _EVAL_22,
  output [2:0]  _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  output [2:0]  _EVAL_27,
  input         _EVAL_28,
  input  [2:0]  _EVAL_29,
  output        _EVAL_30,
  output [24:0] _EVAL_31,
  output [7:0]  _EVAL_32
);
  assign _EVAL_30 = _EVAL_14;
  assign _EVAL_32 = _EVAL_10;
  assign _EVAL_21 = _EVAL_3;
  assign _EVAL_5 = _EVAL_7;
  assign _EVAL_15 = _EVAL_20;
  assign _EVAL_4 = _EVAL_19;
  assign _EVAL_12 = _EVAL_0;
  assign _EVAL_13 = _EVAL_18;
  assign _EVAL_24 = _EVAL_28;
  assign _EVAL_25 = _EVAL_26;
  assign _EVAL_11 = _EVAL_29;
  assign _EVAL_6 = _EVAL_9;
  assign _EVAL_27 = _EVAL_22;
  assign _EVAL_23 = _EVAL_17;
  assign _EVAL_31 = _EVAL_2;
  assign _EVAL = _EVAL_16;
endmodule
