//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_331_assert(
  input        _EVAL_0,
  input        _EVAL_1,
  input        _EVAL_2,
  input  [3:0] currStateReg__EVAL
);
  wire  _EVAL_98;
  wire  _EVAL_71;
  wire  _EVAL_94;
  wire  _EVAL_106;
  wire  _EVAL_109;
  wire  _EVAL_23;
  wire  _EVAL_93;
  wire  _EVAL_64;
  wire  _EVAL_55;
  wire  _EVAL_87;
  wire  _EVAL_12;
  wire  _EVAL_8;
  wire  _EVAL_97;
  wire  _EVAL_11;
  wire  _EVAL_38;
  wire  _EVAL_21;
  wire  _EVAL_83;
  wire  _EVAL_105;
  wire  _EVAL_85;
  wire  _EVAL_5;
  wire  _EVAL_68;
  wire  _EVAL_73;
  wire  _EVAL_32;
  wire  _EVAL_39;
  wire  _EVAL_100;
  wire  _EVAL_102;
  wire  _EVAL_99;
  wire  _EVAL_37;
  wire  _EVAL_52;
  wire  _EVAL_25;
  wire  _EVAL_69;
  wire  _EVAL_60;
  wire  _EVAL_107;
  wire  _EVAL_101;
  wire  _EVAL_67;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_54;
  wire  _EVAL_88;
  wire  _EVAL_81;
  wire  _EVAL_50;
  wire  _EVAL_82;
  wire  _EVAL_15;
  wire  _EVAL_92;
  wire  _EVAL_44;
  wire  _EVAL_59;
  wire  _EVAL_18;
  wire  _EVAL_65;
  wire  _EVAL_45;
  wire  _EVAL_86;
  wire  _EVAL_72;
  wire  _EVAL_40;
  wire  _EVAL_31;
  wire  _EVAL_51;
  wire  _EVAL_63;
  wire  _EVAL_77;
  wire  _EVAL_96;
  wire  _EVAL_36;
  wire  _EVAL_104;
  wire  _EVAL_22;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire  _EVAL_17;
  wire  _EVAL_103;
  wire  _EVAL_66;
  wire  _EVAL_61;
  assign _EVAL_98 = currStateReg__EVAL == 4'h3;
  assign _EVAL_71 = _EVAL_0 == 1'h0;
  assign _EVAL_94 = currStateReg__EVAL == 4'h6;
  assign _EVAL_106 = _EVAL_94 & _EVAL_71;
  assign _EVAL_109 = currStateReg__EVAL == 4'h1;
  assign _EVAL_23 = _EVAL_109 & _EVAL_1;
  assign _EVAL_93 = _EVAL_94 & _EVAL_1;
  assign _EVAL_64 = _EVAL_109 & _EVAL_0;
  assign _EVAL_55 = currStateReg__EVAL == 4'h4;
  assign _EVAL_87 = currStateReg__EVAL == 4'h2;
  assign _EVAL_12 = _EVAL_87 & _EVAL_71;
  assign _EVAL_8 = _EVAL_55 & _EVAL_71;
  assign _EVAL_97 = currStateReg__EVAL == 4'h8;
  assign _EVAL_11 = _EVAL_97 & _EVAL_0;
  assign _EVAL_38 = currStateReg__EVAL == 4'he;
  assign _EVAL_21 = _EVAL_38 & _EVAL_1;
  assign _EVAL_83 = _EVAL_87 & _EVAL_0;
  assign _EVAL_105 = currStateReg__EVAL == 4'hd;
  assign _EVAL_85 = _EVAL_105 & _EVAL_0;
  assign _EVAL_5 = currStateReg__EVAL == 4'h7;
  assign _EVAL_68 = currStateReg__EVAL == 4'h0;
  assign _EVAL_73 = _EVAL_68 & _EVAL_1;
  assign _EVAL_32 = _EVAL_97 & _EVAL_71;
  assign _EVAL_39 = _EVAL_98 & _EVAL_0;
  assign _EVAL_100 = currStateReg__EVAL == 4'h5;
  assign _EVAL_102 = _EVAL_100 & _EVAL_71;
  assign _EVAL_99 = currStateReg__EVAL == 4'h9;
  assign _EVAL_37 = _EVAL_99 & _EVAL_71;
  assign _EVAL_52 = _EVAL_1 == 1'h0;
  assign _EVAL_25 = _EVAL_97 & _EVAL_1;
  assign _EVAL_69 = _EVAL_5 & _EVAL_1;
  assign _EVAL_60 = currStateReg__EVAL == 4'hf;
  assign _EVAL_107 = _EVAL_60 & _EVAL_1;
  assign _EVAL_101 = currStateReg__EVAL == 4'ha;
  assign _EVAL_67 = _EVAL_101 & _EVAL_0;
  assign _EVAL_48 = _EVAL_68 & _EVAL_71;
  assign _EVAL_49 = _EVAL_55 & _EVAL_0;
  assign _EVAL_54 = _EVAL_105 & _EVAL_71;
  assign _EVAL_88 = _EVAL_109 & _EVAL_71;
  assign _EVAL_81 = _EVAL_5 & _EVAL_71;
  assign _EVAL_50 = _EVAL_38 & _EVAL_71;
  assign _EVAL_82 = _EVAL_105 & _EVAL_1;
  assign _EVAL_15 = currStateReg__EVAL == 4'hc;
  assign _EVAL_92 = _EVAL_15 & _EVAL_1;
  assign _EVAL_44 = _EVAL_99 & _EVAL_1;
  assign _EVAL_59 = _EVAL_101 & _EVAL_1;
  assign _EVAL_18 = _EVAL_100 & _EVAL_0;
  assign _EVAL_65 = _EVAL_15 & _EVAL_0;
  assign _EVAL_45 = currStateReg__EVAL == 4'hb;
  assign _EVAL_86 = _EVAL_98 & _EVAL_71;
  assign _EVAL_72 = _EVAL_60 & _EVAL_71;
  assign _EVAL_40 = _EVAL_98 & _EVAL_1;
  assign _EVAL_31 = _EVAL_45 & _EVAL_0;
  assign _EVAL_51 = _EVAL_38 & _EVAL_0;
  assign _EVAL_63 = _EVAL_45 & _EVAL_71;
  assign _EVAL_77 = _EVAL_101 & _EVAL_71;
  assign _EVAL_96 = _EVAL_94 & _EVAL_0;
  assign _EVAL_36 = _EVAL_68 & _EVAL_0;
  assign _EVAL_104 = _EVAL_87 & _EVAL_1;
  assign _EVAL_22 = _EVAL_55 & _EVAL_1;
  assign _EVAL_13 = _EVAL_15 & _EVAL_71;
  assign _EVAL_14 = _EVAL_60 & _EVAL_0;
  assign _EVAL_17 = _EVAL_100 & _EVAL_1;
  assign _EVAL_103 = _EVAL_5 & _EVAL_0;
  assign _EVAL_66 = _EVAL_99 & _EVAL_0;
  assign _EVAL_61 = _EVAL_45 & _EVAL_1;
  always @(posedge _EVAL_2) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc66c66f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(137aad41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(520a3eab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c53aee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(980ab8ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f38dd949)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c6abc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d82be47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f298471b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fec06801)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc55aefe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50aacde2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68d82391)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30399f4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2dd6437)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d2a545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56d8fd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e21f395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14187b10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a41ad91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1551d3d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdd36988)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b132156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(455b87c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8080518a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f2a5445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8a8ea52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(951736b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7b61e6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bec91976)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(299a9313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c52f0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33881c46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c21c23d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a12aaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a6cc042)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54f73c08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63e53b61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f75e0157)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c150c17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c08d59a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f2d3f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e0a8ee6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7132eb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c484752)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9adeae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51d6e326)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cfbd394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
