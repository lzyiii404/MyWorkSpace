//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_316_assert(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [1:0]  _EVAL_3,
  input  [31:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [6:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [2:0]  _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input  [2:0]  _EVAL_22,
  input  [7:0]  _EVAL_23,
  input         _EVAL_24,
  input  [6:0]  _EVAL_25,
  input         _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [1:0]  _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input  [2:0]  _EVAL_31,
  input  [6:0]  _EVAL_32
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_64;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_86;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_87;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_110;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_167;
  reg [31:0] _RAND_4;
  reg [6:0] _EVAL_170;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_187;
  reg [31:0] _RAND_6;
  reg [1:0] _EVAL_226;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_264;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_273;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_293;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_297;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_303;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_318;
  reg [31:0] _RAND_13;
  reg [6:0] _EVAL_337;
  reg [31:0] _RAND_14;
  reg [72:0] _EVAL_338;
  reg [95:0] _RAND_15;
  reg [31:0] _EVAL_394;
  reg [31:0] _RAND_16;
  reg [2:0] _EVAL_421;
  reg [31:0] _RAND_17;
  reg  _EVAL_427;
  reg [31:0] _RAND_18;
  reg [31:0] _EVAL_429;
  reg [31:0] _RAND_19;
  reg [1:0] _EVAL_446;
  reg [31:0] _RAND_20;
  reg [2:0] _EVAL_463;
  reg [31:0] _RAND_21;
  reg  _EVAL_467;
  reg [31:0] _RAND_22;
  reg [31:0] _EVAL_471;
  reg [31:0] _RAND_23;
  reg [2:0] _EVAL_474;
  reg [31:0] _RAND_24;
  reg [2:0] _EVAL_496;
  reg [31:0] _RAND_25;
  reg [2:0] _EVAL_514;
  reg [31:0] _RAND_26;
  reg [2:0] _EVAL_524;
  reg [31:0] _RAND_27;
  wire  _EVAL_74;
  wire  _EVAL_57;
  wire  _EVAL_362;
  wire  _EVAL_360;
  wire  _EVAL_483;
  wire [12:0] _EVAL_98;
  wire [5:0] _EVAL_500;
  wire [5:0] _EVAL_349;
  wire [2:0] _EVAL_133;
  wire [12:0] _EVAL_347;
  wire [5:0] _EVAL_343;
  wire [5:0] _EVAL_140;
  wire [31:0] _EVAL_132;
  wire  _EVAL_218;
  wire  _EVAL_184;
  wire  _EVAL_51;
  wire  _EVAL_71;
  wire  _EVAL_507;
  wire  _EVAL_254;
  wire  _EVAL_185;
  wire [3:0] _EVAL_520;
  wire  _EVAL_215;
  wire [2:0] _EVAL_213;
  wire  _EVAL_450;
  wire  _EVAL_39;
  wire  _EVAL_221;
  wire  _EVAL_91;
  wire  _EVAL_208;
  wire  _EVAL_41;
  wire  _EVAL_313;
  wire  _EVAL_510;
  wire [3:0] _EVAL_171;
  wire  _EVAL_155;
  wire  _EVAL_77;
  wire  _EVAL_212;
  wire  _EVAL_515;
  wire  _EVAL_513;
  wire [31:0] _EVAL_294;
  wire [32:0] _EVAL_419;
  wire  _EVAL_476;
  wire  _EVAL_371;
  wire  _EVAL_528;
  wire  _EVAL_237;
  wire  _EVAL_504;
  wire [127:0] _EVAL_283;
  wire [127:0] _EVAL_298;
  wire [72:0] _EVAL_484;
  wire [72:0] _EVAL_385;
  wire [72:0] _EVAL_61;
  wire [1:0] _EVAL_451;
  wire [3:0] _EVAL_304;
  wire [2:0] _EVAL_162;
  wire [2:0] _EVAL_92;
  wire  _EVAL_404;
  wire  _EVAL_384;
  wire  _EVAL_430;
  wire  _EVAL_280;
  wire  _EVAL_204;
  wire  _EVAL_325;
  wire [2:0] _EVAL_130;
  wire  _EVAL_310;
  wire  _EVAL_75;
  wire  _EVAL_351;
  wire  _EVAL_107;
  wire  _EVAL_222;
  wire  _EVAL_240;
  wire  _EVAL_458;
  wire  _EVAL_248;
  wire  _EVAL_191;
  wire  _EVAL_206;
  wire  _EVAL_411;
  wire  _EVAL_159;
  wire  _EVAL_442;
  wire  _EVAL_529;
  wire  _EVAL_139;
  wire  _EVAL_382;
  wire [31:0] _EVAL_356;
  wire [32:0] _EVAL_327;
  wire [32:0] _EVAL_83;
  wire [32:0] _EVAL_247;
  wire  _EVAL_166;
  wire  _EVAL_284;
  wire  _EVAL_375;
  wire  _EVAL_103;
  wire  _EVAL_420;
  wire  _EVAL_379;
  wire  _EVAL_109;
  wire  _EVAL_258;
  wire  _EVAL_262;
  wire [12:0] _EVAL_486;
  wire [5:0] _EVAL_111;
  wire [5:0] _EVAL_114;
  wire [2:0] _EVAL_506;
  wire [2:0] _EVAL_214;
  wire  _EVAL_516;
  wire  _EVAL_160;
  wire  _EVAL_414;
  wire  _EVAL_174;
  wire  _EVAL_241;
  wire  _EVAL_261;
  wire  _EVAL_134;
  wire  _EVAL_122;
  wire  _EVAL_246;
  wire  _EVAL_54;
  wire [31:0] _EVAL_354;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_59;
  wire  _EVAL_488;
  wire  _EVAL_499;
  wire  _EVAL_196;
  wire  _EVAL_224;
  wire  _EVAL_119;
  wire  _EVAL_357;
  wire  _EVAL_201;
  wire  _EVAL_44;
  wire  _EVAL_50;
  wire  _EVAL_282;
  wire [2:0] _EVAL_372;
  wire  _EVAL_439;
  wire  _EVAL_339;
  wire  _EVAL_152;
  wire  _EVAL_279;
  wire [72:0] _EVAL_120;
  wire  _EVAL_232;
  wire  _EVAL_377;
  wire  _EVAL_186;
  wire  _EVAL_239;
  wire  _EVAL_511;
  wire  _EVAL_126;
  wire [31:0] _EVAL_127;
  wire [32:0] _EVAL_216;
  wire [32:0] _EVAL_129;
  wire  _EVAL_183;
  wire  _EVAL_449;
  wire  _EVAL_154;
  wire  _EVAL_434;
  wire  _EVAL_412;
  wire  _EVAL_276;
  wire  _EVAL_189;
  wire  _EVAL_165;
  wire [127:0] _EVAL_522;
  wire [127:0] _EVAL_243;
  wire  _EVAL_324;
  wire  _EVAL_274;
  wire  _EVAL_457;
  wire  _EVAL_245;
  wire  _EVAL_101;
  wire  _EVAL_334;
  wire  _EVAL_436;
  wire  _EVAL_369;
  wire  _EVAL_518;
  wire  _EVAL_417;
  wire  _EVAL_350;
  wire  _EVAL_113;
  wire  _EVAL_138;
  wire  _EVAL_373;
  wire [1:0] _EVAL_527;
  wire  _EVAL_225;
  wire  _EVAL_381;
  wire  _EVAL_270;
  wire  _EVAL_358;
  wire  _EVAL_301;
  wire [31:0] _EVAL_456;
  wire  _EVAL_426;
  wire  _EVAL_255;
  wire  _EVAL_161;
  wire  _EVAL_33;
  wire  _EVAL_217;
  wire  _EVAL_190;
  wire  _EVAL_517;
  wire  _EVAL_268;
  wire  _EVAL_317;
  wire  _EVAL_141;
  wire  _EVAL_178;
  wire  _EVAL_158;
  wire  _EVAL_437;
  wire  _EVAL_38;
  wire [32:0] _EVAL_157;
  wire  _EVAL_150;
  wire  _EVAL_249;
  wire  _EVAL_195;
  wire  _EVAL_252;
  wire  _EVAL_202;
  wire  _EVAL_387;
  wire  _EVAL_308;
  wire  _EVAL_503;
  wire  _EVAL_169;
  wire  _EVAL_491;
  wire  _EVAL_401;
  wire  _EVAL_300;
  wire  _EVAL_461;
  wire [1:0] _EVAL_142;
  wire [1:0] _EVAL_316;
  wire [1:0] _EVAL_399;
  wire [1:0] _EVAL_532;
  wire  _EVAL_112;
  wire  _EVAL_365;
  wire  _EVAL_392;
  wire  _EVAL_395;
  wire  _EVAL_180;
  wire  _EVAL_331;
  wire [3:0] _EVAL_480;
  wire  _EVAL_521;
  wire  _EVAL_525;
  wire  _EVAL_207;
  wire  _EVAL_79;
  wire  _EVAL_326;
  wire  _EVAL_432;
  wire  _EVAL_231;
  wire  _EVAL_487;
  wire  _EVAL_355;
  wire  _EVAL_320;
  wire  _EVAL_403;
  wire  _EVAL_489;
  wire  _EVAL_335;
  wire  _EVAL_88;
  wire  _EVAL_305;
  wire  _EVAL_275;
  wire  _EVAL_478;
  wire  _EVAL_505;
  wire  _EVAL_497;
  wire  _EVAL_220;
  wire  _EVAL_223;
  wire  _EVAL_415;
  wire  _EVAL_361;
  wire  _EVAL_188;
  wire  _EVAL_100;
  wire  _EVAL_410;
  wire  _EVAL_508;
  wire  _EVAL_228;
  wire [7:0] _EVAL_292;
  wire  _EVAL_163;
  wire  _EVAL_42;
  wire  _EVAL_148;
  wire [7:0] _EVAL_299;
  wire  _EVAL_413;
  wire  _EVAL_182;
  wire  _EVAL_34;
  wire  _EVAL_468;
  wire  _EVAL_43;
  wire [31:0] _EVAL_192;
  wire  _EVAL_250;
  wire [2:0] _EVAL_295;
  wire  _EVAL_49;
  wire  _EVAL_69;
  wire  _EVAL_93;
  wire  _EVAL_63;
  wire  _EVAL_346;
  wire  _EVAL_495;
  wire  _EVAL_393;
  wire  _EVAL_95;
  wire [2:0] _EVAL_374;
  wire  _EVAL_378;
  wire  _EVAL_448;
  wire  _EVAL_259;
  wire  _EVAL_322;
  wire  _EVAL_70;
  wire  _EVAL_37;
  wire  _EVAL_265;
  wire  _EVAL_271;
  wire  _EVAL_323;
  wire  _EVAL_405;
  wire  _EVAL_333;
  wire  _EVAL_80;
  wire  _EVAL_330;
  wire  _EVAL_267;
  wire [1:0] _EVAL_319;
  wire [1:0] _EVAL_156;
  wire  _EVAL_48;
  wire [1:0] _EVAL_376;
  wire  _EVAL_455;
  wire  _EVAL_286;
  wire  _EVAL_153;
  wire  _EVAL_530;
  wire  _EVAL_290;
  wire  _EVAL_453;
  wire  _EVAL_523;
  wire  _EVAL_128;
  wire  _EVAL_433;
  wire  _EVAL_177;
  wire  _EVAL_102;
  wire [7:0] _EVAL_45;
  wire  _EVAL_312;
  wire  _EVAL_210;
  wire  _EVAL_229;
  wire  _EVAL_509;
  wire  _EVAL_199;
  wire  _EVAL_238;
  wire  _EVAL_76;
  wire  _EVAL_454;
  wire  _EVAL_341;
  wire [72:0] _EVAL_78;
  wire  _EVAL_125;
  wire [32:0] _EVAL_473;
  wire  _EVAL_173;
  wire  _EVAL_82;
  wire  _EVAL_251;
  wire  _EVAL_115;
  wire [2:0] _EVAL_340;
  wire  _EVAL_242;
  wire  _EVAL_435;
  wire  _EVAL_368;
  wire  _EVAL_406;
  wire  _EVAL_462;
  wire  _EVAL_197;
  wire [31:0] _EVAL_108;
  wire  _EVAL_408;
  wire  _EVAL_144;
  wire  _EVAL_464;
  wire  _EVAL_172;
  wire [2:0] _EVAL_306;
  wire  _EVAL_391;
  wire  _EVAL_176;
  wire [2:0] _EVAL_475;
  wire  _EVAL_494;
  wire  _EVAL_194;
  wire  _EVAL_502;
  wire  _EVAL_288;
  wire  _EVAL_256;
  wire  _EVAL_400;
  wire  _EVAL_47;
  wire  _EVAL_203;
  wire  _EVAL_307;
  wire  _EVAL_443;
  wire  _EVAL_131;
  wire  _EVAL_135;
  wire  _EVAL_332;
  wire  _EVAL_344;
  wire  _EVAL_418;
  wire  _EVAL_447;
  wire  _EVAL_72;
  wire  _EVAL_84;
  wire  _EVAL_117;
  wire  _EVAL_67;
  wire  _EVAL_440;
  wire  _EVAL_302;
  wire  _EVAL_329;
  wire  _EVAL_263;
  wire  _EVAL_230;
  wire  _EVAL_52;
  wire  _EVAL_470;
  wire  _EVAL_481;
  wire  _EVAL_233;
  wire  _EVAL_367;
  wire  _EVAL_235;
  wire  _EVAL_205;
  wire  _EVAL_227;
  wire  _EVAL_85;
  wire  _EVAL_272;
  wire  _EVAL_136;
  wire  _EVAL_422;
  wire [7:0] _EVAL_118;
  wire  _EVAL_370;
  wire  _EVAL_390;
  wire [2:0] _EVAL_336;
  wire  _EVAL_164;
  wire  _EVAL_168;
  wire  _EVAL_121;
  wire [31:0] _EVAL_266;
  wire  _EVAL_380;
  wire [72:0] _EVAL_423;
  wire  _EVAL_424;
  wire  _EVAL_99;
  wire  _EVAL_402;
  wire  _EVAL_143;
  wire  _EVAL_281;
  wire  _EVAL_465;
  wire  _EVAL_386;
  wire  _EVAL_81;
  wire  _EVAL_219;
  wire  _EVAL_531;
  wire  _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_363;
  wire  _EVAL_311;
  wire [32:0] _EVAL_519;
  wire  _EVAL_342;
  wire  _EVAL_73;
  wire  _EVAL_198;
  wire  _EVAL_89;
  wire  _EVAL_444;
  wire  _EVAL_60;
  wire  _EVAL_460;
  wire  _EVAL_257;
  wire  _EVAL_269;
  wire  _EVAL_431;
  wire  _EVAL_459;
  wire  _EVAL_56;
  wire  _EVAL_35;
  wire [1:0] _EVAL_53;
  wire [1:0] _EVAL_438;
  wire  _EVAL_321;
  wire  _EVAL_277;
  wire  _EVAL_234;
  wire  _EVAL_68;
  wire  _EVAL_46;
  wire  _EVAL_512;
  wire  _EVAL_364;
  wire  _EVAL_441;
  wire  _EVAL_253;
  wire  _EVAL_490;
  wire  _EVAL_62;
  wire  _EVAL_383;
  wire  _EVAL_352;
  wire  _EVAL_501;
  wire  _EVAL_328;
  wire  _EVAL_146;
  wire [2:0] _EVAL_94;
  wire  _EVAL_485;
  wire  _EVAL_285;
  wire  _EVAL_366;
  wire  _EVAL_359;
  wire  _EVAL_97;
  wire  _EVAL_416;
  wire  _EVAL_175;
  wire  _EVAL_493;
  wire  _EVAL_145;
  wire  _EVAL_309;
  wire  _EVAL_236;
  wire  _EVAL_425;
  wire  _EVAL_104;
  wire  _EVAL_181;
  wire  _EVAL_291;
  wire  _EVAL_289;
  wire  _EVAL_482;
  wire  _EVAL_55;
  wire  _EVAL_477;
  wire [72:0] _EVAL_498;
  wire  _EVAL_66;
  wire  _EVAL_123;
  wire  _EVAL_90;
  wire  _EVAL_179;
  wire  _EVAL_389;
  wire  _EVAL_353;
  wire  _EVAL_151;
  wire  _EVAL_200;
  wire [72:0] _EVAL_65;
  wire  _EVAL_278;
  wire  _EVAL_124;
  wire  _EVAL_526;
  wire  _EVAL_193;
  wire  _EVAL_452;
  wire  _EVAL_40;
  wire  _EVAL_315;
  wire  _EVAL_116;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_74 = _EVAL_30 == 1'h0;
  assign _EVAL_57 = _EVAL_5 == _EVAL_463;
  assign _EVAL_362 = _EVAL_57 | _EVAL_30;
  assign _EVAL_360 = _EVAL_22[2];
  assign _EVAL_483 = _EVAL_360 == 1'h0;
  assign _EVAL_98 = 13'h3f << _EVAL_5;
  assign _EVAL_500 = _EVAL_98[5:0];
  assign _EVAL_349 = ~ _EVAL_500;
  assign _EVAL_133 = _EVAL_349[5:3];
  assign _EVAL_347 = 13'h3f << _EVAL_11;
  assign _EVAL_343 = _EVAL_347[5:0];
  assign _EVAL_140 = ~ _EVAL_343;
  assign _EVAL_132 = {{26'd0}, _EVAL_140};
  assign _EVAL_218 = _EVAL_32 == 7'h40;
  assign _EVAL_184 = 3'h6 == _EVAL_5;
  assign _EVAL_51 = _EVAL_218 ? _EVAL_184 : 1'h0;
  assign _EVAL_71 = _EVAL_51 | _EVAL_30;
  assign _EVAL_507 = _EVAL_7 == 7'h48;
  assign _EVAL_254 = _EVAL_7 == 7'h40;
  assign _EVAL_185 = _EVAL_507 | _EVAL_254;
  assign _EVAL_520 = _EVAL_7[6:3];
  assign _EVAL_215 = _EVAL_520 == 4'h8;
  assign _EVAL_213 = _EVAL_7[2:0];
  assign _EVAL_450 = 3'h1 <= _EVAL_213;
  assign _EVAL_39 = _EVAL_215 & _EVAL_450;
  assign _EVAL_221 = _EVAL_185 | _EVAL_39;
  assign _EVAL_91 = _EVAL_7 == 7'h20;
  assign _EVAL_208 = _EVAL_221 | _EVAL_91;
  assign _EVAL_41 = _EVAL_293 == 3'h0;
  assign _EVAL_313 = _EVAL_41 == 1'h0;
  assign _EVAL_510 = _EVAL_0 & _EVAL_313;
  assign _EVAL_171 = _EVAL_25[6:3];
  assign _EVAL_155 = _EVAL_171 == 4'h8;
  assign _EVAL_77 = _EVAL_6 == _EVAL_110;
  assign _EVAL_212 = _EVAL_3 <= 2'h2;
  assign _EVAL_515 = _EVAL_212 | _EVAL_30;
  assign _EVAL_513 = _EVAL_4[2];
  assign _EVAL_294 = _EVAL_4 ^ 32'h80000000;
  assign _EVAL_419 = {1'b0,$signed(_EVAL_294)};
  assign _EVAL_476 = _EVAL_31 <= 3'h4;
  assign _EVAL_371 = _EVAL_476 | _EVAL_30;
  assign _EVAL_528 = _EVAL_24 & _EVAL_9;
  assign _EVAL_237 = _EVAL_187 == 3'h0;
  assign _EVAL_504 = _EVAL_528 & _EVAL_237;
  assign _EVAL_283 = 128'h1 << _EVAL_32;
  assign _EVAL_298 = _EVAL_504 ? _EVAL_283 : 128'h0;
  assign _EVAL_484 = _EVAL_298[72:0];
  assign _EVAL_385 = _EVAL_484 | _EVAL_338;
  assign _EVAL_61 = _EVAL_385 >> _EVAL_25;
  assign _EVAL_451 = _EVAL_5[1:0];
  assign _EVAL_304 = 4'h1 << _EVAL_451;
  assign _EVAL_162 = _EVAL_304[2:0];
  assign _EVAL_92 = _EVAL_162 | 3'h1;
  assign _EVAL_404 = _EVAL_92[2];
  assign _EVAL_384 = _EVAL_513 == 1'h0;
  assign _EVAL_430 = _EVAL_404 & _EVAL_384;
  assign _EVAL_280 = _EVAL_25 == 7'h48;
  assign _EVAL_204 = _EVAL_25 == 7'h40;
  assign _EVAL_325 = _EVAL_280 | _EVAL_204;
  assign _EVAL_130 = _EVAL_25[2:0];
  assign _EVAL_310 = 3'h1 <= _EVAL_130;
  assign _EVAL_75 = _EVAL_155 & _EVAL_310;
  assign _EVAL_351 = _EVAL_325 | _EVAL_75;
  assign _EVAL_107 = _EVAL_25 == 7'h20;
  assign _EVAL_222 = _EVAL_351 | _EVAL_107;
  assign _EVAL_240 = _EVAL_171 == 4'h0;
  assign _EVAL_458 = _EVAL_222 | _EVAL_240;
  assign _EVAL_248 = _EVAL_171 == 4'h1;
  assign _EVAL_191 = _EVAL_458 | _EVAL_248;
  assign _EVAL_206 = _EVAL_171 == 4'h2;
  assign _EVAL_411 = _EVAL_191 | _EVAL_206;
  assign _EVAL_159 = _EVAL_171 == 4'h3;
  assign _EVAL_442 = _EVAL_411 | _EVAL_159;
  assign _EVAL_529 = _EVAL_442 | _EVAL_30;
  assign _EVAL_139 = _EVAL_13 == 1'h0;
  assign _EVAL_382 = _EVAL_338 != 73'h0;
  assign _EVAL_356 = _EVAL ^ 32'h80000000;
  assign _EVAL_327 = {1'b0,$signed(_EVAL_356)};
  assign _EVAL_83 = $signed(_EVAL_327) & $signed(-33'sh20000);
  assign _EVAL_247 = $signed(_EVAL_83);
  assign _EVAL_166 = $signed(_EVAL_247) == $signed(33'sh0);
  assign _EVAL_284 = _EVAL_166 | _EVAL_30;
  assign _EVAL_375 = _EVAL_284 == 1'h0;
  assign _EVAL_103 = _EVAL_529 == 1'h0;
  assign _EVAL_420 = _EVAL_139 | _EVAL_2;
  assign _EVAL_379 = _EVAL_420 | _EVAL_30;
  assign _EVAL_109 = _EVAL_14 & _EVAL_12;
  assign _EVAL_258 = _EVAL_64 == 3'h0;
  assign _EVAL_262 = _EVAL_1[0];
  assign _EVAL_486 = 13'h3f << _EVAL_6;
  assign _EVAL_111 = _EVAL_486[5:0];
  assign _EVAL_114 = ~ _EVAL_111;
  assign _EVAL_506 = _EVAL_114[5:3];
  assign _EVAL_214 = _EVAL_64 - 3'h1;
  assign _EVAL_516 = _EVAL_6 >= 3'h3;
  assign _EVAL_160 = _EVAL_516 | _EVAL_30;
  assign _EVAL_414 = _EVAL_160 == 1'h0;
  assign _EVAL_174 = _EVAL_139 | _EVAL_30;
  assign _EVAL_241 = _EVAL_174 == 1'h0;
  assign _EVAL_261 = _EVAL_474 == 3'h0;
  assign _EVAL_134 = _EVAL_261 == 1'h0;
  assign _EVAL_122 = _EVAL_1 == _EVAL_524;
  assign _EVAL_246 = _EVAL_3 == _EVAL_226;
  assign _EVAL_54 = _EVAL_246 | _EVAL_30;
  assign _EVAL_354 = _EVAL_429 + 32'h1;
  assign _EVAL_105 = _EVAL_167 == 3'h0;
  assign _EVAL_106 = _EVAL_105 == 1'h0;
  assign _EVAL_59 = _EVAL_9 & _EVAL_106;
  assign _EVAL_488 = _EVAL_18 == 3'h1;
  assign _EVAL_499 = _EVAL_21 & _EVAL_488;
  assign _EVAL_196 = _EVAL_1 == 3'h0;
  assign _EVAL_224 = _EVAL_92[1];
  assign _EVAL_119 = _EVAL_4[1];
  assign _EVAL_357 = _EVAL_513 & _EVAL_119;
  assign _EVAL_201 = _EVAL_224 & _EVAL_357;
  assign _EVAL_44 = 3'h6 == _EVAL_11;
  assign _EVAL_50 = _EVAL_254 ? _EVAL_44 : 1'h0;
  assign _EVAL_282 = _EVAL_484 != 73'h0;
  assign _EVAL_372 = _EVAL_87 - 3'h1;
  assign _EVAL_439 = _EVAL_18 == 3'h5;
  assign _EVAL_339 = _EVAL_21 & _EVAL_439;
  assign _EVAL_152 = _EVAL_371 == 1'h0;
  assign _EVAL_279 = _EVAL_528 & _EVAL_105;
  assign _EVAL_120 = _EVAL_338 >> _EVAL_32;
  assign _EVAL_232 = _EVAL_120[0];
  assign _EVAL_377 = _EVAL_232 == 1'h0;
  assign _EVAL_186 = _EVAL_362 == 1'h0;
  assign _EVAL_239 = _EVAL_87 == 3'h0;
  assign _EVAL_511 = _EVAL_1 == 3'h1;
  assign _EVAL_126 = _EVAL_12 & _EVAL_511;
  assign _EVAL_127 = _EVAL_27 ^ 32'h80000000;
  assign _EVAL_216 = {1'b0,$signed(_EVAL_127)};
  assign _EVAL_129 = $signed(_EVAL_216) & $signed(-33'sh20000);
  assign _EVAL_183 = _EVAL_15 == 1'h0;
  assign _EVAL_449 = _EVAL_183 | _EVAL_30;
  assign _EVAL_154 = _EVAL_22 == 3'h0;
  assign _EVAL_434 = _EVAL_9 & _EVAL_154;
  assign _EVAL_412 = _EVAL_109 & _EVAL_258;
  assign _EVAL_276 = _EVAL_1 == 3'h6;
  assign _EVAL_189 = _EVAL_276 == 1'h0;
  assign _EVAL_165 = _EVAL_412 & _EVAL_189;
  assign _EVAL_522 = 128'h1 << _EVAL_25;
  assign _EVAL_243 = _EVAL_165 ? _EVAL_522 : 128'h0;
  assign _EVAL_324 = _EVAL_18 == _EVAL_421;
  assign _EVAL_274 = _EVAL_324 | _EVAL_30;
  assign _EVAL_457 = _EVAL_5 >= 3'h3;
  assign _EVAL_245 = _EVAL_404 & _EVAL_513;
  assign _EVAL_101 = _EVAL_457 | _EVAL_245;
  assign _EVAL_334 = _EVAL_119 == 1'h0;
  assign _EVAL_436 = _EVAL_513 & _EVAL_334;
  assign _EVAL_369 = _EVAL_224 & _EVAL_436;
  assign _EVAL_518 = _EVAL_101 | _EVAL_369;
  assign _EVAL_417 = _EVAL_92[0];
  assign _EVAL_350 = _EVAL_4[0];
  assign _EVAL_113 = _EVAL_436 & _EVAL_350;
  assign _EVAL_138 = _EVAL_417 & _EVAL_113;
  assign _EVAL_373 = _EVAL_518 | _EVAL_138;
  assign _EVAL_527 = 2'h1 << _EVAL_17;
  assign _EVAL_225 = _EVAL_16 == _EVAL_303;
  assign _EVAL_381 = _EVAL_122 | _EVAL_30;
  assign _EVAL_270 = _EVAL_381 == 1'h0;
  assign _EVAL_358 = _EVAL_20 == _EVAL_427;
  assign _EVAL_301 = _EVAL_358 | _EVAL_30;
  assign _EVAL_456 = _EVAL & 32'h3f;
  assign _EVAL_426 = _EVAL_382 == 1'h0;
  assign _EVAL_255 = plusarg_reader_out == 32'h0;
  assign _EVAL_161 = _EVAL_426 | _EVAL_255;
  assign _EVAL_33 = _EVAL_429 < plusarg_reader_out;
  assign _EVAL_217 = _EVAL_161 | _EVAL_33;
  assign _EVAL_190 = _EVAL_217 | _EVAL_30;
  assign _EVAL_517 = _EVAL == _EVAL_394;
  assign _EVAL_268 = _EVAL_22 == 3'h1;
  assign _EVAL_317 = _EVAL_9 & _EVAL_268;
  assign _EVAL_141 = _EVAL_101 | _EVAL_201;
  assign _EVAL_178 = _EVAL_350 == 1'h0;
  assign _EVAL_158 = _EVAL_357 & _EVAL_178;
  assign _EVAL_437 = _EVAL_417 & _EVAL_158;
  assign _EVAL_38 = _EVAL_141 | _EVAL_437;
  assign _EVAL_157 = $signed(_EVAL_419) & $signed(-33'sh20000);
  assign _EVAL_150 = _EVAL_16 <= 3'h5;
  assign _EVAL_249 = _EVAL_150 | _EVAL_30;
  assign _EVAL_195 = _EVAL_249 == 1'h0;
  assign _EVAL_252 = _EVAL_28 == 2'h0;
  assign _EVAL_202 = _EVAL_252 | _EVAL_30;
  assign _EVAL_387 = _EVAL_202 == 1'h0;
  assign _EVAL_308 = _EVAL_514 == 3'h0;
  assign _EVAL_503 = _EVAL_109 & _EVAL_308;
  assign _EVAL_169 = _EVAL_1[2];
  assign _EVAL_491 = _EVAL_1[1];
  assign _EVAL_401 = _EVAL_491 == 1'h0;
  assign _EVAL_300 = _EVAL_169 & _EVAL_401;
  assign _EVAL_461 = _EVAL_503 & _EVAL_300;
  assign _EVAL_142 = 2'h1 << _EVAL_20;
  assign _EVAL_316 = _EVAL_461 ? _EVAL_142 : 2'h0;
  assign _EVAL_399 = _EVAL_316 | _EVAL_297;
  assign _EVAL_532 = _EVAL_399 >> _EVAL_17;
  assign _EVAL_112 = _EVAL_532[0];
  assign _EVAL_365 = _EVAL_112 | _EVAL_30;
  assign _EVAL_392 = _EVAL_365 == 1'h0;
  assign _EVAL_395 = _EVAL_28 == _EVAL_446;
  assign _EVAL_180 = _EVAL_395 | _EVAL_30;
  assign _EVAL_331 = _EVAL_180 == 1'h0;
  assign _EVAL_480 = _EVAL_32[6:3];
  assign _EVAL_521 = _EVAL_480 == 4'h8;
  assign _EVAL_525 = _EVAL_520 == 4'h0;
  assign _EVAL_207 = _EVAL_208 | _EVAL_525;
  assign _EVAL_79 = _EVAL_384 & _EVAL_334;
  assign _EVAL_326 = _EVAL_224 & _EVAL_79;
  assign _EVAL_432 = _EVAL_357 & _EVAL_350;
  assign _EVAL_231 = _EVAL_417 & _EVAL_432;
  assign _EVAL_487 = _EVAL_141 | _EVAL_231;
  assign _EVAL_355 = _EVAL_436 & _EVAL_178;
  assign _EVAL_320 = _EVAL_417 & _EVAL_355;
  assign _EVAL_403 = _EVAL_518 | _EVAL_320;
  assign _EVAL_489 = _EVAL_457 | _EVAL_430;
  assign _EVAL_335 = _EVAL_384 & _EVAL_119;
  assign _EVAL_88 = _EVAL_224 & _EVAL_335;
  assign _EVAL_305 = _EVAL_489 | _EVAL_88;
  assign _EVAL_275 = _EVAL_335 & _EVAL_350;
  assign _EVAL_478 = _EVAL_417 & _EVAL_275;
  assign _EVAL_505 = _EVAL_305 | _EVAL_478;
  assign _EVAL_497 = _EVAL_335 & _EVAL_178;
  assign _EVAL_220 = _EVAL_417 & _EVAL_497;
  assign _EVAL_223 = _EVAL_305 | _EVAL_220;
  assign _EVAL_415 = _EVAL_489 | _EVAL_326;
  assign _EVAL_361 = _EVAL_79 & _EVAL_350;
  assign _EVAL_188 = _EVAL_417 & _EVAL_361;
  assign _EVAL_100 = _EVAL_415 | _EVAL_188;
  assign _EVAL_410 = _EVAL_79 & _EVAL_178;
  assign _EVAL_508 = _EVAL_417 & _EVAL_410;
  assign _EVAL_228 = _EVAL_415 | _EVAL_508;
  assign _EVAL_292 = {_EVAL_487,_EVAL_38,_EVAL_373,_EVAL_403,_EVAL_505,_EVAL_223,_EVAL_100,_EVAL_228};
  assign _EVAL_163 = _EVAL_23 == _EVAL_292;
  assign _EVAL_42 = _EVAL_25 == _EVAL_170;
  assign _EVAL_148 = _EVAL_31 <= 3'h2;
  assign _EVAL_299 = ~ _EVAL_292;
  assign _EVAL_413 = _EVAL_54 == 1'h0;
  assign _EVAL_182 = _EVAL_456 == 32'h0;
  assign _EVAL_34 = _EVAL_182 | _EVAL_30;
  assign _EVAL_468 = _EVAL_16 == 3'h0;
  assign _EVAL_43 = _EVAL_468 | _EVAL_30;
  assign _EVAL_192 = _EVAL_27 & _EVAL_132;
  assign _EVAL_250 = _EVAL_192 == 32'h0;
  assign _EVAL_295 = _EVAL_140[5:3];
  assign _EVAL_49 = _EVAL_31 != 3'h0;
  assign _EVAL_69 = _EVAL_49 | _EVAL_30;
  assign _EVAL_93 = _EVAL_69 == 1'h0;
  assign _EVAL_63 = _EVAL_28 <= 2'h2;
  assign _EVAL_346 = _EVAL_63 | _EVAL_30;
  assign _EVAL_495 = _EVAL_346 == 1'h0;
  assign _EVAL_393 = _EVAL_32 == 7'h48;
  assign _EVAL_95 = _EVAL_393 | _EVAL_218;
  assign _EVAL_374 = _EVAL_32[2:0];
  assign _EVAL_378 = 3'h1 <= _EVAL_374;
  assign _EVAL_448 = _EVAL_521 & _EVAL_378;
  assign _EVAL_259 = _EVAL_95 | _EVAL_448;
  assign _EVAL_322 = _EVAL_32 == 7'h20;
  assign _EVAL_70 = _EVAL_259 | _EVAL_322;
  assign _EVAL_37 = _EVAL_480 == 4'h0;
  assign _EVAL_265 = _EVAL_70 | _EVAL_37;
  assign _EVAL_271 = _EVAL_480 == 4'h1;
  assign _EVAL_323 = _EVAL_265 | _EVAL_271;
  assign _EVAL_405 = _EVAL_480 == 4'h2;
  assign _EVAL_333 = _EVAL_323 | _EVAL_405;
  assign _EVAL_80 = _EVAL_480 == 4'h3;
  assign _EVAL_330 = _EVAL_333 | _EVAL_80;
  assign _EVAL_267 = _EVAL_330 | _EVAL_30;
  assign _EVAL_319 = _EVAL_10 ? _EVAL_527 : 2'h0;
  assign _EVAL_156 = ~ _EVAL_319;
  assign _EVAL_48 = _EVAL_31 == _EVAL_496;
  assign _EVAL_376 = _EVAL_297 >> _EVAL_20;
  assign _EVAL_455 = _EVAL_376[0];
  assign _EVAL_286 = _EVAL_449 == 1'h0;
  assign _EVAL_153 = _EVAL_18 == 3'h4;
  assign _EVAL_530 = _EVAL_12 & _EVAL_196;
  assign _EVAL_290 = _EVAL_520 == 4'h1;
  assign _EVAL_453 = _EVAL_207 | _EVAL_290;
  assign _EVAL_523 = _EVAL_520 == 4'h2;
  assign _EVAL_128 = _EVAL_453 | _EVAL_523;
  assign _EVAL_433 = _EVAL_520 == 4'h3;
  assign _EVAL_177 = _EVAL_128 | _EVAL_433;
  assign _EVAL_102 = _EVAL_177 | _EVAL_30;
  assign _EVAL_45 = ~ _EVAL_23;
  assign _EVAL_312 = _EVAL_45 == 8'h0;
  assign _EVAL_210 = _EVAL_8 & _EVAL_0;
  assign _EVAL_229 = _EVAL_11 >= 3'h3;
  assign _EVAL_509 = _EVAL_229 | _EVAL_30;
  assign _EVAL_199 = _EVAL_509 == 1'h0;
  assign _EVAL_238 = _EVAL_239 == 1'h0;
  assign _EVAL_76 = _EVAL_12 & _EVAL_238;
  assign _EVAL_454 = _EVAL_109 & _EVAL_239;
  assign _EVAL_341 = _EVAL_18 == 3'h6;
  assign _EVAL_78 = _EVAL_243[72:0];
  assign _EVAL_125 = _EVAL_71 == 1'h0;
  assign _EVAL_473 = $signed(_EVAL_129);
  assign _EVAL_173 = $signed(_EVAL_473) == $signed(33'sh0);
  assign _EVAL_82 = _EVAL_173 | _EVAL_30;
  assign _EVAL_251 = _EVAL_82 == 1'h0;
  assign _EVAL_115 = _EVAL_22 == 3'h5;
  assign _EVAL_340 = _EVAL_187 - 3'h1;
  assign _EVAL_242 = _EVAL_31 == 3'h0;
  assign _EVAL_435 = _EVAL_484 != _EVAL_78;
  assign _EVAL_368 = _EVAL_282 == 1'h0;
  assign _EVAL_406 = _EVAL_435 | _EVAL_368;
  assign _EVAL_462 = _EVAL_406 | _EVAL_30;
  assign _EVAL_197 = _EVAL_462 == 1'h0;
  assign _EVAL_108 = {{26'd0}, _EVAL_349};
  assign _EVAL_408 = _EVAL_18 == 3'h0;
  assign _EVAL_144 = _EVAL_250 | _EVAL_30;
  assign _EVAL_464 = _EVAL_144 == 1'h0;
  assign _EVAL_172 = _EVAL_21 & _EVAL_341;
  assign _EVAL_306 = _EVAL_293 - 3'h1;
  assign _EVAL_391 = _EVAL_18 == 3'h7;
  assign _EVAL_176 = _EVAL_21 & _EVAL_391;
  assign _EVAL_475 = _EVAL_167 - 3'h1;
  assign _EVAL_494 = _EVAL_77 | _EVAL_30;
  assign _EVAL_194 = _EVAL_102 == 1'h0;
  assign _EVAL_502 = _EVAL_455 == 1'h0;
  assign _EVAL_288 = _EVAL_502 | _EVAL_30;
  assign _EVAL_256 = _EVAL_288 == 1'h0;
  assign _EVAL_400 = _EVAL_18[0];
  assign _EVAL_47 = _EVAL_515 == 1'h0;
  assign _EVAL_203 = _EVAL_43 == 1'h0;
  assign _EVAL_307 = _EVAL_16 <= 3'h2;
  assign _EVAL_443 = _EVAL_61[0];
  assign _EVAL_131 = _EVAL_443 | _EVAL_30;
  assign _EVAL_135 = _EVAL_131 == 1'h0;
  assign _EVAL_332 = _EVAL_1 <= 3'h6;
  assign _EVAL_344 = _EVAL_332 | _EVAL_30;
  assign _EVAL_418 = _EVAL_344 == 1'h0;
  assign _EVAL_447 = _EVAL_4 == _EVAL_471;
  assign _EVAL_72 = _EVAL_19 & _EVAL_21;
  assign _EVAL_84 = _EVAL_11 <= 3'h6;
  assign _EVAL_117 = _EVAL_84 & _EVAL_173;
  assign _EVAL_67 = _EVAL_117 | _EVAL_30;
  assign _EVAL_440 = _EVAL_2 == 1'h0;
  assign _EVAL_302 = _EVAL_440 | _EVAL_30;
  assign _EVAL_329 = _EVAL_447 | _EVAL_30;
  assign _EVAL_263 = _EVAL_329 == 1'h0;
  assign _EVAL_230 = _EVAL_1 == 3'h4;
  assign _EVAL_52 = _EVAL_22 == 3'h6;
  assign _EVAL_470 = _EVAL_21 & _EVAL_408;
  assign _EVAL_481 = _EVAL_28 != 2'h2;
  assign _EVAL_233 = _EVAL_13 == _EVAL_467;
  assign _EVAL_367 = _EVAL_7 == _EVAL_337;
  assign _EVAL_235 = _EVAL_367 | _EVAL_30;
  assign _EVAL_205 = _EVAL_235 == 1'h0;
  assign _EVAL_227 = _EVAL_27 == _EVAL_318;
  assign _EVAL_85 = _EVAL_227 | _EVAL_30;
  assign _EVAL_272 = _EVAL_85 == 1'h0;
  assign _EVAL_136 = _EVAL_9 & _EVAL_115;
  assign _EVAL_422 = _EVAL_307 | _EVAL_30;
  assign _EVAL_118 = _EVAL_23 & _EVAL_299;
  assign _EVAL_370 = _EVAL_118 == 8'h0;
  assign _EVAL_390 = _EVAL_370 | _EVAL_30;
  assign _EVAL_336 = _EVAL_514 - 3'h1;
  assign _EVAL_164 = _EVAL_32 == _EVAL_86;
  assign _EVAL_168 = _EVAL_164 | _EVAL_30;
  assign _EVAL_121 = _EVAL_168 == 1'h0;
  assign _EVAL_266 = _EVAL_4 & _EVAL_108;
  assign _EVAL_380 = _EVAL_266 == 32'h0;
  assign _EVAL_423 = ~ _EVAL_78;
  assign _EVAL_424 = _EVAL_31 <= 3'h3;
  assign _EVAL_99 = _EVAL_233 | _EVAL_30;
  assign _EVAL_402 = _EVAL_302 == 1'h0;
  assign _EVAL_143 = _EVAL_380 | _EVAL_30;
  assign _EVAL_281 = _EVAL_143 == 1'h0;
  assign _EVAL_465 = _EVAL_1 == 3'h2;
  assign _EVAL_386 = _EVAL_22 == _EVAL_264;
  assign _EVAL_81 = _EVAL_386 | _EVAL_30;
  assign _EVAL_219 = _EVAL_81 == 1'h0;
  assign _EVAL_531 = _EVAL_22 == 3'h7;
  assign _EVAL_396 = _EVAL_9 & _EVAL_531;
  assign _EVAL_397 = _EVAL_12 & _EVAL_230;
  assign _EVAL_363 = _EVAL_190 == 1'h0;
  assign _EVAL_311 = _EVAL_5 <= 3'h6;
  assign _EVAL_519 = $signed(_EVAL_157);
  assign _EVAL_342 = $signed(_EVAL_519) == $signed(33'sh0);
  assign _EVAL_73 = _EVAL_311 & _EVAL_342;
  assign _EVAL_198 = _EVAL_73 | _EVAL_30;
  assign _EVAL_89 = _EVAL_481 | _EVAL_30;
  assign _EVAL_444 = _EVAL_89 == 1'h0;
  assign _EVAL_60 = _EVAL_457 | _EVAL_30;
  assign _EVAL_460 = _EVAL_60 == 1'h0;
  assign _EVAL_257 = _EVAL_42 | _EVAL_30;
  assign _EVAL_269 = _EVAL_528 | _EVAL_109;
  assign _EVAL_431 = _EVAL_225 | _EVAL_30;
  assign _EVAL_459 = _EVAL_431 == 1'h0;
  assign _EVAL_56 = _EVAL_11 == _EVAL_273;
  assign _EVAL_35 = _EVAL_22 == 3'h3;
  assign _EVAL_53 = _EVAL_297 | _EVAL_316;
  assign _EVAL_438 = _EVAL_53 & _EVAL_156;
  assign _EVAL_321 = _EVAL_379 == 1'h0;
  assign _EVAL_277 = _EVAL_50 | _EVAL_30;
  assign _EVAL_234 = _EVAL_277 == 1'h0;
  assign _EVAL_68 = _EVAL_72 & _EVAL_261;
  assign _EVAL_46 = _EVAL_18 == 3'h2;
  assign _EVAL_512 = _EVAL_21 & _EVAL_46;
  assign _EVAL_364 = _EVAL_148 | _EVAL_30;
  assign _EVAL_441 = _EVAL_364 == 1'h0;
  assign _EVAL_253 = _EVAL_424 | _EVAL_30;
  assign _EVAL_490 = _EVAL_422 == 1'h0;
  assign _EVAL_62 = _EVAL_22 == 3'h4;
  assign _EVAL_383 = _EVAL_9 & _EVAL_62;
  assign _EVAL_352 = _EVAL_267 == 1'h0;
  assign _EVAL_501 = _EVAL_29 == 1'h0;
  assign _EVAL_328 = _EVAL_501 | _EVAL_30;
  assign _EVAL_146 = _EVAL_328 == 1'h0;
  assign _EVAL_94 = _EVAL_474 - 3'h1;
  assign _EVAL_485 = _EVAL_1 == 3'h5;
  assign _EVAL_285 = _EVAL_257 == 1'h0;
  assign _EVAL_366 = _EVAL_163 | _EVAL_30;
  assign _EVAL_359 = _EVAL_48 | _EVAL_30;
  assign _EVAL_97 = _EVAL_359 == 1'h0;
  assign _EVAL_416 = _EVAL_242 | _EVAL_30;
  assign _EVAL_175 = _EVAL_416 == 1'h0;
  assign _EVAL_493 = _EVAL_99 == 1'h0;
  assign _EVAL_145 = _EVAL_12 & _EVAL_465;
  assign _EVAL_309 = _EVAL_301 == 1'h0;
  assign _EVAL_236 = _EVAL_56 | _EVAL_30;
  assign _EVAL_425 = _EVAL_236 == 1'h0;
  assign _EVAL_104 = _EVAL_67 == 1'h0;
  assign _EVAL_181 = _EVAL_21 & _EVAL_134;
  assign _EVAL_291 = _EVAL_517 | _EVAL_30;
  assign _EVAL_289 = _EVAL_198 == 1'h0;
  assign _EVAL_482 = _EVAL_9 & _EVAL_52;
  assign _EVAL_55 = _EVAL_253 == 1'h0;
  assign _EVAL_477 = _EVAL_9 & _EVAL_35;
  assign _EVAL_498 = _EVAL_338 | _EVAL_484;
  assign _EVAL_66 = _EVAL_312 | _EVAL_30;
  assign _EVAL_123 = _EVAL_66 == 1'h0;
  assign _EVAL_90 = _EVAL_377 | _EVAL_30;
  assign _EVAL_179 = _EVAL_12 & _EVAL_276;
  assign _EVAL_389 = _EVAL_22 == 3'h2;
  assign _EVAL_353 = _EVAL_494 == 1'h0;
  assign _EVAL_151 = _EVAL_366 == 1'h0;
  assign _EVAL_200 = _EVAL_12 & _EVAL_485;
  assign _EVAL_65 = _EVAL_498 & _EVAL_423;
  assign _EVAL_278 = _EVAL_274 == 1'h0;
  assign _EVAL_124 = _EVAL_21 & _EVAL_153;
  assign _EVAL_526 = _EVAL_390 == 1'h0;
  assign _EVAL_193 = _EVAL_9 & _EVAL_389;
  assign _EVAL_452 = _EVAL_34 == 1'h0;
  assign _EVAL_40 = _EVAL_90 == 1'h0;
  assign _EVAL_315 = _EVAL_210 & _EVAL_41;
  assign _EVAL_116 = _EVAL_291 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_64 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_86 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_87 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_110 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_167 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_170 = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_187 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_226 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_264 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_273 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_293 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_297 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_303 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_318 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_337 = _RAND_14[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {3{`RANDOM}};
  _EVAL_338 = _RAND_15[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_394 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_421 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_427 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_429 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_446 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_463 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_467 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_471 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_474 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_496 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_514 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_524 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_26) begin
    if (_EVAL_30) begin
      _EVAL_64 <= 3'h0;
    end else begin
      if (_EVAL_109) begin
        if (_EVAL_258) begin
          if (_EVAL_262) begin
            _EVAL_64 <= _EVAL_506;
          end else begin
            _EVAL_64 <= 3'h0;
          end
        end else begin
          _EVAL_64 <= _EVAL_214;
        end
      end
    end
    if (_EVAL_279) begin
      _EVAL_86 <= _EVAL_32;
    end
    if (_EVAL_30) begin
      _EVAL_87 <= 3'h0;
    end else begin
      if (_EVAL_109) begin
        if (_EVAL_239) begin
          if (_EVAL_262) begin
            _EVAL_87 <= _EVAL_506;
          end else begin
            _EVAL_87 <= 3'h0;
          end
        end else begin
          _EVAL_87 <= _EVAL_372;
        end
      end
    end
    if (_EVAL_454) begin
      _EVAL_110 <= _EVAL_6;
    end
    if (_EVAL_30) begin
      _EVAL_167 <= 3'h0;
    end else begin
      if (_EVAL_528) begin
        if (_EVAL_105) begin
          if (_EVAL_483) begin
            _EVAL_167 <= _EVAL_133;
          end else begin
            _EVAL_167 <= 3'h0;
          end
        end else begin
          _EVAL_167 <= _EVAL_475;
        end
      end
    end
    if (_EVAL_454) begin
      _EVAL_170 <= _EVAL_25;
    end
    if (_EVAL_30) begin
      _EVAL_187 <= 3'h0;
    end else begin
      if (_EVAL_528) begin
        if (_EVAL_237) begin
          if (_EVAL_483) begin
            _EVAL_187 <= _EVAL_133;
          end else begin
            _EVAL_187 <= 3'h0;
          end
        end else begin
          _EVAL_187 <= _EVAL_340;
        end
      end
    end
    if (_EVAL_315) begin
      _EVAL_226 <= _EVAL_3;
    end
    if (_EVAL_279) begin
      _EVAL_264 <= _EVAL_22;
    end
    if (_EVAL_68) begin
      _EVAL_273 <= _EVAL_11;
    end
    if (_EVAL_30) begin
      _EVAL_293 <= 3'h0;
    end else begin
      if (_EVAL_210) begin
        if (_EVAL_41) begin
          _EVAL_293 <= 3'h0;
        end else begin
          _EVAL_293 <= _EVAL_306;
        end
      end
    end
    if (_EVAL_30) begin
      _EVAL_297 <= 2'h0;
    end else begin
      _EVAL_297 <= _EVAL_438;
    end
    if (_EVAL_68) begin
      _EVAL_303 <= _EVAL_16;
    end
    if (_EVAL_68) begin
      _EVAL_318 <= _EVAL_27;
    end
    if (_EVAL_68) begin
      _EVAL_337 <= _EVAL_7;
    end
    if (_EVAL_30) begin
      _EVAL_338 <= 73'h0;
    end else begin
      _EVAL_338 <= _EVAL_65;
    end
    if (_EVAL_315) begin
      _EVAL_394 <= _EVAL;
    end
    if (_EVAL_68) begin
      _EVAL_421 <= _EVAL_18;
    end
    if (_EVAL_454) begin
      _EVAL_427 <= _EVAL_20;
    end
    if (_EVAL_30) begin
      _EVAL_429 <= 32'h0;
    end else begin
      if (_EVAL_269) begin
        _EVAL_429 <= 32'h0;
      end else begin
        _EVAL_429 <= _EVAL_354;
      end
    end
    if (_EVAL_454) begin
      _EVAL_446 <= _EVAL_28;
    end
    if (_EVAL_279) begin
      _EVAL_463 <= _EVAL_5;
    end
    if (_EVAL_454) begin
      _EVAL_467 <= _EVAL_13;
    end
    if (_EVAL_279) begin
      _EVAL_471 <= _EVAL_4;
    end
    if (_EVAL_30) begin
      _EVAL_474 <= 3'h0;
    end else begin
      if (_EVAL_72) begin
        if (_EVAL_261) begin
          if (_EVAL_400) begin
            _EVAL_474 <= _EVAL_295;
          end else begin
            _EVAL_474 <= 3'h0;
          end
        end else begin
          _EVAL_474 <= _EVAL_94;
        end
      end
    end
    if (_EVAL_279) begin
      _EVAL_496 <= _EVAL_31;
    end
    if (_EVAL_30) begin
      _EVAL_514 <= 3'h0;
    end else begin
      if (_EVAL_109) begin
        if (_EVAL_308) begin
          if (_EVAL_262) begin
            _EVAL_514 <= _EVAL_506;
          end else begin
            _EVAL_514 <= 3'h0;
          end
        end else begin
          _EVAL_514 <= _EVAL_336;
        end
      end
    end
    if (_EVAL_454) begin
      _EVAL_524 <= _EVAL_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_414) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e57bd212)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53ddb67d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aca80f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29b99d32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eae16b50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_495) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6764594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae6aff0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6f3fa55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95643d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e798a54f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5daa2b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a326b3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_414) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(657d278a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_402) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15043e52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_414) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61c8cbc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7384e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_375) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cdda73e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(911070e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6befe919)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_460) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38035396)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_495) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eec92f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a61d7b5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9a70538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40519f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66bcef52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_490) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f61e634a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51a587a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_387) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(958b188e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_452) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f63aea14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d59114c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2aca051)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_402) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4031e19a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac01f130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df8ba527)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(890d636a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_504 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c63bce35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(625a58bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_402) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aa5f1f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5ebfbd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d42942a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ba4103)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c1a99f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_441) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eb92ec2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_452) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14795818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f59debac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_460) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397fe997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_402) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c822545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_414) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe848bfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6511ca9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f4e0e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e07f94fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_375) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3accc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_414) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95e1d9a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57f27c82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d92f2186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_413) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(776a72fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87ee1f6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24eb546b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_460) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92128005)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d51f8d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c7f2d6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d738250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da8c9372)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57397855)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c201020c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d61146)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_413) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6e62bdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74129b24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_495) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44474e55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88c22c61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_493) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ec7c5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81951cb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_441) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a3867f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_402) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fe9a6ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce31e825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6a38ffc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_441) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(947a2593)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9319fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_392) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e1bc6a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddb9f080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25dbaddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fba6389)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_459) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e6aba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afac83bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4a64397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_493) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96eb3b12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab3823f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73c12f5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e606440b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_418) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1f54428)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba7cbfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_495) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e474caa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df2291c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18771d50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb0fc821)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0eb1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_392) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c64455f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_387) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1adb6931)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abaf1da0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f8e76fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0c266f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1545b4e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_460) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b80d9309)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_526) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6da28182)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8a946e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2822d6e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9ff69ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e2c445e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0f92e9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7db7579b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_504 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_402) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c7c4eb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_402) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_414) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_459) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(207c2b71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_387) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9b7fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0b9dad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_402) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(405d698c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4a4cd1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8fd7e50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5330b7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_434 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4f01f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_464) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_490) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(275970ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69f0ddd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd307d6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70012b2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d10f0dd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7563aac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_490) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_425) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(305ce7b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e003a95f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90ed25e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_418) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_363) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5056857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_441) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_526) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4971899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd2231fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191cfef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_387) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc07021f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb402ae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39c1ba7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_490) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_499 & _EVAL_464) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fca129a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_425) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b58e603)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f551c2e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
