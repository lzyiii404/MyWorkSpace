//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_115_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [6:0]  _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [6:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [29:0] _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_0;
  reg  _EVAL_35;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_38;
  reg [31:0] _RAND_2;
  reg [6:0] _EVAL_69;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_148;
  reg [31:0] _RAND_4;
  reg [1:0] _EVAL_149;
  reg [31:0] _RAND_5;
  reg [72:0] _EVAL_158;
  reg [95:0] _RAND_6;
  reg [31:0] _EVAL_164;
  reg [31:0] _RAND_7;
  reg [5:0] _EVAL_172;
  reg [31:0] _RAND_8;
  reg [29:0] _EVAL_174;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_197;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_201;
  reg [31:0] _RAND_11;
  reg  _EVAL_246;
  reg [31:0] _RAND_12;
  reg [6:0] _EVAL_326;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_335;
  reg [31:0] _RAND_14;
  reg [5:0] _EVAL_337;
  reg [31:0] _RAND_15;
  reg [2:0] _EVAL_357;
  reg [31:0] _RAND_16;
  wire  _EVAL_176;
  wire  _EVAL_20;
  wire [1:0] _EVAL_318;
  wire [1:0] _EVAL_235;
  wire  _EVAL_76;
  wire  _EVAL_165;
  wire  _EVAL_282;
  wire  _EVAL_169;
  wire [3:0] _EVAL_256;
  wire  _EVAL_205;
  wire  _EVAL_238;
  wire  _EVAL_138;
  wire  _EVAL_228;
  wire  _EVAL_313;
  wire  _EVAL_258;
  wire  _EVAL_203;
  wire  _EVAL_253;
  wire  _EVAL_28;
  wire  _EVAL_321;
  wire  _EVAL_81;
  wire  _EVAL_54;
  wire  _EVAL_301;
  wire  _EVAL_210;
  wire [2:0] _EVAL_116;
  wire  _EVAL_332;
  wire  _EVAL_274;
  wire  _EVAL_272;
  wire  _EVAL_29;
  wire  _EVAL_93;
  wire  _EVAL_218;
  wire  _EVAL_37;
  wire  _EVAL_56;
  wire  _EVAL_106;
  wire  _EVAL_19;
  wire  _EVAL_168;
  wire  _EVAL_156;
  wire  _EVAL_97;
  wire  _EVAL_227;
  wire  _EVAL_196;
  wire  _EVAL_245;
  wire [22:0] _EVAL_311;
  wire [7:0] _EVAL_239;
  wire [7:0] _EVAL_101;
  wire [29:0] _EVAL_314;
  wire [29:0] _EVAL_45;
  wire  _EVAL_181;
  wire [29:0] _EVAL_202;
  wire [30:0] _EVAL_254;
  wire [30:0] _EVAL_191;
  wire [30:0] _EVAL_113;
  wire  _EVAL_163;
  wire  _EVAL_159;
  wire  _EVAL_251;
  wire  _EVAL_154;
  wire  _EVAL_167;
  wire  _EVAL_281;
  wire [31:0] _EVAL_108;
  wire  _EVAL_298;
  wire [29:0] _EVAL_206;
  wire [30:0] _EVAL_186;
  wire [30:0] _EVAL_85;
  wire [30:0] _EVAL_255;
  wire  _EVAL_360;
  wire [29:0] _EVAL_121;
  wire [30:0] _EVAL_98;
  wire [30:0] _EVAL_128;
  wire [30:0] _EVAL_307;
  wire  _EVAL_316;
  wire  _EVAL_127;
  wire [30:0] _EVAL_139;
  wire [30:0] _EVAL_351;
  wire [30:0] _EVAL_184;
  wire  _EVAL_190;
  wire  _EVAL_25;
  wire  _EVAL_283;
  wire  _EVAL_248;
  wire  _EVAL_278;
  wire  _EVAL_319;
  wire [29:0] _EVAL_322;
  wire [30:0] _EVAL_122;
  wire [30:0] _EVAL_315;
  wire [30:0] _EVAL_308;
  wire  _EVAL_257;
  wire  _EVAL_60;
  wire  _EVAL_275;
  wire  _EVAL_219;
  wire  _EVAL_243;
  wire  _EVAL_207;
  wire  _EVAL_217;
  wire [3:0] _EVAL_162;
  wire  _EVAL_183;
  wire  _EVAL_328;
  wire  _EVAL_72;
  wire  _EVAL_161;
  wire  _EVAL_123;
  wire  _EVAL_55;
  wire  _EVAL_157;
  wire  _EVAL_234;
  wire  _EVAL_216;
  wire  _EVAL_102;
  wire  _EVAL_114;
  wire  _EVAL_136;
  wire  _EVAL_22;
  wire  _EVAL_303;
  wire  _EVAL_64;
  wire  _EVAL_306;
  wire [3:0] _EVAL_170;
  wire [3:0] _EVAL_104;
  wire [3:0] _EVAL_291;
  wire  _EVAL_185;
  wire  _EVAL_226;
  wire [127:0] _EVAL_331;
  wire  _EVAL_324;
  wire  _EVAL_359;
  wire [2:0] _EVAL_92;
  wire  _EVAL_240;
  wire  _EVAL_195;
  wire  _EVAL_21;
  wire  _EVAL_261;
  wire  _EVAL_180;
  wire  _EVAL_208;
  wire  _EVAL_290;
  wire  _EVAL_75;
  wire  _EVAL_317;
  wire [22:0] _EVAL_120;
  wire [7:0] _EVAL_73;
  wire [7:0] _EVAL_339;
  wire [5:0] _EVAL_117;
  wire  _EVAL_353;
  wire  _EVAL_100;
  wire  _EVAL_347;
  wire  _EVAL_27;
  wire  _EVAL_88;
  wire  _EVAL_270;
  wire [29:0] _EVAL_115;
  wire [30:0] _EVAL_31;
  wire [30:0] _EVAL_58;
  wire [30:0] _EVAL_96;
  wire  _EVAL_178;
  wire  _EVAL_271;
  wire  _EVAL_134;
  wire  _EVAL_182;
  wire  _EVAL_329;
  wire [29:0] _EVAL_310;
  wire  _EVAL_279;
  wire  _EVAL_342;
  wire  _EVAL_287;
  wire  _EVAL_350;
  wire  _EVAL_199;
  wire  _EVAL_241;
  wire  _EVAL_212;
  wire  _EVAL_23;
  wire  _EVAL_62;
  wire  _EVAL_348;
  wire  _EVAL_295;
  wire  _EVAL_188;
  wire  _EVAL_53;
  wire  _EVAL_263;
  wire  _EVAL_52;
  wire  _EVAL_70;
  wire  _EVAL_343;
  wire  _EVAL_222;
  wire  _EVAL_211;
  wire  _EVAL_44;
  wire  _EVAL_221;
  wire  _EVAL_302;
  wire [3:0] _EVAL_66;
  wire  _EVAL_68;
  wire  _EVAL_346;
  wire  _EVAL_152;
  wire [127:0] _EVAL_204;
  wire [127:0] _EVAL_173;
  wire [72:0] _EVAL_325;
  wire [72:0] _EVAL_233;
  wire  _EVAL_268;
  wire  _EVAL_83;
  wire  _EVAL_340;
  wire  _EVAL_140;
  wire  _EVAL_250;
  wire  _EVAL_50;
  wire  _EVAL_47;
  wire  _EVAL_71;
  wire  _EVAL_124;
  wire  _EVAL_200;
  wire  _EVAL_79;
  wire  _EVAL_198;
  wire  _EVAL_215;
  wire  _EVAL_82;
  wire  _EVAL_225;
  wire  _EVAL_220;
  wire  _EVAL_141;
  wire [5:0] _EVAL_265;
  wire [30:0] _EVAL_237;
  wire [30:0] _EVAL_135;
  wire [30:0] _EVAL_177;
  wire  _EVAL_252;
  wire  _EVAL_166;
  wire  _EVAL_286;
  wire  _EVAL_297;
  wire  _EVAL_57;
  wire  _EVAL_249;
  wire  _EVAL_118;
  wire  _EVAL_46;
  wire  _EVAL_330;
  wire  _EVAL_260;
  wire  _EVAL_189;
  wire  _EVAL_131;
  wire  _EVAL_300;
  wire [72:0] _EVAL_160;
  wire [72:0] _EVAL_144;
  wire  _EVAL_264;
  wire  _EVAL_267;
  wire  _EVAL_99;
  wire [5:0] _EVAL_276;
  wire [5:0] _EVAL_107;
  wire  _EVAL_320;
  wire  _EVAL_129;
  wire  _EVAL_349;
  wire  _EVAL_284;
  wire  _EVAL_78;
  wire  _EVAL_288;
  wire  _EVAL_231;
  wire  _EVAL_175;
  wire  _EVAL_51;
  wire  _EVAL_91;
  wire  _EVAL_259;
  wire  _EVAL_277;
  wire  _EVAL_262;
  wire  _EVAL_358;
  wire  _EVAL_150;
  wire  _EVAL_305;
  wire  _EVAL_67;
  wire  _EVAL_30;
  wire  _EVAL_294;
  wire  _EVAL_125;
  wire  _EVAL_77;
  wire  _EVAL_119;
  wire  _EVAL_42;
  wire [5:0] _EVAL_48;
  wire  _EVAL_142;
  wire  _EVAL_155;
  wire  _EVAL_145;
  wire  _EVAL_336;
  wire [5:0] _EVAL_90;
  wire  _EVAL_354;
  wire  _EVAL_110;
  wire  _EVAL_179;
  wire  _EVAL_130;
  wire  _EVAL_244;
  wire  _EVAL_61;
  wire  _EVAL_280;
  wire  _EVAL_289;
  wire  _EVAL_153;
  wire  _EVAL_236;
  wire  _EVAL_24;
  wire  _EVAL_312;
  wire  _EVAL_356;
  wire  _EVAL_39;
  wire  _EVAL_112;
  wire  _EVAL_41;
  wire  _EVAL_266;
  wire  _EVAL_194;
  wire  _EVAL_103;
  wire  _EVAL_269;
  wire  _EVAL_49;
  wire  _EVAL_74;
  wire  _EVAL_192;
  wire  _EVAL_355;
  wire  _EVAL_333;
  wire  _EVAL_111;
  wire  _EVAL_323;
  wire  _EVAL_171;
  wire  _EVAL_59;
  wire  _EVAL_345;
  wire  _EVAL_26;
  wire [72:0] _EVAL_33;
  wire [127:0] _EVAL_296;
  wire [72:0] _EVAL_40;
  wire [72:0] _EVAL_137;
  wire [72:0] _EVAL_80;
  wire  _EVAL_341;
  wire  _EVAL_84;
  wire  _EVAL_232;
  wire  _EVAL_334;
  wire  _EVAL_126;
  wire  _EVAL_352;
  wire  _EVAL_193;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_304;
  wire  _EVAL_36;
  wire  _EVAL_87;
  wire  _EVAL_230;
  wire  _EVAL_327;
  wire  _EVAL_209;
  wire  _EVAL_187;
  wire  _EVAL_338;
  wire  _EVAL_247;
  wire  _EVAL_95;
  wire  _EVAL_273;
  wire  _EVAL_223;
  wire  _EVAL_65;
  wire  _EVAL_229;
  wire  _EVAL_344;
  wire  _EVAL_89;
  wire  _EVAL_213;
  wire  _EVAL_133;
  wire  _EVAL_242;
  wire  _EVAL_109;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_176 = _EVAL_4 >= 4'h2;
  assign _EVAL_20 = _EVAL_4[0];
  assign _EVAL_318 = 2'h1 << _EVAL_20;
  assign _EVAL_235 = _EVAL_318 | 2'h1;
  assign _EVAL_76 = _EVAL_235[1];
  assign _EVAL_165 = _EVAL_17[1];
  assign _EVAL_282 = _EVAL_76 & _EVAL_165;
  assign _EVAL_169 = _EVAL_176 | _EVAL_282;
  assign _EVAL_256 = _EVAL_8[6:3];
  assign _EVAL_205 = _EVAL_256 == 4'h3;
  assign _EVAL_238 = _EVAL_15 == _EVAL_35;
  assign _EVAL_138 = _EVAL_238 | _EVAL_18;
  assign _EVAL_228 = _EVAL_10 == _EVAL_69;
  assign _EVAL_313 = _EVAL_228 | _EVAL_18;
  assign _EVAL_258 = _EVAL_1[0];
  assign _EVAL_203 = _EVAL_235[0];
  assign _EVAL_253 = _EVAL_17[0];
  assign _EVAL_28 = _EVAL_165 & _EVAL_253;
  assign _EVAL_321 = _EVAL_203 & _EVAL_28;
  assign _EVAL_81 = _EVAL_8 == 7'h48;
  assign _EVAL_54 = _EVAL_8 == 7'h40;
  assign _EVAL_301 = _EVAL_81 | _EVAL_54;
  assign _EVAL_210 = _EVAL_256 == 4'h8;
  assign _EVAL_116 = _EVAL_8[2:0];
  assign _EVAL_332 = 3'h1 <= _EVAL_116;
  assign _EVAL_274 = _EVAL_210 & _EVAL_332;
  assign _EVAL_272 = _EVAL_301 | _EVAL_274;
  assign _EVAL_29 = _EVAL_8 == 7'h20;
  assign _EVAL_93 = _EVAL_272 | _EVAL_29;
  assign _EVAL_218 = _EVAL_256 == 4'h0;
  assign _EVAL_37 = _EVAL_93 | _EVAL_218;
  assign _EVAL_56 = _EVAL_256 == 4'h1;
  assign _EVAL_106 = _EVAL_37 | _EVAL_56;
  assign _EVAL_19 = _EVAL_256 == 4'h2;
  assign _EVAL_168 = _EVAL_106 | _EVAL_19;
  assign _EVAL_156 = _EVAL_168 | _EVAL_205;
  assign _EVAL_97 = _EVAL_337 == 6'h0;
  assign _EVAL_227 = _EVAL_4 == _EVAL_148;
  assign _EVAL_196 = _EVAL_227 | _EVAL_18;
  assign _EVAL_245 = _EVAL_158 != 73'h0;
  assign _EVAL_311 = 23'hff << _EVAL_4;
  assign _EVAL_239 = _EVAL_311[7:0];
  assign _EVAL_101 = ~ _EVAL_239;
  assign _EVAL_314 = {{22'd0}, _EVAL_101};
  assign _EVAL_45 = _EVAL_17 & _EVAL_314;
  assign _EVAL_181 = _EVAL_45 == 30'h0;
  assign _EVAL_202 = _EVAL_17 ^ 30'h20000000;
  assign _EVAL_254 = {1'b0,$signed(_EVAL_202)};
  assign _EVAL_191 = $signed(_EVAL_254) & $signed(-31'sh2000);
  assign _EVAL_113 = $signed(_EVAL_191);
  assign _EVAL_163 = _EVAL == 3'h0;
  assign _EVAL_159 = _EVAL_163 | _EVAL_18;
  assign _EVAL_251 = _EVAL_159 == 1'h0;
  assign _EVAL_154 = _EVAL_2 & _EVAL_16;
  assign _EVAL_167 = _EVAL_5 & _EVAL_14;
  assign _EVAL_281 = _EVAL_154 | _EVAL_167;
  assign _EVAL_108 = _EVAL_164 + 32'h1;
  assign _EVAL_298 = _EVAL <= 3'h3;
  assign _EVAL_206 = _EVAL_17 ^ 30'hc000000;
  assign _EVAL_186 = {1'b0,$signed(_EVAL_206)};
  assign _EVAL_85 = $signed(_EVAL_186) & $signed(-31'sh4000000);
  assign _EVAL_255 = $signed(_EVAL_85);
  assign _EVAL_360 = $signed(_EVAL_255) == $signed(31'sh0);
  assign _EVAL_121 = _EVAL_17 ^ 30'h2000000;
  assign _EVAL_98 = {1'b0,$signed(_EVAL_121)};
  assign _EVAL_128 = $signed(_EVAL_98) & $signed(-31'sh10000);
  assign _EVAL_307 = $signed(_EVAL_128);
  assign _EVAL_316 = $signed(_EVAL_307) == $signed(31'sh0);
  assign _EVAL_127 = _EVAL_360 | _EVAL_316;
  assign _EVAL_139 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_351 = $signed(_EVAL_139) & $signed(-31'sh5000);
  assign _EVAL_184 = $signed(_EVAL_351);
  assign _EVAL_190 = $signed(_EVAL_184) == $signed(31'sh0);
  assign _EVAL_25 = _EVAL_127 | _EVAL_190;
  assign _EVAL_283 = _EVAL_169 | _EVAL_321;
  assign _EVAL_248 = _EVAL_1 == 3'h4;
  assign _EVAL_278 = _EVAL_14 & _EVAL_248;
  assign _EVAL_319 = _EVAL_4 <= 4'h8;
  assign _EVAL_322 = _EVAL_17 ^ 30'h3000;
  assign _EVAL_122 = {1'b0,$signed(_EVAL_322)};
  assign _EVAL_315 = $signed(_EVAL_122) & $signed(-31'sh1000);
  assign _EVAL_308 = $signed(_EVAL_315);
  assign _EVAL_257 = $signed(_EVAL_308) == $signed(31'sh0);
  assign _EVAL_60 = _EVAL_319 & _EVAL_257;
  assign _EVAL_275 = _EVAL_7 != 2'h2;
  assign _EVAL_219 = _EVAL_172 == 6'h0;
  assign _EVAL_243 = _EVAL_219 == 1'h0;
  assign _EVAL_207 = _EVAL_1 == 3'h2;
  assign _EVAL_217 = _EVAL_14 & _EVAL_207;
  assign _EVAL_162 = _EVAL_10[6:3];
  assign _EVAL_183 = _EVAL_162 == 4'h8;
  assign _EVAL_328 = 4'h6 == _EVAL_4;
  assign _EVAL_72 = _EVAL_3 == 3'h6;
  assign _EVAL_161 = _EVAL_253 == 1'h0;
  assign _EVAL_123 = _EVAL_165 & _EVAL_161;
  assign _EVAL_55 = _EVAL_203 & _EVAL_123;
  assign _EVAL_157 = _EVAL_169 | _EVAL_55;
  assign _EVAL_234 = _EVAL_165 == 1'h0;
  assign _EVAL_216 = _EVAL_76 & _EVAL_234;
  assign _EVAL_102 = _EVAL_176 | _EVAL_216;
  assign _EVAL_114 = _EVAL_234 & _EVAL_253;
  assign _EVAL_136 = _EVAL_203 & _EVAL_114;
  assign _EVAL_22 = _EVAL_102 | _EVAL_136;
  assign _EVAL_303 = _EVAL_234 & _EVAL_161;
  assign _EVAL_64 = _EVAL_203 & _EVAL_303;
  assign _EVAL_306 = _EVAL_102 | _EVAL_64;
  assign _EVAL_170 = {_EVAL_283,_EVAL_157,_EVAL_22,_EVAL_306};
  assign _EVAL_104 = ~ _EVAL_170;
  assign _EVAL_291 = _EVAL_12 & _EVAL_104;
  assign _EVAL_185 = _EVAL_291 == 4'h0;
  assign _EVAL_226 = _EVAL_185 | _EVAL_18;
  assign _EVAL_331 = 128'h1 << _EVAL_10;
  assign _EVAL_324 = _EVAL <= 3'h2;
  assign _EVAL_359 = _EVAL_324 | _EVAL_18;
  assign _EVAL_92 = _EVAL_10[2:0];
  assign _EVAL_240 = 3'h1 <= _EVAL_92;
  assign _EVAL_195 = _EVAL_183 & _EVAL_240;
  assign _EVAL_21 = _EVAL_3[2];
  assign _EVAL_261 = _EVAL_245 == 1'h0;
  assign _EVAL_180 = _EVAL == _EVAL_201;
  assign _EVAL_208 = _EVAL_180 | _EVAL_18;
  assign _EVAL_290 = _EVAL_13 == _EVAL_246;
  assign _EVAL_75 = _EVAL_290 | _EVAL_18;
  assign _EVAL_317 = _EVAL_38 == 6'h0;
  assign _EVAL_120 = 23'hff << _EVAL_9;
  assign _EVAL_73 = _EVAL_120[7:0];
  assign _EVAL_339 = ~ _EVAL_73;
  assign _EVAL_117 = _EVAL_339[7:2];
  assign _EVAL_353 = _EVAL_11 == 1'h0;
  assign _EVAL_100 = _EVAL_1 == 3'h0;
  assign _EVAL_347 = _EVAL_14 & _EVAL_100;
  assign _EVAL_27 = _EVAL_1 <= 3'h6;
  assign _EVAL_88 = _EVAL_27 | _EVAL_18;
  assign _EVAL_270 = _EVAL_88 == 1'h0;
  assign _EVAL_115 = _EVAL_17 ^ 30'h1900000;
  assign _EVAL_31 = {1'b0,$signed(_EVAL_115)};
  assign _EVAL_58 = $signed(_EVAL_31) & $signed(-31'sh2000);
  assign _EVAL_96 = $signed(_EVAL_58);
  assign _EVAL_178 = _EVAL_298 | _EVAL_18;
  assign _EVAL_271 = _EVAL_176 | _EVAL_18;
  assign _EVAL_134 = _EVAL_7 == _EVAL_149;
  assign _EVAL_182 = _EVAL_134 | _EVAL_18;
  assign _EVAL_329 = _EVAL_182 == 1'h0;
  assign _EVAL_310 = _EVAL_17 ^ 30'h1800000;
  assign _EVAL_279 = _EVAL_9 >= 4'h2;
  assign _EVAL_342 = _EVAL_279 | _EVAL_18;
  assign _EVAL_287 = _EVAL_342 == 1'h0;
  assign _EVAL_350 = _EVAL_164 < plusarg_reader_out;
  assign _EVAL_199 = _EVAL_12 == _EVAL_170;
  assign _EVAL_241 = _EVAL_199 | _EVAL_18;
  assign _EVAL_212 = _EVAL_162 == 4'h1;
  assign _EVAL_23 = _EVAL_10 == 7'h48;
  assign _EVAL_62 = _EVAL_10 == 7'h40;
  assign _EVAL_348 = _EVAL_23 | _EVAL_62;
  assign _EVAL_295 = _EVAL_348 | _EVAL_195;
  assign _EVAL_188 = _EVAL_10 == 7'h20;
  assign _EVAL_53 = _EVAL_295 | _EVAL_188;
  assign _EVAL_263 = _EVAL_162 == 4'h0;
  assign _EVAL_52 = _EVAL_53 | _EVAL_263;
  assign _EVAL_70 = _EVAL_52 | _EVAL_212;
  assign _EVAL_343 = _EVAL_162 == 4'h2;
  assign _EVAL_222 = _EVAL_70 | _EVAL_343;
  assign _EVAL_211 = _EVAL_162 == 4'h3;
  assign _EVAL_44 = _EVAL_222 | _EVAL_211;
  assign _EVAL_221 = _EVAL_44 | _EVAL_18;
  assign _EVAL_302 = _EVAL_221 == 1'h0;
  assign _EVAL_66 = ~ _EVAL_12;
  assign _EVAL_68 = _EVAL_317 == 1'h0;
  assign _EVAL_346 = _EVAL_197 == 6'h0;
  assign _EVAL_152 = _EVAL_154 & _EVAL_346;
  assign _EVAL_204 = 128'h1 << _EVAL_8;
  assign _EVAL_173 = _EVAL_152 ? _EVAL_204 : 128'h0;
  assign _EVAL_325 = _EVAL_173[72:0];
  assign _EVAL_233 = _EVAL_158 >> _EVAL_8;
  assign _EVAL_268 = _EVAL_233[0];
  assign _EVAL_83 = _EVAL_268 == 1'h0;
  assign _EVAL_340 = _EVAL_83 | _EVAL_18;
  assign _EVAL_140 = _EVAL_1 == _EVAL_32;
  assign _EVAL_250 = _EVAL_140 | _EVAL_18;
  assign _EVAL_50 = _EVAL_250 == 1'h0;
  assign _EVAL_47 = _EVAL_14 & _EVAL_243;
  assign _EVAL_71 = plusarg_reader_out == 32'h0;
  assign _EVAL_124 = _EVAL_261 | _EVAL_71;
  assign _EVAL_200 = _EVAL_124 | _EVAL_350;
  assign _EVAL_79 = _EVAL_156 | _EVAL_18;
  assign _EVAL_198 = _EVAL != 3'h0;
  assign _EVAL_215 = _EVAL_1 == 3'h6;
  assign _EVAL_82 = _EVAL_14 & _EVAL_215;
  assign _EVAL_225 = _EVAL <= 3'h4;
  assign _EVAL_220 = _EVAL_3 == 3'h0;
  assign _EVAL_141 = _EVAL_16 & _EVAL_220;
  assign _EVAL_265 = _EVAL_38 - 6'h1;
  assign _EVAL_237 = {1'b0,$signed(_EVAL_310)};
  assign _EVAL_135 = $signed(_EVAL_237) & $signed(-31'sh8000);
  assign _EVAL_177 = $signed(_EVAL_135);
  assign _EVAL_252 = $signed(_EVAL_177) == $signed(31'sh0);
  assign _EVAL_166 = _EVAL_4 <= 4'h6;
  assign _EVAL_286 = _EVAL_25 | _EVAL_252;
  assign _EVAL_297 = $signed(_EVAL_96) == $signed(31'sh0);
  assign _EVAL_57 = _EVAL_286 | _EVAL_297;
  assign _EVAL_249 = $signed(_EVAL_113) == $signed(31'sh0);
  assign _EVAL_118 = _EVAL_57 | _EVAL_249;
  assign _EVAL_46 = _EVAL_166 & _EVAL_118;
  assign _EVAL_330 = _EVAL_17 == _EVAL_174;
  assign _EVAL_260 = _EVAL_330 | _EVAL_18;
  assign _EVAL_189 = _EVAL_66 == 4'h0;
  assign _EVAL_131 = _EVAL_189 | _EVAL_18;
  assign _EVAL_300 = _EVAL_131 == 1'h0;
  assign _EVAL_160 = _EVAL_325 | _EVAL_158;
  assign _EVAL_144 = _EVAL_160 >> _EVAL_10;
  assign _EVAL_264 = _EVAL_54 ? _EVAL_328 : 1'h0;
  assign _EVAL_267 = _EVAL_264 | _EVAL_18;
  assign _EVAL_99 = _EVAL_21 == 1'h0;
  assign _EVAL_276 = _EVAL_101[7:2];
  assign _EVAL_107 = _EVAL_197 - 6'h1;
  assign _EVAL_320 = _EVAL_3 == 3'h3;
  assign _EVAL_129 = _EVAL_16 & _EVAL_320;
  assign _EVAL_349 = _EVAL_1 == 3'h1;
  assign _EVAL_284 = _EVAL_14 & _EVAL_349;
  assign _EVAL_78 = _EVAL_4 <= 4'h2;
  assign _EVAL_288 = _EVAL_257 | _EVAL_297;
  assign _EVAL_231 = _EVAL_78 & _EVAL_288;
  assign _EVAL_175 = _EVAL_231 | _EVAL_18;
  assign _EVAL_51 = _EVAL_175 == 1'h0;
  assign _EVAL_91 = _EVAL_3 == 3'h2;
  assign _EVAL_259 = _EVAL_16 & _EVAL_91;
  assign _EVAL_277 = _EVAL_13 == 1'h0;
  assign _EVAL_262 = _EVAL_277 | _EVAL_0;
  assign _EVAL_358 = _EVAL_262 | _EVAL_18;
  assign _EVAL_150 = _EVAL_358 == 1'h0;
  assign _EVAL_305 = _EVAL_3 == 3'h7;
  assign _EVAL_67 = _EVAL_60 | _EVAL_46;
  assign _EVAL_30 = _EVAL_181 | _EVAL_18;
  assign _EVAL_294 = _EVAL_7 == 2'h0;
  assign _EVAL_125 = _EVAL_294 | _EVAL_18;
  assign _EVAL_77 = _EVAL_60 | _EVAL_18;
  assign _EVAL_119 = _EVAL_353 | _EVAL_18;
  assign _EVAL_42 = _EVAL_119 == 1'h0;
  assign _EVAL_48 = _EVAL_337 - 6'h1;
  assign _EVAL_142 = _EVAL_79 == 1'h0;
  assign _EVAL_155 = _EVAL_196 == 1'h0;
  assign _EVAL_145 = _EVAL_0 == 1'h0;
  assign _EVAL_336 = _EVAL_145 | _EVAL_18;
  assign _EVAL_90 = _EVAL_172 - 6'h1;
  assign _EVAL_354 = _EVAL_225 | _EVAL_18;
  assign _EVAL_110 = _EVAL_354 == 1'h0;
  assign _EVAL_179 = _EVAL_144[0];
  assign _EVAL_130 = _EVAL_179 | _EVAL_18;
  assign _EVAL_244 = _EVAL_3 == _EVAL_357;
  assign _EVAL_61 = _EVAL_244 | _EVAL_18;
  assign _EVAL_280 = _EVAL_61 == 1'h0;
  assign _EVAL_289 = _EVAL_313 == 1'h0;
  assign _EVAL_153 = _EVAL_208 == 1'h0;
  assign _EVAL_236 = _EVAL_336 == 1'h0;
  assign _EVAL_24 = _EVAL_9 == _EVAL_335;
  assign _EVAL_312 = _EVAL_24 | _EVAL_18;
  assign _EVAL_356 = _EVAL_7 <= 2'h2;
  assign _EVAL_39 = _EVAL_356 | _EVAL_18;
  assign _EVAL_112 = _EVAL_67 | _EVAL_18;
  assign _EVAL_41 = _EVAL_112 == 1'h0;
  assign _EVAL_266 = _EVAL_16 & _EVAL_68;
  assign _EVAL_194 = _EVAL_167 & _EVAL_97;
  assign _EVAL_103 = _EVAL_215 == 1'h0;
  assign _EVAL_269 = _EVAL_194 & _EVAL_103;
  assign _EVAL_49 = _EVAL_8 == _EVAL_326;
  assign _EVAL_74 = _EVAL_49 | _EVAL_18;
  assign _EVAL_192 = _EVAL_74 == 1'h0;
  assign _EVAL_355 = _EVAL_18 == 1'h0;
  assign _EVAL_333 = _EVAL_3 == 3'h5;
  assign _EVAL_111 = _EVAL_30 == 1'h0;
  assign _EVAL_323 = _EVAL_178 == 1'h0;
  assign _EVAL_171 = _EVAL_200 | _EVAL_18;
  assign _EVAL_59 = _EVAL_171 == 1'h0;
  assign _EVAL_345 = _EVAL_271 == 1'h0;
  assign _EVAL_26 = _EVAL_3 == 3'h1;
  assign _EVAL_33 = _EVAL_158 | _EVAL_325;
  assign _EVAL_296 = _EVAL_269 ? _EVAL_331 : 128'h0;
  assign _EVAL_40 = _EVAL_296[72:0];
  assign _EVAL_137 = ~ _EVAL_40;
  assign _EVAL_80 = _EVAL_33 & _EVAL_137;
  assign _EVAL_341 = _EVAL_198 | _EVAL_18;
  assign _EVAL_84 = _EVAL_3 == 3'h4;
  assign _EVAL_232 = _EVAL_16 & _EVAL_84;
  assign _EVAL_334 = _EVAL_359 == 1'h0;
  assign _EVAL_126 = _EVAL_275 | _EVAL_18;
  assign _EVAL_352 = _EVAL_126 == 1'h0;
  assign _EVAL_193 = _EVAL_277 | _EVAL_18;
  assign _EVAL_292 = _EVAL_193 == 1'h0;
  assign _EVAL_293 = _EVAL_39 == 1'h0;
  assign _EVAL_304 = _EVAL_130 == 1'h0;
  assign _EVAL_36 = _EVAL_167 & _EVAL_219;
  assign _EVAL_87 = _EVAL_341 == 1'h0;
  assign _EVAL_230 = _EVAL_260 == 1'h0;
  assign _EVAL_327 = _EVAL_154 & _EVAL_317;
  assign _EVAL_209 = _EVAL_1 == 3'h5;
  assign _EVAL_187 = _EVAL_14 & _EVAL_209;
  assign _EVAL_338 = _EVAL_16 & _EVAL_26;
  assign _EVAL_247 = _EVAL_138 == 1'h0;
  assign _EVAL_95 = _EVAL_125 == 1'h0;
  assign _EVAL_273 = _EVAL_75 == 1'h0;
  assign _EVAL_223 = _EVAL_16 & _EVAL_333;
  assign _EVAL_65 = _EVAL_241 == 1'h0;
  assign _EVAL_229 = _EVAL_226 == 1'h0;
  assign _EVAL_344 = _EVAL_267 == 1'h0;
  assign _EVAL_89 = _EVAL_312 == 1'h0;
  assign _EVAL_213 = _EVAL_16 & _EVAL_72;
  assign _EVAL_133 = _EVAL_16 & _EVAL_305;
  assign _EVAL_242 = _EVAL_340 == 1'h0;
  assign _EVAL_109 = _EVAL_77 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_38 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_69 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_148 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_149 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  _EVAL_158 = _RAND_6[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_164 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_172 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_174 = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_197 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_201 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_246 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_326 = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_335 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_337 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_357 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_6) begin
    if (_EVAL_36) begin
      _EVAL_32 <= _EVAL_1;
    end
    if (_EVAL_36) begin
      _EVAL_35 <= _EVAL_15;
    end
    if (_EVAL_18) begin
      _EVAL_38 <= 6'h0;
    end else begin
      if (_EVAL_154) begin
        if (_EVAL_317) begin
          if (_EVAL_99) begin
            _EVAL_38 <= _EVAL_276;
          end else begin
            _EVAL_38 <= 6'h0;
          end
        end else begin
          _EVAL_38 <= _EVAL_265;
        end
      end
    end
    if (_EVAL_36) begin
      _EVAL_69 <= _EVAL_10;
    end
    if (_EVAL_327) begin
      _EVAL_148 <= _EVAL_4;
    end
    if (_EVAL_36) begin
      _EVAL_149 <= _EVAL_7;
    end
    if (_EVAL_18) begin
      _EVAL_158 <= 73'h0;
    end else begin
      _EVAL_158 <= _EVAL_80;
    end
    if (_EVAL_18) begin
      _EVAL_164 <= 32'h0;
    end else begin
      if (_EVAL_281) begin
        _EVAL_164 <= 32'h0;
      end else begin
        _EVAL_164 <= _EVAL_108;
      end
    end
    if (_EVAL_18) begin
      _EVAL_172 <= 6'h0;
    end else begin
      if (_EVAL_167) begin
        if (_EVAL_219) begin
          if (_EVAL_258) begin
            _EVAL_172 <= _EVAL_117;
          end else begin
            _EVAL_172 <= 6'h0;
          end
        end else begin
          _EVAL_172 <= _EVAL_90;
        end
      end
    end
    if (_EVAL_327) begin
      _EVAL_174 <= _EVAL_17;
    end
    if (_EVAL_18) begin
      _EVAL_197 <= 6'h0;
    end else begin
      if (_EVAL_154) begin
        if (_EVAL_346) begin
          if (_EVAL_99) begin
            _EVAL_197 <= _EVAL_276;
          end else begin
            _EVAL_197 <= 6'h0;
          end
        end else begin
          _EVAL_197 <= _EVAL_107;
        end
      end
    end
    if (_EVAL_327) begin
      _EVAL_201 <= _EVAL;
    end
    if (_EVAL_36) begin
      _EVAL_246 <= _EVAL_13;
    end
    if (_EVAL_327) begin
      _EVAL_326 <= _EVAL_8;
    end
    if (_EVAL_36) begin
      _EVAL_335 <= _EVAL_9;
    end
    if (_EVAL_18) begin
      _EVAL_337 <= 6'h0;
    end else begin
      if (_EVAL_167) begin
        if (_EVAL_97) begin
          if (_EVAL_258) begin
            _EVAL_337 <= _EVAL_117;
          end else begin
            _EVAL_337 <= 6'h0;
          end
        end else begin
          _EVAL_337 <= _EVAL_48;
        end
      end
    end
    if (_EVAL_327) begin
      _EVAL_357 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdd1af14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93f707d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_329) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5d71ca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26057de7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_345) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918ab113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(264ebb95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3547c264)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8c7c945)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5db932d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16cdc5ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaf5132a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ec209e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_345) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2f4c8eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5669a024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d6fe87f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60fc623a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa8e2c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfa264e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28fb83dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52c0a55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(134f45d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ed667d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ddabab7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6443e310)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9133b0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e551eed5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9702c23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40651ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64f40050)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b621621b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35db4494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f34f466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_334) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1d82c86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_334) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(731c1272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a47d305a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b60b5e7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1baf3536)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e745cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36483e86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa57943b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0948909)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd1d38f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afa525c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_345) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8076d126)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4546bdd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90c0b78c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31bc7e69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(142d9a81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7d4e3ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aefd357b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0181d01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7681a693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64682cb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83940964)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_329) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bf1b9a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf38775c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61950a62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33bfc3aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f4c0576)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ca8532f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27e21020)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a62d785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36959606)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2404683)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ded681)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da685b59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30cc4502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(749eb2dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a9b1384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5073abd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7dff92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d471e5e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af636a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3339824)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37ef0c0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fa7fc71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_345) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acf45559)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(160c0124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76937a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2be2f83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa4db3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1716424)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb1521be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4911462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9f3b811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70f5acbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c2c1429)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d42f9774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d84a833)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
