//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_210(
  input          _EVAL,
  output         _EVAL_0,
  input  [7:0]   _EVAL_1,
  output         _EVAL_2,
  output         _EVAL_3,
  input          _EVAL_4,
  input  [2:0]   _EVAL_5,
  output         _EVAL_6,
  output         _EVAL_7,
  output         _EVAL_8,
  output         _EVAL_9,
  output [31:0]  _EVAL_10,
  input          _EVAL_11,
  output         _EVAL_12,
  output [3:0]   _EVAL_13,
  output [2:0]   _EVAL_14,
  output         _EVAL_15,
  input          _EVAL_16,
  input          _EVAL_17,
  input          _EVAL_18,
  output [7:0]   _EVAL_19,
  input          _EVAL_20,
  input  [127:0] _EVAL_21,
  output         _EVAL_22,
  output [2:0]   _EVAL_23,
  input          _EVAL_24,
  input          _EVAL_25,
  output         _EVAL_26,
  output [7:0]   _EVAL_27,
  input  [127:0] _EVAL_28
);
  wire  d__EVAL;
  wire  d__EVAL_0;
  wire  d__EVAL_1;
  wire  d__EVAL_2;
  wire [7:0] d__EVAL_3;
  wire  d__EVAL_4;
  wire [7:0] d__EVAL_5;
  wire  d__EVAL_6;
  wire  d__EVAL_7;
  wire  d__EVAL_8;
  wire  d__EVAL_9;
  wire  d__EVAL_10;
  reg [2:0] _EVAL_75;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_130;
  reg [31:0] _RAND_1;
  wire [127:0] _EVAL_139;
  wire [128:0] _EVAL_96;
  wire [128:0] _EVAL_99;
  wire [128:0] _EVAL_71;
  wire  _EVAL_78;
  wire [127:0] _EVAL_128;
  wire  _EVAL_44;
  wire [127:0] _EVAL_124;
  wire [128:0] _EVAL_95;
  wire [128:0] _EVAL_111;
  wire [128:0] _EVAL_115;
  wire [128:0] _EVAL_60;
  wire [128:0] _EVAL_109;
  wire [127:0] _EVAL_40;
  wire [128:0] _EVAL_43;
  wire [128:0] _EVAL_45;
  wire  _EVAL_83;
  wire  _EVAL_81;
  wire  _EVAL_69;
  wire  _EVAL_49;
  wire  _EVAL_36;
  wire  _EVAL_125;
  wire  _EVAL_77;
  wire  _EVAL_68;
  wire  _EVAL_110;
  wire  _EVAL_94;
  wire  _EVAL_119;
  wire  _EVAL_118;
  wire [7:0] _EVAL_31;
  wire [7:0] _EVAL_41;
  wire [7:0] _EVAL_142;
  wire  _EVAL_133;
  wire  _EVAL_141;
  wire [2:0] _EVAL_121;
  wire  _EVAL_135;
  wire  _EVAL_97;
  wire [127:0] _EVAL_140;
  wire [128:0] _EVAL_32;
  wire [128:0] _EVAL_87;
  wire [128:0] _EVAL_137;
  wire [128:0] _EVAL_74;
  wire [128:0] _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_84;
  wire  _EVAL_136;
  wire  _EVAL_117;
  wire  _EVAL_123;
  wire  _EVAL_132;
  wire [128:0] _EVAL_42;
  wire  _EVAL_64;
  wire [128:0] _EVAL_67;
  wire  _EVAL_101;
  wire  _EVAL_143;
  wire [127:0] _EVAL_76;
  wire [128:0] _EVAL_91;
  wire [128:0] _EVAL_107;
  wire [128:0] _EVAL_113;
  wire  _EVAL_52;
  wire  _EVAL_104;
  wire [128:0] _EVAL_126;
  wire  _EVAL_98;
  wire  _EVAL_108;
  wire [127:0] _EVAL_80;
  wire [128:0] _EVAL_112;
  wire [128:0] _EVAL_114;
  wire [128:0] _EVAL_88;
  wire  _EVAL_138;
  wire  _EVAL_86;
  wire  _EVAL_103;
  wire  _EVAL_122;
  wire  _EVAL_50;
  wire [1:0] _EVAL_51;
  wire [7:0] _EVAL_35;
  wire [7:0] _EVAL_58;
  wire [7:0] _EVAL_89;
  wire [7:0] _EVAL_39;
  wire [7:0] _EVAL_85;
  wire [7:0] _EVAL_145;
  wire [7:0] _EVAL_90;
  wire [127:0] _EVAL_73;
  wire [128:0] _EVAL_55;
  wire [128:0] _EVAL_62;
  wire [128:0] _EVAL_147;
  wire  _EVAL_120;
  wire  _EVAL_66;
  wire [31:0] _EVAL_47;
  wire  _EVAL_33;
  wire  _EVAL_30;
  wire [3:0] _EVAL_29;
  wire  _EVAL_92;
  SiFive__EVAL_209 d (
    ._EVAL(d__EVAL),
    ._EVAL_0(d__EVAL_0),
    ._EVAL_1(d__EVAL_1),
    ._EVAL_2(d__EVAL_2),
    ._EVAL_3(d__EVAL_3),
    ._EVAL_4(d__EVAL_4),
    ._EVAL_5(d__EVAL_5),
    ._EVAL_6(d__EVAL_6),
    ._EVAL_7(d__EVAL_7),
    ._EVAL_8(d__EVAL_8),
    ._EVAL_9(d__EVAL_9),
    ._EVAL_10(d__EVAL_10)
  );
  assign _EVAL_139 = _EVAL_28 ^ 128'h1900000;
  assign _EVAL_96 = {1'b0,$signed(_EVAL_139)};
  assign _EVAL_99 = $signed(_EVAL_96) & $signed(-129'sh2000);
  assign _EVAL_71 = $signed(_EVAL_99);
  assign _EVAL_78 = d__EVAL_1 & d__EVAL_9;
  assign _EVAL_128 = _EVAL_28 ^ 128'h40000000;
  assign _EVAL_44 = _EVAL_75 == 3'h0;
  assign _EVAL_124 = _EVAL_28 ^ 128'h80000000;
  assign _EVAL_95 = {1'b0,$signed(_EVAL_124)};
  assign _EVAL_111 = $signed(_EVAL_95) & $signed(-129'sh20000);
  assign _EVAL_115 = {1'b0,$signed(_EVAL_28)};
  assign _EVAL_60 = $signed(_EVAL_115) & $signed(-129'sh5000);
  assign _EVAL_109 = $signed(_EVAL_60);
  assign _EVAL_40 = _EVAL_28 ^ 128'hc000000;
  assign _EVAL_43 = {1'b0,$signed(_EVAL_40)};
  assign _EVAL_45 = $signed(_EVAL_43) & $signed(-129'sh4000000);
  assign _EVAL_83 = _EVAL_25 & _EVAL_7;
  assign _EVAL_81 = _EVAL_11 & _EVAL_6;
  assign _EVAL_69 = $signed(_EVAL_71) == $signed(129'sh0);
  assign _EVAL_49 = _EVAL_130 == 3'h2;
  assign _EVAL_36 = _EVAL_130 == 3'h1;
  assign _EVAL_125 = _EVAL_36 | _EVAL_49;
  assign _EVAL_77 = _EVAL_49 & _EVAL_125;
  assign _EVAL_68 = _EVAL_77 & _EVAL_4;
  assign _EVAL_110 = _EVAL_130 == 3'h3;
  assign _EVAL_94 = _EVAL_110 & d__EVAL_1;
  assign _EVAL_119 = _EVAL_94 & d__EVAL_9;
  assign _EVAL_118 = _EVAL_68 | _EVAL_119;
  assign _EVAL_31 = {{5'd0}, _EVAL_75};
  assign _EVAL_41 = 8'h1 << _EVAL_5;
  assign _EVAL_142 = _EVAL_41 - 8'h1;
  assign _EVAL_133 = _EVAL_31 == _EVAL_142;
  assign _EVAL_141 = _EVAL_118 & _EVAL_133;
  assign _EVAL_121 = _EVAL_75 + 3'h1;
  assign _EVAL_135 = _EVAL_119 & _EVAL_133;
  assign _EVAL_97 = _EVAL_130 == 3'h4;
  assign _EVAL_140 = _EVAL_28 ^ 128'h1800000;
  assign _EVAL_32 = {1'b0,$signed(_EVAL_140)};
  assign _EVAL_87 = $signed(_EVAL_32) & $signed(-129'sh8000);
  assign _EVAL_137 = $signed(_EVAL_87);
  assign _EVAL_74 = {1'b0,$signed(_EVAL_128)};
  assign _EVAL_70 = $signed(_EVAL_74) & $signed(-129'sh2000);
  assign _EVAL_72 = $signed(_EVAL_137) == $signed(129'sh0);
  assign _EVAL_84 = _EVAL_75 == 3'h2;
  assign _EVAL_136 = ~ _EVAL_17;
  assign _EVAL_117 = _EVAL_130 == 3'h0;
  assign _EVAL_123 = _EVAL_125 & _EVAL_4;
  assign _EVAL_132 = _EVAL_68 & _EVAL_133;
  assign _EVAL_42 = $signed(_EVAL_70);
  assign _EVAL_64 = $signed(_EVAL_42) == $signed(129'sh0);
  assign _EVAL_67 = $signed(_EVAL_111);
  assign _EVAL_101 = $signed(_EVAL_67) == $signed(129'sh0);
  assign _EVAL_143 = _EVAL_64 | _EVAL_101;
  assign _EVAL_76 = _EVAL_28 ^ 128'h3000;
  assign _EVAL_91 = {1'b0,$signed(_EVAL_76)};
  assign _EVAL_107 = $signed(_EVAL_91) & $signed(-129'sh1000);
  assign _EVAL_113 = $signed(_EVAL_107);
  assign _EVAL_52 = $signed(_EVAL_113) == $signed(129'sh0);
  assign _EVAL_104 = _EVAL_143 | _EVAL_52;
  assign _EVAL_126 = $signed(_EVAL_45);
  assign _EVAL_98 = $signed(_EVAL_126) == $signed(129'sh0);
  assign _EVAL_108 = _EVAL_104 | _EVAL_98;
  assign _EVAL_80 = _EVAL_28 ^ 128'h2000000;
  assign _EVAL_112 = {1'b0,$signed(_EVAL_80)};
  assign _EVAL_114 = $signed(_EVAL_112) & $signed(-129'sh10000);
  assign _EVAL_88 = $signed(_EVAL_114);
  assign _EVAL_138 = $signed(_EVAL_88) == $signed(129'sh0);
  assign _EVAL_86 = _EVAL_108 | _EVAL_138;
  assign _EVAL_103 = $signed(_EVAL_109) == $signed(129'sh0);
  assign _EVAL_122 = _EVAL_86 | _EVAL_103;
  assign _EVAL_50 = _EVAL_122 | _EVAL_72;
  assign _EVAL_51 = _EVAL_75[1:0];
  assign _EVAL_35 = _EVAL_21[31:24];
  assign _EVAL_58 = _EVAL_21[23:16];
  assign _EVAL_89 = _EVAL_21[15:8];
  assign _EVAL_39 = _EVAL_21[7:0];
  assign _EVAL_85 = 2'h1 == _EVAL_51 ? _EVAL_89 : _EVAL_39;
  assign _EVAL_145 = 2'h2 == _EVAL_51 ? _EVAL_58 : _EVAL_85;
  assign _EVAL_90 = 2'h3 == _EVAL_51 ? _EVAL_35 : _EVAL_145;
  assign _EVAL_73 = _EVAL_28 ^ 128'h20000000;
  assign _EVAL_55 = {1'b0,$signed(_EVAL_73)};
  assign _EVAL_62 = $signed(_EVAL_55) & $signed(-129'sh2000);
  assign _EVAL_147 = $signed(_EVAL_62);
  assign _EVAL_120 = _EVAL_75 == 3'h3;
  assign _EVAL_66 = _EVAL_97 & d__EVAL_1;
  assign _EVAL_47 = _EVAL_28[31:0];
  assign _EVAL_33 = _EVAL_50 | _EVAL_69;
  assign _EVAL_30 = _EVAL_75 == 3'h1;
  assign _EVAL_29 = {{1'd0}, _EVAL_5};
  assign _EVAL_92 = $signed(_EVAL_147) == $signed(129'sh0);
  assign _EVAL_13 = _EVAL_36 ? _EVAL_29 : _EVAL_29;
  assign _EVAL_3 = _EVAL_119 & _EVAL_30;
  assign d__EVAL_5 = _EVAL_1;
  assign _EVAL_19 = d__EVAL_3;
  assign d__EVAL_9 = _EVAL_110 | _EVAL_97;
  assign _EVAL_0 = _EVAL_119 & _EVAL_84;
  assign _EVAL_15 = _EVAL_119 & _EVAL_133;
  assign d__EVAL_7 = _EVAL;
  assign _EVAL_9 = _EVAL_66 & d__EVAL_9;
  assign d__EVAL_0 = _EVAL_18;
  assign _EVAL_14 = _EVAL_130;
  assign _EVAL_10 = _EVAL_36 ? _EVAL_47 : _EVAL_47;
  assign d__EVAL_10 = _EVAL_16;
  assign _EVAL_27 = _EVAL_36 ? 8'h0 : _EVAL_90;
  assign _EVAL_22 = _EVAL_119 & _EVAL_120;
  assign _EVAL_8 = d__EVAL | d__EVAL_2;
  assign _EVAL_7 = _EVAL_33 | _EVAL_92;
  assign _EVAL_2 = _EVAL_36 | _EVAL_49;
  assign _EVAL_23 = _EVAL_36 ? 3'h4 : 3'h0;
  assign _EVAL_6 = _EVAL_33 | _EVAL_92;
  assign _EVAL_12 = _EVAL_119 & _EVAL_44;
  assign d__EVAL_6 = _EVAL_20;
  assign d__EVAL_4 = _EVAL_24;
  assign _EVAL_26 = d__EVAL_8;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_75 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_130 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_18) begin
    if (_EVAL_20) begin
      _EVAL_75 <= 3'h0;
    end else begin
      if (_EVAL_141) begin
        _EVAL_75 <= 3'h0;
      end else begin
        if (_EVAL_118) begin
          _EVAL_75 <= _EVAL_121;
        end
      end
    end
    if (_EVAL_20) begin
      _EVAL_130 <= 3'h0;
    end else begin
      if (_EVAL_136) begin
        _EVAL_130 <= 3'h0;
      end else begin
        if (_EVAL_117) begin
          if (_EVAL_83) begin
            _EVAL_130 <= 3'h1;
          end else begin
            if (_EVAL_81) begin
              _EVAL_130 <= 3'h2;
            end
          end
        end else begin
          if (_EVAL_36) begin
            if (_EVAL_123) begin
              _EVAL_130 <= 3'h3;
            end
          end else begin
            if (_EVAL_49) begin
              if (_EVAL_132) begin
                _EVAL_130 <= 3'h4;
              end
            end else begin
              if (_EVAL_110) begin
                if (_EVAL_135) begin
                  _EVAL_130 <= 3'h0;
                end
              end else begin
                if (_EVAL_97) begin
                  if (_EVAL_78) begin
                    _EVAL_130 <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
