//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_323_assert(
  input  [8:0]  _EVAL,
  input  [7:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [8:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input  [31:0] _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_20;
  reg [31:0] _RAND_0;
  reg [31:0] _EVAL_23;
  reg [31:0] _RAND_1;
  reg  _EVAL_25;
  reg [31:0] _RAND_2;
  reg [2:0] _EVAL_26;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_35;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_62;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_104;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_111;
  reg [31:0] _RAND_7;
  reg [2:0] _EVAL_138;
  reg [31:0] _RAND_8;
  reg [511:0] _EVAL_156;
  reg [511:0] _RAND_9;
  reg [2:0] _EVAL_158;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_176;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_185;
  reg [31:0] _RAND_12;
  reg [8:0] _EVAL_268;
  reg [31:0] _RAND_13;
  reg [8:0] _EVAL_273;
  reg [31:0] _RAND_14;
  wire [1:0] _EVAL_114;
  wire [3:0] _EVAL_75;
  wire [2:0] _EVAL_169;
  wire [2:0] _EVAL_44;
  wire  _EVAL_184;
  wire  _EVAL_121;
  wire  _EVAL_237;
  wire  _EVAL_38;
  wire  _EVAL_91;
  wire  _EVAL_202;
  wire  _EVAL_33;
  wire  _EVAL_152;
  wire  _EVAL_76;
  wire  _EVAL_88;
  wire  _EVAL_71;
  wire  _EVAL_145;
  wire  _EVAL_107;
  wire  _EVAL_157;
  wire  _EVAL_190;
  wire  _EVAL_281;
  wire  _EVAL_140;
  wire  _EVAL_163;
  wire  _EVAL_215;
  wire  _EVAL_29;
  wire  _EVAL_68;
  wire  _EVAL_49;
  wire  _EVAL_159;
  wire  _EVAL_103;
  wire  _EVAL_180;
  wire [31:0] _EVAL_51;
  wire [32:0] _EVAL_276;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_108;
  wire  _EVAL_267;
  wire  _EVAL_52;
  wire  _EVAL_124;
  wire  _EVAL_148;
  wire  _EVAL_85;
  wire  _EVAL_133;
  wire  _EVAL_257;
  wire  _EVAL_116;
  wire  _EVAL_222;
  wire  _EVAL_220;
  wire  _EVAL_92;
  wire  _EVAL_197;
  wire  _EVAL_204;
  wire  _EVAL_167;
  wire  _EVAL_66;
  wire  _EVAL_73;
  wire [511:0] _EVAL_235;
  wire [511:0] _EVAL_120;
  wire  _EVAL_149;
  wire  _EVAL_198;
  wire  _EVAL_123;
  wire  _EVAL_41;
  wire  _EVAL_146;
  wire  _EVAL_87;
  wire [511:0] _EVAL_69;
  wire [511:0] _EVAL_48;
  wire  _EVAL_214;
  wire  _EVAL_193;
  wire  _EVAL_126;
  wire  _EVAL_265;
  wire  _EVAL_253;
  wire [12:0] _EVAL_208;
  wire [5:0] _EVAL_53;
  wire [5:0] _EVAL_32;
  wire [31:0] _EVAL_251;
  wire [31:0] _EVAL_275;
  wire  _EVAL_236;
  wire  _EVAL_187;
  wire  _EVAL_117;
  wire  _EVAL_233;
  wire  _EVAL_56;
  wire  _EVAL_72;
  wire  _EVAL_128;
  wire  _EVAL_37;
  wire [2:0] _EVAL_55;
  wire  _EVAL_28;
  wire  _EVAL_80;
  wire [2:0] _EVAL_252;
  wire  _EVAL_224;
  wire  _EVAL_143;
  wire  _EVAL_194;
  wire  _EVAL_263;
  wire  _EVAL_229;
  wire  _EVAL_227;
  wire  _EVAL_39;
  wire  _EVAL_30;
  wire  _EVAL_219;
  wire  _EVAL_186;
  wire  _EVAL_142;
  wire  _EVAL_247;
  wire  _EVAL_188;
  wire  _EVAL_98;
  wire  _EVAL_70;
  wire  _EVAL_199;
  wire  _EVAL_170;
  wire  _EVAL_67;
  wire  _EVAL_31;
  wire  _EVAL_136;
  wire  _EVAL_93;
  wire [7:0] _EVAL_95;
  wire [7:0] _EVAL_105;
  wire [7:0] _EVAL_272;
  wire  _EVAL_261;
  wire  _EVAL_110;
  wire  _EVAL_213;
  wire [2:0] _EVAL_118;
  wire  _EVAL_154;
  wire  _EVAL_231;
  wire [511:0] _EVAL_238;
  wire  _EVAL_97;
  wire  _EVAL_217;
  wire  _EVAL_94;
  wire  _EVAL_239;
  wire  _EVAL_50;
  wire [12:0] _EVAL_40;
  wire [5:0] _EVAL_205;
  wire [5:0] _EVAL_65;
  wire [2:0] _EVAL_135;
  wire  _EVAL_144;
  wire  _EVAL_256;
  wire  _EVAL_280;
  wire  _EVAL_211;
  wire  _EVAL_259;
  wire  _EVAL_209;
  wire  _EVAL_54;
  wire [511:0] _EVAL_89;
  wire  _EVAL_228;
  wire  _EVAL_119;
  wire  _EVAL_109;
  wire  _EVAL_125;
  wire  _EVAL_99;
  wire [511:0] _EVAL_79;
  wire [511:0] _EVAL_221;
  wire  _EVAL_24;
  wire  _EVAL_166;
  wire  _EVAL_250;
  wire  _EVAL_207;
  wire [2:0] _EVAL_153;
  wire  _EVAL_83;
  wire  _EVAL_175;
  wire  _EVAL_61;
  wire  _EVAL_225;
  wire  _EVAL_19;
  wire  _EVAL_74;
  wire  _EVAL_177;
  wire  _EVAL_262;
  wire  _EVAL_226;
  wire  _EVAL_42;
  wire  _EVAL_150;
  wire  _EVAL_36;
  wire  _EVAL_249;
  wire  _EVAL_270;
  wire  _EVAL_246;
  wire [511:0] _EVAL_129;
  wire  _EVAL_200;
  wire  _EVAL_210;
  wire  _EVAL_160;
  wire  _EVAL_203;
  wire  _EVAL_131;
  wire  _EVAL_59;
  wire  _EVAL_134;
  wire  _EVAL_241;
  wire  _EVAL_34;
  wire  _EVAL_63;
  wire  _EVAL_279;
  wire  _EVAL_282;
  wire  _EVAL_277;
  wire  _EVAL_171;
  wire  _EVAL_182;
  wire [7:0] _EVAL_174;
  wire  _EVAL_201;
  wire  _EVAL_27;
  wire  _EVAL_178;
  wire  _EVAL_216;
  wire  _EVAL_84;
  wire  _EVAL_22;
  wire  _EVAL_137;
  wire [2:0] _EVAL_122;
  wire  _EVAL_271;
  wire  _EVAL_243;
  wire  _EVAL_269;
  wire  _EVAL_274;
  wire  _EVAL_248;
  wire  _EVAL_112;
  wire  _EVAL_230;
  wire  _EVAL_130;
  wire  _EVAL_21;
  wire  _EVAL_183;
  wire  _EVAL_283;
  wire  _EVAL_141;
  wire  _EVAL_60;
  wire  _EVAL_223;
  wire  _EVAL_96;
  wire  _EVAL_139;
  wire  _EVAL_161;
  wire  _EVAL_101;
  wire [31:0] _EVAL_82;
  wire  _EVAL_232;
  wire  _EVAL_181;
  wire  _EVAL_255;
  wire  _EVAL_64;
  wire  _EVAL_254;
  wire  _EVAL_58;
  wire  _EVAL_102;
  wire  _EVAL_151;
  wire  _EVAL_278;
  wire  _EVAL_195;
  wire  _EVAL_155;
  wire  _EVAL_264;
  wire  _EVAL_43;
  wire  _EVAL_245;
  wire  _EVAL_189;
  wire  _EVAL_90;
  wire  _EVAL_113;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_78;
  wire  _EVAL_165;
  wire  _EVAL_196;
  wire  _EVAL_206;
  wire  _EVAL_77;
  wire  _EVAL_132;
  wire  _EVAL_18;
  wire  _EVAL_258;
  wire  _EVAL_212;
  wire [511:0] _EVAL_191;
  wire  _EVAL_260;
  wire  _EVAL_168;
  wire  _EVAL_244;
  wire  _EVAL_179;
  wire  _EVAL_266;
  wire  _EVAL_234;
  wire  _EVAL_106;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_114 = _EVAL_1[1:0];
  assign _EVAL_75 = 4'h1 << _EVAL_114;
  assign _EVAL_169 = _EVAL_75[2:0];
  assign _EVAL_44 = _EVAL_169 | 3'h1;
  assign _EVAL_184 = _EVAL_44[1];
  assign _EVAL_121 = _EVAL_176 == 3'h0;
  assign _EVAL_237 = _EVAL_121 == 1'h0;
  assign _EVAL_38 = _EVAL_5 == 3'h4;
  assign _EVAL_91 = _EVAL_1 >= 3'h3;
  assign _EVAL_202 = _EVAL_44[2];
  assign _EVAL_33 = _EVAL_16[2];
  assign _EVAL_152 = _EVAL_33 == 1'h0;
  assign _EVAL_76 = _EVAL_202 & _EVAL_152;
  assign _EVAL_88 = _EVAL_91 | _EVAL_76;
  assign _EVAL_71 = _EVAL_16[1];
  assign _EVAL_145 = _EVAL_152 & _EVAL_71;
  assign _EVAL_107 = _EVAL_184 & _EVAL_145;
  assign _EVAL_157 = _EVAL_88 | _EVAL_107;
  assign _EVAL_190 = _EVAL_12 >= 3'h3;
  assign _EVAL_281 = _EVAL_71 == 1'h0;
  assign _EVAL_140 = _EVAL_152 & _EVAL_281;
  assign _EVAL_163 = _EVAL_184 & _EVAL_140;
  assign _EVAL_215 = _EVAL_88 | _EVAL_163;
  assign _EVAL_29 = _EVAL_44[0];
  assign _EVAL_68 = _EVAL_16[0];
  assign _EVAL_49 = _EVAL_68 == 1'h0;
  assign _EVAL_159 = _EVAL_140 & _EVAL_49;
  assign _EVAL_103 = _EVAL_29 & _EVAL_159;
  assign _EVAL_180 = _EVAL_215 | _EVAL_103;
  assign _EVAL_51 = _EVAL_16 ^ 32'h80000000;
  assign _EVAL_276 = {1'b0,$signed(_EVAL_51)};
  assign _EVAL_172 = $signed(_EVAL_276) & $signed(-33'sh20000);
  assign _EVAL_108 = $signed(_EVAL_172);
  assign _EVAL_267 = $signed(_EVAL_108) == $signed(33'sh0);
  assign _EVAL_52 = _EVAL_1 == _EVAL_35;
  assign _EVAL_124 = _EVAL_52 | _EVAL_8;
  assign _EVAL_148 = _EVAL_124 == 1'h0;
  assign _EVAL_85 = _EVAL_10 == 3'h0;
  assign _EVAL_133 = _EVAL_202 & _EVAL_33;
  assign _EVAL_257 = _EVAL_91 | _EVAL_133;
  assign _EVAL_116 = _EVAL_33 & _EVAL_71;
  assign _EVAL_222 = _EVAL_184 & _EVAL_116;
  assign _EVAL_220 = _EVAL_257 | _EVAL_222;
  assign _EVAL_92 = _EVAL_116 & _EVAL_68;
  assign _EVAL_197 = _EVAL_29 & _EVAL_92;
  assign _EVAL_204 = _EVAL_220 | _EVAL_197;
  assign _EVAL_167 = _EVAL_15 & _EVAL_11;
  assign _EVAL_66 = _EVAL_62 == 3'h0;
  assign _EVAL_73 = _EVAL_167 & _EVAL_66;
  assign _EVAL_235 = 512'h1 << _EVAL;
  assign _EVAL_120 = _EVAL_73 ? _EVAL_235 : 512'h0;
  assign _EVAL_149 = _EVAL_6 & _EVAL_7;
  assign _EVAL_198 = _EVAL_26 == 3'h0;
  assign _EVAL_123 = _EVAL_149 & _EVAL_198;
  assign _EVAL_41 = _EVAL_5 == 3'h6;
  assign _EVAL_146 = _EVAL_41 == 1'h0;
  assign _EVAL_87 = _EVAL_123 & _EVAL_146;
  assign _EVAL_69 = 512'h1 << _EVAL_9;
  assign _EVAL_48 = _EVAL_87 ? _EVAL_69 : 512'h0;
  assign _EVAL_214 = _EVAL_120 != _EVAL_48;
  assign _EVAL_193 = _EVAL_120 != 512'h0;
  assign _EVAL_126 = _EVAL_193 == 1'h0;
  assign _EVAL_265 = _EVAL_214 | _EVAL_126;
  assign _EVAL_253 = _EVAL_265 | _EVAL_8;
  assign _EVAL_208 = 13'h3f << _EVAL_1;
  assign _EVAL_53 = _EVAL_208[5:0];
  assign _EVAL_32 = ~ _EVAL_53;
  assign _EVAL_251 = {{26'd0}, _EVAL_32};
  assign _EVAL_275 = _EVAL_16 & _EVAL_251;
  assign _EVAL_236 = _EVAL_275 == 32'h0;
  assign _EVAL_187 = _EVAL_236 | _EVAL_8;
  assign _EVAL_117 = _EVAL_187 == 1'h0;
  assign _EVAL_233 = _EVAL_10 == 3'h1;
  assign _EVAL_56 = _EVAL_10 == 3'h4;
  assign _EVAL_72 = _EVAL_3 == 1'h0;
  assign _EVAL_128 = _EVAL_156 != 512'h0;
  assign _EVAL_37 = _EVAL_128 == 1'h0;
  assign _EVAL_55 = _EVAL_26 - 3'h1;
  assign _EVAL_28 = _EVAL_10[2];
  assign _EVAL_80 = _EVAL_28 == 1'h0;
  assign _EVAL_252 = _EVAL_32[5:3];
  assign _EVAL_224 = _EVAL_116 & _EVAL_49;
  assign _EVAL_143 = _EVAL_29 & _EVAL_224;
  assign _EVAL_194 = _EVAL_220 | _EVAL_143;
  assign _EVAL_263 = _EVAL_33 & _EVAL_281;
  assign _EVAL_229 = _EVAL_184 & _EVAL_263;
  assign _EVAL_227 = _EVAL_257 | _EVAL_229;
  assign _EVAL_39 = _EVAL_263 & _EVAL_68;
  assign _EVAL_30 = _EVAL_29 & _EVAL_39;
  assign _EVAL_219 = _EVAL_227 | _EVAL_30;
  assign _EVAL_186 = _EVAL_263 & _EVAL_49;
  assign _EVAL_142 = _EVAL_29 & _EVAL_186;
  assign _EVAL_247 = _EVAL_227 | _EVAL_142;
  assign _EVAL_188 = _EVAL_145 & _EVAL_68;
  assign _EVAL_98 = _EVAL_29 & _EVAL_188;
  assign _EVAL_70 = _EVAL_157 | _EVAL_98;
  assign _EVAL_199 = _EVAL_145 & _EVAL_49;
  assign _EVAL_170 = _EVAL_29 & _EVAL_199;
  assign _EVAL_67 = _EVAL_157 | _EVAL_170;
  assign _EVAL_31 = _EVAL_140 & _EVAL_68;
  assign _EVAL_136 = _EVAL_29 & _EVAL_31;
  assign _EVAL_93 = _EVAL_215 | _EVAL_136;
  assign _EVAL_95 = {_EVAL_204,_EVAL_194,_EVAL_219,_EVAL_247,_EVAL_70,_EVAL_67,_EVAL_93,_EVAL_180};
  assign _EVAL_105 = ~ _EVAL_95;
  assign _EVAL_272 = _EVAL_0 & _EVAL_105;
  assign _EVAL_261 = _EVAL_272 == 8'h0;
  assign _EVAL_110 = _EVAL_261 | _EVAL_8;
  assign _EVAL_213 = _EVAL_110 == 1'h0;
  assign _EVAL_118 = _EVAL_138 - 3'h1;
  assign _EVAL_154 = _EVAL_7 & _EVAL_38;
  assign _EVAL_231 = _EVAL_10 == _EVAL_158;
  assign _EVAL_238 = _EVAL_156 | _EVAL_120;
  assign _EVAL_97 = _EVAL_138 == 3'h0;
  assign _EVAL_217 = _EVAL_97 == 1'h0;
  assign _EVAL_94 = _EVAL_11 & _EVAL_217;
  assign _EVAL_239 = _EVAL_13 == 1'h0;
  assign _EVAL_50 = _EVAL_5[0];
  assign _EVAL_40 = 13'h3f << _EVAL_12;
  assign _EVAL_205 = _EVAL_40[5:0];
  assign _EVAL_65 = ~ _EVAL_205;
  assign _EVAL_135 = _EVAL_65[5:3];
  assign _EVAL_144 = _EVAL_1 <= 3'h6;
  assign _EVAL_256 = _EVAL_5 == 3'h5;
  assign _EVAL_280 = _EVAL_2 == _EVAL_25;
  assign _EVAL_211 = _EVAL_280 | _EVAL_8;
  assign _EVAL_259 = _EVAL_5 == _EVAL_185;
  assign _EVAL_209 = _EVAL_259 | _EVAL_8;
  assign _EVAL_54 = _EVAL_209 == 1'h0;
  assign _EVAL_89 = _EVAL_156 >> _EVAL;
  assign _EVAL_228 = _EVAL_89[0];
  assign _EVAL_119 = _EVAL_228 == 1'h0;
  assign _EVAL_109 = _EVAL_14 <= 3'h4;
  assign _EVAL_125 = _EVAL_109 | _EVAL_8;
  assign _EVAL_99 = _EVAL_125 == 1'h0;
  assign _EVAL_79 = _EVAL_120 | _EVAL_156;
  assign _EVAL_221 = _EVAL_79 >> _EVAL_9;
  assign _EVAL_24 = _EVAL_221[0];
  assign _EVAL_166 = _EVAL_24 | _EVAL_8;
  assign _EVAL_250 = _EVAL_5 == 3'h2;
  assign _EVAL_207 = _EVAL_7 & _EVAL_250;
  assign _EVAL_153 = _EVAL_62 - 3'h1;
  assign _EVAL_83 = _EVAL_14 <= 3'h2;
  assign _EVAL_175 = _EVAL_83 | _EVAL_8;
  assign _EVAL_61 = _EVAL_167 | _EVAL_149;
  assign _EVAL_225 = _EVAL_16 == _EVAL_111;
  assign _EVAL_19 = _EVAL_225 | _EVAL_8;
  assign _EVAL_74 = _EVAL_10 == 3'h5;
  assign _EVAL_177 = _EVAL_11 & _EVAL_74;
  assign _EVAL_262 = _EVAL_10 == 3'h2;
  assign _EVAL_226 = _EVAL_9 == _EVAL_273;
  assign _EVAL_42 = _EVAL_226 | _EVAL_8;
  assign _EVAL_150 = _EVAL_42 == 1'h0;
  assign _EVAL_36 = _EVAL_2 == 1'h0;
  assign _EVAL_249 = _EVAL_36 | _EVAL_8;
  assign _EVAL_270 = _EVAL_11 & _EVAL_262;
  assign _EVAL_246 = _EVAL_253 == 1'h0;
  assign _EVAL_129 = ~ _EVAL_48;
  assign _EVAL_200 = _EVAL_14 != 3'h0;
  assign _EVAL_210 = _EVAL_200 | _EVAL_8;
  assign _EVAL_160 = plusarg_reader_out == 32'h0;
  assign _EVAL_203 = _EVAL_37 | _EVAL_160;
  assign _EVAL_131 = _EVAL_23 < plusarg_reader_out;
  assign _EVAL_59 = _EVAL_203 | _EVAL_131;
  assign _EVAL_134 = _EVAL_59 | _EVAL_8;
  assign _EVAL_241 = _EVAL_134 == 1'h0;
  assign _EVAL_34 = _EVAL_7 & _EVAL_237;
  assign _EVAL_63 = _EVAL_5 <= 3'h6;
  assign _EVAL_279 = _EVAL_36 | _EVAL_13;
  assign _EVAL_282 = _EVAL_279 | _EVAL_8;
  assign _EVAL_277 = _EVAL_282 == 1'h0;
  assign _EVAL_171 = _EVAL_239 | _EVAL_8;
  assign _EVAL_182 = _EVAL_171 == 1'h0;
  assign _EVAL_174 = ~ _EVAL_0;
  assign _EVAL_201 = _EVAL_174 == 8'h0;
  assign _EVAL_27 = _EVAL_201 | _EVAL_8;
  assign _EVAL_178 = _EVAL_27 == 1'h0;
  assign _EVAL_216 = _EVAL_10 == 3'h3;
  assign _EVAL_84 = _EVAL_11 & _EVAL_216;
  assign _EVAL_22 = _EVAL == _EVAL_268;
  assign _EVAL_137 = _EVAL_22 | _EVAL_8;
  assign _EVAL_122 = _EVAL_176 - 3'h1;
  assign _EVAL_271 = _EVAL_10 == 3'h6;
  assign _EVAL_243 = _EVAL_249 == 1'h0;
  assign _EVAL_269 = _EVAL_14 == _EVAL_104;
  assign _EVAL_274 = _EVAL_269 | _EVAL_8;
  assign _EVAL_248 = _EVAL_231 | _EVAL_8;
  assign _EVAL_112 = _EVAL_91 | _EVAL_8;
  assign _EVAL_230 = _EVAL_0 == _EVAL_95;
  assign _EVAL_130 = _EVAL_14 <= 3'h3;
  assign _EVAL_21 = _EVAL_130 | _EVAL_8;
  assign _EVAL_183 = _EVAL_21 == 1'h0;
  assign _EVAL_283 = _EVAL_11 & _EVAL_233;
  assign _EVAL_141 = _EVAL_11 & _EVAL_56;
  assign _EVAL_60 = _EVAL_5 == 3'h1;
  assign _EVAL_223 = _EVAL_10 == 3'h7;
  assign _EVAL_96 = _EVAL_11 & _EVAL_223;
  assign _EVAL_139 = _EVAL_175 == 1'h0;
  assign _EVAL_161 = _EVAL_5 == 3'h0;
  assign _EVAL_101 = _EVAL_63 | _EVAL_8;
  assign _EVAL_82 = _EVAL_23 + 32'h1;
  assign _EVAL_232 = _EVAL_19 == 1'h0;
  assign _EVAL_181 = _EVAL_190 | _EVAL_8;
  assign _EVAL_255 = _EVAL_12 == _EVAL_20;
  assign _EVAL_64 = _EVAL_230 | _EVAL_8;
  assign _EVAL_254 = _EVAL_64 == 1'h0;
  assign _EVAL_58 = _EVAL_144 & _EVAL_267;
  assign _EVAL_102 = _EVAL_58 | _EVAL_8;
  assign _EVAL_151 = _EVAL_102 == 1'h0;
  assign _EVAL_278 = _EVAL_11 & _EVAL_271;
  assign _EVAL_195 = _EVAL_14 == 3'h0;
  assign _EVAL_155 = _EVAL_255 | _EVAL_8;
  assign _EVAL_264 = _EVAL_155 == 1'h0;
  assign _EVAL_43 = _EVAL_167 & _EVAL_97;
  assign _EVAL_245 = _EVAL_119 | _EVAL_8;
  assign _EVAL_189 = _EVAL_245 == 1'h0;
  assign _EVAL_90 = _EVAL_7 & _EVAL_161;
  assign _EVAL_113 = _EVAL_72 | _EVAL_8;
  assign _EVAL_46 = _EVAL_113 == 1'h0;
  assign _EVAL_47 = _EVAL_166 == 1'h0;
  assign _EVAL_78 = _EVAL_274 == 1'h0;
  assign _EVAL_165 = _EVAL_8 == 1'h0;
  assign _EVAL_196 = _EVAL_7 & _EVAL_41;
  assign _EVAL_206 = _EVAL_101 == 1'h0;
  assign _EVAL_77 = _EVAL_210 == 1'h0;
  assign _EVAL_132 = _EVAL_195 | _EVAL_8;
  assign _EVAL_18 = _EVAL_11 & _EVAL_85;
  assign _EVAL_258 = _EVAL_248 == 1'h0;
  assign _EVAL_212 = _EVAL_7 & _EVAL_256;
  assign _EVAL_191 = _EVAL_238 & _EVAL_129;
  assign _EVAL_260 = _EVAL_211 == 1'h0;
  assign _EVAL_168 = _EVAL_137 == 1'h0;
  assign _EVAL_244 = _EVAL_112 == 1'h0;
  assign _EVAL_179 = _EVAL_149 & _EVAL_121;
  assign _EVAL_266 = _EVAL_132 == 1'h0;
  assign _EVAL_234 = _EVAL_181 == 1'h0;
  assign _EVAL_106 = _EVAL_7 & _EVAL_60;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_23 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_26 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_35 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_62 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_104 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_111 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_138 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {16{`RANDOM}};
  _EVAL_156 = _RAND_9[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_158 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_176 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_185 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_268 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_273 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_4) begin
    if (_EVAL_179) begin
      _EVAL_20 <= _EVAL_12;
    end
    if (_EVAL_8) begin
      _EVAL_23 <= 32'h0;
    end else begin
      if (_EVAL_61) begin
        _EVAL_23 <= 32'h0;
      end else begin
        _EVAL_23 <= _EVAL_82;
      end
    end
    if (_EVAL_179) begin
      _EVAL_25 <= _EVAL_2;
    end
    if (_EVAL_8) begin
      _EVAL_26 <= 3'h0;
    end else begin
      if (_EVAL_149) begin
        if (_EVAL_198) begin
          if (_EVAL_50) begin
            _EVAL_26 <= _EVAL_135;
          end else begin
            _EVAL_26 <= 3'h0;
          end
        end else begin
          _EVAL_26 <= _EVAL_55;
        end
      end
    end
    if (_EVAL_43) begin
      _EVAL_35 <= _EVAL_1;
    end
    if (_EVAL_8) begin
      _EVAL_62 <= 3'h0;
    end else begin
      if (_EVAL_167) begin
        if (_EVAL_66) begin
          if (_EVAL_80) begin
            _EVAL_62 <= _EVAL_252;
          end else begin
            _EVAL_62 <= 3'h0;
          end
        end else begin
          _EVAL_62 <= _EVAL_153;
        end
      end
    end
    if (_EVAL_43) begin
      _EVAL_104 <= _EVAL_14;
    end
    if (_EVAL_43) begin
      _EVAL_111 <= _EVAL_16;
    end
    if (_EVAL_8) begin
      _EVAL_138 <= 3'h0;
    end else begin
      if (_EVAL_167) begin
        if (_EVAL_97) begin
          if (_EVAL_80) begin
            _EVAL_138 <= _EVAL_252;
          end else begin
            _EVAL_138 <= 3'h0;
          end
        end else begin
          _EVAL_138 <= _EVAL_118;
        end
      end
    end
    if (_EVAL_8) begin
      _EVAL_156 <= 512'h0;
    end else begin
      _EVAL_156 <= _EVAL_191;
    end
    if (_EVAL_43) begin
      _EVAL_158 <= _EVAL_10;
    end
    if (_EVAL_8) begin
      _EVAL_176 <= 3'h0;
    end else begin
      if (_EVAL_149) begin
        if (_EVAL_121) begin
          if (_EVAL_50) begin
            _EVAL_176 <= _EVAL_135;
          end else begin
            _EVAL_176 <= 3'h0;
          end
        end else begin
          _EVAL_176 <= _EVAL_122;
        end
      end
    end
    if (_EVAL_179) begin
      _EVAL_185 <= _EVAL_5;
    end
    if (_EVAL_43) begin
      _EVAL_268 <= _EVAL;
    end
    if (_EVAL_179) begin
      _EVAL_273 <= _EVAL_9;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba9a45d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(521c889d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa4b1171)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1580e5d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30793217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f1c4636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fce97426)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42ce9647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4db7559f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58caf125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854ff628)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5b200fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf646b1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f08fc901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0bac354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aee1d24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da83092d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(137b5f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab80f0e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a64fa00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49543278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5091979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72fc522c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79139b72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(653fde77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380dc372)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d4d5427)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(237cd3e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d151f8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d512f4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cc696b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab59e273)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f88893ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f44da7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c57d068)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4bf4331)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dad4f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc28a13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52fcd8e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a868d0f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a14d02ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(844d226c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(685e7af2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(597c811d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81795b08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31edf4d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5101056a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa546d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(270e9f23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(742cb593)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fd489dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(347e51fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a299eaae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36ac369c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1bb0365)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91bfd4b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bbc8d92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eb96262)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3391ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f080aff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbfc9cd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14b65548)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8689bc70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd2631f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8501a352)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2401901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
