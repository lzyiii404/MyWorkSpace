//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_253(
  input  [63:0] _EVAL,
  input  [2:0]  _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  output [2:0]  _EVAL_3,
  output [63:0] _EVAL_4,
  output        _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  output        _EVAL_10,
  input  [2:0]  _EVAL_11,
  output [7:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [7:0]  _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output [3:0]  _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input  [2:0]  _EVAL_29,
  output        _EVAL_30,
  output [2:0]  _EVAL_31,
  output [31:0] _EVAL_32,
  input  [3:0]  _EVAL_33,
  input  [2:0]  _EVAL_34,
  input  [31:0] _EVAL_35,
  input         _EVAL_36,
  output [63:0] _EVAL_37,
  input  [63:0] _EVAL_38,
  output        _EVAL_39,
  output [2:0]  _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  output [63:0] _EVAL_43,
  output [63:0] _EVAL_44,
  output        _EVAL_45,
  output [3:0]  _EVAL_46,
  output        _EVAL_47,
  input  [63:0] _EVAL_48,
  input  [2:0]  _EVAL_49,
  input  [1:0]  _EVAL_50,
  output        _EVAL_51,
  output [2:0]  _EVAL_52,
  output        _EVAL_53,
  input  [2:0]  _EVAL_54,
  output [7:0]  _EVAL_55,
  input         _EVAL_56,
  output [2:0]  _EVAL_57,
  input         _EVAL_58,
  output        _EVAL_59,
  output        _EVAL_60,
  output [1:0]  _EVAL_61,
  output        _EVAL_62,
  output [1:0]  _EVAL_63,
  output [2:0]  _EVAL_64,
  output [2:0]  _EVAL_65,
  output [2:0]  _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_68,
  output [2:0]  _EVAL_69,
  input  [63:0] _EVAL_70,
  output [31:0] _EVAL_71,
  output        _EVAL_72,
  input  [1:0]  _EVAL_73,
  output [2:0]  _EVAL_74,
  output        _EVAL_75,
  output [24:0] _EVAL_76,
  input         _EVAL_77,
  output [31:0] _EVAL_78,
  input         _EVAL_79,
  output [2:0]  _EVAL_80,
  output [2:0]  _EVAL_81,
  input  [2:0]  _EVAL_82,
  input  [2:0]  _EVAL_83,
  input  [31:0] _EVAL_84,
  output [3:0]  _EVAL_85,
  output        _EVAL_86,
  output        _EVAL_87,
  input         _EVAL_88
);
  reg  _EVAL_98;
  reg [31:0] _RAND_0;
  reg [1:0] _EVAL_123;
  reg [31:0] _RAND_1;
  reg  _EVAL_132;
  reg [31:0] _RAND_2;
  reg [4:0] _EVAL_175;
  reg [31:0] _RAND_3;
  wire [3:0] _EVAL_190;
  wire [22:0] _EVAL_193;
  wire [31:0] _EVAL_152;
  wire [32:0] _EVAL_158;
  wire [32:0] _EVAL_110;
  wire [32:0] _EVAL_146;
  wire [1:0] _EVAL_163;
  wire [31:0] _EVAL_145;
  wire [32:0] _EVAL_149;
  wire [1:0] _EVAL_138;
  wire [1:0] _EVAL_203;
  wire [3:0] _EVAL_113;
  wire [2:0] _EVAL_94;
  wire [3:0] _EVAL_165;
  wire [3:0] _EVAL_99;
  wire [2:0] _EVAL_139;
  wire [3:0] _EVAL_114;
  wire [3:0] _EVAL_121;
  wire [3:0] _EVAL_196;
  wire [1:0] _EVAL_97;
  wire [1:0] _EVAL_185;
  wire [1:0] _EVAL_187;
  wire [1:0] _EVAL_140;
  wire  _EVAL_91;
  wire  _EVAL_172;
  wire  _EVAL_168;
  wire  _EVAL_122;
  wire [20:0] _EVAL_199;
  wire [5:0] _EVAL_181;
  wire [5:0] _EVAL_151;
  wire [2:0] _EVAL_179;
  wire [2:0] _EVAL_200;
  wire [2:0] _EVAL_154;
  wire [32:0] _EVAL_156;
  wire [32:0] _EVAL_89;
  wire  _EVAL_204;
  wire  _EVAL_136;
  wire  _EVAL_195;
  wire [32:0] _EVAL_130;
  wire [32:0] _EVAL_102;
  wire [7:0] _EVAL_184;
  wire [7:0] _EVAL_189;
  wire [32:0] _EVAL_107;
  wire [1:0] _EVAL_117;
  wire [2:0] _EVAL_194;
  wire [31:0] _EVAL_133;
  wire [32:0] _EVAL_171;
  wire [32:0] _EVAL_129;
  wire [32:0] _EVAL_127;
  wire  _EVAL_155;
  wire  _EVAL_182;
  wire  _EVAL_161;
  wire  _EVAL_197;
  wire  _EVAL_119;
  wire  _EVAL_135;
  wire  _EVAL_128;
  wire [31:0] _EVAL_111;
  wire [32:0] _EVAL_131;
  wire [32:0] _EVAL_180;
  wire [32:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_106;
  wire  _EVAL_148;
  wire  _EVAL_104;
  wire [1:0] _EVAL_192;
  wire [1:0] _EVAL_141;
  wire  _EVAL_120;
  wire  _EVAL_126;
  wire  _EVAL_183;
  wire  _EVAL_153;
  wire [4:0] _EVAL_159;
  wire [4:0] _EVAL_116;
  wire [78:0] _EVAL_103;
  wire [4:0] _EVAL_112;
  wire  _EVAL_143;
  wire  _EVAL_92;
  wire  _EVAL_137;
  wire [78:0] _EVAL_96;
  wire  _EVAL_169;
  wire [31:0] _EVAL_142;
  wire  _EVAL_162;
  wire  _EVAL_202;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_157;
  wire [32:0] _EVAL_101;
  wire  _EVAL_173;
  wire  _EVAL_93;
  wire [4:0] _EVAL_100;
  wire [4:0] _EVAL_174;
  wire [78:0] _EVAL_90;
  wire  _EVAL_108;
  wire [78:0] _EVAL_178;
  wire [4:0] _EVAL_144;
  wire [4:0] _EVAL_164;
  wire [78:0] _EVAL_188;
  wire  _EVAL_167;
  assign _EVAL_190 = {{1'd0}, _EVAL_9};
  assign _EVAL_193 = 23'hff << _EVAL_8;
  assign _EVAL_152 = _EVAL_1 ^ 32'h8000000;
  assign _EVAL_158 = {1'b0,$signed(_EVAL_152)};
  assign _EVAL_110 = $signed(_EVAL_158) & $signed(33'she8000000);
  assign _EVAL_146 = $signed(_EVAL_110);
  assign _EVAL_163 = {_EVAL_58,_EVAL_42};
  assign _EVAL_145 = _EVAL_1 ^ 32'h20000000;
  assign _EVAL_149 = {1'b0,$signed(_EVAL_145)};
  assign _EVAL_138 = ~ _EVAL_123;
  assign _EVAL_203 = _EVAL_163 & _EVAL_138;
  assign _EVAL_113 = {_EVAL_203,_EVAL_58,_EVAL_42};
  assign _EVAL_94 = _EVAL_113[3:1];
  assign _EVAL_165 = {{1'd0}, _EVAL_94};
  assign _EVAL_99 = _EVAL_113 | _EVAL_165;
  assign _EVAL_139 = _EVAL_99[3:1];
  assign _EVAL_114 = {{1'd0}, _EVAL_139};
  assign _EVAL_121 = {_EVAL_123, 2'h0};
  assign _EVAL_196 = _EVAL_114 | _EVAL_121;
  assign _EVAL_97 = _EVAL_196[3:2];
  assign _EVAL_185 = _EVAL_196[1:0];
  assign _EVAL_187 = _EVAL_97 & _EVAL_185;
  assign _EVAL_140 = ~ _EVAL_187;
  assign _EVAL_91 = _EVAL_140[0];
  assign _EVAL_172 = _EVAL_132 ? _EVAL_58 : 1'h0;
  assign _EVAL_168 = _EVAL_91 & _EVAL_42;
  assign _EVAL_122 = _EVAL_34[0];
  assign _EVAL_199 = 21'h3f << _EVAL_190;
  assign _EVAL_181 = _EVAL_199[5:0];
  assign _EVAL_151 = ~ _EVAL_181;
  assign _EVAL_179 = _EVAL_151[5:3];
  assign _EVAL_200 = _EVAL_122 ? _EVAL_179 : 3'h0;
  assign _EVAL_154 = _EVAL_168 ? _EVAL_200 : 3'h0;
  assign _EVAL_156 = $signed(_EVAL_149) & $signed(33'she9100000);
  assign _EVAL_89 = $signed(_EVAL_156);
  assign _EVAL_204 = _EVAL_140[1];
  assign _EVAL_136 = _EVAL_204 & _EVAL_58;
  assign _EVAL_195 = _EVAL_42 | _EVAL_58;
  assign _EVAL_130 = {1'b0,$signed(_EVAL_1)};
  assign _EVAL_102 = $signed(_EVAL_130) & $signed(33'sha9100000);
  assign _EVAL_184 = _EVAL_193[7:0];
  assign _EVAL_189 = ~ _EVAL_184;
  assign _EVAL_107 = $signed(_EVAL_102);
  assign _EVAL_117 = _EVAL_140 & _EVAL_163;
  assign _EVAL_194 = {_EVAL_117, 1'h0};
  assign _EVAL_133 = _EVAL_1 ^ 32'h80000000;
  assign _EVAL_171 = {1'b0,$signed(_EVAL_133)};
  assign _EVAL_129 = $signed(_EVAL_171) & $signed(33'she9100000);
  assign _EVAL_127 = $signed(_EVAL_129);
  assign _EVAL_155 = $signed(_EVAL_127) == $signed(33'sh0);
  assign _EVAL_182 = _EVAL_175 == 5'h0;
  assign _EVAL_161 = _EVAL_182 ? _EVAL_91 : _EVAL_98;
  assign _EVAL_197 = $signed(_EVAL_107) == $signed(33'sh0);
  assign _EVAL_119 = _EVAL_197 | _EVAL_155;
  assign _EVAL_135 = $signed(_EVAL_146) == $signed(33'sh0);
  assign _EVAL_128 = _EVAL_119 | _EVAL_135;
  assign _EVAL_111 = _EVAL_1 ^ 32'h1000000;
  assign _EVAL_131 = {1'b0,$signed(_EVAL_111)};
  assign _EVAL_180 = $signed(_EVAL_131) & $signed(33'she9100000);
  assign _EVAL_176 = $signed(_EVAL_180);
  assign _EVAL_177 = $signed(_EVAL_176) == $signed(33'sh0);
  assign _EVAL_106 = _EVAL_128 | _EVAL_177;
  assign _EVAL_148 = $signed(_EVAL_89) == $signed(33'sh0);
  assign _EVAL_104 = _EVAL_106 | _EVAL_148;
  assign _EVAL_192 = _EVAL_194[1:0];
  assign _EVAL_141 = _EVAL_117 | _EVAL_192;
  assign _EVAL_120 = _EVAL_98 ? _EVAL_42 : 1'h0;
  assign _EVAL_126 = _EVAL_120 | _EVAL_172;
  assign _EVAL_183 = _EVAL_182 ? _EVAL_195 : _EVAL_126;
  assign _EVAL_153 = _EVAL_27 & _EVAL_183;
  assign _EVAL_159 = {{4'd0}, _EVAL_153};
  assign _EVAL_116 = _EVAL_175 - _EVAL_159;
  assign _EVAL_103 = {_EVAL_83,_EVAL_73,_EVAL_8,_EVAL_0,_EVAL_68,_EVAL_77,_EVAL_48,_EVAL_26};
  assign _EVAL_112 = _EVAL_189[7:3];
  assign _EVAL_143 = _EVAL_163 != 2'h0;
  assign _EVAL_92 = _EVAL_104 ? _EVAL_36 : 1'h0;
  assign _EVAL_137 = _EVAL_182 ? _EVAL_136 : _EVAL_132;
  assign _EVAL_96 = _EVAL_137 ? _EVAL_103 : 79'h0;
  assign _EVAL_169 = _EVAL_83[0];
  assign _EVAL_142 = _EVAL_1 ^ 32'h1100000;
  assign _EVAL_162 = _EVAL_182 & _EVAL_27;
  assign _EVAL_202 = _EVAL_162 & _EVAL_143;
  assign _EVAL_150 = {1'b0,$signed(_EVAL_142)};
  assign _EVAL_157 = $signed(_EVAL_150) & $signed(33'she9100000);
  assign _EVAL_101 = $signed(_EVAL_157);
  assign _EVAL_173 = $signed(_EVAL_101) == $signed(33'sh0);
  assign _EVAL_93 = _EVAL_173 ? _EVAL_13 : 1'h0;
  assign _EVAL_100 = _EVAL_169 ? _EVAL_112 : 5'h0;
  assign _EVAL_174 = _EVAL_136 ? _EVAL_100 : 5'h0;
  assign _EVAL_90 = {_EVAL_34,2'h0,_EVAL_190,_EVAL_54,2'h0,_EVAL_70,1'h0};
  assign _EVAL_108 = _EVAL_182 ? _EVAL_168 : _EVAL_98;
  assign _EVAL_178 = _EVAL_108 ? _EVAL_90 : 79'h0;
  assign _EVAL_144 = {{2'd0}, _EVAL_154};
  assign _EVAL_164 = _EVAL_144 | _EVAL_174;
  assign _EVAL_188 = _EVAL_178 | _EVAL_96;
  assign _EVAL_167 = _EVAL_182 ? _EVAL_204 : _EVAL_132;
  assign _EVAL_45 = _EVAL_16;
  assign _EVAL_71 = _EVAL_1;
  assign _EVAL_75 = _EVAL_93 | _EVAL_92;
  assign _EVAL_39 = _EVAL_27 & _EVAL_161;
  assign _EVAL_52 = _EVAL_17;
  assign _EVAL_37 = _EVAL;
  assign _EVAL_74 = _EVAL_188[69:67];
  assign _EVAL_5 = _EVAL_2;
  assign _EVAL_81 = _EVAL_33[2:0];
  assign _EVAL_55 = _EVAL_18;
  assign _EVAL_61 = _EVAL_50;
  assign _EVAL_46 = _EVAL_6;
  assign _EVAL_76 = _EVAL_1[24:0];
  assign _EVAL_86 = _EVAL_188[66];
  assign _EVAL_44 = _EVAL;
  assign _EVAL_19 = _EVAL_20 & _EVAL_173;
  assign _EVAL_14 = _EVAL_188[0];
  assign _EVAL_85 = _EVAL_188[73:70];
  assign _EVAL_43 = _EVAL_188[64:1];
  assign _EVAL_32 = _EVAL_35;
  assign _EVAL_51 = _EVAL_20 & _EVAL_104;
  assign _EVAL_40 = _EVAL_29;
  assign _EVAL_10 = _EVAL_21;
  assign _EVAL_62 = _EVAL_79;
  assign _EVAL_66 = _EVAL_11;
  assign _EVAL_15 = _EVAL_27 & _EVAL_167;
  assign _EVAL_4 = _EVAL_38;
  assign _EVAL_53 = _EVAL_88;
  assign _EVAL_65 = _EVAL_49;
  assign _EVAL_60 = _EVAL_67;
  assign _EVAL_63 = _EVAL_188[75:74];
  assign _EVAL_47 = _EVAL_23;
  assign _EVAL_31 = _EVAL_82;
  assign _EVAL_25 = _EVAL_33;
  assign _EVAL_78 = _EVAL_84;
  assign _EVAL_57 = _EVAL_29;
  assign _EVAL_72 = _EVAL_188[65];
  assign _EVAL_30 = _EVAL_28;
  assign _EVAL_80 = _EVAL_17;
  assign _EVAL_12 = _EVAL_18;
  assign _EVAL_64 = _EVAL_22;
  assign _EVAL_41 = _EVAL_182 ? _EVAL_195 : _EVAL_126;
  assign _EVAL_3 = _EVAL_49;
  assign _EVAL_87 = _EVAL_56;
  assign _EVAL_59 = _EVAL_56;
  assign _EVAL_69 = _EVAL_188[78:76];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_98 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_123 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_132 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_175 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_7) begin
    if (_EVAL_24) begin
      _EVAL_98 <= 1'h0;
    end else begin
      if (_EVAL_182) begin
        _EVAL_98 <= _EVAL_168;
      end
    end
    if (_EVAL_24) begin
      _EVAL_123 <= 2'h3;
    end else begin
      if (_EVAL_202) begin
        _EVAL_123 <= _EVAL_141;
      end
    end
    if (_EVAL_24) begin
      _EVAL_132 <= 1'h0;
    end else begin
      if (_EVAL_182) begin
        _EVAL_132 <= _EVAL_136;
      end
    end
    if (_EVAL_24) begin
      _EVAL_175 <= 5'h0;
    end else begin
      if (_EVAL_162) begin
        _EVAL_175 <= _EVAL_164;
      end else begin
        _EVAL_175 <= _EVAL_116;
      end
    end
  end
endmodule
