//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_234(
  input  [31:0]  _EVAL,
  input  [31:0]  _EVAL_0,
  output         _EVAL_1,
  input  [127:0] _EVAL_2,
  input          _EVAL_3,
  input          _EVAL_4,
  input          _EVAL_5,
  input          _EVAL_6,
  input          _EVAL_7,
  input          _EVAL_8,
  input          _EVAL_9,
  input          _EVAL_10,
  input          _EVAL_11,
  input  [2:0]   _EVAL_12,
  input  [31:0]  _EVAL_13,
  output         _EVAL_14,
  input  [1:0]   _EVAL_15,
  input          _EVAL_16,
  output         _EVAL_17,
  input          _EVAL_18,
  input          _EVAL_19,
  input  [2:0]   _EVAL_20,
  input  [31:0]  _EVAL_21,
  output         _EVAL_22,
  input          _EVAL_23,
  input          _EVAL_24,
  output         _EVAL_25,
  output         _EVAL_26,
  input  [29:0]  _EVAL_27,
  input          _EVAL_28,
  input  [1:0]   _EVAL_29,
  input          _EVAL_30,
  output [2:0]   _EVAL_31,
  input  [2:0]   _EVAL_32,
  input          _EVAL_33,
  input          _EVAL_34,
  input          _EVAL_35,
  input          _EVAL_36,
  input          _EVAL_37,
  input          _EVAL_38,
  input          _EVAL_39,
  input          _EVAL_40,
  input          _EVAL_41,
  input  [29:0]  _EVAL_42,
  input  [63:0]  _EVAL_43,
  input          _EVAL_44,
  input          _EVAL_45,
  input          _EVAL_46,
  input          _EVAL_47,
  input          _EVAL_48,
  output [8:0]   _EVAL_49,
  input  [1:0]   _EVAL_50,
  input          _EVAL_51,
  input          _EVAL_52,
  output [63:0]  _EVAL_53,
  input          _EVAL_54,
  input  [31:0]  _EVAL_55,
  output         _EVAL_56,
  input          _EVAL_57,
  input          _EVAL_58,
  input          _EVAL_59,
  input  [1:0]   _EVAL_60,
  output [31:0]  _EVAL_61,
  output [127:0] _EVAL_62,
  input  [63:0]  _EVAL_63,
  input          _EVAL_64,
  input          _EVAL_65,
  output [31:0]  _EVAL_66,
  input          _EVAL_67,
  input  [29:0]  _EVAL_68,
  output [1:0]   _EVAL_69,
  input          _EVAL_70,
  input          _EVAL_71,
  output         _EVAL_72,
  input  [1:0]   _EVAL_73,
  input  [31:0]  _EVAL_74,
  output [1:0]   _EVAL_75,
  output [2:0]   _EVAL_76,
  input          _EVAL_77,
  input  [29:0]  _EVAL_78,
  output         _EVAL_79,
  input          _EVAL_80,
  input  [29:0]  _EVAL_81,
  input  [127:0] _EVAL_82,
  input          _EVAL_83,
  output         _EVAL_84,
  input  [7:0]   _EVAL_85,
  output [2:0]   _EVAL_86,
  input          _EVAL_87,
  input  [1:0]   _EVAL_88,
  input  [31:0]  _EVAL_89,
  input  [1:0]   _EVAL_90,
  output         _EVAL_91,
  input  [31:0]  _EVAL_92,
  input  [29:0]  _EVAL_93,
  input  [31:0]  _EVAL_94,
  input  [31:0]  _EVAL_95,
  output [14:0]  _EVAL_96,
  input  [2:0]   _EVAL_97,
  input  [29:0]  _EVAL_98,
  output         _EVAL_99,
  input          _EVAL_100,
  input  [29:0]  _EVAL_101,
  output [2:0]   _EVAL_102,
  input          _EVAL_103,
  input          _EVAL_104,
  input          _EVAL_105,
  output         _EVAL_106,
  output [11:0]  _EVAL_107,
  output         _EVAL_108,
  input          _EVAL_109,
  output         _EVAL_110,
  output         _EVAL_111,
  input          _EVAL_112,
  input          _EVAL_113,
  input  [1:0]   _EVAL_114,
  input  [1:0]   _EVAL_115,
  input  [1:0]   _EVAL_116,
  input          _EVAL_117,
  input  [14:0]  _EVAL_118,
  input          _EVAL_119,
  output [63:0]  _EVAL_120,
  input  [24:0]  _EVAL_121,
  input  [3:0]   _EVAL_122,
  input          _EVAL_123,
  output         _EVAL_124,
  output         _EVAL_125,
  output         _EVAL_126,
  output         _EVAL_127,
  input  [1:0]   _EVAL_128,
  input  [31:0]  _EVAL_129,
  input  [31:0]  _EVAL_130,
  input          _EVAL_131,
  input          _EVAL_132,
  output         _EVAL_133,
  input          _EVAL_134,
  output         _EVAL_135,
  input          _EVAL_136,
  input  [11:0]  _EVAL_137,
  input          _EVAL_138,
  input  [31:0]  _EVAL_139,
  input          _EVAL_140,
  input          _EVAL_141,
  input          _EVAL_142
);
  wire  packageanon1_3__EVAL;
  wire  packageanon1_3__EVAL_0;
  wire  packageanon1_5__EVAL;
  wire  packageanon1_5__EVAL_0;
  wire  data_arrays_3_0__EVAL;
  wire [63:0] data_arrays_3_0__EVAL_0;
  wire [7:0] data_arrays_3_0__EVAL_1;
  wire  data_arrays_3_0__EVAL_2;
  wire  data_arrays_3_0__EVAL_3;
  wire [63:0] data_arrays_3_0__EVAL_4;
  wire  data_arrays_2_1__EVAL;
  wire [63:0] data_arrays_2_1__EVAL_0;
  wire [7:0] data_arrays_2_1__EVAL_1;
  wire  data_arrays_2_1__EVAL_2;
  wire  data_arrays_2_1__EVAL_3;
  wire [63:0] data_arrays_2_1__EVAL_4;
  wire  data_arrays_1_0__EVAL;
  wire [63:0] data_arrays_1_0__EVAL_0;
  wire [7:0] data_arrays_1_0__EVAL_1;
  wire  data_arrays_1_0__EVAL_2;
  wire  data_arrays_1_0__EVAL_3;
  wire [63:0] data_arrays_1_0__EVAL_4;
  wire  data_arrays_2_0__EVAL;
  wire [63:0] data_arrays_2_0__EVAL_0;
  wire [7:0] data_arrays_2_0__EVAL_1;
  wire  data_arrays_2_0__EVAL_2;
  wire  data_arrays_2_0__EVAL_3;
  wire [63:0] data_arrays_2_0__EVAL_4;
  wire  packageanon1_7__EVAL;
  wire  packageanon1_7__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_1__EVAL;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_0;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_1;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_2;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_3;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_4;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_5;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_6;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_7;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_8;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_9;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_10;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_11;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_12;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_13;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_14;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_15;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_16;
  wire  MaxPeriodFibonacciLFSR_1__EVAL_17;
  wire  predictor_tagged_tables_2__EVAL;
  wire  predictor_tagged_tables_2__EVAL_0;
  wire  predictor_tagged_tables_2__EVAL_1;
  wire  predictor_tagged_tables_2__EVAL_2;
  wire  predictor_tagged_tables_2__EVAL_3;
  wire  predictor_tagged_tables_2__EVAL_4;
  wire  predictor_tagged_tables_2__EVAL_5;
  wire  predictor_tagged_tables_2__EVAL_6;
  wire  predictor_tagged_tables_2__EVAL_7;
  wire  predictor_tagged_tables_2__EVAL_8;
  wire  predictor_tagged_tables_2__EVAL_9;
  wire  predictor_tagged_tables_2__EVAL_10;
  wire  predictor_tagged_tables_2__EVAL_11;
  wire  predictor_tagged_tables_2__EVAL_12;
  wire  predictor_tagged_tables_2__EVAL_13;
  wire  predictor_tagged_tables_2__EVAL_14;
  wire [8:0] predictor_tagged_tables_2__EVAL_15;
  wire  predictor_tagged_tables_2__EVAL_16;
  wire  predictor_tagged_tables_2__EVAL_17;
  wire  predictor_tagged_tables_2__EVAL_18;
  wire  predictor_tagged_tables_2__EVAL_19;
  wire  predictor_tagged_tables_2__EVAL_20;
  wire  predictor_tagged_tables_2__EVAL_21;
  wire  predictor_tagged_tables_2__EVAL_22;
  wire  predictor_tagged_tables_2__EVAL_23;
  wire  predictor_tagged_tables_2__EVAL_24;
  wire  predictor_tagged_tables_2__EVAL_25;
  wire  predictor_tagged_tables_2__EVAL_26;
  wire  predictor_tagged_tables_2__EVAL_27;
  wire  predictor_tagged_tables_2__EVAL_28;
  wire  predictor_tagged_tables_2__EVAL_29;
  wire  predictor_tagged_tables_2__EVAL_30;
  wire  predictor_tagged_tables_2__EVAL_31;
  wire  predictor_tagged_tables_2__EVAL_32;
  wire  predictor_tagged_tables_2__EVAL_33;
  wire  predictor_tagged_tables_2__EVAL_34;
  wire  predictor_tagged_tables_2__EVAL_35;
  wire  predictor_tagged_tables_2__EVAL_36;
  wire  predictor_tagged_tables_2__EVAL_37;
  wire  predictor_tagged_tables_2__EVAL_38;
  wire  predictor_tagged_tables_1__EVAL;
  wire  predictor_tagged_tables_1__EVAL_0;
  wire  predictor_tagged_tables_1__EVAL_1;
  wire  predictor_tagged_tables_1__EVAL_2;
  wire  predictor_tagged_tables_1__EVAL_3;
  wire  predictor_tagged_tables_1__EVAL_4;
  wire  predictor_tagged_tables_1__EVAL_5;
  wire  predictor_tagged_tables_1__EVAL_6;
  wire  predictor_tagged_tables_1__EVAL_7;
  wire  predictor_tagged_tables_1__EVAL_8;
  wire  predictor_tagged_tables_1__EVAL_9;
  wire  predictor_tagged_tables_1__EVAL_10;
  wire  predictor_tagged_tables_1__EVAL_11;
  wire  predictor_tagged_tables_1__EVAL_12;
  wire  predictor_tagged_tables_1__EVAL_13;
  wire  predictor_tagged_tables_1__EVAL_14;
  wire [8:0] predictor_tagged_tables_1__EVAL_15;
  wire  predictor_tagged_tables_1__EVAL_16;
  wire  predictor_tagged_tables_1__EVAL_17;
  wire  predictor_tagged_tables_1__EVAL_18;
  wire  predictor_tagged_tables_1__EVAL_19;
  wire  predictor_tagged_tables_1__EVAL_20;
  wire  predictor_tagged_tables_1__EVAL_21;
  wire  predictor_tagged_tables_1__EVAL_22;
  wire  predictor_tagged_tables_1__EVAL_23;
  wire  predictor_tagged_tables_1__EVAL_24;
  wire  predictor_tagged_tables_1__EVAL_25;
  wire  predictor_tagged_tables_1__EVAL_26;
  wire  predictor_tagged_tables_1__EVAL_27;
  wire  predictor_tagged_tables_1__EVAL_28;
  wire  predictor_tagged_tables_1__EVAL_29;
  wire  predictor_tagged_tables_1__EVAL_30;
  wire  predictor_tagged_tables_1__EVAL_31;
  wire  predictor_tagged_tables_1__EVAL_32;
  wire  predictor_tagged_tables_1__EVAL_33;
  wire  predictor_tagged_tables_1__EVAL_34;
  wire  predictor_tagged_tables_1__EVAL_35;
  wire  predictor_tagged_tables_1__EVAL_36;
  wire  predictor_tagged_tables_1__EVAL_37;
  wire  predictor_tagged_tables_1__EVAL_38;
  wire  icache_clock_gate_in;
  wire  icache_clock_gate_en;
  wire  icache_clock_gate_out;
  wire  data_arrays_1_1__EVAL;
  wire [63:0] data_arrays_1_1__EVAL_0;
  wire [7:0] data_arrays_1_1__EVAL_1;
  wire  data_arrays_1_1__EVAL_2;
  wire  data_arrays_1_1__EVAL_3;
  wire [63:0] data_arrays_1_1__EVAL_4;
  wire  packageanon1_1__EVAL;
  wire  packageanon1_1__EVAL_0;
  wire  packageanon1_2__EVAL;
  wire  packageanon1_2__EVAL_0;
  wire  predictor_tagged_tables_0__EVAL;
  wire  predictor_tagged_tables_0__EVAL_0;
  wire  predictor_tagged_tables_0__EVAL_1;
  wire  predictor_tagged_tables_0__EVAL_2;
  wire  predictor_tagged_tables_0__EVAL_3;
  wire  predictor_tagged_tables_0__EVAL_4;
  wire  predictor_tagged_tables_0__EVAL_5;
  wire  predictor_tagged_tables_0__EVAL_6;
  wire  predictor_tagged_tables_0__EVAL_7;
  wire  predictor_tagged_tables_0__EVAL_8;
  wire  predictor_tagged_tables_0__EVAL_9;
  wire  predictor_tagged_tables_0__EVAL_10;
  wire  predictor_tagged_tables_0__EVAL_11;
  wire  predictor_tagged_tables_0__EVAL_12;
  wire  predictor_tagged_tables_0__EVAL_13;
  wire  predictor_tagged_tables_0__EVAL_14;
  wire [8:0] predictor_tagged_tables_0__EVAL_15;
  wire  predictor_tagged_tables_0__EVAL_16;
  wire  predictor_tagged_tables_0__EVAL_17;
  wire  predictor_tagged_tables_0__EVAL_18;
  wire  predictor_tagged_tables_0__EVAL_19;
  wire  predictor_tagged_tables_0__EVAL_20;
  wire  predictor_tagged_tables_0__EVAL_21;
  wire  predictor_tagged_tables_0__EVAL_22;
  wire  predictor_tagged_tables_0__EVAL_23;
  wire  predictor_tagged_tables_0__EVAL_24;
  wire  predictor_tagged_tables_0__EVAL_25;
  wire  predictor_tagged_tables_0__EVAL_26;
  wire  predictor_tagged_tables_0__EVAL_27;
  wire  predictor_tagged_tables_0__EVAL_28;
  wire  predictor_tagged_tables_0__EVAL_29;
  wire  predictor_tagged_tables_0__EVAL_30;
  wire  predictor_tagged_tables_0__EVAL_31;
  wire  predictor_tagged_tables_0__EVAL_32;
  wire  predictor_tagged_tables_0__EVAL_33;
  wire  predictor_tagged_tables_0__EVAL_34;
  wire  predictor_tagged_tables_0__EVAL_35;
  wire  predictor_tagged_tables_0__EVAL_36;
  wire  predictor_tagged_tables_0__EVAL_37;
  wire  predictor_tagged_tables_0__EVAL_38;
  wire [31:0] predictor_Queue__EVAL;
  wire [31:0] predictor_Queue__EVAL_0;
  wire  predictor_Queue__EVAL_1;
  wire  predictor_Queue__EVAL_2;
  wire  predictor_Queue__EVAL_3;
  wire  predictor_Queue__EVAL_4;
  wire  predictor_Queue__EVAL_5;
  wire [127:0] predictor_Queue__EVAL_6;
  wire  predictor_Queue__EVAL_7;
  wire  predictor_Queue__EVAL_8;
  wire  predictor_Queue__EVAL_9;
  wire  predictor_Queue__EVAL_10;
  wire  predictor_Queue__EVAL_11;
  wire [127:0] predictor_Queue__EVAL_12;
  wire  predictor_Queue__EVAL_13;
  wire  predictor_Queue__EVAL_14;
  wire  packageanon1_8__EVAL;
  wire  packageanon1_8__EVAL_0;
  wire  data_arrays_3_1__EVAL;
  wire [63:0] data_arrays_3_1__EVAL_0;
  wire [7:0] data_arrays_3_1__EVAL_1;
  wire  data_arrays_3_1__EVAL_2;
  wire  data_arrays_3_1__EVAL_3;
  wire [63:0] data_arrays_3_1__EVAL_4;
  wire [5:0] tag_array__EVAL;
  wire [20:0] tag_array__EVAL_0;
  wire [20:0] tag_array__EVAL_1;
  wire [20:0] tag_array__EVAL_2;
  wire [20:0] tag_array__EVAL_3;
  wire  tag_array__EVAL_4;
  wire  tag_array__EVAL_5;
  wire  tag_array__EVAL_6;
  wire [20:0] tag_array__EVAL_7;
  wire  tag_array__EVAL_8;
  wire  tag_array__EVAL_9;
  wire  tag_array__EVAL_10;
  wire [20:0] tag_array__EVAL_11;
  wire [20:0] tag_array__EVAL_12;
  wire  tag_array__EVAL_13;
  wire [20:0] tag_array__EVAL_14;
  wire  packageanon1_6__EVAL;
  wire  packageanon1_6__EVAL_0;
  wire  data_arrays_0_1__EVAL;
  wire [63:0] data_arrays_0_1__EVAL_0;
  wire [7:0] data_arrays_0_1__EVAL_1;
  wire  data_arrays_0_1__EVAL_2;
  wire  data_arrays_0_1__EVAL_3;
  wire [63:0] data_arrays_0_1__EVAL_4;
  wire  predictor_base_table_1__EVAL;
  wire  predictor_base_table_1__EVAL_0;
  wire  predictor_base_table_1__EVAL_1;
  wire  predictor_base_table_1__EVAL_2;
  wire  predictor_base_table_1__EVAL_3;
  wire  predictor_base_table_1__EVAL_4;
  wire  predictor_base_table_1__EVAL_5;
  wire  predictor_base_table_1__EVAL_6;
  wire  predictor_base_table_1__EVAL_7;
  wire [7:0] predictor_base_table_1__EVAL_8;
  wire  predictor_base_table_1__EVAL_9;
  wire  predictor_base_table_1__EVAL_10;
  wire  predictor_base_table_1__EVAL_11;
  wire  predictor_base_table_1__EVAL_12;
  wire  predictor_base_table_1__EVAL_13;
  wire  predictor_base_table_1__EVAL_14;
  wire  predictor_base_table_1__EVAL_15;
  wire  predictor_base_table_1__EVAL_16;
  wire  predictor_base_table_1__EVAL_17;
  wire  predictor_base_table_1__EVAL_18;
  wire  predictor_base_table_1__EVAL_19;
  wire  predictor_base_table_1__EVAL_20;
  wire  predictor_base_table_1__EVAL_21;
  wire  predictor_base_table_1__EVAL_22;
  wire  predictor_base_table_1__EVAL_23;
  wire  predictor_base_table_1__EVAL_24;
  wire  predictor_base_table_1__EVAL_25;
  wire  predictor_base_table_1__EVAL_26;
  wire  predictor_base_table_1__EVAL_27;
  wire  predictor_base_table_1__EVAL_28;
  wire  predictor_base_table_1__EVAL_29;
  wire  MaxPeriodFibonacciLFSR__EVAL;
  wire  MaxPeriodFibonacciLFSR__EVAL_0;
  wire  MaxPeriodFibonacciLFSR__EVAL_1;
  wire  MaxPeriodFibonacciLFSR__EVAL_2;
  wire  MaxPeriodFibonacciLFSR__EVAL_3;
  wire  MaxPeriodFibonacciLFSR__EVAL_4;
  wire  MaxPeriodFibonacciLFSR__EVAL_5;
  wire  MaxPeriodFibonacciLFSR__EVAL_6;
  wire  MaxPeriodFibonacciLFSR__EVAL_7;
  wire  MaxPeriodFibonacciLFSR__EVAL_8;
  wire  MaxPeriodFibonacciLFSR__EVAL_9;
  wire  MaxPeriodFibonacciLFSR__EVAL_10;
  wire  MaxPeriodFibonacciLFSR__EVAL_11;
  wire  MaxPeriodFibonacciLFSR__EVAL_12;
  wire  MaxPeriodFibonacciLFSR__EVAL_13;
  wire  MaxPeriodFibonacciLFSR__EVAL_14;
  wire  MaxPeriodFibonacciLFSR__EVAL_15;
  wire  MaxPeriodFibonacciLFSR__EVAL_16;
  wire  MaxPeriodFibonacciLFSR__EVAL_17;
  wire  predictor_tagged_tables_3__EVAL;
  wire  predictor_tagged_tables_3__EVAL_0;
  wire  predictor_tagged_tables_3__EVAL_1;
  wire  predictor_tagged_tables_3__EVAL_2;
  wire  predictor_tagged_tables_3__EVAL_3;
  wire  predictor_tagged_tables_3__EVAL_4;
  wire  predictor_tagged_tables_3__EVAL_5;
  wire  predictor_tagged_tables_3__EVAL_6;
  wire  predictor_tagged_tables_3__EVAL_7;
  wire  predictor_tagged_tables_3__EVAL_8;
  wire  predictor_tagged_tables_3__EVAL_9;
  wire  predictor_tagged_tables_3__EVAL_10;
  wire  predictor_tagged_tables_3__EVAL_11;
  wire  predictor_tagged_tables_3__EVAL_12;
  wire  predictor_tagged_tables_3__EVAL_13;
  wire  predictor_tagged_tables_3__EVAL_14;
  wire [8:0] predictor_tagged_tables_3__EVAL_15;
  wire  predictor_tagged_tables_3__EVAL_16;
  wire  predictor_tagged_tables_3__EVAL_17;
  wire  predictor_tagged_tables_3__EVAL_18;
  wire  predictor_tagged_tables_3__EVAL_19;
  wire  predictor_tagged_tables_3__EVAL_20;
  wire  predictor_tagged_tables_3__EVAL_21;
  wire  predictor_tagged_tables_3__EVAL_22;
  wire  predictor_tagged_tables_3__EVAL_23;
  wire  predictor_tagged_tables_3__EVAL_24;
  wire  predictor_tagged_tables_3__EVAL_25;
  wire  predictor_tagged_tables_3__EVAL_26;
  wire  predictor_tagged_tables_3__EVAL_27;
  wire  predictor_tagged_tables_3__EVAL_28;
  wire  predictor_tagged_tables_3__EVAL_29;
  wire  predictor_tagged_tables_3__EVAL_30;
  wire  predictor_tagged_tables_3__EVAL_31;
  wire  predictor_tagged_tables_3__EVAL_32;
  wire  predictor_tagged_tables_3__EVAL_33;
  wire  predictor_tagged_tables_3__EVAL_34;
  wire  predictor_tagged_tables_3__EVAL_35;
  wire  predictor_tagged_tables_3__EVAL_36;
  wire  predictor_tagged_tables_3__EVAL_37;
  wire  predictor_tagged_tables_3__EVAL_38;
  wire  data_arrays_0_0__EVAL;
  wire [63:0] data_arrays_0_0__EVAL_0;
  wire [7:0] data_arrays_0_0__EVAL_1;
  wire  data_arrays_0_0__EVAL_2;
  wire  data_arrays_0_0__EVAL_3;
  wire [63:0] data_arrays_0_0__EVAL_4;
  wire  predictor_base_table_0__EVAL;
  wire  predictor_base_table_0__EVAL_0;
  wire  predictor_base_table_0__EVAL_1;
  wire  predictor_base_table_0__EVAL_2;
  wire  predictor_base_table_0__EVAL_3;
  wire  predictor_base_table_0__EVAL_4;
  wire  predictor_base_table_0__EVAL_5;
  wire  predictor_base_table_0__EVAL_6;
  wire  predictor_base_table_0__EVAL_7;
  wire [7:0] predictor_base_table_0__EVAL_8;
  wire  predictor_base_table_0__EVAL_9;
  wire  predictor_base_table_0__EVAL_10;
  wire  predictor_base_table_0__EVAL_11;
  wire  predictor_base_table_0__EVAL_12;
  wire  predictor_base_table_0__EVAL_13;
  wire  predictor_base_table_0__EVAL_14;
  wire  predictor_base_table_0__EVAL_15;
  wire  predictor_base_table_0__EVAL_16;
  wire  predictor_base_table_0__EVAL_17;
  wire  predictor_base_table_0__EVAL_18;
  wire  predictor_base_table_0__EVAL_19;
  wire  predictor_base_table_0__EVAL_20;
  wire  predictor_base_table_0__EVAL_21;
  wire  predictor_base_table_0__EVAL_22;
  wire  predictor_base_table_0__EVAL_23;
  wire  predictor_base_table_0__EVAL_24;
  wire  predictor_base_table_0__EVAL_25;
  wire  predictor_base_table_0__EVAL_26;
  wire  predictor_base_table_0__EVAL_27;
  wire  predictor_base_table_0__EVAL_28;
  wire  predictor_base_table_0__EVAL_29;
  wire  packageanon1_4__EVAL;
  wire  packageanon1_4__EVAL_0;
  wire [1:0] tlb__EVAL;
  wire  tlb__EVAL_0;
  wire [29:0] tlb__EVAL_1;
  wire  tlb__EVAL_2;
  wire  tlb__EVAL_3;
  wire  tlb__EVAL_4;
  wire [1:0] tlb__EVAL_5;
  wire  tlb__EVAL_6;
  wire [1:0] tlb__EVAL_7;
  wire [31:0] tlb__EVAL_8;
  wire [29:0] tlb__EVAL_9;
  wire  tlb__EVAL_10;
  wire  tlb__EVAL_11;
  wire  tlb__EVAL_12;
  wire  tlb__EVAL_13;
  wire  tlb__EVAL_14;
  wire [1:0] tlb__EVAL_15;
  wire [1:0] tlb__EVAL_16;
  wire [31:0] tlb__EVAL_17;
  wire [31:0] tlb__EVAL_18;
  wire  tlb__EVAL_19;
  wire  tlb__EVAL_20;
  wire [29:0] tlb__EVAL_21;
  wire  tlb__EVAL_22;
  wire [29:0] tlb__EVAL_23;
  wire  tlb__EVAL_24;
  wire [1:0] tlb__EVAL_25;
  wire  tlb__EVAL_26;
  wire [29:0] tlb__EVAL_27;
  wire  tlb__EVAL_28;
  wire  tlb__EVAL_29;
  wire  tlb__EVAL_30;
  wire  tlb__EVAL_31;
  wire  tlb__EVAL_32;
  wire  tlb__EVAL_33;
  wire [31:0] tlb__EVAL_34;
  wire  tlb__EVAL_35;
  wire  tlb__EVAL_36;
  wire [31:0] tlb__EVAL_37;
  wire  tlb__EVAL_38;
  wire  tlb__EVAL_39;
  wire [1:0] tlb__EVAL_40;
  wire [29:0] tlb__EVAL_41;
  wire  tlb__EVAL_42;
  wire [29:0] tlb__EVAL_43;
  wire [31:0] tlb__EVAL_44;
  wire  tlb__EVAL_45;
  wire [1:0] tlb__EVAL_46;
  wire [31:0] tlb__EVAL_47;
  wire [31:0] tlb__EVAL_48;
  wire [1:0] tlb__EVAL_49;
  wire [29:0] tlb__EVAL_50;
  wire  tlb__EVAL_51;
  wire  tlb__EVAL_52;
  wire  tlb__EVAL_53;
  wire  tlb__EVAL_54;
  wire  tlb__EVAL_55;
  wire  tlb__EVAL_56;
  wire [31:0] tlb__EVAL_57;
  wire  tlb__EVAL_58;
  wire [31:0] tlb__EVAL_59;
  wire  tlb__EVAL_60;
  wire  tlb__EVAL_61;
  wire  tlb__EVAL_62;
  wire  itim_array__EVAL;
  wire  itim_array__EVAL_0;
  wire [11:0] itim_array__EVAL_1;
  wire [63:0] itim_array__EVAL_2;
  wire  itim_array__EVAL_3;
  wire [63:0] itim_array__EVAL_4;
  wire [31:0] packageanon1__EVAL;
  wire [31:0] packageanon1__EVAL_0;
  reg  _EVAL_215 [0:3];
  reg [31:0] _RAND_0;
  wire  _EVAL_215__EVAL_216_data;
  wire [1:0] _EVAL_215__EVAL_216_addr;
  wire  _EVAL_215__EVAL_217_data;
  wire [1:0] _EVAL_215__EVAL_217_addr;
  wire  _EVAL_215__EVAL_217_mask;
  wire  _EVAL_215__EVAL_217_en;
  reg  _EVAL_319 [0:0];
  reg [31:0] _RAND_1;
  wire  _EVAL_319__EVAL_320_data;
  wire  _EVAL_319__EVAL_320_addr;
  wire  _EVAL_319__EVAL_321_data;
  wire  _EVAL_319__EVAL_321_addr;
  wire  _EVAL_319__EVAL_321_mask;
  wire  _EVAL_319__EVAL_321_en;
  reg  _EVAL_363 [0:3];
  reg [31:0] _RAND_2;
  wire  _EVAL_363__EVAL_364_data;
  wire [1:0] _EVAL_363__EVAL_364_addr;
  wire  _EVAL_363__EVAL_365_data;
  wire [1:0] _EVAL_363__EVAL_365_addr;
  wire  _EVAL_363__EVAL_365_mask;
  wire  _EVAL_363__EVAL_365_en;
  reg [2:0] _EVAL_386 [0:3];
  reg [31:0] _RAND_3;
  wire [2:0] _EVAL_386__EVAL_387_data;
  wire [1:0] _EVAL_386__EVAL_387_addr;
  wire [2:0] _EVAL_386__EVAL_388_data;
  wire [1:0] _EVAL_386__EVAL_388_addr;
  wire  _EVAL_386__EVAL_388_mask;
  wire  _EVAL_386__EVAL_388_en;
  reg  _EVAL_394 [0:0];
  reg [31:0] _RAND_4;
  wire  _EVAL_394__EVAL_395_data;
  wire  _EVAL_394__EVAL_395_addr;
  wire  _EVAL_394__EVAL_396_data;
  wire  _EVAL_394__EVAL_396_addr;
  wire  _EVAL_394__EVAL_396_mask;
  wire  _EVAL_394__EVAL_396_en;
  reg  _EVAL_403 [0:0];
  reg [31:0] _RAND_5;
  wire  _EVAL_403__EVAL_404_data;
  wire  _EVAL_403__EVAL_404_addr;
  wire  _EVAL_403__EVAL_405_data;
  wire  _EVAL_403__EVAL_405_addr;
  wire  _EVAL_403__EVAL_405_mask;
  wire  _EVAL_403__EVAL_405_en;
  reg [127:0] _EVAL_489 [0:3];
  reg [127:0] _RAND_6;
  wire [127:0] _EVAL_489__EVAL_490_data;
  wire [1:0] _EVAL_489__EVAL_490_addr;
  wire [127:0] _EVAL_489__EVAL_491_data;
  wire [1:0] _EVAL_489__EVAL_491_addr;
  wire  _EVAL_489__EVAL_491_mask;
  wire  _EVAL_489__EVAL_491_en;
  reg [2:0] _EVAL_530 [0:0];
  reg [31:0] _RAND_7;
  wire [2:0] _EVAL_530__EVAL_531_data;
  wire  _EVAL_530__EVAL_531_addr;
  wire [2:0] _EVAL_530__EVAL_532_data;
  wire  _EVAL_530__EVAL_532_addr;
  wire  _EVAL_530__EVAL_532_mask;
  wire  _EVAL_530__EVAL_532_en;
  reg  _EVAL_548 [0:3];
  reg [31:0] _RAND_8;
  wire  _EVAL_548__EVAL_549_data;
  wire [1:0] _EVAL_548__EVAL_549_addr;
  wire  _EVAL_548__EVAL_550_data;
  wire [1:0] _EVAL_548__EVAL_550_addr;
  wire  _EVAL_548__EVAL_550_mask;
  wire  _EVAL_548__EVAL_550_en;
  reg  _EVAL_658 [0:0];
  reg [31:0] _RAND_9;
  wire  _EVAL_658__EVAL_659_data;
  wire  _EVAL_658__EVAL_659_addr;
  wire  _EVAL_658__EVAL_660_data;
  wire  _EVAL_658__EVAL_660_addr;
  wire  _EVAL_658__EVAL_660_mask;
  wire  _EVAL_658__EVAL_660_en;
  reg [63:0] _EVAL_719 [0:3];
  reg [63:0] _RAND_10;
  wire [63:0] _EVAL_719__EVAL_720_data;
  wire [1:0] _EVAL_719__EVAL_720_addr;
  wire [63:0] _EVAL_719__EVAL_721_data;
  wire [1:0] _EVAL_719__EVAL_721_addr;
  wire  _EVAL_719__EVAL_721_mask;
  wire  _EVAL_719__EVAL_721_en;
  reg  _EVAL_725 [0:0];
  reg [31:0] _RAND_11;
  wire  _EVAL_725__EVAL_726_data;
  wire  _EVAL_725__EVAL_726_addr;
  wire  _EVAL_725__EVAL_727_data;
  wire  _EVAL_725__EVAL_727_addr;
  wire  _EVAL_725__EVAL_727_mask;
  wire  _EVAL_725__EVAL_727_en;
  reg  _EVAL_744 [0:3];
  reg [31:0] _RAND_12;
  wire  _EVAL_744__EVAL_745_data;
  wire [1:0] _EVAL_744__EVAL_745_addr;
  wire  _EVAL_744__EVAL_746_data;
  wire [1:0] _EVAL_744__EVAL_746_addr;
  wire  _EVAL_744__EVAL_746_mask;
  wire  _EVAL_744__EVAL_746_en;
  reg  _EVAL_931 [0:3];
  reg [31:0] _RAND_13;
  wire  _EVAL_931__EVAL_932_data;
  wire [1:0] _EVAL_931__EVAL_932_addr;
  wire  _EVAL_931__EVAL_933_data;
  wire [1:0] _EVAL_931__EVAL_933_addr;
  wire  _EVAL_931__EVAL_933_mask;
  wire  _EVAL_931__EVAL_933_en;
  reg  _EVAL_949 [0:0];
  reg [31:0] _RAND_14;
  wire  _EVAL_949__EVAL_950_data;
  wire  _EVAL_949__EVAL_950_addr;
  wire  _EVAL_949__EVAL_951_data;
  wire  _EVAL_949__EVAL_951_addr;
  wire  _EVAL_949__EVAL_951_mask;
  wire  _EVAL_949__EVAL_951_en;
  reg [8:0] _EVAL_961 [0:3];
  reg [31:0] _RAND_15;
  wire [8:0] _EVAL_961__EVAL_962_data;
  wire [1:0] _EVAL_961__EVAL_962_addr;
  wire [8:0] _EVAL_961__EVAL_963_data;
  wire [1:0] _EVAL_961__EVAL_963_addr;
  wire  _EVAL_961__EVAL_963_mask;
  wire  _EVAL_961__EVAL_963_en;
  reg [2:0] _EVAL_982 [0:0];
  reg [31:0] _RAND_16;
  wire [2:0] _EVAL_982__EVAL_983_data;
  wire  _EVAL_982__EVAL_983_addr;
  wire [2:0] _EVAL_982__EVAL_984_data;
  wire  _EVAL_982__EVAL_984_addr;
  wire  _EVAL_982__EVAL_984_mask;
  wire  _EVAL_982__EVAL_984_en;
  reg  _EVAL_1119 [0:0];
  reg [31:0] _RAND_17;
  wire  _EVAL_1119__EVAL_1120_data;
  wire  _EVAL_1119__EVAL_1120_addr;
  wire  _EVAL_1119__EVAL_1121_data;
  wire  _EVAL_1119__EVAL_1121_addr;
  wire  _EVAL_1119__EVAL_1121_mask;
  wire  _EVAL_1119__EVAL_1121_en;
  reg  _EVAL_1140 [0:3];
  reg [31:0] _RAND_18;
  wire  _EVAL_1140__EVAL_1141_data;
  wire [1:0] _EVAL_1140__EVAL_1141_addr;
  wire  _EVAL_1140__EVAL_1142_data;
  wire [1:0] _EVAL_1140__EVAL_1142_addr;
  wire  _EVAL_1140__EVAL_1142_mask;
  wire  _EVAL_1140__EVAL_1142_en;
  reg [8:0] _EVAL_1147 [0:0];
  reg [31:0] _RAND_19;
  wire [8:0] _EVAL_1147__EVAL_1148_data;
  wire  _EVAL_1147__EVAL_1148_addr;
  wire [8:0] _EVAL_1147__EVAL_1149_data;
  wire  _EVAL_1147__EVAL_1149_addr;
  wire  _EVAL_1147__EVAL_1149_mask;
  wire  _EVAL_1147__EVAL_1149_en;
  reg  _EVAL_1440 [0:3];
  reg [31:0] _RAND_20;
  wire  _EVAL_1440__EVAL_1441_data;
  wire [1:0] _EVAL_1440__EVAL_1441_addr;
  wire  _EVAL_1440__EVAL_1442_data;
  wire [1:0] _EVAL_1440__EVAL_1442_addr;
  wire  _EVAL_1440__EVAL_1442_mask;
  wire  _EVAL_1440__EVAL_1442_en;
  reg [127:0] _EVAL_1465 [0:0];
  reg [127:0] _RAND_21;
  wire [127:0] _EVAL_1465__EVAL_1466_data;
  wire  _EVAL_1465__EVAL_1466_addr;
  wire [127:0] _EVAL_1465__EVAL_1467_data;
  wire  _EVAL_1465__EVAL_1467_addr;
  wire  _EVAL_1465__EVAL_1467_mask;
  wire  _EVAL_1465__EVAL_1467_en;
  reg [2:0] _EVAL_1481 [0:0];
  reg [31:0] _RAND_22;
  wire [2:0] _EVAL_1481__EVAL_1482_data;
  wire  _EVAL_1481__EVAL_1482_addr;
  wire [2:0] _EVAL_1481__EVAL_1483_data;
  wire  _EVAL_1481__EVAL_1483_addr;
  wire  _EVAL_1481__EVAL_1483_mask;
  wire  _EVAL_1481__EVAL_1483_en;
  reg [31:0] _EVAL_1518 [0:3];
  reg [31:0] _RAND_23;
  wire [31:0] _EVAL_1518__EVAL_1519_data;
  wire [1:0] _EVAL_1518__EVAL_1519_addr;
  wire [31:0] _EVAL_1518__EVAL_1520_data;
  wire [1:0] _EVAL_1518__EVAL_1520_addr;
  wire  _EVAL_1518__EVAL_1520_mask;
  wire  _EVAL_1518__EVAL_1520_en;
  reg  _EVAL_1652 [0:0];
  reg [31:0] _RAND_24;
  wire  _EVAL_1652__EVAL_1653_data;
  wire  _EVAL_1652__EVAL_1653_addr;
  wire  _EVAL_1652__EVAL_1654_data;
  wire  _EVAL_1652__EVAL_1654_addr;
  wire  _EVAL_1652__EVAL_1654_mask;
  wire  _EVAL_1652__EVAL_1654_en;
  reg  _EVAL_1716 [0:0];
  reg [31:0] _RAND_25;
  wire  _EVAL_1716__EVAL_1717_data;
  wire  _EVAL_1716__EVAL_1717_addr;
  wire  _EVAL_1716__EVAL_1718_data;
  wire  _EVAL_1716__EVAL_1718_addr;
  wire  _EVAL_1716__EVAL_1718_mask;
  wire  _EVAL_1716__EVAL_1718_en;
  reg [31:0] _EVAL_1767 [0:5];
  reg [31:0] _RAND_26;
  wire [31:0] _EVAL_1767__EVAL_1768_data;
  wire [2:0] _EVAL_1767__EVAL_1768_addr;
  reg [31:0] _RAND_27;
  wire [31:0] _EVAL_1767__EVAL_1769_data;
  wire [2:0] _EVAL_1767__EVAL_1769_addr;
  wire  _EVAL_1767__EVAL_1769_mask;
  wire  _EVAL_1767__EVAL_1769_en;
  reg [39:0] _EVAL_1859 [0:7];
  reg [63:0] _RAND_28;
  wire [39:0] _EVAL_1859__EVAL_1860_data;
  wire [2:0] _EVAL_1859__EVAL_1860_addr;
  wire [39:0] _EVAL_1859__EVAL_1861_data;
  wire [2:0] _EVAL_1859__EVAL_1861_addr;
  wire [39:0] _EVAL_1859__EVAL_1862_data;
  wire [2:0] _EVAL_1859__EVAL_1862_addr;
  wire  _EVAL_1859__EVAL_1862_mask;
  wire  _EVAL_1859__EVAL_1862_en;
  reg  _EVAL_1895 [0:0];
  reg [31:0] _RAND_29;
  wire  _EVAL_1895__EVAL_1896_data;
  wire  _EVAL_1895__EVAL_1896_addr;
  wire  _EVAL_1895__EVAL_1897_data;
  wire  _EVAL_1895__EVAL_1897_addr;
  wire  _EVAL_1895__EVAL_1897_mask;
  wire  _EVAL_1895__EVAL_1897_en;
  reg  _EVAL_1986 [0:3];
  reg [31:0] _RAND_30;
  wire  _EVAL_1986__EVAL_1987_data;
  wire [1:0] _EVAL_1986__EVAL_1987_addr;
  wire  _EVAL_1986__EVAL_1988_data;
  wire [1:0] _EVAL_1986__EVAL_1988_addr;
  wire  _EVAL_1986__EVAL_1988_mask;
  wire  _EVAL_1986__EVAL_1988_en;
  reg  _EVAL_2023 [0:0];
  reg [31:0] _RAND_31;
  wire  _EVAL_2023__EVAL_2024_data;
  wire  _EVAL_2023__EVAL_2024_addr;
  wire  _EVAL_2023__EVAL_2025_data;
  wire  _EVAL_2023__EVAL_2025_addr;
  wire  _EVAL_2023__EVAL_2025_mask;
  wire  _EVAL_2023__EVAL_2025_en;
  reg [1:0] _EVAL_2073 [0:3];
  reg [31:0] _RAND_32;
  wire [1:0] _EVAL_2073__EVAL_2074_data;
  wire [1:0] _EVAL_2073__EVAL_2074_addr;
  wire [1:0] _EVAL_2073__EVAL_2075_data;
  wire [1:0] _EVAL_2073__EVAL_2075_addr;
  wire  _EVAL_2073__EVAL_2075_mask;
  wire  _EVAL_2073__EVAL_2075_en;
  reg  _EVAL_2081 [0:3];
  reg [31:0] _RAND_33;
  wire  _EVAL_2081__EVAL_2082_data;
  wire [1:0] _EVAL_2081__EVAL_2082_addr;
  wire  _EVAL_2081__EVAL_2083_data;
  wire [1:0] _EVAL_2081__EVAL_2083_addr;
  wire  _EVAL_2081__EVAL_2083_mask;
  wire  _EVAL_2081__EVAL_2083_en;
  reg  _EVAL_2177 [0:3];
  reg [31:0] _RAND_34;
  wire  _EVAL_2177__EVAL_2178_data;
  wire [1:0] _EVAL_2177__EVAL_2178_addr;
  wire  _EVAL_2177__EVAL_2179_data;
  wire [1:0] _EVAL_2177__EVAL_2179_addr;
  wire  _EVAL_2177__EVAL_2179_mask;
  wire  _EVAL_2177__EVAL_2179_en;
  reg [63:0] _EVAL_2229 [0:0];
  reg [63:0] _RAND_35;
  wire [63:0] _EVAL_2229__EVAL_2230_data;
  wire  _EVAL_2229__EVAL_2230_addr;
  wire [63:0] _EVAL_2229__EVAL_2231_data;
  wire  _EVAL_2229__EVAL_2231_addr;
  wire  _EVAL_2229__EVAL_2231_mask;
  wire  _EVAL_2229__EVAL_2231_en;
  reg [31:0] _EVAL_2337 [0:0];
  reg [31:0] _RAND_36;
  wire [31:0] _EVAL_2337__EVAL_2338_data;
  wire  _EVAL_2337__EVAL_2338_addr;
  wire [31:0] _EVAL_2337__EVAL_2339_data;
  wire  _EVAL_2337__EVAL_2339_addr;
  wire  _EVAL_2337__EVAL_2339_mask;
  wire  _EVAL_2337__EVAL_2339_en;
  reg [14:0] _EVAL_2478 [0:0];
  reg [31:0] _RAND_37;
  wire [14:0] _EVAL_2478__EVAL_2479_data;
  wire  _EVAL_2478__EVAL_2479_addr;
  wire [14:0] _EVAL_2478__EVAL_2480_data;
  wire  _EVAL_2478__EVAL_2480_addr;
  wire  _EVAL_2478__EVAL_2480_mask;
  wire  _EVAL_2478__EVAL_2480_en;
  reg  _EVAL_2542 [0:0];
  reg [31:0] _RAND_38;
  wire  _EVAL_2542__EVAL_2543_data;
  wire  _EVAL_2542__EVAL_2543_addr;
  wire  _EVAL_2542__EVAL_2544_data;
  wire  _EVAL_2542__EVAL_2544_addr;
  wire  _EVAL_2542__EVAL_2544_mask;
  wire  _EVAL_2542__EVAL_2544_en;
  reg [14:0] _EVAL_2573 [0:3];
  reg [31:0] _RAND_39;
  wire [14:0] _EVAL_2573__EVAL_2574_data;
  wire [1:0] _EVAL_2573__EVAL_2574_addr;
  wire [14:0] _EVAL_2573__EVAL_2575_data;
  wire [1:0] _EVAL_2573__EVAL_2575_addr;
  wire  _EVAL_2573__EVAL_2575_mask;
  wire  _EVAL_2573__EVAL_2575_en;
  reg  _EVAL_2580 [0:3];
  reg [31:0] _RAND_40;
  wire  _EVAL_2580__EVAL_2581_data;
  wire [1:0] _EVAL_2580__EVAL_2581_addr;
  wire  _EVAL_2580__EVAL_2582_data;
  wire [1:0] _EVAL_2580__EVAL_2582_addr;
  wire  _EVAL_2580__EVAL_2582_mask;
  wire  _EVAL_2580__EVAL_2582_en;
  reg [2:0] _EVAL_2591 [0:3];
  reg [31:0] _RAND_41;
  wire [2:0] _EVAL_2591__EVAL_2592_data;
  wire [1:0] _EVAL_2591__EVAL_2592_addr;
  wire [2:0] _EVAL_2591__EVAL_2593_data;
  wire [1:0] _EVAL_2591__EVAL_2593_addr;
  wire  _EVAL_2591__EVAL_2593_mask;
  wire  _EVAL_2591__EVAL_2593_en;
  reg  _EVAL_2712 [0:0];
  reg [31:0] _RAND_42;
  wire  _EVAL_2712__EVAL_2713_data;
  wire  _EVAL_2712__EVAL_2713_addr;
  wire  _EVAL_2712__EVAL_2714_data;
  wire  _EVAL_2712__EVAL_2714_addr;
  wire  _EVAL_2712__EVAL_2714_mask;
  wire  _EVAL_2712__EVAL_2714_en;
  reg  _EVAL_2773 [0:3];
  reg [31:0] _RAND_43;
  wire  _EVAL_2773__EVAL_2774_data;
  wire [1:0] _EVAL_2773__EVAL_2774_addr;
  wire  _EVAL_2773__EVAL_2775_data;
  wire [1:0] _EVAL_2773__EVAL_2775_addr;
  wire  _EVAL_2773__EVAL_2775_mask;
  wire  _EVAL_2773__EVAL_2775_en;
  reg  _EVAL_2852 [0:3];
  reg [31:0] _RAND_44;
  wire  _EVAL_2852__EVAL_2853_data;
  wire [1:0] _EVAL_2852__EVAL_2853_addr;
  wire  _EVAL_2852__EVAL_2854_data;
  wire [1:0] _EVAL_2852__EVAL_2854_addr;
  wire  _EVAL_2852__EVAL_2854_mask;
  wire  _EVAL_2852__EVAL_2854_en;
  reg  _EVAL_3001 [0:0];
  reg [31:0] _RAND_45;
  wire  _EVAL_3001__EVAL_3002_data;
  wire  _EVAL_3001__EVAL_3002_addr;
  wire  _EVAL_3001__EVAL_3003_data;
  wire  _EVAL_3001__EVAL_3003_addr;
  wire  _EVAL_3001__EVAL_3003_mask;
  wire  _EVAL_3001__EVAL_3003_en;
  reg [1:0] _EVAL_3082 [0:0];
  reg [31:0] _RAND_46;
  wire [1:0] _EVAL_3082__EVAL_3083_data;
  wire  _EVAL_3082__EVAL_3083_addr;
  wire [1:0] _EVAL_3082__EVAL_3084_data;
  wire  _EVAL_3082__EVAL_3084_addr;
  wire  _EVAL_3082__EVAL_3084_mask;
  wire  _EVAL_3082__EVAL_3084_en;
  reg [2:0] _EVAL_3112 [0:3];
  reg [31:0] _RAND_47;
  wire [2:0] _EVAL_3112__EVAL_3113_data;
  wire [1:0] _EVAL_3112__EVAL_3113_addr;
  wire [2:0] _EVAL_3112__EVAL_3114_data;
  wire [1:0] _EVAL_3112__EVAL_3114_addr;
  wire  _EVAL_3112__EVAL_3114_mask;
  wire  _EVAL_3112__EVAL_3114_en;
  reg  _EVAL_3335 [0:3];
  reg [31:0] _RAND_48;
  wire  _EVAL_3335__EVAL_3336_data;
  wire [1:0] _EVAL_3335__EVAL_3336_addr;
  wire  _EVAL_3335__EVAL_3337_data;
  wire [1:0] _EVAL_3335__EVAL_3337_addr;
  wire  _EVAL_3335__EVAL_3337_mask;
  wire  _EVAL_3335__EVAL_3337_en;
  reg  _EVAL_155;
  reg [31:0] _RAND_49;
  wire  _EVAL_228;
  reg  _EVAL_227;
  reg [31:0] _RAND_50;
  reg [51:0] _EVAL_253;
  reg [63:0] _RAND_51;
  wire  _EVAL_751;
  wire  _EVAL_255;
  reg [1:0] _EVAL_254;
  reg [31:0] _RAND_52;
  reg  _EVAL_271;
  reg [31:0] _RAND_53;
  reg  _EVAL_287;
  reg [31:0] _RAND_54;
  reg [2:0] _EVAL_306;
  reg [31:0] _RAND_55;
  reg [7:0] _EVAL_314;
  reg [31:0] _RAND_56;
  reg  _EVAL_339;
  reg [31:0] _RAND_57;
  reg  _EVAL_344;
  reg [31:0] _RAND_58;
  reg [8:0] _EVAL_352;
  reg [31:0] _RAND_59;
  reg  _EVAL_374;
  reg [31:0] _RAND_60;
  reg [51:0] _EVAL_397;
  reg [63:0] _RAND_61;
  reg  _EVAL_430;
  reg [31:0] _RAND_62;
  reg [51:0] _EVAL_446;
  reg [63:0] _RAND_63;
  reg [7:0] _EVAL_454;
  reg [31:0] _RAND_64;
  reg [2:0] _EVAL_481;
  reg [31:0] _RAND_65;
  reg [51:0] _EVAL_492;
  reg [63:0] _RAND_66;
  reg  _EVAL_591;
  reg [31:0] _RAND_67;
  reg  _EVAL_664;
  reg [31:0] _RAND_68;
  reg  _EVAL_700;
  reg [31:0] _RAND_69;
  reg [51:0] _EVAL_722;
  reg [63:0] _RAND_70;
  reg  _EVAL_731;
  reg [31:0] _RAND_71;
  reg [51:0] _EVAL_794;
  reg [63:0] _RAND_72;
  reg [127:0] _EVAL_837;
  reg [127:0] _RAND_73;
  reg  _EVAL_839;
  reg [31:0] _RAND_74;
  reg [20:0] _EVAL_849;
  reg [31:0] _RAND_75;
  reg [51:0] _EVAL_856;
  reg [63:0] _RAND_76;
  reg  _EVAL_865;
  reg [31:0] _RAND_77;
  reg  _EVAL_900;
  reg [31:0] _RAND_78;
  reg  _EVAL_927;
  reg [31:0] _RAND_79;
  reg  _EVAL_928;
  reg [31:0] _RAND_80;
  reg  _EVAL_947;
  reg [31:0] _RAND_81;
  reg [8:0] _EVAL_954;
  reg [31:0] _RAND_82;
  reg  _EVAL_957;
  reg [31:0] _RAND_83;
  reg  _EVAL_959;
  reg [31:0] _RAND_84;
  wire  _EVAL_973;
  reg  _EVAL_972;
  reg [31:0] _RAND_85;
  reg  _EVAL_975;
  reg [31:0] _RAND_86;
  reg  _EVAL_1004;
  reg [31:0] _RAND_87;
  reg [20:0] _EVAL_1023;
  reg [31:0] _RAND_88;
  reg  _EVAL_1031;
  reg [31:0] _RAND_89;
  reg  _EVAL_1085;
  reg [31:0] _RAND_90;
  reg [2:0] _EVAL_1102;
  reg [31:0] _RAND_91;
  reg [8:0] _EVAL_1128;
  reg [31:0] _RAND_92;
  reg [51:0] _EVAL_1152;
  reg [63:0] _RAND_93;
  reg [31:0] _EVAL_1163;
  reg [31:0] _RAND_94;
  reg  _EVAL_1165;
  reg [31:0] _RAND_95;
  reg [63:0] _EVAL_1168;
  reg [63:0] _RAND_96;
  reg [51:0] _EVAL_1175;
  reg [63:0] _RAND_97;
  reg  _EVAL_1176;
  reg [31:0] _RAND_98;
  reg  _EVAL_1199;
  reg [31:0] _RAND_99;
  reg [31:0] _EVAL_1243;
  reg [31:0] _RAND_100;
  reg  _EVAL_1244;
  reg [31:0] _RAND_101;
  reg [8:0] _EVAL_1259;
  reg [31:0] _RAND_102;
  reg  _EVAL_1269;
  reg [31:0] _RAND_103;
  reg  _EVAL_1272;
  reg [31:0] _RAND_104;
  reg  _EVAL_1303;
  reg [31:0] _RAND_105;
  reg  _EVAL_1344;
  reg [31:0] _RAND_106;
  reg [51:0] _EVAL_1352;
  reg [63:0] _RAND_107;
  reg  _EVAL_1372;
  reg [31:0] _RAND_108;
  reg  _EVAL_1386;
  reg [31:0] _RAND_109;
  reg [6:0] _EVAL_1387;
  reg [31:0] _RAND_110;
  reg [8:0] _EVAL_1394;
  reg [31:0] _RAND_111;
  reg  _EVAL_1412;
  reg [31:0] _RAND_112;
  reg  _EVAL_1415;
  reg [31:0] _RAND_113;
  reg [63:0] _EVAL_1434;
  reg [63:0] _RAND_114;
  reg [51:0] _EVAL_1487;
  reg [63:0] _RAND_115;
  reg [11:0] _EVAL_1522;
  reg [31:0] _RAND_116;
  reg  _EVAL_1523;
  reg [31:0] _RAND_117;
  reg  _EVAL_1529;
  reg [31:0] _RAND_118;
  reg [63:0] _EVAL_1544;
  reg [63:0] _RAND_119;
  reg  _EVAL_1591;
  reg [31:0] _RAND_120;
  reg  _EVAL_1649;
  reg [31:0] _RAND_121;
  reg  _EVAL_1663;
  reg [31:0] _RAND_122;
  reg  _EVAL_1673;
  reg [31:0] _RAND_123;
  reg  _EVAL_1692;
  reg [31:0] _RAND_124;
  reg [3:0] _EVAL_1706;
  reg [31:0] _RAND_125;
  reg [127:0] _EVAL_1714;
  reg [127:0] _RAND_126;
  reg  _EVAL_1731;
  reg [31:0] _RAND_127;
  reg [8:0] _EVAL_1746;
  reg [31:0] _RAND_128;
  reg  _EVAL_1748;
  reg [31:0] _RAND_129;
  reg [8:0] _EVAL_1755;
  reg [31:0] _RAND_130;
  reg  _EVAL_1762;
  reg [31:0] _RAND_131;
  reg [20:0] _EVAL_1785;
  reg [31:0] _RAND_132;
  reg  _EVAL_1807;
  reg [31:0] _RAND_133;
  reg  _EVAL_1836;
  reg [31:0] _RAND_134;
  reg [24:0] _EVAL_1846;
  reg [31:0] _RAND_135;
  reg  _EVAL_1848;
  reg [31:0] _RAND_136;
  reg [14:0] _EVAL_1886;
  reg [31:0] _RAND_137;
  reg  _EVAL_1953;
  reg [31:0] _RAND_138;
  reg  _EVAL_1954;
  reg [31:0] _RAND_139;
  reg  _EVAL_1957;
  reg [31:0] _RAND_140;
  reg [4:0] _EVAL_1993;
  reg [31:0] _RAND_141;
  reg [255:0] _EVAL_2031;
  reg [255:0] _RAND_142;
  reg  _EVAL_2053;
  reg [31:0] _RAND_143;
  reg [63:0] _EVAL_2062;
  reg [63:0] _RAND_144;
  reg [63:0] _EVAL_2078;
  reg [63:0] _RAND_145;
  reg  _EVAL_2084;
  reg [31:0] _RAND_146;
  reg [51:0] _EVAL_2170;
  reg [63:0] _RAND_147;
  reg  _EVAL_2189;
  reg [31:0] _RAND_148;
  reg [1:0] _EVAL_2212;
  reg [31:0] _RAND_149;
  reg [31:0] _EVAL_2235;
  reg [31:0] _RAND_150;
  reg [1:0] _EVAL_2248;
  reg [31:0] _RAND_151;
  reg  _EVAL_2252;
  reg [31:0] _RAND_152;
  reg [51:0] _EVAL_2270;
  reg [63:0] _RAND_153;
  reg [31:0] _EVAL_2273;
  reg [31:0] _RAND_154;
  reg  _EVAL_2274;
  reg [31:0] _RAND_155;
  reg  _EVAL_2292;
  reg [31:0] _RAND_156;
  reg  _EVAL_2294;
  reg [31:0] _RAND_157;
  reg  _EVAL_2304;
  reg [31:0] _RAND_158;
  reg  _EVAL_2347;
  reg [31:0] _RAND_159;
  reg  _EVAL_2378;
  reg [31:0] _RAND_160;
  reg [63:0] _EVAL_2383;
  reg [63:0] _RAND_161;
  reg [31:0] _EVAL_2392;
  reg [31:0] _RAND_162;
  reg  _EVAL_2398;
  reg [31:0] _RAND_163;
  reg  _EVAL_2399;
  reg [31:0] _RAND_164;
  reg [31:0] _EVAL_2402;
  reg [31:0] _RAND_165;
  reg  _EVAL_2413;
  reg [31:0] _RAND_166;
  reg  _EVAL_2447;
  reg [31:0] _RAND_167;
  reg  _EVAL_2518;
  reg [31:0] _RAND_168;
  reg [1:0] _EVAL_2528;
  reg [31:0] _RAND_169;
  reg [63:0] _EVAL_2534;
  reg [63:0] _RAND_170;
  reg [31:0] _EVAL_2549;
  reg [31:0] _RAND_171;
  reg  _EVAL_2550;
  reg [31:0] _RAND_172;
  reg  _EVAL_2629;
  reg [31:0] _RAND_173;
  reg  _EVAL_2640;
  reg [31:0] _RAND_174;
  reg [63:0] _EVAL_2655;
  reg [63:0] _RAND_175;
  reg  _EVAL_2663;
  reg [31:0] _RAND_176;
  reg [31:0] _EVAL_2686;
  reg [31:0] _RAND_177;
  reg [8:0] _EVAL_2721;
  reg [31:0] _RAND_178;
  reg [51:0] _EVAL_2746;
  reg [63:0] _RAND_179;
  reg [63:0] _EVAL_2785;
  reg [63:0] _RAND_180;
  reg  _EVAL_2799;
  reg [31:0] _RAND_181;
  reg  _EVAL_2806;
  reg [31:0] _RAND_182;
  reg  _EVAL_2808;
  reg [31:0] _RAND_183;
  reg  _EVAL_2880;
  reg [31:0] _RAND_184;
  reg  _EVAL_2882;
  reg [31:0] _RAND_185;
  reg  _EVAL_2887;
  reg [31:0] _RAND_186;
  reg  _EVAL_2888;
  reg [31:0] _RAND_187;
  reg  _EVAL_2915;
  reg [31:0] _RAND_188;
  reg [127:0] _EVAL_2928;
  reg [127:0] _RAND_189;
  reg [127:0] _EVAL_2950;
  reg [127:0] _RAND_190;
  reg [63:0] _EVAL_2971;
  reg [63:0] _RAND_191;
  reg  _EVAL_3019;
  reg [31:0] _RAND_192;
  reg [6:0] _EVAL_3050;
  reg [31:0] _RAND_193;
  reg  _EVAL_3054;
  reg [31:0] _RAND_194;
  reg  _EVAL_3089;
  reg [31:0] _RAND_195;
  reg [1:0] _EVAL_3143;
  reg [31:0] _RAND_196;
  reg  _EVAL_3173;
  reg [31:0] _RAND_197;
  reg [51:0] _EVAL_3187;
  reg [63:0] _RAND_198;
  reg [51:0] _EVAL_3198;
  reg [63:0] _RAND_199;
  reg  _EVAL_3220;
  reg [31:0] _RAND_200;
  reg [20:0] _EVAL_3225;
  reg [31:0] _RAND_201;
  reg  _EVAL_3261;
  reg [31:0] _RAND_202;
  reg  _EVAL_3284;
  reg [31:0] _RAND_203;
  reg [1:0] _EVAL_3292;
  reg [31:0] _RAND_204;
  reg [15:0] _EVAL_3338;
  reg [31:0] _RAND_205;
  reg  _EVAL_3340;
  reg [31:0] _RAND_206;
  reg  _EVAL_3370;
  reg [31:0] _RAND_207;
  reg [15:0] _EVAL_3376;
  reg [31:0] _RAND_208;
  reg  _EVAL_3394;
  reg [31:0] _RAND_209;
  reg  _EVAL_3402;
  reg [31:0] _RAND_210;
  reg [7:0] _EVAL_3406;
  reg [31:0] _RAND_211;
  wire  _EVAL_1981;
  wire  _EVAL_3080;
  wire  _EVAL_1781;
  wire  _EVAL_2472;
  wire  _EVAL_2092;
  wire [8:0] _EVAL_2897;
  wire  _EVAL_1677;
  wire  _EVAL_1751;
  wire  _EVAL_1192;
  wire  _EVAL_1636;
  wire [11:0] _EVAL_1980;
  wire  _EVAL_1215;
  wire  _EVAL_3321;
  wire  _EVAL_1955;
  wire  _EVAL_362;
  wire  _EVAL_3076;
  wire  _EVAL_1983;
  wire  _EVAL_1365;
  wire  _EVAL_1589;
  wire  _EVAL_1841;
  wire  _EVAL_2288;
  wire  _EVAL_1797;
  wire  _EVAL_3092;
  wire  _EVAL_542;
  wire  _EVAL_182;
  wire  _EVAL_3181;
  wire  _EVAL_645;
  wire  _EVAL_956;
  wire [1:0] _EVAL_169;
  wire  _EVAL_2191;
  wire [2:0] _EVAL_2658;
  wire  _EVAL_518;
  wire  _EVAL_2969;
  wire  _EVAL_2018;
  wire  _EVAL_159;
  wire [1:0] _EVAL_724;
  wire  _EVAL_786;
  wire  _EVAL_1313;
  wire  _EVAL_282;
  wire  _EVAL_1605;
  wire  _EVAL_2723;
  wire  _EVAL_2465;
  wire  _EVAL_1426;
  wire  _EVAL_2133;
  wire  _EVAL_769;
  wire  _EVAL_1930;
  wire  _EVAL_2443;
  wire  _EVAL_2366;
  wire [63:0] _EVAL_1295;
  wire [63:0] _EVAL_1271;
  wire [63:0] _EVAL_2668;
  wire [63:0] _EVAL_2618;
  wire [63:0] _EVAL_1214;
  wire [63:0] _EVAL_1402;
  wire [63:0] _EVAL_3203;
  wire [63:0] _EVAL_164;
  wire [63:0] _EVAL_442;
  wire [63:0] _EVAL_993;
  wire [63:0] _EVAL_1550;
  wire [63:0] _EVAL_342;
  wire [63:0] _EVAL_502;
  wire [63:0] _EVAL_1613;
  wire [63:0] _EVAL_2947;
  wire [63:0] _EVAL_2761;
  wire [63:0] _EVAL_1504;
  wire [15:0] _EVAL_2227;
  wire [1:0] _EVAL_2168;
  wire  _EVAL_3211;
  wire  _EVAL_2327;
  wire  _EVAL_315;
  wire  _EVAL_2980;
  wire  _EVAL_2621;
  wire [6:0] _EVAL_2728;
  wire [6:0] _EVAL_3276;
  wire  _EVAL_1245;
  wire  _EVAL_1719;
  wire  _EVAL_194;
  wire [15:0] _EVAL_995;
  wire [1:0] _EVAL_1545;
  wire  _EVAL_2645;
  wire  _EVAL_1610;
  wire  _EVAL_3071;
  wire  _EVAL_1607;
  wire  _EVAL_2012;
  wire [6:0] _EVAL_3281;
  wire [6:0] _EVAL_2326;
  wire  _EVAL_684;
  wire  _EVAL_942;
  wire  _EVAL_1114;
  wire [15:0] _EVAL_2291;
  wire [1:0] _EVAL_1952;
  wire  _EVAL_1934;
  wire  _EVAL_1642;
  wire  _EVAL_1557;
  wire  _EVAL_1008;
  wire  _EVAL_902;
  wire [6:0] _EVAL_174;
  wire [6:0] _EVAL_1221;
  wire  _EVAL_393;
  wire  _EVAL_740;
  wire  _EVAL_1078;
  wire [15:0] _EVAL_1336;
  wire [1:0] _EVAL_3064;
  wire  _EVAL_1867;
  wire  _EVAL_2103;
  wire  _EVAL_2557;
  wire  _EVAL_381;
  wire  _EVAL_1035;
  wire  _EVAL_3000;
  wire  _EVAL_336;
  wire  _EVAL_1091;
  wire  _EVAL_1209;
  wire  _EVAL_1967;
  wire  _EVAL_2336;
  wire  _EVAL_1100;
  wire  _EVAL_1732;
  wire  _EVAL_2030;
  wire  _EVAL_2173;
  wire  _EVAL_3348;
  wire  _EVAL_3039;
  wire  _EVAL_402;
  wire  _EVAL_3107;
  wire  _EVAL_1226;
  wire  _EVAL_3303;
  wire  _EVAL_230;
  wire  _EVAL_2458;
  wire  _EVAL_1996;
  wire [126:0] _EVAL_2066;
  wire [127:0] _EVAL_3155;
  wire [127:0] _EVAL_2115;
  wire [1:0] _EVAL_1502;
  wire [125:0] _EVAL_295;
  wire [127:0] _EVAL_1305;
  wire [127:0] _EVAL_349;
  wire [3:0] _EVAL_1893;
  wire [123:0] _EVAL_3038;
  wire [127:0] _EVAL_1358;
  wire [127:0] _EVAL_1772;
  wire [7:0] _EVAL_699;
  wire [119:0] _EVAL_3308;
  wire [127:0] _EVAL_1916;
  wire [127:0] _EVAL_2286;
  wire [15:0] _EVAL_1978;
  wire [111:0] _EVAL_2160;
  wire [127:0] _EVAL_2899;
  wire [127:0] _EVAL_1491;
  wire [31:0] _EVAL_2426;
  wire [95:0] _EVAL_247;
  wire [127:0] _EVAL_1292;
  wire [127:0] _EVAL_2100;
  wire [63:0] _EVAL_2569;
  wire [63:0] _EVAL_2464;
  wire [127:0] _EVAL_2436;
  wire [127:0] _EVAL_1670;
  wire [128:0] _EVAL_691;
  wire  _EVAL_3405;
  wire  _EVAL_2218;
  wire  _EVAL_325;
  wire  _EVAL_2120;
  wire  _EVAL_761;
  wire  _EVAL_187;
  wire  _EVAL_1377;
  wire [128:0] _EVAL_2059;
  wire [127:0] _EVAL_3265;
  wire [128:0] _EVAL_2765;
  wire  _EVAL_892;
  wire [6:0] _EVAL_1592;
  wire [6:0] _EVAL_520;
  wire  _EVAL_2330;
  wire  _EVAL_2486;
  wire  _EVAL_2293;
  wire  _EVAL_178;
  wire [6:0] _EVAL_2365;
  wire  _EVAL_713;
  wire  _EVAL_3075;
  wire  _EVAL_3186;
  wire  _EVAL_3179;
  wire  _EVAL_3006;
  wire  _EVAL_204;
  wire  _EVAL_2794;
  wire [1:0] _EVAL_304;
  wire  _EVAL_3135;
  wire  _EVAL_2384;
  wire [2:0] _EVAL_2068;
  wire  _EVAL_773;
  wire  _EVAL_858;
  wire [1:0] _EVAL_2877;
  wire  _EVAL_2940;
  wire  _EVAL_1851;
  wire  _EVAL_1855;
  wire  _EVAL_2973;
  wire  _EVAL_3016;
  wire  _EVAL_2410;
  wire  _EVAL_2613;
  wire  _EVAL_1143;
  wire  _EVAL_1154;
  wire  _EVAL_2014;
  wire [6:0] _EVAL_1976;
  wire  _EVAL_3106;
  wire  _EVAL_2499;
  wire  _EVAL_1631;
  wire  _EVAL_300;
  wire  _EVAL_249;
  wire  _EVAL_1070;
  wire  _EVAL_2972;
  wire  _EVAL_2975;
  wire  _EVAL_2044;
  wire  _EVAL_867;
  wire  _EVAL_3133;
  wire  _EVAL_2158;
  wire [2:0] _EVAL_779;
  wire  _EVAL_369;
  wire  _EVAL_1343;
  wire [1:0] _EVAL_3258;
  wire  _EVAL_2556;
  wire  _EVAL_2363;
  wire  _EVAL_1025;
  wire  _EVAL_2289;
  wire  _EVAL_735;
  wire  _EVAL_1686;
  wire  _EVAL_2697;
  wire  _EVAL_1159;
  wire  _EVAL_3323;
  wire  _EVAL_1011;
  wire [6:0] _EVAL_2692;
  wire  _EVAL_970;
  wire  _EVAL_2756;
  wire  _EVAL_1564;
  wire  _EVAL_515;
  wire  _EVAL_378;
  wire  _EVAL_2306;
  wire  _EVAL_3163;
  wire  _EVAL_1051;
  wire  _EVAL_2885;
  wire  _EVAL_868;
  wire  _EVAL_3117;
  wire  _EVAL_1276;
  wire [2:0] _EVAL_2755;
  wire  _EVAL_238;
  wire  _EVAL_2431;
  wire [1:0] _EVAL_920;
  wire  _EVAL_1758;
  wire  _EVAL_2043;
  wire  _EVAL_641;
  wire  _EVAL_1400;
  wire  _EVAL_771;
  wire  _EVAL_3063;
  wire  _EVAL_231;
  wire  _EVAL_2020;
  wire  _EVAL_1032;
  wire  _EVAL_1883;
  wire [6:0] _EVAL_989;
  wire  _EVAL_2742;
  wire  _EVAL_1965;
  wire  _EVAL_3319;
  wire  _EVAL_3250;
  wire  _EVAL_184;
  wire  _EVAL_3398;
  wire  _EVAL_2816;
  wire  _EVAL_3169;
  wire  _EVAL_607;
  wire  _EVAL_3105;
  wire [2:0] _EVAL_1580;
  wire  _EVAL_1733;
  wire  _EVAL_2396;
  wire [1:0] _EVAL_3364;
  wire  _EVAL_2451;
  wire  _EVAL_748;
  wire  _EVAL_1193;
  wire  _EVAL_874;
  wire  _EVAL_309;
  wire  _EVAL_1537;
  wire  _EVAL_2353;
  wire  _EVAL_1439;
  wire  _EVAL_1827;
  wire  _EVAL_2198;
  wire  _EVAL_1995;
  wire  _EVAL_935;
  wire  _EVAL_316;
  wire [128:0] _EVAL_2284;
  wire [126:0] _EVAL_2538;
  wire [128:0] _EVAL_166;
  wire [127:0] _EVAL_2531;
  wire  _EVAL_1500;
  wire  _EVAL_624;
  wire  _EVAL_667;
  wire  _EVAL_1311;
  wire  _EVAL_2810;
  wire  _EVAL_3266;
  wire  _EVAL_2049;
  wire  _EVAL_3299;
  wire  _EVAL_1443;
  wire  _EVAL_2521;
  wire  _EVAL_3139;
  wire  _EVAL_2387;
  wire  _EVAL_3264;
  wire  _EVAL_1129;
  wire  _EVAL_3388;
  wire  _EVAL_1711;
  wire  _EVAL_1927;
  wire  _EVAL_2553;
  wire [8:0] _EVAL_2283;
  wire [17:0] _EVAL_2172;
  wire  _EVAL_1195;
  wire  _EVAL_861;
  wire  _EVAL_1804;
  wire  _EVAL_2029;
  wire  _EVAL_145;
  wire  _EVAL_3033;
  wire  _EVAL_3053;
  wire  _EVAL_1475;
  wire  _EVAL_1312;
  wire  _EVAL_419;
  wire  _EVAL_1077;
  wire  _EVAL_2860;
  wire  _EVAL_1640;
  wire  _EVAL_2843;
  wire  _EVAL_273;
  wire  _EVAL_1366;
  wire  _EVAL_3296;
  wire  _EVAL_1463;
  wire  _EVAL_2789;
  wire  _EVAL_1991;
  wire  _EVAL_1375;
  wire  _EVAL_2900;
  wire  _EVAL_2139;
  wire  _EVAL_1169;
  wire  _EVAL_919;
  wire  _EVAL_2394;
  wire  _EVAL_377;
  wire  _EVAL_1036;
  wire  _EVAL_758;
  wire  _EVAL_2671;
  wire  _EVAL_1407;
  wire  _EVAL_474;
  wire [31:0] _EVAL_930;
  wire [31:0] _EVAL_158;
  wire [31:0] _EVAL_1492;
  wire  _EVAL_777;
  wire [15:0] _EVAL_1633;
  wire [13:0] _EVAL_1678;
  wire [2:0] _EVAL_622;
  wire  _EVAL_818;
  wire [4:0] _EVAL_1779;
  wire  _EVAL_1618;
  wire [1:0] _EVAL_305;
  wire  _EVAL_1136;
  wire  _EVAL_553;
  wire  _EVAL_937;
  wire  _EVAL_1469;
  wire [1:0] _EVAL_1870;
  wire [1:0] _EVAL_318;
  wire [15:0] _EVAL_1189;
  wire [13:0] _EVAL_1517;
  wire [2:0] _EVAL_1556;
  wire  _EVAL_3234;
  wire [4:0] _EVAL_1021;
  wire  _EVAL_235;
  wire [1:0] _EVAL_1721;
  wire  _EVAL_2351;
  wire  _EVAL_657;
  wire  _EVAL_1045;
  wire  _EVAL_2099;
  wire [1:0] _EVAL_2833;
  wire [1:0] _EVAL_2085;
  wire [31:0] _EVAL_876;
  wire  _EVAL_2342;
  wire  _EVAL_2646;
  wire  _EVAL_2913;
  wire  _EVAL_2165;
  wire [10:0] _EVAL_2867;
  wire [10:0] _EVAL_3278;
  wire [7:0] _EVAL_1948;
  wire [7:0] _EVAL_882;
  wire [7:0] _EVAL_1079;
  wire  _EVAL_2493;
  wire  _EVAL_1274;
  wire  _EVAL_1056;
  wire [5:0] _EVAL_3248;
  wire [3:0] _EVAL_3014;
  wire [31:0] _EVAL_2876;
  wire [31:0] _EVAL_860;
  wire [7:0] _EVAL_445;
  wire [7:0] _EVAL_2105;
  wire  _EVAL_331;
  wire  _EVAL_2101;
  wire  _EVAL_829;
  wire [3:0] _EVAL_3061;
  wire [31:0] _EVAL_1219;
  wire [31:0] _EVAL_1014;
  wire [31:0] _EVAL_1743;
  wire  _EVAL_2134;
  wire  _EVAL_3361;
  wire [4:0] _EVAL_2540;
  wire [1:0] _EVAL_2709;
  wire  _EVAL_3159;
  wire [1:0] _EVAL_756;
  wire [1:0] _EVAL_1588;
  wire [12:0] _EVAL_3212;
  wire [12:0] _EVAL_2367;
  wire [9:0] _EVAL_1551;
  wire  _EVAL_2673;
  wire [1:0] _EVAL_1575;
  wire  _EVAL_156;
  wire  _EVAL_2904;
  wire  _EVAL_511;
  wire [2:0] _EVAL_527;
  wire [20:0] _EVAL_1038;
  wire [20:0] _EVAL_604;
  wire [20:0] _EVAL_1362;
  wire [31:0] _EVAL_1534;
  wire [31:0] _EVAL_817;
  wire [31:0] _EVAL_2890;
  wire [31:0] _EVAL_2257;
  wire [31:0] _EVAL_922;
  wire [31:0] _EVAL_2233;
  wire [31:0] _EVAL_3009;
  wire [32:0] _EVAL_1096;
  wire [31:0] _EVAL_462;
  wire [31:0] _EVAL_650;
  wire [31:0] _EVAL_1627;
  wire [4:0] _EVAL_2051;
  wire [4:0] _EVAL_189;
  wire  _EVAL_1926;
  wire  _EVAL_3324;
  wire  _EVAL_2411;
  wire  _EVAL_925;
  wire [3:0] _EVAL_578;
  wire [3:0] _EVAL_2264;
  wire  _EVAL_2701;
  wire  _EVAL_3210;
  wire  _EVAL_272;
  wire [31:0] _EVAL_2977;
  wire [31:0] _EVAL_803;
  wire [31:0] _EVAL_1130;
  wire  _EVAL_1847;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_2504;
  wire  _EVAL_683;
  wire  _EVAL_1111;
  wire  _EVAL_1374;
  wire  _EVAL_1029;
  wire  _EVAL_1281;
  wire  _EVAL_2046;
  wire  _EVAL_1621;
  wire  _EVAL_3333;
  wire  _EVAL_955;
  wire  _EVAL_343;
  wire  _EVAL_1413;
  wire [31:0] _EVAL_477;
  wire [31:0] _EVAL_3178;
  wire  _EVAL_830;
  wire [15:0] _EVAL_3068;
  wire [13:0] _EVAL_540;
  wire [2:0] _EVAL_2921;
  wire  _EVAL_1759;
  wire [4:0] _EVAL_2266;
  wire  _EVAL_1828;
  wire [1:0] _EVAL_1028;
  wire  _EVAL_2425;
  wire  _EVAL_1217;
  wire  _EVAL_2603;
  wire  _EVAL_2533;
  wire [1:0] _EVAL_3282;
  wire [1:0] _EVAL_896;
  wire [15:0] _EVAL_1756;
  wire [13:0] _EVAL_3127;
  wire [2:0] _EVAL_835;
  wire  _EVAL_1146;
  wire [4:0] _EVAL_2878;
  wire  _EVAL_2599;
  wire [1:0] _EVAL_3341;
  wire  _EVAL_3136;
  wire  _EVAL_2174;
  wire  _EVAL_2314;
  wire  _EVAL_766;
  wire [1:0] _EVAL_1211;
  wire [1:0] _EVAL_1735;
  wire [31:0] _EVAL_1144;
  wire  _EVAL_1834;
  wire  _EVAL_1069;
  wire  _EVAL_648;
  wire  _EVAL_2258;
  wire [10:0] _EVAL_2991;
  wire [10:0] _EVAL_384;
  wire [7:0] _EVAL_3395;
  wire [7:0] _EVAL_1929;
  wire [7:0] _EVAL_2130;
  wire  _EVAL_535;
  wire  _EVAL_1567;
  wire  _EVAL_3352;
  wire [5:0] _EVAL_1041;
  wire [3:0] _EVAL_680;
  wire [31:0] _EVAL_1643;
  wire [31:0] _EVAL_1720;
  wire [7:0] _EVAL_3238;
  wire [7:0] _EVAL_2666;
  wire  _EVAL_2088;
  wire  _EVAL_2041;
  wire  _EVAL_2832;
  wire [3:0] _EVAL_1210;
  wire [31:0] _EVAL_1266;
  wire [31:0] _EVAL_1962;
  wire [31:0] _EVAL_360;
  wire  _EVAL_2335;
  wire  _EVAL_1829;
  wire [4:0] _EVAL_763;
  wire [1:0] _EVAL_2171;
  wire  _EVAL_3399;
  wire [1:0] _EVAL_1975;
  wire [1:0] _EVAL_256;
  wire [12:0] _EVAL_755;
  wire [12:0] _EVAL_2834;
  wire [9:0] _EVAL_3379;
  wire  _EVAL_1116;
  wire [1:0] _EVAL_313;
  wire  _EVAL_284;
  wire  _EVAL_1346;
  wire  _EVAL_1960;
  wire [2:0] _EVAL_898;
  wire [20:0] _EVAL_1345;
  wire [20:0] _EVAL_485;
  wire [20:0] _EVAL_2369;
  wire [31:0] _EVAL_1204;
  wire [31:0] _EVAL_573;
  wire [31:0] _EVAL_1672;
  wire [31:0] _EVAL_391;
  wire [31:0] _EVAL_1205;
  wire [31:0] _EVAL_1411;
  wire [4:0] _EVAL_2187;
  wire [4:0] _EVAL_2220;
  wire  _EVAL_1528;
  wire  _EVAL_2060;
  wire  _EVAL_1424;
  wire  _EVAL_416;
  wire [3:0] _EVAL_2872;
  wire [3:0] _EVAL_168;
  wire  _EVAL_1109;
  wire  _EVAL_3056;
  wire  _EVAL_2236;
  wire [31:0] _EVAL_566;
  wire [31:0] _EVAL_302;
  wire [31:0] _EVAL_1602;
  wire  _EVAL_3372;
  wire  _EVAL_1688;
  wire  _EVAL_310;
  wire  _EVAL_1907;
  wire  _EVAL_1308;
  wire  _EVAL_1257;
  wire  _EVAL_2930;
  wire  _EVAL_2938;
  wire  _EVAL_3196;
  wire  _EVAL_1805;
  wire  _EVAL_1300;
  wire  _EVAL_3098;
  wire  _EVAL_431;
  wire  _EVAL_2966;
  wire  _EVAL_2623;
  wire [31:0] _EVAL_2419;
  wire [31:0] _EVAL_581;
  wire  _EVAL_3015;
  wire [15:0] _EVAL_2108;
  wire [13:0] _EVAL_1799;
  wire [2:0] _EVAL_3285;
  wire  _EVAL_2590;
  wire [4:0] _EVAL_939;
  wire  _EVAL_329;
  wire [1:0] _EVAL_1490;
  wire  _EVAL_473;
  wire  _EVAL_2874;
  wire  _EVAL_432;
  wire  _EVAL_2333;
  wire [1:0] _EVAL_2140;
  wire [1:0] _EVAL_2745;
  wire [15:0] _EVAL_1680;
  wire [13:0] _EVAL_884;
  wire [2:0] _EVAL_1830;
  wire  _EVAL_2561;
  wire [4:0] _EVAL_1554;
  wire  _EVAL_2155;
  wire [1:0] _EVAL_1232;
  wire  _EVAL_2512;
  wire  _EVAL_210;
  wire  _EVAL_2644;
  wire  _EVAL_2837;
  wire [1:0] _EVAL_1187;
  wire [1:0] _EVAL_3312;
  wire [31:0] _EVAL_2798;
  wire  _EVAL_1373;
  wire  _EVAL_2551;
  wire  _EVAL_968;
  wire  _EVAL_1979;
  wire [10:0] _EVAL_638;
  wire [10:0] _EVAL_768;
  wire [7:0] _EVAL_3100;
  wire [7:0] _EVAL_1538;
  wire [7:0] _EVAL_2356;
  wire  _EVAL_3294;
  wire  _EVAL_3334;
  wire  _EVAL_244;
  wire [5:0] _EVAL_514;
  wire [3:0] _EVAL_2281;
  wire [31:0] _EVAL_3293;
  wire [31:0] _EVAL_3286;
  wire [7:0] _EVAL_1059;
  wire [7:0] _EVAL_3102;
  wire  _EVAL_3152;
  wire  _EVAL_2287;
  wire  _EVAL_1309;
  wire [3:0] _EVAL_1330;
  wire [31:0] _EVAL_1177;
  wire [31:0] _EVAL_2954;
  wire [31:0] _EVAL_2205;
  wire  _EVAL_1155;
  wire  _EVAL_423;
  wire [4:0] _EVAL_2523;
  wire [1:0] _EVAL_1115;
  wire  _EVAL_2530;
  wire [1:0] _EVAL_1868;
  wire [1:0] _EVAL_1455;
  wire [12:0] _EVAL_754;
  wire [12:0] _EVAL_1752;
  wire [9:0] _EVAL_1275;
  wire  _EVAL_3255;
  wire [1:0] _EVAL_555;
  wire  _EVAL_400;
  wire  _EVAL_863;
  wire  _EVAL_2290;
  wire [2:0] _EVAL_1082;
  wire [20:0] _EVAL_2263;
  wire [20:0] _EVAL_2439;
  wire [20:0] _EVAL_2822;
  wire [31:0] _EVAL_3008;
  wire [31:0] _EVAL_687;
  wire [31:0] _EVAL_1549;
  wire [31:0] _EVAL_2490;
  wire [31:0] _EVAL_2232;
  wire [31:0] _EVAL_2766;
  wire [4:0] _EVAL_2323;
  wire [4:0] _EVAL_2965;
  wire  _EVAL_3208;
  wire  _EVAL_1310;
  wire  _EVAL_1453;
  wire  _EVAL_203;
  wire [3:0] _EVAL_2964;
  wire [3:0] _EVAL_833;
  wire  _EVAL_2718;
  wire  _EVAL_1882;
  wire  _EVAL_3410;
  wire [31:0] _EVAL_1290;
  wire [31:0] _EVAL_1134;
  wire [31:0] _EVAL_3407;
  wire  _EVAL_2516;
  wire  _EVAL_2520;
  wire  _EVAL_3262;
  wire  _EVAL_1572;
  wire  _EVAL_2309;
  wire  _EVAL_2163;
  wire  _EVAL_2866;
  wire  _EVAL_3161;
  wire  _EVAL_2208;
  wire  _EVAL_3141;
  wire  _EVAL_192;
  wire  _EVAL_3209;
  wire  _EVAL_618;
  wire  _EVAL_1315;
  wire [31:0] _EVAL_1097;
  wire [31:0] _EVAL_1773;
  wire  _EVAL_3342;
  wire [15:0] _EVAL_245;
  wire [13:0] _EVAL_598;
  wire [2:0] _EVAL_2895;
  wire  _EVAL_2579;
  wire [4:0] _EVAL_2678;
  wire  _EVAL_3289;
  wire [1:0] _EVAL_2881;
  wire  _EVAL_2702;
  wire  _EVAL_1206;
  wire  _EVAL_1002;
  wire  _EVAL_1318;
  wire [1:0] _EVAL_229;
  wire [1:0] _EVAL_3277;
  wire [15:0] _EVAL_1355;
  wire [13:0] _EVAL_2219;
  wire [2:0] _EVAL_1648;
  wire  _EVAL_1959;
  wire [4:0] _EVAL_1604;
  wire  _EVAL_3290;
  wire [1:0] _EVAL_2272;
  wire  _EVAL_1397;
  wire  _EVAL_2840;
  wire  _EVAL_2909;
  wire  _EVAL_1888;
  wire [1:0] _EVAL_1816;
  wire [1:0] _EVAL_3409;
  wire [31:0] _EVAL_2681;
  wire  _EVAL_150;
  wire  _EVAL_2382;
  wire  _EVAL_870;
  wire  _EVAL_3041;
  wire [10:0] _EVAL_2352;
  wire [10:0] _EVAL_2355;
  wire [7:0] _EVAL_2240;
  wire [7:0] _EVAL_213;
  wire [7:0] _EVAL_1559;
  wire  _EVAL_2423;
  wire  _EVAL_163;
  wire  _EVAL_2738;
  wire [5:0] _EVAL_2960;
  wire [3:0] _EVAL_565;
  wire [31:0] _EVAL_2129;
  wire [31:0] _EVAL_782;
  wire [7:0] _EVAL_1630;
  wire [7:0] _EVAL_1823;
  wire  _EVAL_3185;
  wire  _EVAL_1461;
  wire  _EVAL_276;
  wire [3:0] _EVAL_625;
  wire [31:0] _EVAL_1060;
  wire [31:0] _EVAL_3018;
  wire [31:0] _EVAL_3166;
  wire  _EVAL_653;
  wire  _EVAL_875;
  wire [4:0] _EVAL_3396;
  wire [1:0] _EVAL_2433;
  wire  _EVAL_2262;
  wire [1:0] _EVAL_1495;
  wire [1:0] _EVAL_3060;
  wire [12:0] _EVAL_185;
  wire [12:0] _EVAL_1162;
  wire [9:0] _EVAL_2009;
  wire  _EVAL_2389;
  wire [1:0] _EVAL_819;
  wire  _EVAL_1327;
  wire  _EVAL_1969;
  wire  _EVAL_2814;
  wire [2:0] _EVAL_2583;
  wire [20:0] _EVAL_3087;
  wire [20:0] _EVAL_525;
  wire [20:0] _EVAL_3384;
  wire [31:0] _EVAL_2156;
  wire [31:0] _EVAL_3326;
  wire [31:0] _EVAL_2803;
  wire [31:0] _EVAL_2079;
  wire [31:0] _EVAL_2175;
  wire [31:0] _EVAL_191;
  wire [4:0] _EVAL_2376;
  wire [4:0] _EVAL_3377;
  wire  _EVAL_842;
  wire  _EVAL_1887;
  wire  _EVAL_1478;
  wire  _EVAL_1508;
  wire [3:0] _EVAL_2142;
  wire [3:0] _EVAL_2968;
  wire  _EVAL_3267;
  wire  _EVAL_2546;
  wire  _EVAL_1644;
  wire [31:0] _EVAL_161;
  wire [31:0] _EVAL_1579;
  wire [31:0] _EVAL_233;
  wire  _EVAL_1236;
  wire  _EVAL_3221;
  wire [31:0] _EVAL_1742;
  wire [15:0] _EVAL_696;
  wire [15:0] _EVAL_1662;
  wire [15:0] _EVAL_197;
  wire [31:0] _EVAL_1657;
  wire  _EVAL_3316;
  wire [15:0] _EVAL_605;
  wire [13:0] _EVAL_1183;
  wire [2:0] _EVAL_347;
  wire  _EVAL_193;
  wire [4:0] _EVAL_2317;
  wire  _EVAL_546;
  wire [1:0] _EVAL_3142;
  wire  _EVAL_2036;
  wire  _EVAL_2585;
  wire  _EVAL_1815;
  wire  _EVAL_2350;
  wire [1:0] _EVAL_311;
  wire [1:0] _EVAL_2176;
  wire [15:0] _EVAL_1885;
  wire [13:0] _EVAL_2986;
  wire [2:0] _EVAL_2996;
  wire  _EVAL_517;
  wire [4:0] _EVAL_407;
  wire  _EVAL_1421;
  wire [1:0] _EVAL_3360;
  wire  _EVAL_2689;
  wire  _EVAL_1174;
  wire  _EVAL_469;
  wire  _EVAL_1433;
  wire [1:0] _EVAL_307;
  wire [1:0] _EVAL_1570;
  wire [31:0] _EVAL_998;
  wire  _EVAL_2334;
  wire  _EVAL_2097;
  wire  _EVAL_1831;
  wire  _EVAL_1821;
  wire [10:0] _EVAL_2871;
  wire [10:0] _EVAL_1361;
  wire [7:0] _EVAL_2597;
  wire [7:0] _EVAL_268;
  wire [7:0] _EVAL_3260;
  wire  _EVAL_3020;
  wire  _EVAL_188;
  wire  _EVAL_332;
  wire [5:0] _EVAL_1027;
  wire [3:0] _EVAL_853;
  wire [31:0] _EVAL_3193;
  wire [31:0] _EVAL_1444;
  wire [7:0] _EVAL_2739;
  wire [7:0] _EVAL_1098;
  wire  _EVAL_375;
  wire  _EVAL_2095;
  wire  _EVAL_2606;
  wire [3:0] _EVAL_1220;
  wire [31:0] _EVAL_2498;
  wire [31:0] _EVAL_3382;
  wire [31:0] _EVAL_1367;
  wire  _EVAL_2733;
  wire  _EVAL_358;
  wire [4:0] _EVAL_3130;
  wire [1:0] _EVAL_554;
  wire  _EVAL_296;
  wire [1:0] _EVAL_3263;
  wire [1:0] _EVAL_2344;
  wire [12:0] _EVAL_1200;
  wire [12:0] _EVAL_199;
  wire [9:0] _EVAL_3109;
  wire  _EVAL_1818;
  wire [1:0] _EVAL_2167;
  wire  _EVAL_2957;
  wire  _EVAL_2244;
  wire  _EVAL_2650;
  wire [2:0] _EVAL_615;
  wire [20:0] _EVAL_749;
  wire [20:0] _EVAL_2328;
  wire [20:0] _EVAL_1796;
  wire [31:0] _EVAL_646;
  wire [31:0] _EVAL_859;
  wire [31:0] _EVAL_2788;
  wire [31:0] _EVAL_2605;
  wire [4:0] _EVAL_2223;
  wire [4:0] _EVAL_1760;
  wire  _EVAL_1596;
  wire [31:0] _EVAL_2061;
  wire [31:0] _EVAL_3201;
  wire [31:0] _EVAL_1780;
  wire [31:0] _EVAL_757;
  wire [31:0] _EVAL_1510;
  wire [31:0] _EVAL_2136;
  wire [31:0] _EVAL_690;
  wire  _EVAL_1260;
  wire  _EVAL_820;
  wire  _EVAL_997;
  wire [14:0] _EVAL_417;
  wire [14:0] _EVAL_647;
  wire  _EVAL_2894;
  wire  _EVAL_572;
  wire  _EVAL_2388;
  wire  _EVAL_907;
  wire [14:0] _EVAL_2662;
  wire  _EVAL_889;
  wire  _EVAL_1909;
  wire  _EVAL_2424;
  wire  _EVAL_3287;
  wire [14:0] _EVAL_341;
  wire  _EVAL_2898;
  wire  _EVAL_335;
  wire  _EVAL_3153;
  wire  _EVAL_2994;
  wire [14:0] _EVAL_2724;
  wire  _EVAL_243;
  wire  _EVAL_2135;
  wire  _EVAL_3128;
  wire  _EVAL_3346;
  wire [14:0] _EVAL_1946;
  wire  _EVAL_1705;
  wire  _EVAL_3048;
  wire  _EVAL_2370;
  wire  _EVAL_1617;
  wire [14:0] _EVAL_2400;
  wire  _EVAL_270;
  wire  _EVAL_1094;
  wire  _EVAL_753;
  wire  _EVAL_1218;
  wire [14:0] _EVAL_1687;
  wire  _EVAL_1354;
  wire  _EVAL_2405;
  wire  _EVAL_3373;
  wire  _EVAL_815;
  wire [14:0] _EVAL_2757;
  wire  _EVAL_149;
  wire  _EVAL_1436;
  wire  _EVAL_2444;
  wire  _EVAL_816;
  wire [14:0] _EVAL_2936;
  wire  _EVAL_1428;
  wire  _EVAL_3030;
  wire  _EVAL_1974;
  wire  _EVAL_2507;
  wire [14:0] _EVAL_1026;
  wire  _EVAL_1524;
  wire  _EVAL_569;
  wire  _EVAL_1691;
  wire  _EVAL_594;
  wire [14:0] _EVAL_977;
  wire  _EVAL_3218;
  wire  _EVAL_2146;
  wire  _EVAL_2297;
  wire  _EVAL_2217;
  wire [14:0] _EVAL_221;
  wire  _EVAL_678;
  wire  _EVAL_3275;
  wire  _EVAL_2607;
  wire  _EVAL_2839;
  wire [14:0] _EVAL_2277;
  wire  _EVAL_767;
  wire  _EVAL_2740;
  wire  _EVAL_2111;
  wire  _EVAL_2541;
  wire [14:0] _EVAL_1539;
  wire  _EVAL_479;
  wire  _EVAL_420;
  wire  _EVAL_990;
  wire  _EVAL_2427;
  wire [14:0] _EVAL_1729;
  wire  _EVAL_2373;
  wire  _EVAL_2495;
  wire  _EVAL_2261;
  wire  _EVAL_1734;
  wire [14:0] _EVAL_2005;
  wire  _EVAL_1808;
  wire  _EVAL_3189;
  wire [7:0] _EVAL_439;
  wire [15:0] _EVAL_3329;
  wire  _EVAL_2063;
  wire  _EVAL_1503;
  wire [51:0] _EVAL_3230;
  wire [51:0] _EVAL_1363;
  wire [51:0] _EVAL_3274;
  wire [51:0] _EVAL_1863;
  wire [51:0] _EVAL_3116;
  wire [51:0] _EVAL_1766;
  wire [51:0] _EVAL_2729;
  wire [51:0] _EVAL_2948;
  wire [51:0] _EVAL_1599;
  wire [51:0] _EVAL_3245;
  wire [51:0] _EVAL_3151;
  wire [51:0] _EVAL_1940;
  wire [51:0] _EVAL_1937;
  wire [51:0] _EVAL_2857;
  wire [51:0] _EVAL_552;
  wire [51:0] _EVAL_176;
  wire [51:0] _EVAL_1178;
  wire [51:0] _EVAL_1197;
  wire [51:0] _EVAL_2162;
  wire [51:0] _EVAL_2343;
  wire [51:0] _EVAL_1561;
  wire [51:0] _EVAL_654;
  wire [51:0] _EVAL_936;
  wire [51:0] _EVAL_3025;
  wire [51:0] _EVAL_2896;
  wire [51:0] _EVAL_2253;
  wire [51:0] _EVAL_1963;
  wire [51:0] _EVAL_389;
  wire [51:0] _EVAL_941;
  wire [51:0] _EVAL_1679;
  wire [51:0] _EVAL_1540;
  wire [31:0] _EVAL_1933;
  wire  _EVAL_183;
  wire  _EVAL_3049;
  wire  _EVAL_413;
  wire [10:0] _EVAL_1007;
  wire  _EVAL_1634;
  wire  _EVAL_2552;
  wire  _EVAL_2519;
  wire  _EVAL_541;
  wire [10:0] _EVAL_1289;
  wire [10:0] _EVAL_1396;
  wire [10:0] _EVAL_2403;
  wire [10:0] _EVAL_2159;
  wire [10:0] _EVAL_2301;
  wire [20:0] _EVAL_241;
  wire [31:0] _EVAL_1432;
  wire [31:0] _EVAL_519;
  wire [31:0] _EVAL_895;
  wire [31:0] _EVAL_617;
  wire [31:0] _EVAL_811;
  wire [31:0] _EVAL_710;
  wire [31:0] _EVAL_3356;
  wire [31:0] _EVAL_1099;
  wire [31:0] _EVAL_175;
  wire [30:0] _EVAL_2690;
  wire [14:0] _EVAL_2754;
  wire [8:0] _EVAL_791;
  wire [26:0] _EVAL_3259;
  wire [8:0] _EVAL_2131;
  wire [3:0] _EVAL_2660;
  wire [4:0] _EVAL_436;
  wire [8:0] _EVAL_3301;
  wire [8:0] _EVAL_770;
  wire [4:0] _EVAL_2704;
  wire [3:0] _EVAL_408;
  wire [8:0] _EVAL_2985;
  wire [8:0] _EVAL_1123;
  wire  _EVAL_2958;
  wire  _EVAL_3028;
  wire  _EVAL_1536;
  wire  _EVAL_1230;
  wire  _EVAL_3012;
  wire  _EVAL_2166;
  wire  _EVAL_1695;
  wire  _EVAL_1353;
  wire  _EVAL_846;
  wire  _EVAL_2612;
  wire  _EVAL_1117;
  wire [4:0] _EVAL_380;
  wire  _EVAL_2907;
  wire  _EVAL_1273;
  wire  _EVAL_2782;
  wire  _EVAL_695;
  wire  _EVAL_698;
  wire  _EVAL_1087;
  wire  _EVAL_2595;
  wire  _EVAL_3057;
  wire  _EVAL_810;
  wire  _EVAL_2657;
  wire [9:0] _EVAL_1628;
  wire [14:0] _EVAL_878;
  wire [35:0] _EVAL_3026;
  wire [8:0] _EVAL_484;
  wire [4:0] _EVAL_2107;
  wire [3:0] _EVAL_1403;
  wire [8:0] _EVAL_1782;
  wire [8:0] _EVAL_2604;
  wire [5:0] _EVAL_1898;
  wire [2:0] _EVAL_157;
  wire [8:0] _EVAL_2641;
  wire [8:0] _EVAL_1891;
  wire  _EVAL_2511;
  wire  _EVAL_2967;
  wire [7:0] _EVAL_1068;
  wire [15:0] _EVAL_1172;
  wire  _EVAL_822;
  wire  _EVAL_672;
  wire  _EVAL_493;
  wire  _EVAL_3272;
  wire  _EVAL_3157;
  wire  _EVAL_2194;
  wire  _EVAL_299;
  wire  _EVAL_1489;
  wire  _EVAL_686;
  wire  _EVAL_2414;
  wire  _EVAL_200;
  wire  _EVAL_1016;
  wire  _EVAL_1089;
  wire  _EVAL_2000;
  wire  _EVAL_2316;
  wire  _EVAL_2779;
  wire [7:0] _EVAL_2380;
  wire [15:0] _EVAL_2359;
  wire [3:0] _EVAL_1317;
  wire [15:0] _EVAL_616;
  wire  _EVAL_3188;
  wire  _EVAL_844;
  wire  _EVAL_2412;
  wire  _EVAL_996;
  wire  _EVAL_2039;
  wire  _EVAL_275;
  wire  _EVAL_1113;
  wire  _EVAL_522;
  wire  _EVAL_632;
  wire  _EVAL_1184;
  wire  _EVAL_1049;
  wire  _EVAL_1689;
  wire  _EVAL_716;
  wire  _EVAL_960;
  wire  _EVAL_437;
  wire  _EVAL_2995;
  wire  _EVAL_805;
  wire  _EVAL_1081;
  wire  _EVAL_715;
  wire  _EVAL_2150;
  wire  _EVAL_2193;
  wire  _EVAL_2824;
  wire  _EVAL_2652;
  wire  _EVAL_966;
  wire  _EVAL_373;
  wire  _EVAL_2572;
  wire [4:0] _EVAL_2345;
  wire  _EVAL_3115;
  wire  _EVAL_1435;
  wire  _EVAL_1044;
  wire  _EVAL_2037;
  wire  _EVAL_2256;
  wire  _EVAL_917;
  wire  _EVAL_2239;
  wire [9:0] _EVAL_1238;
  wire [35:0] _EVAL_1864;
  wire [8:0] _EVAL_453;
  wire [4:0] _EVAL_3097;
  wire [3:0] _EVAL_845;
  wire [8:0] _EVAL_2477;
  wire [8:0] _EVAL_1075;
  wire [5:0] _EVAL_712;
  wire [2:0] _EVAL_3347;
  wire [8:0] _EVAL_2787;
  wire [8:0] _EVAL_288;
  wire [8:0] _EVAL_560;
  wire [6:0] _EVAL_2903;
  wire [1:0] _EVAL_2161;
  wire [8:0] _EVAL_2500;
  wire [8:0] _EVAL_2048;
  wire [8:0] _EVAL_1131;
  wire [7:0] _EVAL_2125;
  wire  _EVAL_2186;
  wire [8:0] _EVAL_261;
  wire [8:0] _EVAL_2564;
  wire  _EVAL_1213;
  wire  _EVAL_1160;
  wire  _EVAL_2711;
  wire  _EVAL_1763;
  wire  _EVAL_2949;
  wire  _EVAL_2797;
  wire  _EVAL_2993;
  wire  _EVAL_165;
  wire  _EVAL_2559;
  wire  _EVAL_1822;
  wire  _EVAL_3236;
  wire  _EVAL_1379;
  wire  _EVAL_543;
  wire [15:0] _EVAL_2554;
  wire [13:0] _EVAL_368;
  wire [2:0] _EVAL_703;
  wire  _EVAL_994;
  wire [4:0] _EVAL_2147;
  wire  _EVAL_1800;
  wire [1:0] _EVAL_3239;
  wire  _EVAL_827;
  wire  _EVAL_427;
  wire  _EVAL_2706;
  wire  _EVAL_2616;
  wire [1:0] _EVAL_1249;
  wire [1:0] _EVAL_3034;
  wire [15:0] _EVAL_781;
  wire [13:0] _EVAL_237;
  wire [2:0] _EVAL_190;
  wire  _EVAL_836;
  wire [4:0] _EVAL_2951;
  wire  _EVAL_3244;
  wire [1:0] _EVAL_504;
  wire  _EVAL_1126;
  wire  _EVAL_1104;
  wire  _EVAL_3297;
  wire  _EVAL_269;
  wire [1:0] _EVAL_3223;
  wire [1:0] _EVAL_265;
  wire [15:0] _EVAL_1431;
  wire [13:0] _EVAL_1598;
  wire [2:0] _EVAL_1063;
  wire  _EVAL_2687;
  wire [4:0] _EVAL_2418;
  wire  _EVAL_1294;
  wire [1:0] _EVAL_1658;
  wire  _EVAL_915;
  wire  _EVAL_1383;
  wire  _EVAL_929;
  wire  _EVAL_2567;
  wire [1:0] _EVAL_2254;
  wire [1:0] _EVAL_913;
  wire [15:0] _EVAL_3197;
  wire [13:0] _EVAL_2237;
  wire [2:0] _EVAL_3369;
  wire  _EVAL_3242;
  wire [4:0] _EVAL_670;
  wire  _EVAL_2199;
  wire [1:0] _EVAL_3389;
  wire  _EVAL_2675;
  wire  _EVAL_3090;
  wire  _EVAL_1669;
  wire  _EVAL_862;
  wire [1:0] _EVAL_472;
  wire [1:0] _EVAL_2688;
  wire [63:0] _EVAL_1641;
  wire [63:0] _EVAL_3247;
  wire [7:0] _EVAL_2826;
  wire  _EVAL_2271;
  wire [2:0] _EVAL_575;
  wire  _EVAL_965;
  wire  _EVAL_2741;
  wire  _EVAL_3381;
  wire  _EVAL_222;
  wire  _EVAL_3021;
  wire  _EVAL_2614;
  wire  _EVAL_1645;
  wire  _EVAL_3029;
  wire  _EVAL_2008;
  wire  _EVAL_635;
  wire  _EVAL_2829;
  wire  _EVAL_2064;
  wire  _EVAL_1037;
  wire  _EVAL_1794;
  wire  _EVAL_219;
  wire  _EVAL_487;
  wire  _EVAL_2911;
  wire [8:0] _EVAL_2568;
  wire [17:0] _EVAL_2143;
  wire [8:0] _EVAL_1006;
  wire [26:0] _EVAL_326;
  wire [8:0] _EVAL_717;
  wire  _EVAL_1376;
  wire  _EVAL_2434;
  wire  _EVAL_1931;
  wire [4:0] _EVAL_843;
  wire  _EVAL_711;
  wire  _EVAL_2508;
  wire  _EVAL_2922;
  wire  _EVAL_1616;
  wire  _EVAL_2138;
  wire  _EVAL_1697;
  wire  _EVAL_2279;
  wire  _EVAL_441;
  wire  _EVAL_2879;
  wire  _EVAL_1694;
  wire  _EVAL_623;
  wire  _EVAL_587;
  wire  _EVAL_2211;
  wire  _EVAL_153;
  wire  _EVAL_3380;
  wire [8:0] _EVAL_2635;
  wire [17:0] _EVAL_676;
  wire [26:0] _EVAL_1990;
  wire [8:0] _EVAL_1019;
  wire [5:0] _EVAL_590;
  wire [2:0] _EVAL_1739;
  wire [8:0] _EVAL_2496;
  wire [8:0] _EVAL_1404;
  wire [6:0] _EVAL_1683;
  wire [1:0] _EVAL_2463;
  wire [8:0] _EVAL_629;
  wire [8:0] _EVAL_729;
  wire  _EVAL_1708;
  wire  _EVAL_976;
  wire  _EVAL_3004;
  wire  _EVAL_460;
  wire  _EVAL_147;
  wire  _EVAL_2636;
  wire  _EVAL_813;
  wire [2:0] _EVAL_626;
  wire [1:0] _EVAL_2584;
  wire [2:0] _EVAL_1468;
  wire [2:0] _EVAL_223;
  wire [3:0] _EVAL_1778;
  wire [3:0] _EVAL_1306;
  wire  _EVAL_350;
  wire  _EVAL_759;
  wire [3:0] _EVAL_2747;
  wire [3:0] _EVAL_495;
  wire [3:0] _EVAL_1297;
  wire [2:0] _EVAL_2743;
  wire  _EVAL_3302;
  wire  _EVAL_2071;
  wire  _EVAL_1514;
  wire  _EVAL_851;
  wire  _EVAL_444;
  wire  _EVAL_901;
  wire  _EVAL_3066;
  wire  _EVAL_665;
  wire  _EVAL_2255;
  wire  _EVAL_2188;
  wire  _EVAL_945;
  wire  _EVAL_2360;
  wire  _EVAL_2783;
  wire [15:0] _EVAL_693;
  wire  _EVAL_814;
  wire  _EVAL_1369;
  wire [15:0] _EVAL_2804;
  wire [15:0] _EVAL_606;
  wire [15:0] _EVAL_3146;
  wire [1:0] _EVAL_399;
  wire  _EVAL_1994;
  wire [11:0] _EVAL_523;
  wire [13:0] _EVAL_671;
  wire  _EVAL_601;
  wire  _EVAL_1793;
  wire  _EVAL_2796;
  wire  _EVAL_248;
  wire  _EVAL_2407;
  wire  _EVAL_2276;
  wire  _EVAL_2295;
  wire  _EVAL_944;
  wire  _EVAL_3408;
  wire  _EVAL_2959;
  wire  _EVAL_728;
  wire  _EVAL_1961;
  wire  _EVAL_2659;
  wire  _EVAL_1384;
  wire  _EVAL_3232;
  wire  _EVAL_2035;
  wire  _EVAL_2238;
  wire  _EVAL_2625;
  wire  _EVAL_885;
  wire  _EVAL_2484;
  wire  _EVAL_2385;
  wire  _EVAL_613;
  wire  _EVAL_3047;
  wire  _EVAL_2719;
  wire  _EVAL_2241;
  wire  _EVAL_1910;
  wire  _EVAL_2132;
  wire  _EVAL_3168;
  wire  _EVAL_1749;
  wire [7:0] _EVAL_796;
  wire [7:0] _EVAL_682;
  wire [6:0] _EVAL_3386;
  wire [6:0] _EVAL_1414;
  wire [6:0] _EVAL_2988;
  wire  _EVAL_737;
  wire  _EVAL_2268;
  wire [1:0] _EVAL_938;
  wire [1:0] _EVAL_1825;
  wire  _EVAL_3231;
  wire  _EVAL_2216;
  wire [1:0] _EVAL_3121;
  wire [1:0] _EVAL_2767;
  wire  _EVAL_2251;
  wire  _EVAL_2157;
  wire  _EVAL_1700;
  wire  _EVAL_3177;
  wire  _EVAL_2807;
  wire  _EVAL_1790;
  wire  _EVAL_666;
  wire  _EVAL_804;
  wire  _EVAL_2934;
  wire  _EVAL_2821;
  wire  _EVAL_1390;
  wire  _EVAL_1535;
  wire [2:0] _EVAL_2642;
  wire [2:0] _EVAL_571;
  wire [2:0] _EVAL_1342;
  wire [2:0] _EVAL_1638;
  wire [5:0] _EVAL_880;
  wire [11:0] _EVAL_2452;
  wire  _EVAL_2467;
  wire [1:0] _EVAL_1382;
  wire [13:0] _EVAL_2610;
  wire [13:0] _EVAL_3172;
  wire [10:0] _EVAL_2016;
  wire [2:0] _EVAL_2121;
  wire [10:0] _EVAL_3119;
  wire [10:0] _EVAL_433;
  wire [138:0] _EVAL_1083;
  wire [138:0] _EVAL_2570;
  wire [138:0] _EVAL_797;
  wire [2:0] _EVAL_1279;
  wire  _EVAL_2210;
  wire  _EVAL_258;
  wire  _EVAL_1423;
  wire  _EVAL_750;
  wire  _EVAL_2468;
  wire  _EVAL_1753;
  wire  _EVAL_181;
  wire  _EVAL_1188;
  wire  _EVAL_1419;
  wire  _EVAL_1922;
  wire  _EVAL_2052;
  wire  _EVAL_707;
  wire  _EVAL_1062;
  wire  _EVAL_1299;
  wire  _EVAL_2999;
  wire  _EVAL_3270;
  wire  _EVAL_366;
  wire  _EVAL_3154;
  wire  _EVAL_576;
  wire  _EVAL_513;
  wire  _EVAL_1584;
  wire  _EVAL_1685;
  wire  _EVAL_2707;
  wire  _EVAL_1371;
  wire  _EVAL_274;
  wire  _EVAL_563;
  wire  _EVAL_1145;
  wire  _EVAL_1736;
  wire  _EVAL_1889;
  wire  _EVAL_1569;
  wire  _EVAL_2446;
  wire  _EVAL_866;
  wire  _EVAL_894;
  wire  _EVAL_2040;
  wire  _EVAL_206;
  wire  _EVAL_883;
  wire  _EVAL_2440;
  wire  _EVAL_466;
  wire  _EVAL_201;
  wire  _EVAL_906;
  wire  _EVAL_2748;
  wire  _EVAL_1603;
  wire  _EVAL_2001;
  wire  _EVAL_2299;
  wire [8:0] _EVAL_2054;
  wire  _EVAL_3167;
  wire  _EVAL_2902;
  wire [1:0] _EVAL_428;
  wire [2:0] _EVAL_3200;
  wire [3:0] _EVAL_2851;
  wire [2:0] _EVAL_3110;
  wire  _EVAL_3044;
  wire  _EVAL_3327;
  wire  _EVAL_1255;
  wire  _EVAL_1237;
  wire  _EVAL_2070;
  wire  _EVAL_1445;
  wire [5:0] _EVAL_1899;
  wire  _EVAL_1553;
  wire  _EVAL_1787;
  wire  _EVAL_2801;
  wire  _EVAL_2905;
  wire [14:0] _EVAL_1857;
  wire  _EVAL_1964;
  wire  _EVAL_3318;
  wire  _EVAL_1932;
  wire  _EVAL_3011;
  wire  _EVAL_1709;
  wire  _EVAL_1010;
  wire  _EVAL_834;
  wire [15:0] _EVAL_1786;
  wire [2:0] _EVAL_1263;
  wire  _EVAL_1552;
  wire  _EVAL_3040;
  wire  _EVAL_1151;
  wire  _EVAL_2893;
  wire  _EVAL_3183;
  wire  _EVAL_589;
  wire  _EVAL_709;
  wire  _EVAL_1340;
  wire  _EVAL_855;
  wire  _EVAL_2087;
  wire  _EVAL_2974;
  wire  _EVAL_251;
  wire [4:0] _EVAL_461;
  wire  _EVAL_2828;
  wire [1:0] _EVAL_1639;
  wire  _EVAL_2282;
  wire  _EVAL_3237;
  wire  _EVAL_1844;
  wire [4:0] _EVAL_333;
  wire [4:0] _EVAL_528;
  wire  _EVAL_3215;
  wire [28:0] _EVAL_2910;
  wire [30:0] _EVAL_2397;
  wire [1:0] _EVAL_841;
  wire [30:0] _EVAL_1186;
  wire [30:0] _EVAL_1915;
  wire [2:0] _EVAL_2015;
  wire [10:0] _EVAL_2633;
  wire [7:0] _EVAL_2278;
  wire [15:0] _EVAL_614;
  wire  _EVAL_1138;
  wire  _EVAL_2615;
  wire  _EVAL_3070;
  wire  _EVAL_943;
  wire  _EVAL_1325;
  wire  _EVAL_2430;
  wire  _EVAL_958;
  wire  _EVAL_1626;
  wire  _EVAL_583;
  wire  _EVAL_3317;
  wire  _EVAL_3219;
  wire  _EVAL_1167;
  wire  _EVAL_2768;
  wire  _EVAL_628;
  wire  _EVAL_1233;
  wire  _EVAL_3132;
  wire [7:0] _EVAL_356;
  wire [15:0] _EVAL_2393;
  wire [1:0] _EVAL_2918;
  wire  _EVAL_979;
  wire [5:0] _EVAL_708;
  wire [8:0] _EVAL_1880;
  wire  _EVAL_2003;
  wire [22:0] _EVAL_1456;
  wire [7:0] _EVAL_2537;
  wire [7:0] _EVAL_2267;
  wire [4:0] _EVAL_1494;
  wire [4:0] _EVAL_639;
  wire [4:0] _EVAL_3144;
  wire [8:0] _EVAL_2106;
  wire [8:0] _EVAL_2122;
  wire  _EVAL_903;
  wire  _EVAL_2705;
  wire [31:0] _EVAL_1357;
  wire [31:0] _EVAL_2437;
  wire [15:0] _EVAL_1810;
  wire [2:0] _EVAL_1458;
  wire  _EVAL_1989;
  wire  _EVAL_179;
  wire  _EVAL_2331;
  wire  _EVAL_2626;
  wire  _EVAL_2539;
  wire  _EVAL_2285;
  wire  _EVAL_904;
  wire  _EVAL_3332;
  wire [9:0] _EVAL_1335;
  wire [35:0] _EVAL_656;
  wire [8:0] _EVAL_1224;
  wire  _EVAL_1585;
  wire [7:0] _EVAL_1998;
  wire [8:0] _EVAL_1972;
  wire  _EVAL_1873;
  wire  _EVAL_2149;
  wire  _EVAL_739;
  wire  _EVAL_1750;
  wire  _EVAL_293;
  wire  _EVAL_2817;
  wire  _EVAL_2944;
  wire [1:0] _EVAL_3206;
  wire  _EVAL_850;
  wire [6:0] _EVAL_1071;
  wire  _EVAL_2422;
  wire  _EVAL_264;
  wire  _EVAL_2485;
  wire  _EVAL_3401;
  wire  _EVAL_1001;
  wire  _EVAL_3072;
  wire  _EVAL_3344;
  wire  _EVAL_609;
  wire  _EVAL_1727;
  wire  _EVAL_3067;
  wire  _EVAL_3311;
  wire  _EVAL_2197;
  wire  _EVAL_1856;
  wire  _EVAL_1106;
  wire  _EVAL_2119;
  wire  _EVAL_1939;
  wire  _EVAL_494;
  wire  _EVAL_2815;
  wire  _EVAL_1582;
  wire  _EVAL_1901;
  wire  _EVAL_3123;
  wire  _EVAL_1280;
  wire  _EVAL_1427;
  wire  _EVAL_2777;
  wire  _EVAL_2677;
  wire  _EVAL_2013;
  wire  _EVAL_2448;
  wire  _EVAL_2250;
  wire  _EVAL_1947;
  wire  _EVAL_1332;
  wire  _EVAL_2303;
  wire  _EVAL_694;
  wire  _EVAL_3378;
  wire  _EVAL_2925;
  wire  _EVAL_1676;
  wire  _EVAL_981;
  wire  _EVAL_3240;
  wire  _EVAL_697;
  wire  _EVAL_2152;
  wire  _EVAL_1632;
  wire  _EVAL_2676;
  wire  _EVAL_577;
  wire  _EVAL_1242;
  wire  _EVAL_689;
  wire  _EVAL_2093;
  wire  _EVAL_832;
  wire [2:0] _EVAL_2202;
  wire  _EVAL_809;
  wire  _EVAL_1460;
  wire [4:0] _EVAL_2933;
  wire  _EVAL_3022;
  wire  _EVAL_1878;
  wire [9:0] _EVAL_3055;
  wire [35:0] _EVAL_260;
  wire [8:0] _EVAL_1093;
  wire [2:0] _EVAL_3404;
  wire  _EVAL_2164;
  wire  _EVAL_1170;
  wire  _EVAL_1359;
  wire  _EVAL_250;
  wire  _EVAL_536;
  wire  _EVAL_1328;
  wire  _EVAL_1715;
  wire  _EVAL_2809;
  wire  _EVAL_1425;
  wire  _EVAL_1370;
  wire  _EVAL_1405;
  wire  _EVAL_3184;
  wire  _EVAL_1659;
  wire  _EVAL_2325;
  wire  _EVAL_1984;
  wire  _EVAL_3217;
  wire  _EVAL_3351;
  wire  _EVAL_1803;
  wire  _EVAL_226;
  wire  _EVAL_1533;
  wire  _EVAL_2260;
  wire  _EVAL_783;
  wire  _EVAL_1977;
  wire  _EVAL_2154;
  wire  _EVAL_3031;
  wire  _EVAL_286;
  wire [15:0] _EVAL_2151;
  wire [4:0] _EVAL_649;
  wire  _EVAL_3058;
  wire  _EVAL_2050;
  wire  _EVAL_2275;
  wire  _EVAL_1018;
  wire  _EVAL_2790;
  wire  _EVAL_3032;
  wire [25:0] _EVAL_916;
  wire  _EVAL_2067;
  wire  _EVAL_1479;
  wire  _EVAL_1173;
  wire  _EVAL_567;
  wire  _EVAL_1282;
  wire  _EVAL_2916;
  wire  _EVAL_1612;
  wire  _EVAL_556;
  wire  _EVAL_1420;
  wire [4:0] _EVAL_1783;
  wire [9:0] _EVAL_760;
  wire [35:0] _EVAL_2868;
  wire  _EVAL_914;
  wire  _EVAL_1430;
  wire  _EVAL_2474;
  wire  _EVAL_2535;
  wire  _EVAL_1437;
  wire  _EVAL_3283;
  wire  _EVAL_2145;
  wire  _EVAL_1712;
  wire  _EVAL_3288;
  wire [4:0] _EVAL_2835;
  wire  _EVAL_1917;
  wire  _EVAL_1307;
  wire  _EVAL_1042;
  wire  _EVAL_2245;
  wire [9:0] _EVAL_3358;
  wire [35:0] _EVAL_3138;
  wire [8:0] _EVAL_2578;
  wire  _EVAL_1565;
  wire [7:0] _EVAL_1270;
  wire [8:0] _EVAL_2823;
  wire [1:0] _EVAL_2664;
  wire  _EVAL_730;
  wire  _EVAL_1105;
  wire  _EVAL_790;
  wire  _EVAL_148;
  wire  _EVAL_2144;
  wire  _EVAL_2760;
  wire  _EVAL_2771;
  wire  _EVAL_651;
  wire  _EVAL_3156;
  wire  _EVAL_338;
  wire  _EVAL_470;
  wire  _EVAL_1664;
  wire  _EVAL_2560;
  wire [1:0] _EVAL_1956;
  wire [1:0] _EVAL_1728;
  wire [1:0] _EVAL_376;
  wire [1:0] _EVAL_1331;
  wire [1:0] _EVAL_266;
  wire  _EVAL_580;
  wire  _EVAL_1824;
  wire [1:0] _EVAL_2608;
  wire  _EVAL_1593;
  wire  _EVAL_2683;
  wire [1:0] _EVAL_1945;
  wire [1:0] _EVAL_2221;
  wire [1:0] _EVAL_2307;
  wire [1:0] _EVAL_636;
  wire [1:0] _EVAL_787;
  wire [1:0] _EVAL_561;
  wire  _EVAL_1511;
  wire  _EVAL_1157;
  wire  _EVAL_3129;
  wire  _EVAL_2010;
  wire  _EVAL_146;
  wire  _EVAL_1248;
  wire [8:0] _EVAL_278;
  wire  _EVAL_2349;
  wire  _EVAL_1410;
  wire [8:0] _EVAL_2080;
  wire [17:0] _EVAL_1067;
  wire [26:0] _EVAL_3387;
  wire [8:0] _EVAL_568;
  wire [7:0] _EVAL_946;
  wire [1:0] _EVAL_2825;
  wire  _EVAL_2180;
  wire  _EVAL_2929;
  wire  _EVAL_2931;
  wire  _EVAL_1725;
  wire  _EVAL_3043;
  wire  _EVAL_785;
  wire  _EVAL_854;
  wire  _EVAL_1894;
  wire  _EVAL_1562;
  wire  _EVAL_2492;
  wire [4:0] _EVAL_1858;
  wire [9:0] _EVAL_2002;
  wire [35:0] _EVAL_234;
  wire [8:0] _EVAL_1936;
  wire [4:0] _EVAL_2588;
  wire [7:0] _EVAL_2791;
  wire [7:0] _EVAL_1103;
  wire [6:0] _EVAL_1158;
  wire  _EVAL_1448;
  wire  _EVAL_999;
  wire  _EVAL_1837;
  wire  _EVAL_2566;
  wire  _EVAL_2487;
  wire  _EVAL_1806;
  wire  _EVAL_3307;
  wire  _EVAL_172;
  wire  _EVAL_1301;
  wire  _EVAL_2609;
  wire  _EVAL_2466;
  wire  _EVAL_220;
  wire  _EVAL_2805;
  wire  _EVAL_2698;
  wire  _EVAL_2891;
  wire  _EVAL_1908;
  wire [63:0] _EVAL_1350;
  wire  _EVAL_2296;
  wire  _EVAL_2845;
  wire  _EVAL_456;
  wire  _EVAL_2886;
  wire  _EVAL_2482;
  wire [15:0] _EVAL_3304;
  wire [2:0] _EVAL_2269;
  wire  _EVAL_2181;
  wire [15:0] _EVAL_2846;
  wire [1:0] _EVAL_308;
  wire  _EVAL_1629;
  wire [5:0] _EVAL_1459;
  wire [11:0] _EVAL_741;
  wire [8:0] _EVAL_637;
  wire [8:0] _EVAL_2601;
  wire  _EVAL_3213;
  wire [8:0] _EVAL_3088;
  wire [8:0] _EVAL_1497;
  wire  _EVAL_1635;
  wire  _EVAL_357;
  wire  _EVAL_1826;
  wire  _EVAL_3069;
  wire  _EVAL_1110;
  wire  _EVAL_1543;
  wire  _EVAL_2200;
  wire  _EVAL_3233;
  wire  _EVAL_2182;
  wire  _EVAL_3013;
  wire  _EVAL_1227;
  wire [2:0] _EVAL_1973;
  wire  _EVAL_312;
  wire [128:0] _EVAL_764;
  wire [128:0] _EVAL_1854;
  wire [15:0] _EVAL_298;
  wire [4:0] _EVAL_1185;
  wire  _EVAL_3345;
  wire [3:0] _EVAL_912;
  wire [8:0] _EVAL_170;
  wire [3:0] _EVAL_2778;
  wire [4:0] _EVAL_2375;
  wire [8:0] _EVAL_2875;
  wire  _EVAL_655;
  wire [127:0] _EVAL_1583;
  wire [1:0] _EVAL_1928;
  wire [125:0] _EVAL_465;
  wire [127:0] _EVAL_2432;
  wire [127:0] _EVAL_524;
  wire [123:0] _EVAL_733;
  wire  _EVAL_2716;
  wire  _EVAL_2090;
  wire  _EVAL_1356;
  wire  _EVAL_1622;
  wire  _EVAL_1581;
  wire [8:0] _EVAL_236;
  wire [17:0] _EVAL_2190;
  wire [26:0] _EVAL_1161;
  wire [8:0] _EVAL_429;
  wire [4:0] _EVAL_1095;
  wire  _EVAL_346;
  wire  _EVAL_1997;
  wire [1:0] _EVAL_1278;
  wire [1:0] _EVAL_499;
  wire  _EVAL_2450;
  wire  _EVAL_2617;
  wire [20:0] _EVAL_1268;
  wire  _EVAL_2420;
  wire [15:0] _EVAL_1968;
  wire [8:0] _EVAL_3295;
  wire [1:0] _EVAL_586;
  wire [5:0] _EVAL_2406;
  wire [7:0] _EVAL_881;
  wire [19:0] _EVAL_2602;
  wire  _EVAL_2892;
  wire  _EVAL_475;
  wire  _EVAL_2114;
  wire  _EVAL_2204;
  wire  _EVAL_1938;
  wire  _EVAL_1418;
  wire  _EVAL_303;
  wire [8:0] _EVAL_2672;
  wire [17:0] _EVAL_1839;
  wire [26:0] _EVAL_1057;
  wire [8:0] _EVAL_2997;
  wire  _EVAL_2332;
  wire  _EVAL_2571;
  wire  _EVAL_1501;
  wire  _EVAL_534;
  wire [28:0] _EVAL_808;
  wire [2:0] _EVAL_2312;
  wire [7:0] _EVAL_1817;
  wire  _EVAL_644;
  wire [7:0] _EVAL_2992;
  wire  _EVAL_1471;
  wire  _EVAL_2442;
  wire  _EVAL_257;
  wire [20:0] _EVAL_2725;
  wire  _EVAL_143;
  wire [7:0] _EVAL_418;
  wire [4:0] _EVAL_1515;
  wire  _EVAL_1698;
  wire  _EVAL_2224;
  wire  _EVAL_934;
  wire  _EVAL_1925;
  wire  _EVAL_1526;
  wire  _EVAL_372;
  wire  _EVAL_1288;
  wire  _EVAL_1388;
  wire  _EVAL_1507;
  wire  _EVAL_3126;
  wire  _EVAL_450;
  wire  _EVAL_2700;
  wire  _EVAL_738;
  wire  _EVAL_1235;
  wire  _EVAL_2863;
  wire [14:0] _EVAL_2653;
  wire [1:0] _EVAL_831;
  wire  _EVAL_788;
  wire [31:0] _EVAL_1054;
  wire [14:0] _EVAL_2941;
  wire  _EVAL_2935;
  wire [51:0] _EVAL_2377;
  wire  _EVAL_864;
  wire  _EVAL_2038;
  wire  _EVAL_3363;
  wire  _EVAL_1139;
  wire  _EVAL_778;
  wire  _EVAL_1682;
  wire [4:0] _EVAL_3094;
  wire  _EVAL_1879;
  wire  _EVAL_621;
  wire  _EVAL_879;
  wire [9:0] _EVAL_2979;
  wire [35:0] _EVAL_3257;
  wire [8:0] _EVAL_2831;
  wire [31:0] _EVAL_2717;
  wire [25:0] _EVAL_3162;
  wire  _EVAL_2749;
  wire [4:0] _EVAL_467;
  wire  _EVAL_2056;
  wire [2:0] _EVAL_2818;
  wire  _EVAL_1222;
  wire [1:0] _EVAL_1696;
  wire  _EVAL_2981;
  wire  _EVAL_847;
  wire [8:0] _EVAL_3325;
  wire [5:0] _EVAL_2184;
  wire  _EVAL_798;
  wire  _EVAL_348;
  wire  _EVAL_1496;
  wire  _EVAL_1577;
  wire  _EVAL_2515;
  wire  _EVAL_792;
  wire  _EVAL_160;
  wire [4:0] _EVAL_2762;
  wire  _EVAL_2736;
  wire  _EVAL_705;
  wire  _EVAL_2622;
  wire  _EVAL_1256;
  wire  _EVAL_196;
  wire [1:0] _EVAL_1137;
  wire [31:0] _EVAL_2576;
  wire [30:0] _EVAL_3095;
  wire [14:0] _EVAL_1090;
  wire [11:0] _EVAL_1665;
  wire [13:0] _EVAL_3204;
  wire [1:0] _EVAL_1262;
  wire [13:0] _EVAL_620;
  wire [13:0] _EVAL_1050;
  wire [4:0] _EVAL_242;
  wire  _EVAL_2183;
  wire [1:0] _EVAL_496;
  wire  _EVAL_322;
  wire  _EVAL_2726;
  wire  _EVAL_2415;
  wire  _EVAL_3081;
  wire [1:0] _EVAL_214;
  wire [5:0] _EVAL_1066;
  wire [11:0] _EVAL_1924;
  wire [8:0] _EVAL_2032;
  wire  _EVAL_2148;
  wire  _EVAL_2927;
  wire  _EVAL_2454;
  wire [8:0] _EVAL_468;
  wire [17:0] _EVAL_1876;
  wire [26:0] _EVAL_1684;
  wire [8:0] _EVAL_152;
  wire [28:0] _EVAL_464;
  wire  _EVAL_1203;
  wire  _EVAL_3191;
  wire  _EVAL_2441;
  wire  _EVAL_3192;
  wire  _EVAL_3079;
  wire  _EVAL_1261;
  wire  _EVAL_1578;
  wire [15:0] _EVAL_1774;
  wire [1:0] _EVAL_1853;
  wire [3:0] _EVAL_2028;
  wire  _EVAL_1771;
  wire [127:0] _EVAL_2529;
  wire  _EVAL_2404;
  wire  _EVAL_1234;
  wire  _EVAL_2368;
  wire [8:0] _EVAL_478;
  wire [1:0] _EVAL_2358;
  wire [6:0] _EVAL_3313;
  wire [8:0] _EVAL_412;
  wire [8:0] _EVAL_2737;
  wire  _EVAL_3391;
  wire  _EVAL_551;
  wire [63:0] _EVAL_1546;
  wire  _EVAL_1513;
  wire  _EVAL_2207;
  wire  _EVAL_2319;
  wire  _EVAL_1935;
  wire  _EVAL_2792;
  wire  _EVAL_564;
  wire  _EVAL_1866;
  wire  _EVAL_3268;
  wire  _EVAL_1108;
  wire [8:0] _EVAL_1323;
  wire  _EVAL_3241;
  wire [8:0] _EVAL_177;
  wire [4:0] _EVAL_3051;
  wire  _EVAL_1902;
  wire [4:0] _EVAL_2196;
  wire  _EVAL_2864;
  wire  _EVAL_2558;
  wire  _EVAL_1904;
  wire  _EVAL_1022;
  wire  _EVAL_463;
  wire  _EVAL_2638;
  wire  _EVAL_3120;
  wire  _EVAL_1462;
  wire [10:0] _EVAL_3343;
  wire [10:0] _EVAL_1474;
  wire [138:0] _EVAL_599;
  wire [138:0] _EVAL_1180;
  wire [138:0] _EVAL_2732;
  wire [135:0] _EVAL_246;
  wire [7:0] _EVAL_2619;
  wire [2:0] _EVAL_1765;
  wire  _EVAL_2226;
  wire  _EVAL_1784;
  wire  _EVAL_3042;
  wire  _EVAL_2361;
  wire  _EVAL_1171;
  wire  _EVAL_1164;
  wire  _EVAL_3149;
  wire  _EVAL_2962;
  wire  _EVAL_2536;
  wire  _EVAL_455;
  wire  _EVAL_367;
  wire  _EVAL_277;
  wire  _EVAL_2475;
  wire  _EVAL_3291;
  wire  _EVAL_3096;
  wire  _EVAL_1499;
  wire [3:0] _EVAL_1558;
  wire [127:0] _EVAL_2547;
  wire [127:0] _EVAL_452;
  wire [7:0] _EVAL_872;
  wire [119:0] _EVAL_2417;
  wire [127:0] _EVAL_2734;
  wire [127:0] _EVAL_2983;
  wire [15:0] _EVAL_2620;
  wire [111:0] _EVAL_1009;
  wire [127:0] _EVAL_1877;
  wire [127:0] _EVAL_3007;
  wire [31:0] _EVAL_2476;
  wire [95:0] _EVAL_2545;
  wire [127:0] _EVAL_2703;
  wire [127:0] _EVAL_2594;
  wire [63:0] _EVAL_2813;
  wire [63:0] _EVAL_500;
  wire [127:0] _EVAL_533;
  wire  _EVAL_2109;
  wire  _EVAL_3227;
  wire  _EVAL_3315;
  wire  _EVAL_1250;
  wire [5:0] _EVAL_2058;
  wire [11:0] _EVAL_2192;
  wire  _EVAL_1133;
  wire  _EVAL_211;
  wire  _EVAL_825;
  wire [8:0] _EVAL_826;
  wire [7:0] _EVAL_3062;
  wire [63:0] _EVAL_1788;
  wire [7:0] _EVAL_1498;
  wire  _EVAL_2710;
  wire [31:0] _EVAL_1754;
  wire [5:0] _EVAL_1324;
  wire [8:0] _EVAL_424;
  wire  _EVAL_2069;
  wire  _EVAL_2859;
  wire  _EVAL_1911;
  wire  _EVAL_2390;
  wire  _EVAL_2242;
  wire  _EVAL_1619;
  wire  _EVAL_2937;
  wire  _EVAL_2661;
  wire  _EVAL_1982;
  wire  _EVAL_2042;
  wire [25:0] _EVAL_2491;
  wire  _EVAL_1024;
  wire  _EVAL_899;
  wire [10:0] _EVAL_1291;
  wire [8:0] _EVAL_2524;
  wire [7:0] _EVAL_1971;
  wire  _EVAL_3331;
  wire  _EVAL_501;
  wire [3:0] _EVAL_2525;
  wire [3:0] _EVAL_449;
  wire  _EVAL_2708;
  wire  _EVAL_848;
  wire  _EVAL_3010;
  wire [1:0] _EVAL_1216;
  wire  _EVAL_2259;
  wire  _EVAL_1777;
  wire  _EVAL_2027;
  wire [8:0] _EVAL_1391;
  wire [6:0] _EVAL_1321;
  wire [8:0] _EVAL_723;
  wire [3:0] _EVAL_2065;
  wire [4:0] _EVAL_252;
  wire [8:0] _EVAL_205;
  wire  _EVAL_2481;
  wire [4:0] _EVAL_1398;
  wire  _EVAL_406;
  wire  _EVAL_1065;
  wire  _EVAL_497;
  wire  _EVAL_3368;
  wire  _EVAL_1681;
  wire [1:0] _EVAL_2870;
  wire [1:0] _EVAL_2630;
  wire  _EVAL_1741;
  wire [1:0] _EVAL_1048;
  wire  _EVAL_421;
  wire [8:0] _EVAL_1486;
  wire  _EVAL_281;
  wire  _EVAL_1576;
  wire  _EVAL_2007;
  wire  _EVAL_1127;
  wire  _EVAL_3216;
  wire  _EVAL_602;
  wire  _EVAL_926;
  wire  _EVAL_162;
  wire  _EVAL_1625;
  wire  _EVAL_267;
  wire  _EVAL_3309;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [3:0] _EVAL_323;
  wire [8:0] _EVAL_3214;
  wire  _EVAL_2006;
  wire  _EVAL_1874;
  wire  _EVAL_2827;
  wire  _EVAL_2924;
  wire  _EVAL_280;
  wire  _EVAL_1484;
  wire  _EVAL_2694;
  wire  _EVAL_2989;
  wire  _EVAL_1667;
  wire [19:0] _EVAL_2364;
  wire [19:0] _EVAL_588;
  wire  _EVAL_3349;
  wire  _EVAL_743;
  wire  _EVAL_1944;
  wire [4:0] _EVAL_2932;
  wire  _EVAL_1905;
  wire  _EVAL_3205;
  wire  _EVAL_2695;
  wire  _EVAL_3322;
  wire  _EVAL_1608;
  wire [1:0] _EVAL_1298;
  wire [14:0] _EVAL_2648;
  wire [31:0] _EVAL_1941;
  wire [31:0] _EVAL_3164;
  wire [31:0] _EVAL_451;
  wire  _EVAL_2124;
  wire  _EVAL_2455;
  wire [28:0] _EVAL_688;
  wire [8:0] _EVAL_869;
  wire [17:0] _EVAL_1820;
  wire [26:0] _EVAL_3353;
  wire [8:0] _EVAL_1416;
  wire [1:0] _EVAL_752;
  wire [6:0] _EVAL_1493;
  wire [8:0] _EVAL_1000;
  wire  _EVAL_359;
  wire  _EVAL_2750;
  wire  _EVAL_633;
  wire  _EVAL_986;
  wire  _EVAL_2811;
  wire [8:0] _EVAL_652;
  wire  _EVAL_1422;
  wire [7:0] _EVAL_486;
  wire [8:0] _EVAL_1597;
  wire [6:0] _EVAL_2195;
  wire [8:0] _EVAL_3150;
  wire [8:0] _EVAL_574;
  wire [5:0] _EVAL_1015;
  wire [8:0] _EVAL_1166;
  wire [8:0] _EVAL_775;
  wire [8:0] _EVAL_3366;
  wire [11:0] _EVAL_3397;
  wire [8:0] _EVAL_3310;
  wire  _EVAL_2300;
  wire  _EVAL_3375;
  wire  _EVAL_2639;
  wire  _EVAL_1231;
  wire  _EVAL_806;
  wire [8:0] _EVAL_2565;
  wire  _EVAL_1179;
  wire  _EVAL_1393;
  wire [127:0] _EVAL_1871;
  wire [125:0] _EVAL_1809;
  wire  _EVAL_1473;
  wire  _EVAL_1568;
  wire [3:0] _EVAL_2324;
  wire [7:0] _EVAL_2600;
  wire [7:0] _EVAL_2116;
  wire [7:0] _EVAL_3256;
  wire [7:0] _EVAL_3350;
  wire  _EVAL_3091;
  wire [13:0] _EVAL_353;
  wire  _EVAL_3108;
  wire  _EVAL_3111;
  wire  _EVAL_2998;
  wire  _EVAL_2856;
  wire  _EVAL_1347;
  wire  _EVAL_3371;
  wire [63:0] _EVAL_2506;
  wire  _EVAL_2912;
  wire [4:0] _EVAL_2628;
  wire  _EVAL_2632;
  wire  _EVAL_1464;
  wire  _EVAL_978;
  wire  _EVAL_1675;
  wire  _EVAL_2842;
  wire [1:0] _EVAL_2722;
  wire [1:0] _EVAL_886;
  wire [13:0] _EVAL_1395;
  wire  _EVAL_1623;
  wire [1:0] _EVAL_663;
  wire [31:0] _EVAL_2371;
  wire [13:0] _EVAL_1587;
  wire [13:0] _EVAL_2459;
  wire  _EVAL_2072;
  wire  _EVAL_1086;
  wire [1:0] _EVAL_714;
  wire [1:0] _EVAL_2117;
  wire [31:0] _EVAL_1013;
  wire [63:0] _EVAL_2011;
  wire [63:0] _EVAL_823;
  wire  _EVAL_1594;
  wire  _EVAL_2990;
  wire  _EVAL_202;
  wire [8:0] _EVAL_1951;
  wire [6:0] _EVAL_2841;
  wire [1:0] _EVAL_1912;
  wire [8:0] _EVAL_3158;
  wire [8:0] _EVAL_2470;
  wire [13:0] _EVAL_2680;
  wire  _EVAL_2691;
  wire  _EVAL_1881;
  wire [1:0] _EVAL_1671;
  wire [1:0] _EVAL_1101;
  wire [13:0] _EVAL_1918;
  wire [2:0] _EVAL_1064;
  wire  _EVAL_1251;
  wire  _EVAL_2318;
  wire [1:0] _EVAL_2469;
  wire [1:0] _EVAL_1451;
  wire [31:0] _EVAL_747;
  wire [63:0] _EVAL_3269;
  wire [7:0] _EVAL_2471;
  wire  _EVAL_1304;
  wire  _EVAL_1560;
  wire [2:0] _EVAL_2670;
  wire [8:0] _EVAL_2169;
  wire [8:0] _EVAL_2735;
  wire [3:0] _EVAL_2812;
  wire [4:0] _EVAL_3199;
  wire [8:0] _EVAL_440;
  wire [8:0] _EVAL_1033;
  wire [3:0] _EVAL_1884;
  wire [8:0] _EVAL_1723;
  wire [8:0] _EVAL_2838;
  wire [8:0] _EVAL_1446;
  wire [5:0] _EVAL_2473;
  wire [2:0] _EVAL_2769;
  wire [8:0] _EVAL_2883;
  wire [8:0] _EVAL_1950;
  wire [8:0] _EVAL_802;
  wire [6:0] _EVAL_887;
  wire [255:0] _EVAL_1775;
  wire  _EVAL_2329;
  wire  _EVAL_2679;
  wire  _EVAL_1737;
  wire  _EVAL_225;
  wire  _EVAL_603;
  wire  _EVAL_1872;
  wire  _EVAL_3125;
  wire  _EVAL_2770;
  wire  _EVAL_2311;
  wire  _EVAL_2128;
  wire  _EVAL_457;
  wire  _EVAL_2715;
  wire [3:0] _EVAL_1875;
  wire [3:0] _EVAL_3195;
  wire [7:0] _EVAL_2920;
  wire [255:0] _EVAL_1378;
  wire  _EVAL_1624;
  wire [8:0] _EVAL_1958;
  wire [3:0] _EVAL_410;
  wire [4:0] _EVAL_661;
  wire [8:0] _EVAL_422;
  wire [8:0] _EVAL_2094;
  wire [8:0] _EVAL_2577;
  wire  _EVAL_1392;
  wire  _EVAL_186;
  wire  _EVAL_2946;
  wire  _EVAL_1970;
  wire  _EVAL_3101;
  wire [8:0] _EVAL_1707;
  wire [8:0] _EVAL_2780;
  wire [2:0] _EVAL_3330;
  wire [5:0] _EVAL_2086;
  wire [8:0] _EVAL_212;
  wire [8:0] _EVAL_742;
  wire [4:0] _EVAL_2699;
  wire  _EVAL_3131;
  wire  _EVAL_2033;
  wire  _EVAL_2869;
  wire  _EVAL_1409;
  wire  _EVAL_1740;
  wire [28:0] _EVAL_871;
  wire [2:0] _EVAL_2110;
  wire [7:0] _EVAL_3074;
  wire  _EVAL_1296;
  wire  _EVAL_2497;
  wire  _EVAL_908;
  wire  _EVAL_510;
  wire  _EVAL_2381;
  wire  _EVAL_1322;
  wire  _EVAL_2752;
  wire  _EVAL_762;
  wire  _EVAL_2315;
  wire  _EVAL_2246;
  wire  _EVAL_1196;
  wire  _EVAL_1850;
  wire  _EVAL_2901;
  wire [8:0] _EVAL_596;
  wire  _EVAL_3037;
  wire  _EVAL_1586;
  wire [8:0] _EVAL_1302;
  wire  _EVAL_2089;
  wire [13:0] _EVAL_3145;
  wire  _EVAL_897;
  wire [2:0] _EVAL_2836;
  wire [2:0] _EVAL_1744;
  wire [2:0] _EVAL_2096;
  wire  _EVAL_1334;
  wire  _EVAL_351;
  wire  _EVAL_789;
  wire  _EVAL_969;
  wire  _EVAL_673;
  wire  _EVAL_807;
  wire  _EVAL_967;
  wire  _EVAL_1314;
  wire  _EVAL_627;
  wire  _EVAL_1385;
  wire  _EVAL_704;
  wire  _EVAL_2214;
  wire  _EVAL_2637;
  wire  _EVAL_1043;
  wire  _EVAL_232;
  wire  _EVAL_2213;
  wire  _EVAL_2763;
  wire  _EVAL_209;
  wire  _EVAL_1701;
  wire [1:0] _EVAL_987;
  wire  _EVAL_471;
  wire  _EVAL_2249;
  wire  _EVAL_1548;
  wire  _EVAL_3229;
  wire  _EVAL_1842;
  wire [4:0] _EVAL_390;
  wire  _EVAL_1074;
  wire [31:0] _EVAL_1795;
  wire [31:0] _EVAL_544;
  wire  _EVAL_1949;
  wire [7:0] _EVAL_1381;
  wire [255:0] _EVAL_3065;
  wire  _EVAL_1764;
  wire [20:0] _EVAL_2098;
  wire [19:0] _EVAL_1865;
  wire  _EVAL_1417;
  wire  _EVAL_1811;
  wire  _EVAL_2978;
  wire  _EVAL_3280;
  wire  _EVAL_354;
  wire  _EVAL_3365;
  wire [6:0] _EVAL_776;
  wire [255:0] _EVAL_921;
  wire  _EVAL_2243;
  wire [20:0] _EVAL_2939;
  wire [19:0] _EVAL_334;
  wire  _EVAL_3357;
  wire  _EVAL_1088;
  wire  _EVAL_1985;
  wire  _EVAL_2505;
  wire [4:0] _EVAL_991;
  wire [2:0] _EVAL_3140;
  wire [5:0] _EVAL_401;
  wire [8:0] _EVAL_1722;
  wire [8:0] _EVAL_2984;
  wire [3:0] _EVAL_3228;
  wire [8:0] _EVAL_1030;
  wire [8:0] _EVAL_2201;
  wire [8:0] _EVAL_2926;
  wire  _EVAL_1999;
  wire [1:0] _EVAL_1247;
  wire [30:0] _EVAL_1555;
  wire [31:0] _EVAL_3253;
  wire [8:0] _EVAL_2555;
  wire [2:0] _EVAL_674;
  wire [5:0] _EVAL_3086;
  wire [8:0] _EVAL_1449;
  wire [8:0] _EVAL_1005;
  wire [8:0] _EVAL_482;
  wire [3:0] _EVAL_585;
  wire [4:0] _EVAL_1316;
  wire [8:0] _EVAL_340;
  wire [8:0] _EVAL_3354;
  wire [7:0] _EVAL_1207;
  wire [8:0] _EVAL_294;
  wire [8:0] _EVAL_1757;
  wire  _EVAL_669;
  wire  _EVAL_610;
  wire  _EVAL_3046;
  wire  _EVAL_1531;
  wire  _EVAL_1812;
  wire  _EVAL_2976;
  wire [255:0] _EVAL_488;
  wire [255:0] _EVAL_285;
  wire [255:0] _EVAL_1802;
  wire [255:0] _EVAL_1406;
  wire [255:0] _EVAL_734;
  wire  _EVAL_2889;
  wire  _EVAL_317;
  wire  _EVAL_595;
  wire [63:0] _EVAL_701;
  wire  _EVAL_985;
  wire  _EVAL_2457;
  wire  _EVAL_2720;
  wire  _EVAL_3165;
  wire  _EVAL_1693;
  wire  _EVAL_2961;
  wire  _EVAL_3254;
  wire  _EVAL_2057;
  wire [8:0] _EVAL_3222;
  wire  _EVAL_1337;
  wire [7:0] _EVAL_1704;
  wire  _EVAL_2265;
  wire  _EVAL_718;
  wire [3:0] _EVAL_3300;
  wire [3:0] _EVAL_1606;
  wire  _EVAL_2987;
  wire  _EVAL_2669;
  wire  _EVAL_799;
  wire  _EVAL_801;
  wire  _EVAL_2395;
  wire  _EVAL_2982;
  wire  _EVAL_630;
  wire  _EVAL_1341;
  wire [1:0] _EVAL_558;
  wire  _EVAL_1601;
  wire  _EVAL_1265;
  wire  _EVAL_2322;
  wire  _EVAL_980;
  wire  _EVAL_3359;
  wire  _EVAL_2203;
  wire  _EVAL_1194;
  wire  _EVAL_3362;
  wire  _EVAL_1339;
  wire  _EVAL_3190;
  wire [7:0] _EVAL_3298;
  wire [8:0] _EVAL_3374;
  wire [2:0] _EVAL_1703;
  wire  _EVAL_2772;
  wire  _EVAL_1191;
  wire  _EVAL_795;
  wire [7:0] _EVAL_2379;
  wire [7:0] _EVAL_507;
  wire [6:0] _EVAL_2461;
  wire [8:0] _EVAL_2206;
  wire [1:0] _EVAL_2449;
  wire  _EVAL_1182;
  wire  _EVAL_1319;
  wire  _EVAL_685;
  wire  _EVAL_1776;
  wire  _EVAL_425;
  wire  _EVAL_2004;
  wire  _EVAL_662;
  wire  _EVAL_2906;
  wire [1:0] _EVAL_2501;
  wire  _EVAL_2017;
  wire  _EVAL_1254;
  wire  _EVAL_1472;
  wire  _EVAL_345;
  wire [1:0] _EVAL_1401;
  wire [1:0] _EVAL_1246;
  wire [7:0] _EVAL_1849;
  wire [6:0] _EVAL_1055;
  wire [2:0] _EVAL_2884;
  wire  _EVAL_1223;
  wire  _EVAL_2308;
  wire [2:0] _EVAL_459;
  wire [10:0] _EVAL_940;
  wire [10:0] _EVAL_1034;
  wire  _EVAL_2386;
  wire  _EVAL_592;
  wire [13:0] _EVAL_1747;
  wire [1:0] _EVAL_1710;
  wire [31:0] _EVAL_1992;
  wire  _EVAL_337;
  wire  _EVAL_1132;
  wire  _EVAL_1477;
  wire  _EVAL_905;
  wire  _EVAL_3273;
  wire  _EVAL_3174;
  wire  _EVAL_1080;
  wire  _EVAL_173;
  wire  _EVAL_411;
  wire [6:0] _EVAL_1485;
  wire [1:0] _EVAL_370;
  wire [8:0] _EVAL_3147;
  wire [8:0] _EVAL_2855;
  wire [7:0] _EVAL_1092;
  wire  _EVAL_1920;
  wire [8:0] _EVAL_2527;
  wire [8:0] _EVAL_1943;
  wire [8:0] _EVAL_330;
  wire [8:0] _EVAL_1293;
  wire [25:0] _EVAL_2861;
  wire [31:0] _EVAL_1942;
  wire  _EVAL_2586;
  wire  _EVAL_2126;
  wire  _EVAL_3104;
  wire  _EVAL_1512;
  wire [31:0] _EVAL_1333;
  wire [31:0] _EVAL_2113;
  wire [31:0] _EVAL_1061;
  wire  _EVAL_774;
  wire  _EVAL_2280;
  wire  _EVAL_890;
  wire  _EVAL_1509;
  wire  _EVAL_1258;
  wire [8:0] _EVAL_2489;
  wire [2:0] _EVAL_383;
  wire  _EVAL_392;
  wire  _EVAL_2908;
  wire [11:0] _EVAL_1228;
  wire [7:0] _EVAL_385;
  wire  _EVAL_2123;
  wire  _EVAL_1201;
  wire  _EVAL_2858;
  wire [31:0] _EVAL_1615;
  wire [127:0] _EVAL_2963;
  wire [138:0] _EVAL_582;
  wire [138:0] _EVAL_3182;
  wire [138:0] _EVAL_2409;
  wire [135:0] _EVAL_171;
  wire [7:0] _EVAL_2526;
  wire  _EVAL_198;
  wire  _EVAL_1646;
  wire  _EVAL_2429;
  wire  _EVAL_1229;
  wire  _EVAL_3392;
  wire  _EVAL_600;
  wire [5:0] _EVAL_702;
  wire [8:0] _EVAL_679;
  wire [8:0] _EVAL_2408;
  wire  _EVAL_3383;
  wire  _EVAL_1900;
  wire  _EVAL_3052;
  wire [8:0] _EVAL_1726;
  wire [5:0] _EVAL_2656;
  wire  _EVAL_765;
  wire  _EVAL_448;
  wire [6:0] _EVAL_2026;
  wire [127:0] _EVAL_1135;
  wire  _EVAL_2153;
  wire  _EVAL_2759;
  wire  _EVAL_283;
  wire  _EVAL_3170;
  wire  _EVAL_873;
  wire  _EVAL_1107;
  wire  _EVAL_824;
  wire  _EVAL_1264;
  wire [8:0] _EVAL_2647;
  wire [19:0] _EVAL_643;
  wire [2:0] _EVAL_328;
  wire [2:0] _EVAL_1017;
  wire [2:0] _EVAL_974;
  wire [2:0] _EVAL_3085;
  wire [2:0] _EVAL_2127;
  wire [2:0] _EVAL_1480;
  wire [2:0] _EVAL_1713;
  wire  _EVAL_1845;
  wire  _EVAL_910;
  wire [8:0] _EVAL_784;
  wire [6:0] _EVAL_2634;
  wire [1:0] _EVAL_1505;
  wire [8:0] _EVAL_327;
  wire [8:0] _EVAL_2952;
  wire [8:0] _EVAL_2624;
  wire [8:0] _EVAL_1084;
  wire [8:0] _EVAL_3175;
  wire [8:0] _EVAL_1349;
  wire [11:0] _EVAL_1253;
  wire  _EVAL_1532;
  wire  _EVAL_382;
  wire  _EVAL_1320;
  wire [13:0] _EVAL_434;
  wire [2:0] _EVAL_2764;
  wire  _EVAL_2305;
  wire  _EVAL_971;
  wire [2:0] _EVAL_301;
  wire [2:0] _EVAL_426;
  wire  _EVAL_1738;
  wire  _EVAL_2104;
  wire  _EVAL_1789;
  wire  _EVAL_2019;
  wire  _EVAL_1819;
  wire [2:0] _EVAL_1541;
  wire [2:0] _EVAL_1914;
  wire [2:0] _EVAL_2222;
  wire  _EVAL_1450;
  wire  _EVAL_924;
  wire [5:0] _EVAL_3118;
  wire  _EVAL_988;
  wire  _EVAL_2850;
  wire  _EVAL_1656;
  wire  _EVAL_3390;
  wire [2:0] _EVAL_2914;
  wire [8:0] _EVAL_2022;
  wire  _EVAL_1840;
  wire [7:0] _EVAL_1364;
  wire [8:0] _EVAL_2302;
  wire [8:0] _EVAL_2532;
  wire  _EVAL_2460;
  wire  _EVAL_1267;
  wire  _EVAL_2654;
  wire  _EVAL_3355;
  wire [2:0] _EVAL_151;
  wire  _EVAL_1835;
  wire  _EVAL_195;
  wire  _EVAL_2684;
  wire [8:0] _EVAL_2598;
  wire [5:0] _EVAL_640;
  wire [2:0] _EVAL_1438;
  wire [3:0] _EVAL_2548;
  wire  _EVAL_2091;
  wire [31:0] _EVAL_3148;
  wire [8:0] _EVAL_1053;
  wire [8:0] _EVAL_2800;
  wire [8:0] _EVAL_2955;
  wire [8:0] _EVAL_692;
  wire [8:0] _EVAL_2456;
  wire [2:0] _EVAL_435;
  wire [8:0] _EVAL_1906;
  wire [8:0] _EVAL_2428;
  wire [31:0] _EVAL_1674;
  wire  _EVAL_2234;
  wire  _EVAL_2494;
  wire [8:0] _EVAL_1285;
  wire [1:0] _EVAL_3226;
  wire  _EVAL_1650;
  wire  _EVAL_1890;
  wire  _EVAL_2674;
  wire  _EVAL_2667;
  wire  _EVAL_1351;
  wire  _EVAL_800;
  wire  _EVAL_1770;
  wire  _EVAL_263;
  wire  _EVAL_2517;
  wire  _EVAL_911;
  wire  _EVAL_677;
  wire [63:0] _EVAL_458;
  wire [7:0] _EVAL_3271;
  wire [63:0] _EVAL_1198;
  wire [63:0] _EVAL_1153;
  wire  _EVAL_1530;
  wire  _EVAL_398;
  wire [63:0] _EVAL_2784;
  wire [7:0] _EVAL_1124;
  wire  _EVAL_2310;
  wire  _EVAL_224;
  wire [2:0] _EVAL_2346;
  wire  _EVAL_1590;
  wire [2:0] _EVAL_1571;
  wire [2:0] _EVAL_1903;
  wire  _EVAL_2753;
  wire  _EVAL_3235;
  wire [6:0] _EVAL_1150;
  wire [8:0] _EVAL_891;
  wire [5:0] _EVAL_3073;
  wire [8:0] _EVAL_1012;
  wire [8:0] _EVAL_508;
  wire [3:0] _EVAL_2953;
  wire [4:0] _EVAL_447;
  wire [8:0] _EVAL_1225;
  wire [8:0] _EVAL_852;
  wire  _EVAL_2696;
  wire  _EVAL_1286;
  wire  _EVAL_2665;
  wire  _EVAL_1833;
  wire [31:0] _EVAL_1329;
  wire  _EVAL_2627;
  wire [7:0] _EVAL_2372;
  wire [7:0] _EVAL_2919;
  wire  _EVAL_2228;
  wire  _EVAL_3103;
  wire  _EVAL_2502;
  wire  _EVAL_1212;
  wire [2:0] _EVAL_1360;
  wire [2:0] _EVAL_483;
  wire  _EVAL_409;
  wire [13:0] _EVAL_1573;
  wire  _EVAL_668;
  wire [127:0] _EVAL_1156;
  wire  _EVAL_291;
  wire  _EVAL_1620;
  wire  _EVAL_2247;
  wire  _EVAL_675;
  wire  _EVAL_3176;
  wire  _EVAL_1852;
  wire  _EVAL_1542;
  wire  _EVAL_1020;
  wire [1:0] _EVAL_877;
  wire [8:0] _EVAL_2786;
  wire  _EVAL_2682;
  wire  _EVAL_2793;
  wire [6:0] _EVAL_3249;
  wire [127:0] _EVAL_1730;
  wire [8:0] _EVAL_1046;
  wire [8:0] _EVAL_2917;
  wire [7:0] _EVAL_1832;
  wire  _EVAL_1702;
  wire  _EVAL_3078;
  wire [63:0] _EVAL_559;
  wire [7:0] _EVAL_2209;
  wire [63:0] _EVAL_964;
  wire  _EVAL_1287;
  wire  _EVAL_2141;
  wire [2:0] _EVAL_1389;
  wire [31:0] _EVAL_1040;
  wire  _EVAL_2076;
  wire [8:0] _EVAL_2438;
  wire  _EVAL_1072;
  wire  _EVAL_2401;
  wire [1:0] _EVAL_1284;
  wire [8:0] _EVAL_2589;
  wire [127:0] _EVAL_167;
  wire [127:0] _EVAL_1666;
  wire [127:0] _EVAL_2225;
  wire  _EVAL_1724;
  wire [24:0] _EVAL_2215;
  wire [31:0] _EVAL_1112;
  wire  _EVAL_1919;
  wire  _EVAL_2374;
  wire  _EVAL_3305;
  wire [2:0] _EVAL_2942;
  wire [8:0] _EVAL_480;
  wire [6:0] _EVAL_207;
  wire [8:0] _EVAL_498;
  wire [8:0] _EVAL_2357;
  wire [8:0] _EVAL_1699;
  wire [8:0] _EVAL_2802;
  wire [11:0] _EVAL_1792;
  wire  _EVAL_579;
  wire [2:0] _EVAL_2483;
  wire  _EVAL_3202;
  wire  _EVAL_557;
  wire  _EVAL_3367;
  wire [19:0] _EVAL_608;
  wire [31:0] _EVAL_443;
  wire  _EVAL_3246;
  wire  _EVAL_1563;
  wire  _EVAL_2820;
  wire [8:0] _EVAL_3224;
  wire [13:0] _EVAL_3385;
  wire [63:0] _EVAL_539;
  wire  _EVAL_1647;
  wire  _EVAL_1181;
  wire [1:0] _EVAL_838;
  wire  _EVAL_918;
  wire [8:0] _EVAL_2923;
  wire [1:0] _EVAL_732;
  wire  _EVAL_2685;
  wire [11:0] _EVAL_379;
  wire  _EVAL_1338;
  wire  _EVAL_3045;
  wire  _EVAL_948;
  wire  _EVAL_218;
  wire  _EVAL_992;
  wire [13:0] _EVAL_1869;
  wire [1:0] _EVAL_1452;
  wire [31:0] _EVAL_3252;
  wire [8:0] _EVAL_2340;
  wire  _EVAL_1326;
  wire  _EVAL_1447;
  wire [7:0] _EVAL_262;
  wire  _EVAL_923;
  wire  _EVAL_1609;
  wire [127:0] _EVAL_292;
  wire [127:0] _EVAL_1380;
  wire [7:0] _EVAL_154;
  wire [2:0] _EVAL_3306;
  wire  _EVAL_2862;
  wire  _EVAL_1506;
  wire  _EVAL_537;
  wire [1:0] _EVAL_840;
  wire [31:0] _EVAL_780;
  wire [2:0] _EVAL_3393;
  wire  _EVAL_516;
  wire  _EVAL_634;
  wire  _EVAL_3036;
  wire [31:0] _EVAL_593;
  wire [31:0] _EVAL_570;
  wire [1:0] _EVAL_821;
  wire  _EVAL_1814;
  wire  _EVAL_1660;
  wire  _EVAL_1637;
  wire  _EVAL_2354;
  wire  _EVAL_1801;
  wire [14:0] _EVAL_2776;
  wire [14:0] _EVAL_545;
  wire [2:0] _EVAL_2956;
  wire  _EVAL_642;
  wire [1:0] _EVAL_1600;
  wire [127:0] _EVAL_2118;
  wire  _EVAL_2445;
  wire  _EVAL_1454;
  wire  _EVAL_2587;
  wire  _EVAL_1429;
  wire  _EVAL_1348;
  wire  _EVAL_2416;
  wire  _EVAL_3194;
  wire  _EVAL_3134;
  wire  _EVAL_2021;
  wire  _EVAL_3160;
  wire [8:0] _EVAL_3243;
  wire  _EVAL_2513;
  wire  _EVAL_1761;
  wire [1:0] _EVAL_1047;
  wire  _EVAL_681;
  wire  _EVAL_3328;
  wire  _EVAL_772;
  wire [15:0] _EVAL_2509;
  wire [8:0] _EVAL_2522;
  wire [14:0] _EVAL_1838;
  wire  _EVAL_2348;
  wire  _EVAL_952;
  wire  _EVAL_909;
  wire  _EVAL_828;
  wire  _EVAL_2643;
  wire  _EVAL_2847;
  wire  _EVAL_1003;
  wire  _EVAL_3124;
  wire [31:0] _EVAL_2651;
  wire [127:0] _EVAL_2873;
  wire  _EVAL_812;
  wire  _EVAL_1574;
  wire  _EVAL_438;
  wire  _EVAL_505;
  wire  _EVAL_2034;
  wire  _EVAL_1521;
  wire  _EVAL_361;
  wire  _EVAL_3024;
  wire [127:0] _EVAL_1843;
  wire [6:0] _EVAL_3279;
  wire [6:0] _EVAL_415;
  wire  _EVAL_2298;
  wire [127:0] _EVAL_2562;
  wire [8:0] _EVAL_1745;
  wire  _EVAL_2421;
  wire [2:0] _EVAL_2731;
  wire [8:0] _EVAL_509;
  wire [14:0] _EVAL_3339;
  wire [14:0] _EVAL_1457;
  wire  _EVAL_2055;
  wire [31:0] _EVAL_3403;
  wire  _EVAL_1408;
  wire  _EVAL_2945;
  wire  _EVAL_2819;
  wire  _EVAL_2435;
  wire  _EVAL_893;
  wire  _EVAL_2488;
  wire  _EVAL_1239;
  wire  _EVAL_736;
  wire  _EVAL_612;
  wire  _EVAL_2611;
  wire  _EVAL_2830;
  wire [8:0] _EVAL_631;
  wire  _EVAL_1690;
  wire  _EVAL_208;
  wire  _EVAL_1470;
  wire  _EVAL_2102;
  wire [8:0] _EVAL_3077;
  wire [8:0] _EVAL_526;
  wire [11:0] _EVAL_2844;
  wire  _EVAL_1892;
  wire [2:0] _EVAL_597;
  wire [2:0] _EVAL_2313;
  wire [11:0] _EVAL_2362;
  wire  _EVAL_793;
  wire  _EVAL_611;
  SiFive__EVAL_233 packageanon1_3 (
    ._EVAL(packageanon1_3__EVAL),
    ._EVAL_0(packageanon1_3__EVAL_0)
  );
  SiFive__EVAL_233 packageanon1_5 (
    ._EVAL(packageanon1_5__EVAL),
    ._EVAL_0(packageanon1_5__EVAL_0)
  );
  SiFive__EVAL_340 data_arrays_3_0 (
    ._EVAL(data_arrays_3_0__EVAL),
    ._EVAL_0(data_arrays_3_0__EVAL_0),
    ._EVAL_1(data_arrays_3_0__EVAL_1),
    ._EVAL_2(data_arrays_3_0__EVAL_2),
    ._EVAL_3(data_arrays_3_0__EVAL_3),
    ._EVAL_4(data_arrays_3_0__EVAL_4)
  );
  SiFive__EVAL_340 data_arrays_2_1 (
    ._EVAL(data_arrays_2_1__EVAL),
    ._EVAL_0(data_arrays_2_1__EVAL_0),
    ._EVAL_1(data_arrays_2_1__EVAL_1),
    ._EVAL_2(data_arrays_2_1__EVAL_2),
    ._EVAL_3(data_arrays_2_1__EVAL_3),
    ._EVAL_4(data_arrays_2_1__EVAL_4)
  );
  SiFive__EVAL_340 data_arrays_1_0 (
    ._EVAL(data_arrays_1_0__EVAL),
    ._EVAL_0(data_arrays_1_0__EVAL_0),
    ._EVAL_1(data_arrays_1_0__EVAL_1),
    ._EVAL_2(data_arrays_1_0__EVAL_2),
    ._EVAL_3(data_arrays_1_0__EVAL_3),
    ._EVAL_4(data_arrays_1_0__EVAL_4)
  );
  SiFive__EVAL_340 data_arrays_2_0 (
    ._EVAL(data_arrays_2_0__EVAL),
    ._EVAL_0(data_arrays_2_0__EVAL_0),
    ._EVAL_1(data_arrays_2_0__EVAL_1),
    ._EVAL_2(data_arrays_2_0__EVAL_2),
    ._EVAL_3(data_arrays_2_0__EVAL_3),
    ._EVAL_4(data_arrays_2_0__EVAL_4)
  );
  SiFive__EVAL_233 packageanon1_7 (
    ._EVAL(packageanon1_7__EVAL),
    ._EVAL_0(packageanon1_7__EVAL_0)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR_1 (
    ._EVAL(MaxPeriodFibonacciLFSR_1__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR_1__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR_1__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR_1__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR_1__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR_1__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR_1__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR_1__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR_1__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR_1__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR_1__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR_1__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR_1__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR_1__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR_1__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR_1__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR_1__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR_1__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR_1__EVAL_17)
  );
  SiFive__EVAL_338 predictor_tagged_tables_2 (
    ._EVAL(predictor_tagged_tables_2__EVAL),
    ._EVAL_0(predictor_tagged_tables_2__EVAL_0),
    ._EVAL_1(predictor_tagged_tables_2__EVAL_1),
    ._EVAL_2(predictor_tagged_tables_2__EVAL_2),
    ._EVAL_3(predictor_tagged_tables_2__EVAL_3),
    ._EVAL_4(predictor_tagged_tables_2__EVAL_4),
    ._EVAL_5(predictor_tagged_tables_2__EVAL_5),
    ._EVAL_6(predictor_tagged_tables_2__EVAL_6),
    ._EVAL_7(predictor_tagged_tables_2__EVAL_7),
    ._EVAL_8(predictor_tagged_tables_2__EVAL_8),
    ._EVAL_9(predictor_tagged_tables_2__EVAL_9),
    ._EVAL_10(predictor_tagged_tables_2__EVAL_10),
    ._EVAL_11(predictor_tagged_tables_2__EVAL_11),
    ._EVAL_12(predictor_tagged_tables_2__EVAL_12),
    ._EVAL_13(predictor_tagged_tables_2__EVAL_13),
    ._EVAL_14(predictor_tagged_tables_2__EVAL_14),
    ._EVAL_15(predictor_tagged_tables_2__EVAL_15),
    ._EVAL_16(predictor_tagged_tables_2__EVAL_16),
    ._EVAL_17(predictor_tagged_tables_2__EVAL_17),
    ._EVAL_18(predictor_tagged_tables_2__EVAL_18),
    ._EVAL_19(predictor_tagged_tables_2__EVAL_19),
    ._EVAL_20(predictor_tagged_tables_2__EVAL_20),
    ._EVAL_21(predictor_tagged_tables_2__EVAL_21),
    ._EVAL_22(predictor_tagged_tables_2__EVAL_22),
    ._EVAL_23(predictor_tagged_tables_2__EVAL_23),
    ._EVAL_24(predictor_tagged_tables_2__EVAL_24),
    ._EVAL_25(predictor_tagged_tables_2__EVAL_25),
    ._EVAL_26(predictor_tagged_tables_2__EVAL_26),
    ._EVAL_27(predictor_tagged_tables_2__EVAL_27),
    ._EVAL_28(predictor_tagged_tables_2__EVAL_28),
    ._EVAL_29(predictor_tagged_tables_2__EVAL_29),
    ._EVAL_30(predictor_tagged_tables_2__EVAL_30),
    ._EVAL_31(predictor_tagged_tables_2__EVAL_31),
    ._EVAL_32(predictor_tagged_tables_2__EVAL_32),
    ._EVAL_33(predictor_tagged_tables_2__EVAL_33),
    ._EVAL_34(predictor_tagged_tables_2__EVAL_34),
    ._EVAL_35(predictor_tagged_tables_2__EVAL_35),
    ._EVAL_36(predictor_tagged_tables_2__EVAL_36),
    ._EVAL_37(predictor_tagged_tables_2__EVAL_37),
    ._EVAL_38(predictor_tagged_tables_2__EVAL_38)
  );
  SiFive__EVAL_338 predictor_tagged_tables_1 (
    ._EVAL(predictor_tagged_tables_1__EVAL),
    ._EVAL_0(predictor_tagged_tables_1__EVAL_0),
    ._EVAL_1(predictor_tagged_tables_1__EVAL_1),
    ._EVAL_2(predictor_tagged_tables_1__EVAL_2),
    ._EVAL_3(predictor_tagged_tables_1__EVAL_3),
    ._EVAL_4(predictor_tagged_tables_1__EVAL_4),
    ._EVAL_5(predictor_tagged_tables_1__EVAL_5),
    ._EVAL_6(predictor_tagged_tables_1__EVAL_6),
    ._EVAL_7(predictor_tagged_tables_1__EVAL_7),
    ._EVAL_8(predictor_tagged_tables_1__EVAL_8),
    ._EVAL_9(predictor_tagged_tables_1__EVAL_9),
    ._EVAL_10(predictor_tagged_tables_1__EVAL_10),
    ._EVAL_11(predictor_tagged_tables_1__EVAL_11),
    ._EVAL_12(predictor_tagged_tables_1__EVAL_12),
    ._EVAL_13(predictor_tagged_tables_1__EVAL_13),
    ._EVAL_14(predictor_tagged_tables_1__EVAL_14),
    ._EVAL_15(predictor_tagged_tables_1__EVAL_15),
    ._EVAL_16(predictor_tagged_tables_1__EVAL_16),
    ._EVAL_17(predictor_tagged_tables_1__EVAL_17),
    ._EVAL_18(predictor_tagged_tables_1__EVAL_18),
    ._EVAL_19(predictor_tagged_tables_1__EVAL_19),
    ._EVAL_20(predictor_tagged_tables_1__EVAL_20),
    ._EVAL_21(predictor_tagged_tables_1__EVAL_21),
    ._EVAL_22(predictor_tagged_tables_1__EVAL_22),
    ._EVAL_23(predictor_tagged_tables_1__EVAL_23),
    ._EVAL_24(predictor_tagged_tables_1__EVAL_24),
    ._EVAL_25(predictor_tagged_tables_1__EVAL_25),
    ._EVAL_26(predictor_tagged_tables_1__EVAL_26),
    ._EVAL_27(predictor_tagged_tables_1__EVAL_27),
    ._EVAL_28(predictor_tagged_tables_1__EVAL_28),
    ._EVAL_29(predictor_tagged_tables_1__EVAL_29),
    ._EVAL_30(predictor_tagged_tables_1__EVAL_30),
    ._EVAL_31(predictor_tagged_tables_1__EVAL_31),
    ._EVAL_32(predictor_tagged_tables_1__EVAL_32),
    ._EVAL_33(predictor_tagged_tables_1__EVAL_33),
    ._EVAL_34(predictor_tagged_tables_1__EVAL_34),
    ._EVAL_35(predictor_tagged_tables_1__EVAL_35),
    ._EVAL_36(predictor_tagged_tables_1__EVAL_36),
    ._EVAL_37(predictor_tagged_tables_1__EVAL_37),
    ._EVAL_38(predictor_tagged_tables_1__EVAL_38)
  );
  EICG_wrapper icache_clock_gate (
    .in(icache_clock_gate_in),
    .en(icache_clock_gate_en),
    .out(icache_clock_gate_out)
  );
  SiFive__EVAL_340 data_arrays_1_1 (
    ._EVAL(data_arrays_1_1__EVAL),
    ._EVAL_0(data_arrays_1_1__EVAL_0),
    ._EVAL_1(data_arrays_1_1__EVAL_1),
    ._EVAL_2(data_arrays_1_1__EVAL_2),
    ._EVAL_3(data_arrays_1_1__EVAL_3),
    ._EVAL_4(data_arrays_1_1__EVAL_4)
  );
  SiFive__EVAL_233 packageanon1_1 (
    ._EVAL(packageanon1_1__EVAL),
    ._EVAL_0(packageanon1_1__EVAL_0)
  );
  SiFive__EVAL_233 packageanon1_2 (
    ._EVAL(packageanon1_2__EVAL),
    ._EVAL_0(packageanon1_2__EVAL_0)
  );
  SiFive__EVAL_338 predictor_tagged_tables_0 (
    ._EVAL(predictor_tagged_tables_0__EVAL),
    ._EVAL_0(predictor_tagged_tables_0__EVAL_0),
    ._EVAL_1(predictor_tagged_tables_0__EVAL_1),
    ._EVAL_2(predictor_tagged_tables_0__EVAL_2),
    ._EVAL_3(predictor_tagged_tables_0__EVAL_3),
    ._EVAL_4(predictor_tagged_tables_0__EVAL_4),
    ._EVAL_5(predictor_tagged_tables_0__EVAL_5),
    ._EVAL_6(predictor_tagged_tables_0__EVAL_6),
    ._EVAL_7(predictor_tagged_tables_0__EVAL_7),
    ._EVAL_8(predictor_tagged_tables_0__EVAL_8),
    ._EVAL_9(predictor_tagged_tables_0__EVAL_9),
    ._EVAL_10(predictor_tagged_tables_0__EVAL_10),
    ._EVAL_11(predictor_tagged_tables_0__EVAL_11),
    ._EVAL_12(predictor_tagged_tables_0__EVAL_12),
    ._EVAL_13(predictor_tagged_tables_0__EVAL_13),
    ._EVAL_14(predictor_tagged_tables_0__EVAL_14),
    ._EVAL_15(predictor_tagged_tables_0__EVAL_15),
    ._EVAL_16(predictor_tagged_tables_0__EVAL_16),
    ._EVAL_17(predictor_tagged_tables_0__EVAL_17),
    ._EVAL_18(predictor_tagged_tables_0__EVAL_18),
    ._EVAL_19(predictor_tagged_tables_0__EVAL_19),
    ._EVAL_20(predictor_tagged_tables_0__EVAL_20),
    ._EVAL_21(predictor_tagged_tables_0__EVAL_21),
    ._EVAL_22(predictor_tagged_tables_0__EVAL_22),
    ._EVAL_23(predictor_tagged_tables_0__EVAL_23),
    ._EVAL_24(predictor_tagged_tables_0__EVAL_24),
    ._EVAL_25(predictor_tagged_tables_0__EVAL_25),
    ._EVAL_26(predictor_tagged_tables_0__EVAL_26),
    ._EVAL_27(predictor_tagged_tables_0__EVAL_27),
    ._EVAL_28(predictor_tagged_tables_0__EVAL_28),
    ._EVAL_29(predictor_tagged_tables_0__EVAL_29),
    ._EVAL_30(predictor_tagged_tables_0__EVAL_30),
    ._EVAL_31(predictor_tagged_tables_0__EVAL_31),
    ._EVAL_32(predictor_tagged_tables_0__EVAL_32),
    ._EVAL_33(predictor_tagged_tables_0__EVAL_33),
    ._EVAL_34(predictor_tagged_tables_0__EVAL_34),
    ._EVAL_35(predictor_tagged_tables_0__EVAL_35),
    ._EVAL_36(predictor_tagged_tables_0__EVAL_36),
    ._EVAL_37(predictor_tagged_tables_0__EVAL_37),
    ._EVAL_38(predictor_tagged_tables_0__EVAL_38)
  );
  SiFive__EVAL_231 predictor_Queue (
    ._EVAL(predictor_Queue__EVAL),
    ._EVAL_0(predictor_Queue__EVAL_0),
    ._EVAL_1(predictor_Queue__EVAL_1),
    ._EVAL_2(predictor_Queue__EVAL_2),
    ._EVAL_3(predictor_Queue__EVAL_3),
    ._EVAL_4(predictor_Queue__EVAL_4),
    ._EVAL_5(predictor_Queue__EVAL_5),
    ._EVAL_6(predictor_Queue__EVAL_6),
    ._EVAL_7(predictor_Queue__EVAL_7),
    ._EVAL_8(predictor_Queue__EVAL_8),
    ._EVAL_9(predictor_Queue__EVAL_9),
    ._EVAL_10(predictor_Queue__EVAL_10),
    ._EVAL_11(predictor_Queue__EVAL_11),
    ._EVAL_12(predictor_Queue__EVAL_12),
    ._EVAL_13(predictor_Queue__EVAL_13),
    ._EVAL_14(predictor_Queue__EVAL_14)
  );
  SiFive__EVAL_233 packageanon1_8 (
    ._EVAL(packageanon1_8__EVAL),
    ._EVAL_0(packageanon1_8__EVAL_0)
  );
  SiFive__EVAL_340 data_arrays_3_1 (
    ._EVAL(data_arrays_3_1__EVAL),
    ._EVAL_0(data_arrays_3_1__EVAL_0),
    ._EVAL_1(data_arrays_3_1__EVAL_1),
    ._EVAL_2(data_arrays_3_1__EVAL_2),
    ._EVAL_3(data_arrays_3_1__EVAL_3),
    ._EVAL_4(data_arrays_3_1__EVAL_4)
  );
  SiFive__EVAL_339 tag_array (
    ._EVAL(tag_array__EVAL),
    ._EVAL_0(tag_array__EVAL_0),
    ._EVAL_1(tag_array__EVAL_1),
    ._EVAL_2(tag_array__EVAL_2),
    ._EVAL_3(tag_array__EVAL_3),
    ._EVAL_4(tag_array__EVAL_4),
    ._EVAL_5(tag_array__EVAL_5),
    ._EVAL_6(tag_array__EVAL_6),
    ._EVAL_7(tag_array__EVAL_7),
    ._EVAL_8(tag_array__EVAL_8),
    ._EVAL_9(tag_array__EVAL_9),
    ._EVAL_10(tag_array__EVAL_10),
    ._EVAL_11(tag_array__EVAL_11),
    ._EVAL_12(tag_array__EVAL_12),
    ._EVAL_13(tag_array__EVAL_13),
    ._EVAL_14(tag_array__EVAL_14)
  );
  SiFive__EVAL_233 packageanon1_6 (
    ._EVAL(packageanon1_6__EVAL),
    ._EVAL_0(packageanon1_6__EVAL_0)
  );
  SiFive__EVAL_340 data_arrays_0_1 (
    ._EVAL(data_arrays_0_1__EVAL),
    ._EVAL_0(data_arrays_0_1__EVAL_0),
    ._EVAL_1(data_arrays_0_1__EVAL_1),
    ._EVAL_2(data_arrays_0_1__EVAL_2),
    ._EVAL_3(data_arrays_0_1__EVAL_3),
    ._EVAL_4(data_arrays_0_1__EVAL_4)
  );
  SiFive__EVAL_337 predictor_base_table_1 (
    ._EVAL(predictor_base_table_1__EVAL),
    ._EVAL_0(predictor_base_table_1__EVAL_0),
    ._EVAL_1(predictor_base_table_1__EVAL_1),
    ._EVAL_2(predictor_base_table_1__EVAL_2),
    ._EVAL_3(predictor_base_table_1__EVAL_3),
    ._EVAL_4(predictor_base_table_1__EVAL_4),
    ._EVAL_5(predictor_base_table_1__EVAL_5),
    ._EVAL_6(predictor_base_table_1__EVAL_6),
    ._EVAL_7(predictor_base_table_1__EVAL_7),
    ._EVAL_8(predictor_base_table_1__EVAL_8),
    ._EVAL_9(predictor_base_table_1__EVAL_9),
    ._EVAL_10(predictor_base_table_1__EVAL_10),
    ._EVAL_11(predictor_base_table_1__EVAL_11),
    ._EVAL_12(predictor_base_table_1__EVAL_12),
    ._EVAL_13(predictor_base_table_1__EVAL_13),
    ._EVAL_14(predictor_base_table_1__EVAL_14),
    ._EVAL_15(predictor_base_table_1__EVAL_15),
    ._EVAL_16(predictor_base_table_1__EVAL_16),
    ._EVAL_17(predictor_base_table_1__EVAL_17),
    ._EVAL_18(predictor_base_table_1__EVAL_18),
    ._EVAL_19(predictor_base_table_1__EVAL_19),
    ._EVAL_20(predictor_base_table_1__EVAL_20),
    ._EVAL_21(predictor_base_table_1__EVAL_21),
    ._EVAL_22(predictor_base_table_1__EVAL_22),
    ._EVAL_23(predictor_base_table_1__EVAL_23),
    ._EVAL_24(predictor_base_table_1__EVAL_24),
    ._EVAL_25(predictor_base_table_1__EVAL_25),
    ._EVAL_26(predictor_base_table_1__EVAL_26),
    ._EVAL_27(predictor_base_table_1__EVAL_27),
    ._EVAL_28(predictor_base_table_1__EVAL_28),
    ._EVAL_29(predictor_base_table_1__EVAL_29)
  );
  SiFive__EVAL_232 MaxPeriodFibonacciLFSR (
    ._EVAL(MaxPeriodFibonacciLFSR__EVAL),
    ._EVAL_0(MaxPeriodFibonacciLFSR__EVAL_0),
    ._EVAL_1(MaxPeriodFibonacciLFSR__EVAL_1),
    ._EVAL_2(MaxPeriodFibonacciLFSR__EVAL_2),
    ._EVAL_3(MaxPeriodFibonacciLFSR__EVAL_3),
    ._EVAL_4(MaxPeriodFibonacciLFSR__EVAL_4),
    ._EVAL_5(MaxPeriodFibonacciLFSR__EVAL_5),
    ._EVAL_6(MaxPeriodFibonacciLFSR__EVAL_6),
    ._EVAL_7(MaxPeriodFibonacciLFSR__EVAL_7),
    ._EVAL_8(MaxPeriodFibonacciLFSR__EVAL_8),
    ._EVAL_9(MaxPeriodFibonacciLFSR__EVAL_9),
    ._EVAL_10(MaxPeriodFibonacciLFSR__EVAL_10),
    ._EVAL_11(MaxPeriodFibonacciLFSR__EVAL_11),
    ._EVAL_12(MaxPeriodFibonacciLFSR__EVAL_12),
    ._EVAL_13(MaxPeriodFibonacciLFSR__EVAL_13),
    ._EVAL_14(MaxPeriodFibonacciLFSR__EVAL_14),
    ._EVAL_15(MaxPeriodFibonacciLFSR__EVAL_15),
    ._EVAL_16(MaxPeriodFibonacciLFSR__EVAL_16),
    ._EVAL_17(MaxPeriodFibonacciLFSR__EVAL_17)
  );
  SiFive__EVAL_338 predictor_tagged_tables_3 (
    ._EVAL(predictor_tagged_tables_3__EVAL),
    ._EVAL_0(predictor_tagged_tables_3__EVAL_0),
    ._EVAL_1(predictor_tagged_tables_3__EVAL_1),
    ._EVAL_2(predictor_tagged_tables_3__EVAL_2),
    ._EVAL_3(predictor_tagged_tables_3__EVAL_3),
    ._EVAL_4(predictor_tagged_tables_3__EVAL_4),
    ._EVAL_5(predictor_tagged_tables_3__EVAL_5),
    ._EVAL_6(predictor_tagged_tables_3__EVAL_6),
    ._EVAL_7(predictor_tagged_tables_3__EVAL_7),
    ._EVAL_8(predictor_tagged_tables_3__EVAL_8),
    ._EVAL_9(predictor_tagged_tables_3__EVAL_9),
    ._EVAL_10(predictor_tagged_tables_3__EVAL_10),
    ._EVAL_11(predictor_tagged_tables_3__EVAL_11),
    ._EVAL_12(predictor_tagged_tables_3__EVAL_12),
    ._EVAL_13(predictor_tagged_tables_3__EVAL_13),
    ._EVAL_14(predictor_tagged_tables_3__EVAL_14),
    ._EVAL_15(predictor_tagged_tables_3__EVAL_15),
    ._EVAL_16(predictor_tagged_tables_3__EVAL_16),
    ._EVAL_17(predictor_tagged_tables_3__EVAL_17),
    ._EVAL_18(predictor_tagged_tables_3__EVAL_18),
    ._EVAL_19(predictor_tagged_tables_3__EVAL_19),
    ._EVAL_20(predictor_tagged_tables_3__EVAL_20),
    ._EVAL_21(predictor_tagged_tables_3__EVAL_21),
    ._EVAL_22(predictor_tagged_tables_3__EVAL_22),
    ._EVAL_23(predictor_tagged_tables_3__EVAL_23),
    ._EVAL_24(predictor_tagged_tables_3__EVAL_24),
    ._EVAL_25(predictor_tagged_tables_3__EVAL_25),
    ._EVAL_26(predictor_tagged_tables_3__EVAL_26),
    ._EVAL_27(predictor_tagged_tables_3__EVAL_27),
    ._EVAL_28(predictor_tagged_tables_3__EVAL_28),
    ._EVAL_29(predictor_tagged_tables_3__EVAL_29),
    ._EVAL_30(predictor_tagged_tables_3__EVAL_30),
    ._EVAL_31(predictor_tagged_tables_3__EVAL_31),
    ._EVAL_32(predictor_tagged_tables_3__EVAL_32),
    ._EVAL_33(predictor_tagged_tables_3__EVAL_33),
    ._EVAL_34(predictor_tagged_tables_3__EVAL_34),
    ._EVAL_35(predictor_tagged_tables_3__EVAL_35),
    ._EVAL_36(predictor_tagged_tables_3__EVAL_36),
    ._EVAL_37(predictor_tagged_tables_3__EVAL_37),
    ._EVAL_38(predictor_tagged_tables_3__EVAL_38)
  );
  SiFive__EVAL_340 data_arrays_0_0 (
    ._EVAL(data_arrays_0_0__EVAL),
    ._EVAL_0(data_arrays_0_0__EVAL_0),
    ._EVAL_1(data_arrays_0_0__EVAL_1),
    ._EVAL_2(data_arrays_0_0__EVAL_2),
    ._EVAL_3(data_arrays_0_0__EVAL_3),
    ._EVAL_4(data_arrays_0_0__EVAL_4)
  );
  SiFive__EVAL_337 predictor_base_table_0 (
    ._EVAL(predictor_base_table_0__EVAL),
    ._EVAL_0(predictor_base_table_0__EVAL_0),
    ._EVAL_1(predictor_base_table_0__EVAL_1),
    ._EVAL_2(predictor_base_table_0__EVAL_2),
    ._EVAL_3(predictor_base_table_0__EVAL_3),
    ._EVAL_4(predictor_base_table_0__EVAL_4),
    ._EVAL_5(predictor_base_table_0__EVAL_5),
    ._EVAL_6(predictor_base_table_0__EVAL_6),
    ._EVAL_7(predictor_base_table_0__EVAL_7),
    ._EVAL_8(predictor_base_table_0__EVAL_8),
    ._EVAL_9(predictor_base_table_0__EVAL_9),
    ._EVAL_10(predictor_base_table_0__EVAL_10),
    ._EVAL_11(predictor_base_table_0__EVAL_11),
    ._EVAL_12(predictor_base_table_0__EVAL_12),
    ._EVAL_13(predictor_base_table_0__EVAL_13),
    ._EVAL_14(predictor_base_table_0__EVAL_14),
    ._EVAL_15(predictor_base_table_0__EVAL_15),
    ._EVAL_16(predictor_base_table_0__EVAL_16),
    ._EVAL_17(predictor_base_table_0__EVAL_17),
    ._EVAL_18(predictor_base_table_0__EVAL_18),
    ._EVAL_19(predictor_base_table_0__EVAL_19),
    ._EVAL_20(predictor_base_table_0__EVAL_20),
    ._EVAL_21(predictor_base_table_0__EVAL_21),
    ._EVAL_22(predictor_base_table_0__EVAL_22),
    ._EVAL_23(predictor_base_table_0__EVAL_23),
    ._EVAL_24(predictor_base_table_0__EVAL_24),
    ._EVAL_25(predictor_base_table_0__EVAL_25),
    ._EVAL_26(predictor_base_table_0__EVAL_26),
    ._EVAL_27(predictor_base_table_0__EVAL_27),
    ._EVAL_28(predictor_base_table_0__EVAL_28),
    ._EVAL_29(predictor_base_table_0__EVAL_29)
  );
  SiFive__EVAL_233 packageanon1_4 (
    ._EVAL(packageanon1_4__EVAL),
    ._EVAL_0(packageanon1_4__EVAL_0)
  );
  SiFive__EVAL_229 tlb (
    ._EVAL(tlb__EVAL),
    ._EVAL_0(tlb__EVAL_0),
    ._EVAL_1(tlb__EVAL_1),
    ._EVAL_2(tlb__EVAL_2),
    ._EVAL_3(tlb__EVAL_3),
    ._EVAL_4(tlb__EVAL_4),
    ._EVAL_5(tlb__EVAL_5),
    ._EVAL_6(tlb__EVAL_6),
    ._EVAL_7(tlb__EVAL_7),
    ._EVAL_8(tlb__EVAL_8),
    ._EVAL_9(tlb__EVAL_9),
    ._EVAL_10(tlb__EVAL_10),
    ._EVAL_11(tlb__EVAL_11),
    ._EVAL_12(tlb__EVAL_12),
    ._EVAL_13(tlb__EVAL_13),
    ._EVAL_14(tlb__EVAL_14),
    ._EVAL_15(tlb__EVAL_15),
    ._EVAL_16(tlb__EVAL_16),
    ._EVAL_17(tlb__EVAL_17),
    ._EVAL_18(tlb__EVAL_18),
    ._EVAL_19(tlb__EVAL_19),
    ._EVAL_20(tlb__EVAL_20),
    ._EVAL_21(tlb__EVAL_21),
    ._EVAL_22(tlb__EVAL_22),
    ._EVAL_23(tlb__EVAL_23),
    ._EVAL_24(tlb__EVAL_24),
    ._EVAL_25(tlb__EVAL_25),
    ._EVAL_26(tlb__EVAL_26),
    ._EVAL_27(tlb__EVAL_27),
    ._EVAL_28(tlb__EVAL_28),
    ._EVAL_29(tlb__EVAL_29),
    ._EVAL_30(tlb__EVAL_30),
    ._EVAL_31(tlb__EVAL_31),
    ._EVAL_32(tlb__EVAL_32),
    ._EVAL_33(tlb__EVAL_33),
    ._EVAL_34(tlb__EVAL_34),
    ._EVAL_35(tlb__EVAL_35),
    ._EVAL_36(tlb__EVAL_36),
    ._EVAL_37(tlb__EVAL_37),
    ._EVAL_38(tlb__EVAL_38),
    ._EVAL_39(tlb__EVAL_39),
    ._EVAL_40(tlb__EVAL_40),
    ._EVAL_41(tlb__EVAL_41),
    ._EVAL_42(tlb__EVAL_42),
    ._EVAL_43(tlb__EVAL_43),
    ._EVAL_44(tlb__EVAL_44),
    ._EVAL_45(tlb__EVAL_45),
    ._EVAL_46(tlb__EVAL_46),
    ._EVAL_47(tlb__EVAL_47),
    ._EVAL_48(tlb__EVAL_48),
    ._EVAL_49(tlb__EVAL_49),
    ._EVAL_50(tlb__EVAL_50),
    ._EVAL_51(tlb__EVAL_51),
    ._EVAL_52(tlb__EVAL_52),
    ._EVAL_53(tlb__EVAL_53),
    ._EVAL_54(tlb__EVAL_54),
    ._EVAL_55(tlb__EVAL_55),
    ._EVAL_56(tlb__EVAL_56),
    ._EVAL_57(tlb__EVAL_57),
    ._EVAL_58(tlb__EVAL_58),
    ._EVAL_59(tlb__EVAL_59),
    ._EVAL_60(tlb__EVAL_60),
    ._EVAL_61(tlb__EVAL_61),
    ._EVAL_62(tlb__EVAL_62)
  );
  SiFive__EVAL_341 itim_array (
    ._EVAL(itim_array__EVAL),
    ._EVAL_0(itim_array__EVAL_0),
    ._EVAL_1(itim_array__EVAL_1),
    ._EVAL_2(itim_array__EVAL_2),
    ._EVAL_3(itim_array__EVAL_3),
    ._EVAL_4(itim_array__EVAL_4)
  );
  SiFive__EVAL_230 packageanon1 (
    ._EVAL(packageanon1__EVAL),
    ._EVAL_0(packageanon1__EVAL_0)
  );
  assign _EVAL_215__EVAL_216_addr = _EVAL_2248;
  assign _EVAL_215__EVAL_216_data = _EVAL_215[_EVAL_215__EVAL_216_addr];
  assign _EVAL_215__EVAL_217_data = _EVAL_2034;
  assign _EVAL_215__EVAL_217_addr = _EVAL_254;
  assign _EVAL_215__EVAL_217_mask = 1'h1;
  assign _EVAL_215__EVAL_217_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_319__EVAL_320_addr = 1'h0;
  assign _EVAL_319__EVAL_320_data = _EVAL_319[_EVAL_319__EVAL_320_addr];
  assign _EVAL_319__EVAL_321_data = _EVAL_1560;
  assign _EVAL_319__EVAL_321_addr = 1'h0;
  assign _EVAL_319__EVAL_321_mask = 1'h1;
  assign _EVAL_319__EVAL_321_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_363__EVAL_364_addr = _EVAL_2248;
  assign _EVAL_363__EVAL_364_data = _EVAL_363[_EVAL_363__EVAL_364_addr];
  assign _EVAL_363__EVAL_365_data = _EVAL_1337;
  assign _EVAL_363__EVAL_365_addr = _EVAL_254;
  assign _EVAL_363__EVAL_365_mask = 1'h1;
  assign _EVAL_363__EVAL_365_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_386__EVAL_387_addr = _EVAL_2248;
  assign _EVAL_386__EVAL_387_data = _EVAL_386[_EVAL_386__EVAL_387_addr];
  assign _EVAL_386__EVAL_388_data = _EVAL_3306;
  assign _EVAL_386__EVAL_388_addr = _EVAL_254;
  assign _EVAL_386__EVAL_388_mask = 1'h1;
  assign _EVAL_386__EVAL_388_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_394__EVAL_395_addr = 1'h0;
  assign _EVAL_394__EVAL_395_data = _EVAL_394[_EVAL_394__EVAL_395_addr];
  assign _EVAL_394__EVAL_396_data = _EVAL_1234;
  assign _EVAL_394__EVAL_396_addr = 1'h0;
  assign _EVAL_394__EVAL_396_mask = 1'h1;
  assign _EVAL_394__EVAL_396_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_403__EVAL_404_addr = 1'h0;
  assign _EVAL_403__EVAL_404_data = _EVAL_403[_EVAL_403__EVAL_404_addr];
  assign _EVAL_403__EVAL_405_data = _EVAL_224;
  assign _EVAL_403__EVAL_405_addr = 1'h0;
  assign _EVAL_403__EVAL_405_mask = 1'h1;
  assign _EVAL_403__EVAL_405_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_489__EVAL_490_addr = _EVAL_2248;
  assign _EVAL_489__EVAL_490_data = _EVAL_489[_EVAL_489__EVAL_490_addr];
  assign _EVAL_489__EVAL_491_data = _EVAL_2118;
  assign _EVAL_489__EVAL_491_addr = _EVAL_254;
  assign _EVAL_489__EVAL_491_mask = 1'h1;
  assign _EVAL_489__EVAL_491_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_530__EVAL_531_addr = 1'h0;
  assign _EVAL_530__EVAL_531_data = _EVAL_530[_EVAL_530__EVAL_531_addr];
  assign _EVAL_530__EVAL_532_data = _EVAL_597;
  assign _EVAL_530__EVAL_532_addr = 1'h0;
  assign _EVAL_530__EVAL_532_mask = 1'h1;
  assign _EVAL_530__EVAL_532_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_548__EVAL_549_addr = _EVAL_2248;
  assign _EVAL_548__EVAL_549_data = _EVAL_548[_EVAL_548__EVAL_549_addr];
  assign _EVAL_548__EVAL_550_data = _EVAL_3160;
  assign _EVAL_548__EVAL_550_addr = _EVAL_254;
  assign _EVAL_548__EVAL_550_mask = 1'h1;
  assign _EVAL_548__EVAL_550_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_658__EVAL_659_addr = 1'h0;
  assign _EVAL_658__EVAL_659_data = _EVAL_658[_EVAL_658__EVAL_659_addr];
  assign _EVAL_658__EVAL_660_data = _EVAL_2586;
  assign _EVAL_658__EVAL_660_addr = 1'h0;
  assign _EVAL_658__EVAL_660_mask = 1'h1;
  assign _EVAL_658__EVAL_660_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_719__EVAL_720_addr = _EVAL_2248;
  assign _EVAL_719__EVAL_720_data = _EVAL_719[_EVAL_719__EVAL_720_addr];
  assign _EVAL_719__EVAL_721_data = _EVAL_701;
  assign _EVAL_719__EVAL_721_addr = _EVAL_254;
  assign _EVAL_719__EVAL_721_mask = 1'h1;
  assign _EVAL_719__EVAL_721_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_725__EVAL_726_addr = 1'h0;
  assign _EVAL_725__EVAL_726_data = _EVAL_725[_EVAL_725__EVAL_726_addr];
  assign _EVAL_725__EVAL_727_data = _EVAL_2247;
  assign _EVAL_725__EVAL_727_addr = 1'h0;
  assign _EVAL_725__EVAL_727_mask = 1'h1;
  assign _EVAL_725__EVAL_727_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_744__EVAL_745_addr = _EVAL_2248;
  assign _EVAL_744__EVAL_745_data = _EVAL_744[_EVAL_744__EVAL_745_addr];
  assign _EVAL_744__EVAL_746_data = _EVAL_772;
  assign _EVAL_744__EVAL_746_addr = _EVAL_254;
  assign _EVAL_744__EVAL_746_mask = 1'h1;
  assign _EVAL_744__EVAL_746_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_931__EVAL_932_addr = _EVAL_2248;
  assign _EVAL_931__EVAL_932_data = _EVAL_931[_EVAL_931__EVAL_932_addr];
  assign _EVAL_931__EVAL_933_data = _EVAL_675;
  assign _EVAL_931__EVAL_933_addr = _EVAL_254;
  assign _EVAL_931__EVAL_933_mask = 1'h1;
  assign _EVAL_931__EVAL_933_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_949__EVAL_950_addr = 1'h0;
  assign _EVAL_949__EVAL_950_data = _EVAL_949[_EVAL_949__EVAL_950_addr];
  assign _EVAL_949__EVAL_951_data = _EVAL_218;
  assign _EVAL_949__EVAL_951_addr = 1'h0;
  assign _EVAL_949__EVAL_951_mask = 1'h1;
  assign _EVAL_949__EVAL_951_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_961__EVAL_962_addr = _EVAL_2248;
  assign _EVAL_961__EVAL_962_data = _EVAL_961[_EVAL_961__EVAL_962_addr];
  assign _EVAL_961__EVAL_963_data = _EVAL_526;
  assign _EVAL_961__EVAL_963_addr = _EVAL_254;
  assign _EVAL_961__EVAL_963_mask = 1'h1;
  assign _EVAL_961__EVAL_963_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_982__EVAL_983_addr = 1'h0;
  assign _EVAL_982__EVAL_983_data = _EVAL_982[_EVAL_982__EVAL_983_addr];
  assign _EVAL_982__EVAL_984_data = _EVAL_1713;
  assign _EVAL_982__EVAL_984_addr = 1'h0;
  assign _EVAL_982__EVAL_984_mask = 1'h1;
  assign _EVAL_982__EVAL_984_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1119__EVAL_1120_addr = 1'h0;
  assign _EVAL_1119__EVAL_1120_data = _EVAL_1119[_EVAL_1119__EVAL_1120_addr];
  assign _EVAL_1119__EVAL_1121_data = _EVAL_1890;
  assign _EVAL_1119__EVAL_1121_addr = 1'h0;
  assign _EVAL_1119__EVAL_1121_mask = 1'h1;
  assign _EVAL_1119__EVAL_1121_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1140__EVAL_1141_addr = _EVAL_2248;
  assign _EVAL_1140__EVAL_1141_data = _EVAL_1140[_EVAL_1140__EVAL_1141_addr];
  assign _EVAL_1140__EVAL_1142_data = _EVAL_589;
  assign _EVAL_1140__EVAL_1142_addr = _EVAL_254;
  assign _EVAL_1140__EVAL_1142_mask = 1'h1;
  assign _EVAL_1140__EVAL_1142_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_1147__EVAL_1148_addr = 1'h0;
  assign _EVAL_1147__EVAL_1148_data = _EVAL_1147[_EVAL_1147__EVAL_1148_addr];
  assign _EVAL_1147__EVAL_1149_data = _EVAL_692;
  assign _EVAL_1147__EVAL_1149_addr = 1'h0;
  assign _EVAL_1147__EVAL_1149_mask = 1'h1;
  assign _EVAL_1147__EVAL_1149_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1440__EVAL_1441_addr = _EVAL_2248;
  assign _EVAL_1440__EVAL_1441_data = _EVAL_1440[_EVAL_1440__EVAL_1441_addr];
  assign _EVAL_1440__EVAL_1442_data = _EVAL_2856;
  assign _EVAL_1440__EVAL_1442_addr = _EVAL_254;
  assign _EVAL_1440__EVAL_1442_mask = 1'h1;
  assign _EVAL_1440__EVAL_1442_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_1465__EVAL_1466_addr = 1'h0;
  assign _EVAL_1465__EVAL_1466_data = _EVAL_1465[_EVAL_1465__EVAL_1466_addr];
  assign _EVAL_1465__EVAL_1467_data = _EVAL_1843;
  assign _EVAL_1465__EVAL_1467_addr = 1'h0;
  assign _EVAL_1465__EVAL_1467_mask = 1'h1;
  assign _EVAL_1465__EVAL_1467_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1481__EVAL_1482_addr = 1'h0;
  assign _EVAL_1481__EVAL_1482_data = _EVAL_1481[_EVAL_1481__EVAL_1482_addr];
  assign _EVAL_1481__EVAL_1483_data = _EVAL_151;
  assign _EVAL_1481__EVAL_1483_addr = 1'h0;
  assign _EVAL_1481__EVAL_1483_mask = 1'h1;
  assign _EVAL_1481__EVAL_1483_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1518__EVAL_1519_addr = _EVAL_2248;
  assign _EVAL_1518__EVAL_1519_data = _EVAL_1518[_EVAL_1518__EVAL_1519_addr];
  assign _EVAL_1518__EVAL_1520_data = _EVAL_593;
  assign _EVAL_1518__EVAL_1520_addr = _EVAL_254;
  assign _EVAL_1518__EVAL_1520_mask = 1'h1;
  assign _EVAL_1518__EVAL_1520_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_1652__EVAL_1653_addr = 1'h0;
  assign _EVAL_1652__EVAL_1653_data = _EVAL_1652[_EVAL_1652__EVAL_1653_addr];
  assign _EVAL_1652__EVAL_1654_data = _EVAL_812;
  assign _EVAL_1652__EVAL_1654_addr = 1'h0;
  assign _EVAL_1652__EVAL_1654_mask = 1'h1;
  assign _EVAL_1652__EVAL_1654_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1716__EVAL_1717_addr = 1'h0;
  assign _EVAL_1716__EVAL_1717_data = _EVAL_1716[_EVAL_1716__EVAL_1717_addr];
  assign _EVAL_1716__EVAL_1718_data = _EVAL_883;
  assign _EVAL_1716__EVAL_1718_addr = 1'h0;
  assign _EVAL_1716__EVAL_1718_mask = 1'h1;
  assign _EVAL_1716__EVAL_1718_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1767__EVAL_1768_addr = _EVAL_1102;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_1767__EVAL_1768_data = _EVAL_1767[_EVAL_1767__EVAL_1768_addr];
  `else
  assign _EVAL_1767__EVAL_1768_data = _EVAL_1767__EVAL_1768_addr >= 3'h6 ? _RAND_27[31:0] : _EVAL_1767[_EVAL_1767__EVAL_1768_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_1767__EVAL_1769_data = _EVAL_3148 | _EVAL_570;
  assign _EVAL_1767__EVAL_1769_addr = _EVAL_1606[2:0];
  assign _EVAL_1767__EVAL_1769_mask = 1'h1;
  assign _EVAL_1767__EVAL_1769_en = _EVAL_1077 ? _EVAL_971 : 1'h0;
  assign _EVAL_1859__EVAL_1860_addr = _EVAL_871[2:0];
  assign _EVAL_1859__EVAL_1860_data = _EVAL_1859[_EVAL_1859__EVAL_1860_addr];
  assign _EVAL_1859__EVAL_1861_addr = _EVAL_808[2:0];
  assign _EVAL_1859__EVAL_1861_data = _EVAL_1859[_EVAL_1859__EVAL_1861_addr];
  assign _EVAL_1859__EVAL_1862_data = {_EVAL_129,_EVAL_385};
  assign _EVAL_1859__EVAL_1862_addr = _EVAL_808[2:0];
  assign _EVAL_1859__EVAL_1862_mask = 1'h1;
  assign _EVAL_1859__EVAL_1862_en = _EVAL_77 ? _EVAL_257 : 1'h0;
  assign _EVAL_1895__EVAL_1896_addr = 1'h0;
  assign _EVAL_1895__EVAL_1896_data = _EVAL_1895[_EVAL_1895__EVAL_1896_addr];
  assign _EVAL_1895__EVAL_1897_data = _EVAL_2643;
  assign _EVAL_1895__EVAL_1897_addr = 1'h0;
  assign _EVAL_1895__EVAL_1897_mask = 1'h1;
  assign _EVAL_1895__EVAL_1897_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1986__EVAL_1987_addr = _EVAL_2248;
  assign _EVAL_1986__EVAL_1987_data = _EVAL_1986[_EVAL_1986__EVAL_1987_addr];
  assign _EVAL_1986__EVAL_1988_data = _EVAL_2055;
  assign _EVAL_1986__EVAL_1988_addr = _EVAL_254;
  assign _EVAL_1986__EVAL_1988_mask = 1'h1;
  assign _EVAL_1986__EVAL_1988_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2023__EVAL_2024_addr = 1'h0;
  assign _EVAL_2023__EVAL_2024_data = _EVAL_2023[_EVAL_2023__EVAL_2024_addr];
  assign _EVAL_2023__EVAL_2025_data = _EVAL_1385;
  assign _EVAL_2023__EVAL_2025_addr = 1'h0;
  assign _EVAL_2023__EVAL_2025_mask = 1'h1;
  assign _EVAL_2023__EVAL_2025_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_2073__EVAL_2074_addr = _EVAL_2248;
  assign _EVAL_2073__EVAL_2074_data = _EVAL_2073[_EVAL_2073__EVAL_2074_addr];
  assign _EVAL_2073__EVAL_2075_data = _EVAL_732;
  assign _EVAL_2073__EVAL_2075_addr = _EVAL_254;
  assign _EVAL_2073__EVAL_2075_mask = 1'h1;
  assign _EVAL_2073__EVAL_2075_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2081__EVAL_2082_addr = _EVAL_2248;
  assign _EVAL_2081__EVAL_2082_data = _EVAL_2081[_EVAL_2081__EVAL_2082_addr];
  assign _EVAL_2081__EVAL_2083_data = _EVAL_2057;
  assign _EVAL_2081__EVAL_2083_addr = _EVAL_254;
  assign _EVAL_2081__EVAL_2083_mask = 1'h1;
  assign _EVAL_2081__EVAL_2083_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2177__EVAL_2178_addr = _EVAL_2248;
  assign _EVAL_2177__EVAL_2178_data = _EVAL_2177[_EVAL_2177__EVAL_2178_addr];
  assign _EVAL_2177__EVAL_2179_data = _EVAL_1647;
  assign _EVAL_2177__EVAL_2179_addr = _EVAL_254;
  assign _EVAL_2177__EVAL_2179_mask = 1'h1;
  assign _EVAL_2177__EVAL_2179_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2229__EVAL_2230_addr = 1'h0;
  assign _EVAL_2229__EVAL_2230_data = _EVAL_2229[_EVAL_2229__EVAL_2230_addr];
  assign _EVAL_2229__EVAL_2231_data = _EVAL_823;
  assign _EVAL_2229__EVAL_2231_addr = 1'h0;
  assign _EVAL_2229__EVAL_2231_mask = 1'h1;
  assign _EVAL_2229__EVAL_2231_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_2337__EVAL_2338_addr = 1'h0;
  assign _EVAL_2337__EVAL_2338_data = _EVAL_2337[_EVAL_2337__EVAL_2338_addr];
  assign _EVAL_2337__EVAL_2339_data = _EVAL_2651;
  assign _EVAL_2337__EVAL_2339_addr = 1'h0;
  assign _EVAL_2337__EVAL_2339_mask = 1'h1;
  assign _EVAL_2337__EVAL_2339_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_2478__EVAL_2479_addr = 1'h0;
  assign _EVAL_2478__EVAL_2479_data = _EVAL_2478[_EVAL_2478__EVAL_2479_addr];
  assign _EVAL_2478__EVAL_2480_data = _EVAL_545;
  assign _EVAL_2478__EVAL_2480_addr = 1'h0;
  assign _EVAL_2478__EVAL_2480_mask = 1'h1;
  assign _EVAL_2478__EVAL_2480_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_2542__EVAL_2543_addr = 1'h0;
  assign _EVAL_2542__EVAL_2543_data = _EVAL_2542[_EVAL_2542__EVAL_2543_addr];
  assign _EVAL_2542__EVAL_2544_data = _EVAL_1020;
  assign _EVAL_2542__EVAL_2544_addr = 1'h0;
  assign _EVAL_2542__EVAL_2544_mask = 1'h1;
  assign _EVAL_2542__EVAL_2544_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_2573__EVAL_2574_addr = _EVAL_2248;
  assign _EVAL_2573__EVAL_2574_data = _EVAL_2573[_EVAL_2573__EVAL_2574_addr];
  assign _EVAL_2573__EVAL_2575_data = _EVAL_1838;
  assign _EVAL_2573__EVAL_2575_addr = _EVAL_254;
  assign _EVAL_2573__EVAL_2575_mask = 1'h1;
  assign _EVAL_2573__EVAL_2575_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2580__EVAL_2581_addr = _EVAL_2248;
  assign _EVAL_2580__EVAL_2581_data = _EVAL_2580[_EVAL_2580__EVAL_2581_addr];
  assign _EVAL_2580__EVAL_2582_data = _EVAL_2617;
  assign _EVAL_2580__EVAL_2582_addr = _EVAL_254;
  assign _EVAL_2580__EVAL_2582_mask = 1'h1;
  assign _EVAL_2580__EVAL_2582_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2591__EVAL_2592_addr = _EVAL_2248;
  assign _EVAL_2591__EVAL_2592_data = _EVAL_2591[_EVAL_2591__EVAL_2592_addr];
  assign _EVAL_2591__EVAL_2593_data = _EVAL_2313;
  assign _EVAL_2591__EVAL_2593_addr = _EVAL_254;
  assign _EVAL_2591__EVAL_2593_mask = 1'h1;
  assign _EVAL_2591__EVAL_2593_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2712__EVAL_2713_addr = 1'h0;
  assign _EVAL_2712__EVAL_2713_data = _EVAL_2712[_EVAL_2712__EVAL_2713_addr];
  assign _EVAL_2712__EVAL_2714_data = _EVAL_3024;
  assign _EVAL_2712__EVAL_2714_addr = 1'h0;
  assign _EVAL_2712__EVAL_2714_mask = 1'h1;
  assign _EVAL_2712__EVAL_2714_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_2773__EVAL_2774_addr = _EVAL_2248;
  assign _EVAL_2773__EVAL_2774_data = _EVAL_2773[_EVAL_2773__EVAL_2774_addr];
  assign _EVAL_2773__EVAL_2775_data = _EVAL_595;
  assign _EVAL_2773__EVAL_2775_addr = _EVAL_254;
  assign _EVAL_2773__EVAL_2775_mask = 1'h1;
  assign _EVAL_2773__EVAL_2775_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2852__EVAL_2853_addr = _EVAL_2248;
  assign _EVAL_2852__EVAL_2853_data = _EVAL_2852[_EVAL_2852__EVAL_2853_addr];
  assign _EVAL_2852__EVAL_2854_data = _EVAL_909;
  assign _EVAL_2852__EVAL_2854_addr = _EVAL_254;
  assign _EVAL_2852__EVAL_2854_mask = 1'h1;
  assign _EVAL_2852__EVAL_2854_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_3001__EVAL_3002_addr = 1'h0;
  assign _EVAL_3001__EVAL_3002_data = _EVAL_3001[_EVAL_3001__EVAL_3002_addr];
  assign _EVAL_3001__EVAL_3003_data = _EVAL_1072;
  assign _EVAL_3001__EVAL_3003_addr = 1'h0;
  assign _EVAL_3001__EVAL_3003_mask = 1'h1;
  assign _EVAL_3001__EVAL_3003_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_3082__EVAL_3083_addr = 1'h0;
  assign _EVAL_3082__EVAL_3083_data = _EVAL_3082[_EVAL_3082__EVAL_3083_addr];
  assign _EVAL_3082__EVAL_3084_data = _EVAL_1047;
  assign _EVAL_3082__EVAL_3084_addr = 1'h0;
  assign _EVAL_3082__EVAL_3084_mask = 1'h1;
  assign _EVAL_3082__EVAL_3084_en = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_3112__EVAL_3113_addr = _EVAL_2248;
  assign _EVAL_3112__EVAL_3113_data = _EVAL_3112[_EVAL_3112__EVAL_3113_addr];
  assign _EVAL_3112__EVAL_3114_data = _EVAL_3393;
  assign _EVAL_3112__EVAL_3114_addr = _EVAL_254;
  assign _EVAL_3112__EVAL_3114_mask = 1'h1;
  assign _EVAL_3112__EVAL_3114_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_3335__EVAL_3336_addr = _EVAL_2248;
  assign _EVAL_3335__EVAL_3336_data = _EVAL_3335[_EVAL_3335__EVAL_3336_addr];
  assign _EVAL_3335__EVAL_3337_data = 1'h0;
  assign _EVAL_3335__EVAL_3337_addr = _EVAL_254;
  assign _EVAL_3335__EVAL_3337_mask = 1'h1;
  assign _EVAL_3335__EVAL_3337_en = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_228 = icache_clock_gate_out;
  assign _EVAL_751 = _EVAL_57;
  assign _EVAL_255 = _EVAL_751;
  assign _EVAL_973 = _EVAL_751;
  assign _EVAL_1981 = _EVAL_481 == 3'h3;
  assign _EVAL_3080 = _EVAL_1981 == 1'h0;
  assign _EVAL_1781 = _EVAL_1836 == 1'h0;
  assign _EVAL_2472 = _EVAL_3080 & _EVAL_1781;
  assign _EVAL_2092 = _EVAL_2472 ? 1'h0 : 1'h1;
  assign _EVAL_2897 = _EVAL_2472 ? 9'h0 : 9'h1ff;
  assign _EVAL_1677 = _EVAL_2880 != _EVAL_2413;
  assign _EVAL_1751 = _EVAL_1677 == 1'h0;
  assign _EVAL_1192 = _EVAL_1751 & _EVAL_900;
  assign _EVAL_1636 = _EVAL_3080 | _EVAL_1192;
  assign _EVAL_1980 = {_EVAL_2092,_EVAL_2092,_EVAL_2897,_EVAL_1636};
  assign _EVAL_1215 = _EVAL_3261 == 1'h0;
  assign _EVAL_3321 = _EVAL_1386 == 1'h0;
  assign _EVAL_1955 = _EVAL_2629 == 1'h0;
  assign _EVAL_362 = _EVAL_1954 == 1'h0;
  assign _EVAL_3076 = _EVAL_3089;
  assign _EVAL_1983 = _EVAL_362 & _EVAL_3076;
  assign _EVAL_1365 = _EVAL_3019 | _EVAL_1983;
  assign _EVAL_1589 = _EVAL_1955 & _EVAL_1365;
  assign _EVAL_1841 = _EVAL_1244 | _EVAL_1589;
  assign _EVAL_2288 = _EVAL_3321 & _EVAL_1841;
  assign _EVAL_1797 = _EVAL_928 | _EVAL_2288;
  assign _EVAL_3092 = _EVAL_1215 & _EVAL_1797;
  assign _EVAL_542 = _EVAL_1415 | _EVAL_3092;
  assign _EVAL_182 = _EVAL_542 == 1'h0;
  assign _EVAL_3181 = _EVAL_1412 == 1'h0;
  assign _EVAL_645 = _EVAL_182 & _EVAL_3181;
  assign _EVAL_956 = _EVAL_645 == 1'h0;
  assign _EVAL_169 = _EVAL_3376[1:0];
  assign _EVAL_2191 = _EVAL_169 == 2'h1;
  assign _EVAL_2658 = _EVAL_3376[15:13];
  assign _EVAL_518 = _EVAL_2658 == 3'h1;
  assign _EVAL_2969 = _EVAL_2191 & _EVAL_518;
  assign _EVAL_2018 = _EVAL_3376[15];
  assign _EVAL_159 = _EVAL_2191 & _EVAL_2018;
  assign _EVAL_724 = _EVAL_3376[14:13];
  assign _EVAL_786 = _EVAL_724 == 2'h1;
  assign _EVAL_1313 = _EVAL_159 & _EVAL_786;
  assign _EVAL_282 = _EVAL_2969 | _EVAL_1313;
  assign _EVAL_1605 = _EVAL_2084 & _EVAL_3181;
  assign _EVAL_2723 = _EVAL_1605 == 1'h0;
  assign _EVAL_2465 = _EVAL_282 & _EVAL_2723;
  assign _EVAL_1426 = _EVAL_724 == 2'h0;
  assign _EVAL_2133 = _EVAL_159 & _EVAL_1426;
  assign _EVAL_769 = _EVAL_2465 | _EVAL_2133;
  assign _EVAL_1930 = _EVAL_3376[14];
  assign _EVAL_2443 = _EVAL_159 & _EVAL_1930;
  assign _EVAL_2366 = _EVAL_542 != _EVAL_1412;
  assign _EVAL_1295 = _EVAL_1004 ? _EVAL_1544 : 64'h0;
  assign _EVAL_1271 = _EVAL_2799 ? _EVAL_2971 : 64'h0;
  assign _EVAL_2668 = _EVAL_1295 | _EVAL_1271;
  assign _EVAL_2618 = _EVAL_1344 ? _EVAL_1168 : 64'h0;
  assign _EVAL_1214 = _EVAL_839 ? _EVAL_1434 : 64'h0;
  assign _EVAL_1402 = _EVAL_2618 | _EVAL_1214;
  assign _EVAL_3203 = _EVAL_2668 | _EVAL_1402;
  assign _EVAL_164 = _EVAL_1085 ? _EVAL_2062 : 64'h0;
  assign _EVAL_442 = _EVAL_2888 ? _EVAL_2383 : 64'h0;
  assign _EVAL_993 = _EVAL_164 | _EVAL_442;
  assign _EVAL_1550 = _EVAL_3203 | _EVAL_993;
  assign _EVAL_342 = _EVAL_3220 ? _EVAL_2078 : 64'h0;
  assign _EVAL_502 = _EVAL_1807 ? _EVAL_2655 : 64'h0;
  assign _EVAL_1613 = _EVAL_342 | _EVAL_502;
  assign _EVAL_2947 = _EVAL_1550 | _EVAL_1613;
  assign _EVAL_2761 = _EVAL_731 ? _EVAL_2785 : 64'h0;
  assign _EVAL_1504 = _EVAL_2947 | _EVAL_2761;
  assign _EVAL_2227 = _EVAL_1504[15:0];
  assign _EVAL_2168 = _EVAL_2227[1:0];
  assign _EVAL_3211 = _EVAL_2168 == 2'h1;
  assign _EVAL_2327 = _EVAL_2227[15];
  assign _EVAL_315 = _EVAL_3211 & _EVAL_2327;
  assign _EVAL_2980 = _EVAL_2227[14];
  assign _EVAL_2621 = _EVAL_315 & _EVAL_2980;
  assign _EVAL_2728 = _EVAL_2227[6:0];
  assign _EVAL_3276 = _EVAL_2728 & 7'h77;
  assign _EVAL_1245 = _EVAL_3276 == 7'h63;
  assign _EVAL_1719 = _EVAL_2621 | _EVAL_1245;
  assign _EVAL_194 = _EVAL_2168 < 2'h3;
  assign _EVAL_995 = _EVAL_1504[31:16];
  assign _EVAL_1545 = _EVAL_995[1:0];
  assign _EVAL_2645 = _EVAL_1545 == 2'h1;
  assign _EVAL_1610 = _EVAL_995[15];
  assign _EVAL_3071 = _EVAL_2645 & _EVAL_1610;
  assign _EVAL_1607 = _EVAL_995[14];
  assign _EVAL_2012 = _EVAL_3071 & _EVAL_1607;
  assign _EVAL_3281 = _EVAL_995[6:0];
  assign _EVAL_2326 = _EVAL_3281 & 7'h77;
  assign _EVAL_684 = _EVAL_2326 == 7'h63;
  assign _EVAL_942 = _EVAL_2012 | _EVAL_684;
  assign _EVAL_1114 = _EVAL_1545 < 2'h3;
  assign _EVAL_2291 = _EVAL_1504[47:32];
  assign _EVAL_1952 = _EVAL_2291[1:0];
  assign _EVAL_1934 = _EVAL_1952 == 2'h1;
  assign _EVAL_1642 = _EVAL_2291[15];
  assign _EVAL_1557 = _EVAL_1934 & _EVAL_1642;
  assign _EVAL_1008 = _EVAL_2291[14];
  assign _EVAL_902 = _EVAL_1557 & _EVAL_1008;
  assign _EVAL_174 = _EVAL_2291[6:0];
  assign _EVAL_1221 = _EVAL_174 & 7'h77;
  assign _EVAL_393 = _EVAL_1221 == 7'h63;
  assign _EVAL_740 = _EVAL_902 | _EVAL_393;
  assign _EVAL_1078 = _EVAL_1952 < 2'h3;
  assign _EVAL_1336 = _EVAL_1504[63:48];
  assign _EVAL_3064 = _EVAL_1336[1:0];
  assign _EVAL_1867 = _EVAL_3064 == 2'h1;
  assign _EVAL_2103 = _EVAL_1336[15];
  assign _EVAL_2557 = _EVAL_1867 & _EVAL_2103;
  assign _EVAL_381 = _EVAL_1336[14];
  assign _EVAL_1035 = _EVAL_2557 & _EVAL_381;
  assign _EVAL_3000 = _EVAL_1078 ? _EVAL_1035 : 1'h0;
  assign _EVAL_336 = _EVAL_740 | _EVAL_3000;
  assign _EVAL_1091 = _EVAL_1114 ? _EVAL_336 : _EVAL_1035;
  assign _EVAL_1209 = _EVAL_942 | _EVAL_1091;
  assign _EVAL_1967 = _EVAL_194 ? _EVAL_1209 : _EVAL_336;
  assign _EVAL_2336 = _EVAL_1719 | _EVAL_1967;
  assign _EVAL_1100 = _EVAL_2366 | _EVAL_2336;
  assign _EVAL_1732 = _EVAL_2443 & _EVAL_1100;
  assign _EVAL_2030 = _EVAL_769 | _EVAL_1732;
  assign _EVAL_2173 = _EVAL_2518 & _EVAL_2030;
  assign _EVAL_3348 = _EVAL_2950[2];
  assign _EVAL_3039 = _EVAL_1387[6];
  assign _EVAL_402 = _EVAL_1387[5];
  assign _EVAL_3107 = _EVAL_1387[4];
  assign _EVAL_1226 = _EVAL_1387[3];
  assign _EVAL_3303 = _EVAL_1387[2];
  assign _EVAL_230 = _EVAL_1387[1];
  assign _EVAL_2458 = _EVAL_1387[0];
  assign _EVAL_1996 = _EVAL_837[0];
  assign _EVAL_2066 = _EVAL_837[127:1];
  assign _EVAL_3155 = {_EVAL_1996,_EVAL_2066};
  assign _EVAL_2115 = _EVAL_2458 ? _EVAL_3155 : _EVAL_837;
  assign _EVAL_1502 = _EVAL_2115[1:0];
  assign _EVAL_295 = _EVAL_2115[127:2];
  assign _EVAL_1305 = {_EVAL_1502,_EVAL_295};
  assign _EVAL_349 = _EVAL_230 ? _EVAL_1305 : _EVAL_2115;
  assign _EVAL_1893 = _EVAL_349[3:0];
  assign _EVAL_3038 = _EVAL_349[127:4];
  assign _EVAL_1358 = {_EVAL_1893,_EVAL_3038};
  assign _EVAL_1772 = _EVAL_3303 ? _EVAL_1358 : _EVAL_349;
  assign _EVAL_699 = _EVAL_1772[7:0];
  assign _EVAL_3308 = _EVAL_1772[127:8];
  assign _EVAL_1916 = {_EVAL_699,_EVAL_3308};
  assign _EVAL_2286 = _EVAL_1226 ? _EVAL_1916 : _EVAL_1772;
  assign _EVAL_1978 = _EVAL_2286[15:0];
  assign _EVAL_2160 = _EVAL_2286[127:16];
  assign _EVAL_2899 = {_EVAL_1978,_EVAL_2160};
  assign _EVAL_1491 = _EVAL_3107 ? _EVAL_2899 : _EVAL_2286;
  assign _EVAL_2426 = _EVAL_1491[31:0];
  assign _EVAL_247 = _EVAL_1491[127:32];
  assign _EVAL_1292 = {_EVAL_2426,_EVAL_247};
  assign _EVAL_2100 = _EVAL_402 ? _EVAL_1292 : _EVAL_1491;
  assign _EVAL_2569 = _EVAL_2100[63:0];
  assign _EVAL_2464 = _EVAL_2100[127:64];
  assign _EVAL_2436 = {_EVAL_2569,_EVAL_2464};
  assign _EVAL_1670 = _EVAL_3039 ? _EVAL_2436 : _EVAL_2100;
  assign _EVAL_691 = {{1'd0}, _EVAL_1670};
  assign _EVAL_3405 = _EVAL_927 == 1'h0;
  assign _EVAL_2218 = _EVAL_1412 & _EVAL_3405;
  assign _EVAL_325 = _EVAL_2218 & _EVAL_182;
  assign _EVAL_2120 = _EVAL_325 == 1'h0;
  assign _EVAL_761 = _EVAL_2252 == 1'h0;
  assign _EVAL_187 = _EVAL_344 & _EVAL_761;
  assign _EVAL_1377 = _EVAL_1529 ? _EVAL_2120 : _EVAL_187;
  assign _EVAL_2059 = _EVAL_691 << _EVAL_1377;
  assign _EVAL_3265 = _EVAL_2059[127:0];
  assign _EVAL_2765 = {{1'd0}, _EVAL_3265};
  assign _EVAL_892 = _EVAL_344 & _EVAL_1529;
  assign _EVAL_1592 = _EVAL_3376[6:0];
  assign _EVAL_520 = _EVAL_1592 & 7'h7b;
  assign _EVAL_2330 = _EVAL_520 == 7'h6b;
  assign _EVAL_2486 = _EVAL_2330 & _EVAL_2723;
  assign _EVAL_2293 = _EVAL_1592 == 7'h67;
  assign _EVAL_178 = _EVAL_2486 | _EVAL_2293;
  assign _EVAL_2365 = _EVAL_1592 & 7'h77;
  assign _EVAL_713 = _EVAL_2365 == 7'h63;
  assign _EVAL_3075 = _EVAL_2366 | _EVAL_1209;
  assign _EVAL_3186 = _EVAL_713 & _EVAL_3075;
  assign _EVAL_3179 = _EVAL_178 | _EVAL_3186;
  assign _EVAL_3006 = _EVAL_2518 & _EVAL_3179;
  assign _EVAL_204 = _EVAL_2173 | _EVAL_3006;
  assign _EVAL_2794 = _EVAL_169 < 2'h3;
  assign _EVAL_304 = _EVAL_2392[2:1];
  assign _EVAL_3135 = 2'h0 >= _EVAL_304;
  assign _EVAL_2384 = _EVAL_2518 ? _EVAL_2794 : _EVAL_3135;
  assign _EVAL_2068 = _EVAL_2227[15:13];
  assign _EVAL_773 = _EVAL_2068 == 3'h1;
  assign _EVAL_858 = _EVAL_3211 & _EVAL_773;
  assign _EVAL_2877 = _EVAL_2227[14:13];
  assign _EVAL_2940 = _EVAL_2877 == 2'h1;
  assign _EVAL_1851 = _EVAL_315 & _EVAL_2940;
  assign _EVAL_1855 = _EVAL_858 | _EVAL_1851;
  assign _EVAL_2973 = _EVAL_1855 & _EVAL_2723;
  assign _EVAL_3016 = _EVAL_2877 == 2'h0;
  assign _EVAL_2410 = _EVAL_315 & _EVAL_3016;
  assign _EVAL_2613 = _EVAL_2973 | _EVAL_2410;
  assign _EVAL_1143 = _EVAL_2621 & _EVAL_3075;
  assign _EVAL_1154 = _EVAL_2613 | _EVAL_1143;
  assign _EVAL_2014 = _EVAL_2384 & _EVAL_1154;
  assign _EVAL_1976 = _EVAL_2728 & 7'h7b;
  assign _EVAL_3106 = _EVAL_1976 == 7'h6b;
  assign _EVAL_2499 = _EVAL_3106 & _EVAL_2723;
  assign _EVAL_1631 = _EVAL_2728 == 7'h67;
  assign _EVAL_300 = _EVAL_2499 | _EVAL_1631;
  assign _EVAL_249 = _EVAL_2366 | _EVAL_336;
  assign _EVAL_1070 = _EVAL_1245 & _EVAL_249;
  assign _EVAL_2972 = _EVAL_300 | _EVAL_1070;
  assign _EVAL_2975 = _EVAL_2384 & _EVAL_2972;
  assign _EVAL_2044 = _EVAL_2014 | _EVAL_2975;
  assign _EVAL_867 = _EVAL_204 | _EVAL_2044;
  assign _EVAL_3133 = 2'h1 >= _EVAL_304;
  assign _EVAL_2158 = _EVAL_2384 ? _EVAL_194 : _EVAL_3133;
  assign _EVAL_779 = _EVAL_995[15:13];
  assign _EVAL_369 = _EVAL_779 == 3'h1;
  assign _EVAL_1343 = _EVAL_2645 & _EVAL_369;
  assign _EVAL_3258 = _EVAL_995[14:13];
  assign _EVAL_2556 = _EVAL_3258 == 2'h1;
  assign _EVAL_2363 = _EVAL_3071 & _EVAL_2556;
  assign _EVAL_1025 = _EVAL_1343 | _EVAL_2363;
  assign _EVAL_2289 = _EVAL_1025 & _EVAL_2723;
  assign _EVAL_735 = _EVAL_3258 == 2'h0;
  assign _EVAL_1686 = _EVAL_3071 & _EVAL_735;
  assign _EVAL_2697 = _EVAL_2289 | _EVAL_1686;
  assign _EVAL_1159 = _EVAL_2012 & _EVAL_249;
  assign _EVAL_3323 = _EVAL_2697 | _EVAL_1159;
  assign _EVAL_1011 = _EVAL_2158 & _EVAL_3323;
  assign _EVAL_2692 = _EVAL_3281 & 7'h7b;
  assign _EVAL_970 = _EVAL_2692 == 7'h6b;
  assign _EVAL_2756 = _EVAL_970 & _EVAL_2723;
  assign _EVAL_1564 = _EVAL_3281 == 7'h67;
  assign _EVAL_515 = _EVAL_2756 | _EVAL_1564;
  assign _EVAL_378 = _EVAL_2366 | _EVAL_1035;
  assign _EVAL_2306 = _EVAL_684 & _EVAL_378;
  assign _EVAL_3163 = _EVAL_515 | _EVAL_2306;
  assign _EVAL_1051 = _EVAL_2158 & _EVAL_3163;
  assign _EVAL_2885 = _EVAL_1011 | _EVAL_1051;
  assign _EVAL_868 = _EVAL_867 | _EVAL_2885;
  assign _EVAL_3117 = 2'h2 >= _EVAL_304;
  assign _EVAL_1276 = _EVAL_2158 ? _EVAL_1114 : _EVAL_3117;
  assign _EVAL_2755 = _EVAL_2291[15:13];
  assign _EVAL_238 = _EVAL_2755 == 3'h1;
  assign _EVAL_2431 = _EVAL_1934 & _EVAL_238;
  assign _EVAL_920 = _EVAL_2291[14:13];
  assign _EVAL_1758 = _EVAL_920 == 2'h1;
  assign _EVAL_2043 = _EVAL_1557 & _EVAL_1758;
  assign _EVAL_641 = _EVAL_2431 | _EVAL_2043;
  assign _EVAL_1400 = _EVAL_641 & _EVAL_2723;
  assign _EVAL_771 = _EVAL_920 == 2'h0;
  assign _EVAL_3063 = _EVAL_1557 & _EVAL_771;
  assign _EVAL_231 = _EVAL_1400 | _EVAL_3063;
  assign _EVAL_2020 = _EVAL_902 & _EVAL_378;
  assign _EVAL_1032 = _EVAL_231 | _EVAL_2020;
  assign _EVAL_1883 = _EVAL_1276 & _EVAL_1032;
  assign _EVAL_989 = _EVAL_174 & 7'h7b;
  assign _EVAL_2742 = _EVAL_989 == 7'h6b;
  assign _EVAL_1965 = _EVAL_2742 & _EVAL_2723;
  assign _EVAL_3319 = _EVAL_174 == 7'h67;
  assign _EVAL_3250 = _EVAL_1965 | _EVAL_3319;
  assign _EVAL_184 = _EVAL_393 & _EVAL_2366;
  assign _EVAL_3398 = _EVAL_3250 | _EVAL_184;
  assign _EVAL_2816 = _EVAL_1276 & _EVAL_3398;
  assign _EVAL_3169 = _EVAL_1883 | _EVAL_2816;
  assign _EVAL_607 = _EVAL_868 | _EVAL_3169;
  assign _EVAL_3105 = _EVAL_1276 ? _EVAL_1078 : 1'h1;
  assign _EVAL_1580 = _EVAL_1336[15:13];
  assign _EVAL_1733 = _EVAL_1580 == 3'h1;
  assign _EVAL_2396 = _EVAL_1867 & _EVAL_1733;
  assign _EVAL_3364 = _EVAL_1336[14:13];
  assign _EVAL_2451 = _EVAL_3364 == 2'h1;
  assign _EVAL_748 = _EVAL_2557 & _EVAL_2451;
  assign _EVAL_1193 = _EVAL_2396 | _EVAL_748;
  assign _EVAL_874 = _EVAL_1193 & _EVAL_2723;
  assign _EVAL_309 = _EVAL_3364 == 2'h0;
  assign _EVAL_1537 = _EVAL_2557 & _EVAL_309;
  assign _EVAL_2353 = _EVAL_874 | _EVAL_1537;
  assign _EVAL_1439 = _EVAL_1035 & _EVAL_2366;
  assign _EVAL_1827 = _EVAL_2353 | _EVAL_1439;
  assign _EVAL_2198 = _EVAL_3105 & _EVAL_1827;
  assign _EVAL_1995 = _EVAL_607 | _EVAL_2198;
  assign _EVAL_935 = _EVAL_1995 == 1'h0;
  assign _EVAL_316 = _EVAL_892 & _EVAL_935;
  assign _EVAL_2284 = _EVAL_2765 << _EVAL_316;
  assign _EVAL_2538 = _EVAL_2284[128:2];
  assign _EVAL_166 = {_EVAL_2538, 2'h0};
  assign _EVAL_2531 = _EVAL_166[127:0];
  assign _EVAL_1500 = _EVAL_2531[70];
  assign _EVAL_624 = _EVAL_2531[65];
  assign _EVAL_667 = _EVAL_2531[61];
  assign _EVAL_1311 = _EVAL_2531[57];
  assign _EVAL_2810 = _EVAL_2531[53];
  assign _EVAL_3266 = _EVAL_2531[49];
  assign _EVAL_2049 = _EVAL_2531[45];
  assign _EVAL_3299 = _EVAL_2531[41];
  assign _EVAL_1443 = _EVAL_2531[37];
  assign _EVAL_2521 = _EVAL_2531[32];
  assign _EVAL_3139 = _EVAL_2531[28];
  assign _EVAL_2387 = _EVAL_2531[24];
  assign _EVAL_3264 = _EVAL_2531[20];
  assign _EVAL_1129 = _EVAL_2531[16];
  assign _EVAL_3388 = _EVAL_2531[12];
  assign _EVAL_1711 = _EVAL_2531[8];
  assign _EVAL_1927 = _EVAL_2531[4];
  assign _EVAL_2553 = _EVAL_2531[0];
  assign _EVAL_2283 = {_EVAL_2521,_EVAL_3139,_EVAL_2387,_EVAL_3264,_EVAL_1129,_EVAL_3388,_EVAL_1711,_EVAL_1927,_EVAL_2553};
  assign _EVAL_2172 = {_EVAL_1500,_EVAL_624,_EVAL_667,_EVAL_1311,_EVAL_2810,_EVAL_3266,_EVAL_2049,_EVAL_3299,_EVAL_1443,_EVAL_2283};
  assign _EVAL_1195 = _EVAL_1523 | _EVAL_1272;
  assign _EVAL_861 = _EVAL_1195 | _EVAL_2399;
  assign _EVAL_1804 = _EVAL_861 | _EVAL_664;
  assign _EVAL_2029 = _EVAL_1804 | _EVAL_731;
  assign _EVAL_145 = _EVAL_2029 == 1'h0;
  assign _EVAL_3033 = _EVAL_145 & _EVAL_1591;
  assign _EVAL_3053 = _EVAL_1731 == 1'h0;
  assign _EVAL_1475 = _EVAL_3033 & _EVAL_3053;
  assign _EVAL_1312 = _EVAL_2029 | _EVAL_1475;
  assign _EVAL_419 = _EVAL_1312 | _EVAL_957;
  assign _EVAL_1077 = _EVAL_1529 & _EVAL_419;
  assign _EVAL_2860 = _EVAL_1077 == 1'h0;
  assign _EVAL_1640 = _EVAL_2252 & _EVAL_2860;
  assign _EVAL_2843 = _EVAL_1640 | _EVAL_3370;
  assign _EVAL_273 = _EVAL_2843 == 1'h0;
  assign _EVAL_1366 = _EVAL_273 & _EVAL_2252;
  assign _EVAL_3296 = _EVAL_1366 & _EVAL_1995;
  assign _EVAL_1463 = _EVAL_2133 | _EVAL_2293;
  assign _EVAL_2789 = _EVAL_282 | _EVAL_2330;
  assign _EVAL_1991 = _EVAL_1463 | _EVAL_2789;
  assign _EVAL_1375 = _EVAL_1991 | _EVAL_1732;
  assign _EVAL_2900 = _EVAL_1375 | _EVAL_3186;
  assign _EVAL_2139 = _EVAL_2518 & _EVAL_2900;
  assign _EVAL_1169 = _EVAL_3376[1];
  assign _EVAL_919 = _EVAL_1169 == 1'h0;
  assign _EVAL_2394 = _EVAL_3376[3];
  assign _EVAL_377 = _EVAL_919 ? _EVAL_786 : _EVAL_2394;
  assign _EVAL_1036 = _EVAL_3376[2];
  assign _EVAL_758 = _EVAL_1036 == 1'h0;
  assign _EVAL_2671 = _EVAL_919 ? _EVAL_1930 : _EVAL_758;
  assign _EVAL_1407 = _EVAL_2671 & _EVAL_542;
  assign _EVAL_474 = _EVAL_377 | _EVAL_1407;
  assign _EVAL_930 = _EVAL_2273 | 32'h6;
  assign _EVAL_158 = $signed(_EVAL_930);
  assign _EVAL_1492 = {_EVAL_2227,_EVAL_3376};
  assign _EVAL_777 = _EVAL_1492[1];
  assign _EVAL_1633 = _EVAL_1492[31:16];
  assign _EVAL_1678 = _EVAL_1633[15:2];
  assign _EVAL_622 = _EVAL_1633[15:13];
  assign _EVAL_818 = _EVAL_622 == 3'h4;
  assign _EVAL_1779 = _EVAL_1633[6:2];
  assign _EVAL_1618 = _EVAL_1779 == 5'h0;
  assign _EVAL_305 = _EVAL_1633[1:0];
  assign _EVAL_1136 = _EVAL_305[0];
  assign _EVAL_553 = _EVAL_305[1];
  assign _EVAL_937 = _EVAL_1618 ? _EVAL_1136 : _EVAL_553;
  assign _EVAL_1469 = _EVAL_553 == _EVAL_1136;
  assign _EVAL_1870 = {_EVAL_937,_EVAL_1469};
  assign _EVAL_318 = _EVAL_818 ? _EVAL_1870 : _EVAL_305;
  assign _EVAL_1189 = _EVAL_1492[15:0];
  assign _EVAL_1517 = _EVAL_1189[15:2];
  assign _EVAL_1556 = _EVAL_1189[15:13];
  assign _EVAL_3234 = _EVAL_1556 == 3'h4;
  assign _EVAL_1021 = _EVAL_1189[6:2];
  assign _EVAL_235 = _EVAL_1021 == 5'h0;
  assign _EVAL_1721 = _EVAL_1189[1:0];
  assign _EVAL_2351 = _EVAL_1721[0];
  assign _EVAL_657 = _EVAL_1721[1];
  assign _EVAL_1045 = _EVAL_235 ? _EVAL_2351 : _EVAL_657;
  assign _EVAL_2099 = _EVAL_657 == _EVAL_2351;
  assign _EVAL_2833 = {_EVAL_1045,_EVAL_2099};
  assign _EVAL_2085 = _EVAL_3234 ? _EVAL_2833 : _EVAL_1721;
  assign _EVAL_876 = {_EVAL_1678,_EVAL_318,_EVAL_1517,_EVAL_2085};
  assign _EVAL_2342 = _EVAL_876[3];
  assign _EVAL_2646 = _EVAL_876[31];
  assign _EVAL_2913 = $signed(_EVAL_2646);
  assign _EVAL_2165 = $unsigned(_EVAL_2913);
  assign _EVAL_2867 = {11{_EVAL_2913}};
  assign _EVAL_3278 = $unsigned(_EVAL_2867);
  assign _EVAL_1948 = _EVAL_876[19:12];
  assign _EVAL_882 = $signed(_EVAL_1948);
  assign _EVAL_1079 = $unsigned(_EVAL_882);
  assign _EVAL_2493 = _EVAL_876[20];
  assign _EVAL_1274 = $signed(_EVAL_2493);
  assign _EVAL_1056 = $unsigned(_EVAL_1274);
  assign _EVAL_3248 = _EVAL_876[30:25];
  assign _EVAL_3014 = _EVAL_876[24:21];
  assign _EVAL_2876 = {_EVAL_2165,_EVAL_3278,_EVAL_1079,_EVAL_1056,_EVAL_3248,_EVAL_3014,1'h0};
  assign _EVAL_860 = $signed(_EVAL_2876);
  assign _EVAL_445 = {8{_EVAL_2913}};
  assign _EVAL_2105 = $unsigned(_EVAL_445);
  assign _EVAL_331 = _EVAL_876[7];
  assign _EVAL_2101 = $signed(_EVAL_331);
  assign _EVAL_829 = $unsigned(_EVAL_2101);
  assign _EVAL_3061 = _EVAL_876[11:8];
  assign _EVAL_1219 = {_EVAL_2165,_EVAL_3278,_EVAL_2105,_EVAL_829,_EVAL_3248,_EVAL_3061,1'h0};
  assign _EVAL_1014 = $signed(_EVAL_1219);
  assign _EVAL_1743 = _EVAL_2342 ? $signed(_EVAL_860) : $signed(_EVAL_1014);
  assign _EVAL_2134 = _EVAL_1492[14];
  assign _EVAL_3361 = _EVAL_1492[12];
  assign _EVAL_2540 = _EVAL_3361 ? 5'h1f : 5'h0;
  assign _EVAL_2709 = _EVAL_1492[6:5];
  assign _EVAL_3159 = _EVAL_1492[2];
  assign _EVAL_756 = _EVAL_1492[11:10];
  assign _EVAL_1588 = _EVAL_1492[4:3];
  assign _EVAL_3212 = {_EVAL_2540,_EVAL_2709,_EVAL_3159,_EVAL_756,_EVAL_1588,1'h0};
  assign _EVAL_2367 = $signed(_EVAL_3212);
  assign _EVAL_1551 = _EVAL_3361 ? 10'h3ff : 10'h0;
  assign _EVAL_2673 = _EVAL_1492[8];
  assign _EVAL_1575 = _EVAL_1492[10:9];
  assign _EVAL_156 = _EVAL_1492[6];
  assign _EVAL_2904 = _EVAL_1492[7];
  assign _EVAL_511 = _EVAL_1492[11];
  assign _EVAL_527 = _EVAL_1492[5:3];
  assign _EVAL_1038 = {_EVAL_1551,_EVAL_2673,_EVAL_1575,_EVAL_156,_EVAL_2904,_EVAL_3159,_EVAL_511,_EVAL_527,1'h0};
  assign _EVAL_604 = $signed(_EVAL_1038);
  assign _EVAL_1362 = _EVAL_2134 ? $signed({{8{_EVAL_2367[12]}},_EVAL_2367}) : $signed(_EVAL_604);
  assign _EVAL_1534 = _EVAL_777 ? $signed(_EVAL_1743) : $signed({{11{_EVAL_1362[20]}},_EVAL_1362});
  assign _EVAL_817 = $signed(_EVAL_158) + $signed(_EVAL_1534);
  assign _EVAL_2890 = $signed(_EVAL_817);
  assign _EVAL_2257 = $unsigned(_EVAL_2890);
  assign _EVAL_922 = ~ _EVAL_2392;
  assign _EVAL_2233 = _EVAL_922 | 32'h7;
  assign _EVAL_3009 = ~ _EVAL_2233;
  assign _EVAL_1096 = {{1'd0}, _EVAL_3009};
  assign _EVAL_462 = _EVAL_1096[31:0];
  assign _EVAL_650 = _EVAL_3009 + 32'h2;
  assign _EVAL_1627 = _EVAL_919 ? _EVAL_462 : _EVAL_650;
  assign _EVAL_2051 = _EVAL_3376[11:7];
  assign _EVAL_189 = _EVAL_2051 & 5'h1b;
  assign _EVAL_1926 = 5'h1 == _EVAL_189;
  assign _EVAL_3324 = _EVAL_3376[7];
  assign _EVAL_2411 = _EVAL_3324 == 1'h0;
  assign _EVAL_925 = _EVAL_2411 & _EVAL_2018;
  assign _EVAL_578 = _EVAL_2227[3:0];
  assign _EVAL_2264 = _EVAL_578 & 4'hd;
  assign _EVAL_2701 = 4'h0 == _EVAL_2264;
  assign _EVAL_3210 = _EVAL_925 & _EVAL_2701;
  assign _EVAL_272 = _EVAL_919 ? _EVAL_1926 : _EVAL_3210;
  assign _EVAL_2977 = _EVAL_272 ? _EVAL_1163 : _EVAL_1243;
  assign _EVAL_803 = _EVAL_2671 ? _EVAL_1627 : _EVAL_2977;
  assign _EVAL_1130 = _EVAL_474 ? _EVAL_2257 : _EVAL_803;
  assign _EVAL_1847 = _EVAL_2410 | _EVAL_1631;
  assign _EVAL_239 = _EVAL_1855 | _EVAL_3106;
  assign _EVAL_240 = _EVAL_1847 | _EVAL_239;
  assign _EVAL_2504 = _EVAL_240 | _EVAL_1143;
  assign _EVAL_683 = _EVAL_2504 | _EVAL_1070;
  assign _EVAL_1111 = _EVAL_2384 & _EVAL_683;
  assign _EVAL_1374 = _EVAL_2227[1];
  assign _EVAL_1029 = _EVAL_1374 == 1'h0;
  assign _EVAL_1281 = _EVAL_2227[3];
  assign _EVAL_2046 = _EVAL_1029 ? _EVAL_2940 : _EVAL_1281;
  assign _EVAL_1621 = _EVAL_2227[2];
  assign _EVAL_3333 = _EVAL_1621 == 1'h0;
  assign _EVAL_955 = _EVAL_1029 ? _EVAL_2980 : _EVAL_3333;
  assign _EVAL_343 = _EVAL_955 & _EVAL_542;
  assign _EVAL_1413 = _EVAL_2046 | _EVAL_343;
  assign _EVAL_477 = $signed(_EVAL_462);
  assign _EVAL_3178 = {_EVAL_995,_EVAL_2227};
  assign _EVAL_830 = _EVAL_3178[1];
  assign _EVAL_3068 = _EVAL_3178[31:16];
  assign _EVAL_540 = _EVAL_3068[15:2];
  assign _EVAL_2921 = _EVAL_3068[15:13];
  assign _EVAL_1759 = _EVAL_2921 == 3'h4;
  assign _EVAL_2266 = _EVAL_3068[6:2];
  assign _EVAL_1828 = _EVAL_2266 == 5'h0;
  assign _EVAL_1028 = _EVAL_3068[1:0];
  assign _EVAL_2425 = _EVAL_1028[0];
  assign _EVAL_1217 = _EVAL_1028[1];
  assign _EVAL_2603 = _EVAL_1828 ? _EVAL_2425 : _EVAL_1217;
  assign _EVAL_2533 = _EVAL_1217 == _EVAL_2425;
  assign _EVAL_3282 = {_EVAL_2603,_EVAL_2533};
  assign _EVAL_896 = _EVAL_1759 ? _EVAL_3282 : _EVAL_1028;
  assign _EVAL_1756 = _EVAL_3178[15:0];
  assign _EVAL_3127 = _EVAL_1756[15:2];
  assign _EVAL_835 = _EVAL_1756[15:13];
  assign _EVAL_1146 = _EVAL_835 == 3'h4;
  assign _EVAL_2878 = _EVAL_1756[6:2];
  assign _EVAL_2599 = _EVAL_2878 == 5'h0;
  assign _EVAL_3341 = _EVAL_1756[1:0];
  assign _EVAL_3136 = _EVAL_3341[0];
  assign _EVAL_2174 = _EVAL_3341[1];
  assign _EVAL_2314 = _EVAL_2599 ? _EVAL_3136 : _EVAL_2174;
  assign _EVAL_766 = _EVAL_2174 == _EVAL_3136;
  assign _EVAL_1211 = {_EVAL_2314,_EVAL_766};
  assign _EVAL_1735 = _EVAL_1146 ? _EVAL_1211 : _EVAL_3341;
  assign _EVAL_1144 = {_EVAL_540,_EVAL_896,_EVAL_3127,_EVAL_1735};
  assign _EVAL_1834 = _EVAL_1144[3];
  assign _EVAL_1069 = _EVAL_1144[31];
  assign _EVAL_648 = $signed(_EVAL_1069);
  assign _EVAL_2258 = $unsigned(_EVAL_648);
  assign _EVAL_2991 = {11{_EVAL_648}};
  assign _EVAL_384 = $unsigned(_EVAL_2991);
  assign _EVAL_3395 = _EVAL_1144[19:12];
  assign _EVAL_1929 = $signed(_EVAL_3395);
  assign _EVAL_2130 = $unsigned(_EVAL_1929);
  assign _EVAL_535 = _EVAL_1144[20];
  assign _EVAL_1567 = $signed(_EVAL_535);
  assign _EVAL_3352 = $unsigned(_EVAL_1567);
  assign _EVAL_1041 = _EVAL_1144[30:25];
  assign _EVAL_680 = _EVAL_1144[24:21];
  assign _EVAL_1643 = {_EVAL_2258,_EVAL_384,_EVAL_2130,_EVAL_3352,_EVAL_1041,_EVAL_680,1'h0};
  assign _EVAL_1720 = $signed(_EVAL_1643);
  assign _EVAL_3238 = {8{_EVAL_648}};
  assign _EVAL_2666 = $unsigned(_EVAL_3238);
  assign _EVAL_2088 = _EVAL_1144[7];
  assign _EVAL_2041 = $signed(_EVAL_2088);
  assign _EVAL_2832 = $unsigned(_EVAL_2041);
  assign _EVAL_1210 = _EVAL_1144[11:8];
  assign _EVAL_1266 = {_EVAL_2258,_EVAL_384,_EVAL_2666,_EVAL_2832,_EVAL_1041,_EVAL_1210,1'h0};
  assign _EVAL_1962 = $signed(_EVAL_1266);
  assign _EVAL_360 = _EVAL_1834 ? $signed(_EVAL_1720) : $signed(_EVAL_1962);
  assign _EVAL_2335 = _EVAL_3178[14];
  assign _EVAL_1829 = _EVAL_3178[12];
  assign _EVAL_763 = _EVAL_1829 ? 5'h1f : 5'h0;
  assign _EVAL_2171 = _EVAL_3178[6:5];
  assign _EVAL_3399 = _EVAL_3178[2];
  assign _EVAL_1975 = _EVAL_3178[11:10];
  assign _EVAL_256 = _EVAL_3178[4:3];
  assign _EVAL_755 = {_EVAL_763,_EVAL_2171,_EVAL_3399,_EVAL_1975,_EVAL_256,1'h0};
  assign _EVAL_2834 = $signed(_EVAL_755);
  assign _EVAL_3379 = _EVAL_1829 ? 10'h3ff : 10'h0;
  assign _EVAL_1116 = _EVAL_3178[8];
  assign _EVAL_313 = _EVAL_3178[10:9];
  assign _EVAL_284 = _EVAL_3178[6];
  assign _EVAL_1346 = _EVAL_3178[7];
  assign _EVAL_1960 = _EVAL_3178[11];
  assign _EVAL_898 = _EVAL_3178[5:3];
  assign _EVAL_1345 = {_EVAL_3379,_EVAL_1116,_EVAL_313,_EVAL_284,_EVAL_1346,_EVAL_3399,_EVAL_1960,_EVAL_898,1'h0};
  assign _EVAL_485 = $signed(_EVAL_1345);
  assign _EVAL_2369 = _EVAL_2335 ? $signed({{8{_EVAL_2834[12]}},_EVAL_2834}) : $signed(_EVAL_485);
  assign _EVAL_1204 = _EVAL_830 ? $signed(_EVAL_360) : $signed({{11{_EVAL_2369[20]}},_EVAL_2369});
  assign _EVAL_573 = $signed(_EVAL_477) + $signed(_EVAL_1204);
  assign _EVAL_1672 = $signed(_EVAL_573);
  assign _EVAL_391 = $unsigned(_EVAL_1672);
  assign _EVAL_1205 = _EVAL_3009 + 32'h4;
  assign _EVAL_1411 = _EVAL_1029 ? _EVAL_650 : _EVAL_1205;
  assign _EVAL_2187 = _EVAL_2227[11:7];
  assign _EVAL_2220 = _EVAL_2187 & 5'h1b;
  assign _EVAL_1528 = 5'h1 == _EVAL_2220;
  assign _EVAL_2060 = _EVAL_2227[7];
  assign _EVAL_1424 = _EVAL_2060 == 1'h0;
  assign _EVAL_416 = _EVAL_1424 & _EVAL_2327;
  assign _EVAL_2872 = _EVAL_995[3:0];
  assign _EVAL_168 = _EVAL_2872 & 4'hd;
  assign _EVAL_1109 = 4'h0 == _EVAL_168;
  assign _EVAL_3056 = _EVAL_416 & _EVAL_1109;
  assign _EVAL_2236 = _EVAL_1029 ? _EVAL_1528 : _EVAL_3056;
  assign _EVAL_566 = _EVAL_2236 ? _EVAL_1163 : _EVAL_1243;
  assign _EVAL_302 = _EVAL_955 ? _EVAL_1411 : _EVAL_566;
  assign _EVAL_1602 = _EVAL_1413 ? _EVAL_391 : _EVAL_302;
  assign _EVAL_3372 = _EVAL_1686 | _EVAL_1564;
  assign _EVAL_1688 = _EVAL_1025 | _EVAL_970;
  assign _EVAL_310 = _EVAL_3372 | _EVAL_1688;
  assign _EVAL_1907 = _EVAL_310 | _EVAL_1159;
  assign _EVAL_1308 = _EVAL_1907 | _EVAL_2306;
  assign _EVAL_1257 = _EVAL_2158 & _EVAL_1308;
  assign _EVAL_2930 = _EVAL_995[1];
  assign _EVAL_2938 = _EVAL_2930 == 1'h0;
  assign _EVAL_3196 = _EVAL_995[3];
  assign _EVAL_1805 = _EVAL_2938 ? _EVAL_2556 : _EVAL_3196;
  assign _EVAL_1300 = _EVAL_995[2];
  assign _EVAL_3098 = _EVAL_1300 == 1'h0;
  assign _EVAL_431 = _EVAL_2938 ? _EVAL_1607 : _EVAL_3098;
  assign _EVAL_2966 = _EVAL_431 & _EVAL_542;
  assign _EVAL_2623 = _EVAL_1805 | _EVAL_2966;
  assign _EVAL_2419 = $signed(_EVAL_650);
  assign _EVAL_581 = {_EVAL_2291,_EVAL_995};
  assign _EVAL_3015 = _EVAL_581[1];
  assign _EVAL_2108 = _EVAL_581[31:16];
  assign _EVAL_1799 = _EVAL_2108[15:2];
  assign _EVAL_3285 = _EVAL_2108[15:13];
  assign _EVAL_2590 = _EVAL_3285 == 3'h4;
  assign _EVAL_939 = _EVAL_2108[6:2];
  assign _EVAL_329 = _EVAL_939 == 5'h0;
  assign _EVAL_1490 = _EVAL_2108[1:0];
  assign _EVAL_473 = _EVAL_1490[0];
  assign _EVAL_2874 = _EVAL_1490[1];
  assign _EVAL_432 = _EVAL_329 ? _EVAL_473 : _EVAL_2874;
  assign _EVAL_2333 = _EVAL_2874 == _EVAL_473;
  assign _EVAL_2140 = {_EVAL_432,_EVAL_2333};
  assign _EVAL_2745 = _EVAL_2590 ? _EVAL_2140 : _EVAL_1490;
  assign _EVAL_1680 = _EVAL_581[15:0];
  assign _EVAL_884 = _EVAL_1680[15:2];
  assign _EVAL_1830 = _EVAL_1680[15:13];
  assign _EVAL_2561 = _EVAL_1830 == 3'h4;
  assign _EVAL_1554 = _EVAL_1680[6:2];
  assign _EVAL_2155 = _EVAL_1554 == 5'h0;
  assign _EVAL_1232 = _EVAL_1680[1:0];
  assign _EVAL_2512 = _EVAL_1232[0];
  assign _EVAL_210 = _EVAL_1232[1];
  assign _EVAL_2644 = _EVAL_2155 ? _EVAL_2512 : _EVAL_210;
  assign _EVAL_2837 = _EVAL_210 == _EVAL_2512;
  assign _EVAL_1187 = {_EVAL_2644,_EVAL_2837};
  assign _EVAL_3312 = _EVAL_2561 ? _EVAL_1187 : _EVAL_1232;
  assign _EVAL_2798 = {_EVAL_1799,_EVAL_2745,_EVAL_884,_EVAL_3312};
  assign _EVAL_1373 = _EVAL_2798[3];
  assign _EVAL_2551 = _EVAL_2798[31];
  assign _EVAL_968 = $signed(_EVAL_2551);
  assign _EVAL_1979 = $unsigned(_EVAL_968);
  assign _EVAL_638 = {11{_EVAL_968}};
  assign _EVAL_768 = $unsigned(_EVAL_638);
  assign _EVAL_3100 = _EVAL_2798[19:12];
  assign _EVAL_1538 = $signed(_EVAL_3100);
  assign _EVAL_2356 = $unsigned(_EVAL_1538);
  assign _EVAL_3294 = _EVAL_2798[20];
  assign _EVAL_3334 = $signed(_EVAL_3294);
  assign _EVAL_244 = $unsigned(_EVAL_3334);
  assign _EVAL_514 = _EVAL_2798[30:25];
  assign _EVAL_2281 = _EVAL_2798[24:21];
  assign _EVAL_3293 = {_EVAL_1979,_EVAL_768,_EVAL_2356,_EVAL_244,_EVAL_514,_EVAL_2281,1'h0};
  assign _EVAL_3286 = $signed(_EVAL_3293);
  assign _EVAL_1059 = {8{_EVAL_968}};
  assign _EVAL_3102 = $unsigned(_EVAL_1059);
  assign _EVAL_3152 = _EVAL_2798[7];
  assign _EVAL_2287 = $signed(_EVAL_3152);
  assign _EVAL_1309 = $unsigned(_EVAL_2287);
  assign _EVAL_1330 = _EVAL_2798[11:8];
  assign _EVAL_1177 = {_EVAL_1979,_EVAL_768,_EVAL_3102,_EVAL_1309,_EVAL_514,_EVAL_1330,1'h0};
  assign _EVAL_2954 = $signed(_EVAL_1177);
  assign _EVAL_2205 = _EVAL_1373 ? $signed(_EVAL_3286) : $signed(_EVAL_2954);
  assign _EVAL_1155 = _EVAL_581[14];
  assign _EVAL_423 = _EVAL_581[12];
  assign _EVAL_2523 = _EVAL_423 ? 5'h1f : 5'h0;
  assign _EVAL_1115 = _EVAL_581[6:5];
  assign _EVAL_2530 = _EVAL_581[2];
  assign _EVAL_1868 = _EVAL_581[11:10];
  assign _EVAL_1455 = _EVAL_581[4:3];
  assign _EVAL_754 = {_EVAL_2523,_EVAL_1115,_EVAL_2530,_EVAL_1868,_EVAL_1455,1'h0};
  assign _EVAL_1752 = $signed(_EVAL_754);
  assign _EVAL_1275 = _EVAL_423 ? 10'h3ff : 10'h0;
  assign _EVAL_3255 = _EVAL_581[8];
  assign _EVAL_555 = _EVAL_581[10:9];
  assign _EVAL_400 = _EVAL_581[6];
  assign _EVAL_863 = _EVAL_581[7];
  assign _EVAL_2290 = _EVAL_581[11];
  assign _EVAL_1082 = _EVAL_581[5:3];
  assign _EVAL_2263 = {_EVAL_1275,_EVAL_3255,_EVAL_555,_EVAL_400,_EVAL_863,_EVAL_2530,_EVAL_2290,_EVAL_1082,1'h0};
  assign _EVAL_2439 = $signed(_EVAL_2263);
  assign _EVAL_2822 = _EVAL_1155 ? $signed({{8{_EVAL_1752[12]}},_EVAL_1752}) : $signed(_EVAL_2439);
  assign _EVAL_3008 = _EVAL_3015 ? $signed(_EVAL_2205) : $signed({{11{_EVAL_2822[20]}},_EVAL_2822});
  assign _EVAL_687 = $signed(_EVAL_2419) + $signed(_EVAL_3008);
  assign _EVAL_1549 = $signed(_EVAL_687);
  assign _EVAL_2490 = $unsigned(_EVAL_1549);
  assign _EVAL_2232 = _EVAL_3009 + 32'h6;
  assign _EVAL_2766 = _EVAL_2938 ? _EVAL_1205 : _EVAL_2232;
  assign _EVAL_2323 = _EVAL_995[11:7];
  assign _EVAL_2965 = _EVAL_2323 & 5'h1b;
  assign _EVAL_3208 = 5'h1 == _EVAL_2965;
  assign _EVAL_1310 = _EVAL_995[7];
  assign _EVAL_1453 = _EVAL_1310 == 1'h0;
  assign _EVAL_203 = _EVAL_1453 & _EVAL_1610;
  assign _EVAL_2964 = _EVAL_2291[3:0];
  assign _EVAL_833 = _EVAL_2964 & 4'hd;
  assign _EVAL_2718 = 4'h0 == _EVAL_833;
  assign _EVAL_1882 = _EVAL_203 & _EVAL_2718;
  assign _EVAL_3410 = _EVAL_2938 ? _EVAL_3208 : _EVAL_1882;
  assign _EVAL_1290 = _EVAL_3410 ? _EVAL_1163 : _EVAL_1243;
  assign _EVAL_1134 = _EVAL_431 ? _EVAL_2766 : _EVAL_1290;
  assign _EVAL_3407 = _EVAL_2623 ? _EVAL_2490 : _EVAL_1134;
  assign _EVAL_2516 = _EVAL_1078 == 1'h0;
  assign _EVAL_2520 = _EVAL_2516 | _EVAL_3063;
  assign _EVAL_3262 = _EVAL_2520 | _EVAL_641;
  assign _EVAL_1572 = _EVAL_3262 | _EVAL_2020;
  assign _EVAL_2309 = _EVAL_1276 & _EVAL_1572;
  assign _EVAL_2163 = _EVAL_2291[1];
  assign _EVAL_2866 = _EVAL_2163 == 1'h0;
  assign _EVAL_3161 = _EVAL_2291[3];
  assign _EVAL_2208 = _EVAL_2866 ? _EVAL_1758 : _EVAL_3161;
  assign _EVAL_3141 = _EVAL_2291[2];
  assign _EVAL_192 = _EVAL_3141 == 1'h0;
  assign _EVAL_3209 = _EVAL_2866 ? _EVAL_1008 : _EVAL_192;
  assign _EVAL_618 = _EVAL_3209 & _EVAL_542;
  assign _EVAL_1315 = _EVAL_2208 | _EVAL_618;
  assign _EVAL_1097 = $signed(_EVAL_1205);
  assign _EVAL_1773 = {_EVAL_1336,_EVAL_2291};
  assign _EVAL_3342 = _EVAL_1773[1];
  assign _EVAL_245 = _EVAL_1773[31:16];
  assign _EVAL_598 = _EVAL_245[15:2];
  assign _EVAL_2895 = _EVAL_245[15:13];
  assign _EVAL_2579 = _EVAL_2895 == 3'h4;
  assign _EVAL_2678 = _EVAL_245[6:2];
  assign _EVAL_3289 = _EVAL_2678 == 5'h0;
  assign _EVAL_2881 = _EVAL_245[1:0];
  assign _EVAL_2702 = _EVAL_2881[0];
  assign _EVAL_1206 = _EVAL_2881[1];
  assign _EVAL_1002 = _EVAL_3289 ? _EVAL_2702 : _EVAL_1206;
  assign _EVAL_1318 = _EVAL_1206 == _EVAL_2702;
  assign _EVAL_229 = {_EVAL_1002,_EVAL_1318};
  assign _EVAL_3277 = _EVAL_2579 ? _EVAL_229 : _EVAL_2881;
  assign _EVAL_1355 = _EVAL_1773[15:0];
  assign _EVAL_2219 = _EVAL_1355[15:2];
  assign _EVAL_1648 = _EVAL_1355[15:13];
  assign _EVAL_1959 = _EVAL_1648 == 3'h4;
  assign _EVAL_1604 = _EVAL_1355[6:2];
  assign _EVAL_3290 = _EVAL_1604 == 5'h0;
  assign _EVAL_2272 = _EVAL_1355[1:0];
  assign _EVAL_1397 = _EVAL_2272[0];
  assign _EVAL_2840 = _EVAL_2272[1];
  assign _EVAL_2909 = _EVAL_3290 ? _EVAL_1397 : _EVAL_2840;
  assign _EVAL_1888 = _EVAL_2840 == _EVAL_1397;
  assign _EVAL_1816 = {_EVAL_2909,_EVAL_1888};
  assign _EVAL_3409 = _EVAL_1959 ? _EVAL_1816 : _EVAL_2272;
  assign _EVAL_2681 = {_EVAL_598,_EVAL_3277,_EVAL_2219,_EVAL_3409};
  assign _EVAL_150 = _EVAL_2681[3];
  assign _EVAL_2382 = _EVAL_2681[31];
  assign _EVAL_870 = $signed(_EVAL_2382);
  assign _EVAL_3041 = $unsigned(_EVAL_870);
  assign _EVAL_2352 = {11{_EVAL_870}};
  assign _EVAL_2355 = $unsigned(_EVAL_2352);
  assign _EVAL_2240 = _EVAL_2681[19:12];
  assign _EVAL_213 = $signed(_EVAL_2240);
  assign _EVAL_1559 = $unsigned(_EVAL_213);
  assign _EVAL_2423 = _EVAL_2681[20];
  assign _EVAL_163 = $signed(_EVAL_2423);
  assign _EVAL_2738 = $unsigned(_EVAL_163);
  assign _EVAL_2960 = _EVAL_2681[30:25];
  assign _EVAL_565 = _EVAL_2681[24:21];
  assign _EVAL_2129 = {_EVAL_3041,_EVAL_2355,_EVAL_1559,_EVAL_2738,_EVAL_2960,_EVAL_565,1'h0};
  assign _EVAL_782 = $signed(_EVAL_2129);
  assign _EVAL_1630 = {8{_EVAL_870}};
  assign _EVAL_1823 = $unsigned(_EVAL_1630);
  assign _EVAL_3185 = _EVAL_2681[7];
  assign _EVAL_1461 = $signed(_EVAL_3185);
  assign _EVAL_276 = $unsigned(_EVAL_1461);
  assign _EVAL_625 = _EVAL_2681[11:8];
  assign _EVAL_1060 = {_EVAL_3041,_EVAL_2355,_EVAL_1823,_EVAL_276,_EVAL_2960,_EVAL_625,1'h0};
  assign _EVAL_3018 = $signed(_EVAL_1060);
  assign _EVAL_3166 = _EVAL_150 ? $signed(_EVAL_782) : $signed(_EVAL_3018);
  assign _EVAL_653 = _EVAL_1773[14];
  assign _EVAL_875 = _EVAL_1773[12];
  assign _EVAL_3396 = _EVAL_875 ? 5'h1f : 5'h0;
  assign _EVAL_2433 = _EVAL_1773[6:5];
  assign _EVAL_2262 = _EVAL_1773[2];
  assign _EVAL_1495 = _EVAL_1773[11:10];
  assign _EVAL_3060 = _EVAL_1773[4:3];
  assign _EVAL_185 = {_EVAL_3396,_EVAL_2433,_EVAL_2262,_EVAL_1495,_EVAL_3060,1'h0};
  assign _EVAL_1162 = $signed(_EVAL_185);
  assign _EVAL_2009 = _EVAL_875 ? 10'h3ff : 10'h0;
  assign _EVAL_2389 = _EVAL_1773[8];
  assign _EVAL_819 = _EVAL_1773[10:9];
  assign _EVAL_1327 = _EVAL_1773[6];
  assign _EVAL_1969 = _EVAL_1773[7];
  assign _EVAL_2814 = _EVAL_1773[11];
  assign _EVAL_2583 = _EVAL_1773[5:3];
  assign _EVAL_3087 = {_EVAL_2009,_EVAL_2389,_EVAL_819,_EVAL_1327,_EVAL_1969,_EVAL_2262,_EVAL_2814,_EVAL_2583,1'h0};
  assign _EVAL_525 = $signed(_EVAL_3087);
  assign _EVAL_3384 = _EVAL_653 ? $signed({{8{_EVAL_1162[12]}},_EVAL_1162}) : $signed(_EVAL_525);
  assign _EVAL_2156 = _EVAL_3342 ? $signed(_EVAL_3166) : $signed({{11{_EVAL_3384[20]}},_EVAL_3384});
  assign _EVAL_3326 = $signed(_EVAL_1097) + $signed(_EVAL_2156);
  assign _EVAL_2803 = $signed(_EVAL_3326);
  assign _EVAL_2079 = $unsigned(_EVAL_2803);
  assign _EVAL_2175 = _EVAL_3009 + 32'h8;
  assign _EVAL_191 = _EVAL_2866 ? _EVAL_2232 : _EVAL_2175;
  assign _EVAL_2376 = _EVAL_2291[11:7];
  assign _EVAL_3377 = _EVAL_2376 & 5'h1b;
  assign _EVAL_842 = 5'h1 == _EVAL_3377;
  assign _EVAL_1887 = _EVAL_2291[7];
  assign _EVAL_1478 = _EVAL_1887 == 1'h0;
  assign _EVAL_1508 = _EVAL_1478 & _EVAL_1642;
  assign _EVAL_2142 = _EVAL_1336[3:0];
  assign _EVAL_2968 = _EVAL_2142 & 4'hd;
  assign _EVAL_3267 = 4'h0 == _EVAL_2968;
  assign _EVAL_2546 = _EVAL_1508 & _EVAL_3267;
  assign _EVAL_1644 = _EVAL_2866 ? _EVAL_842 : _EVAL_2546;
  assign _EVAL_161 = _EVAL_1644 ? _EVAL_1163 : _EVAL_1243;
  assign _EVAL_1579 = _EVAL_3209 ? _EVAL_191 : _EVAL_161;
  assign _EVAL_233 = _EVAL_1315 ? _EVAL_2079 : _EVAL_1579;
  assign _EVAL_1236 = _EVAL_381 & _EVAL_542;
  assign _EVAL_3221 = _EVAL_2451 | _EVAL_1236;
  assign _EVAL_1742 = $signed(_EVAL_2232);
  assign _EVAL_696 = ~ _EVAL_1336;
  assign _EVAL_1662 = _EVAL_696 | 16'h3;
  assign _EVAL_197 = ~ _EVAL_1662;
  assign _EVAL_1657 = {16'h0,_EVAL_197};
  assign _EVAL_3316 = _EVAL_1657[1];
  assign _EVAL_605 = _EVAL_1657[31:16];
  assign _EVAL_1183 = _EVAL_605[15:2];
  assign _EVAL_347 = _EVAL_605[15:13];
  assign _EVAL_193 = _EVAL_347 == 3'h4;
  assign _EVAL_2317 = _EVAL_605[6:2];
  assign _EVAL_546 = _EVAL_2317 == 5'h0;
  assign _EVAL_3142 = _EVAL_605[1:0];
  assign _EVAL_2036 = _EVAL_3142[0];
  assign _EVAL_2585 = _EVAL_3142[1];
  assign _EVAL_1815 = _EVAL_546 ? _EVAL_2036 : _EVAL_2585;
  assign _EVAL_2350 = _EVAL_2585 == _EVAL_2036;
  assign _EVAL_311 = {_EVAL_1815,_EVAL_2350};
  assign _EVAL_2176 = _EVAL_193 ? _EVAL_311 : _EVAL_3142;
  assign _EVAL_1885 = _EVAL_1657[15:0];
  assign _EVAL_2986 = _EVAL_1885[15:2];
  assign _EVAL_2996 = _EVAL_1885[15:13];
  assign _EVAL_517 = _EVAL_2996 == 3'h4;
  assign _EVAL_407 = _EVAL_1885[6:2];
  assign _EVAL_1421 = _EVAL_407 == 5'h0;
  assign _EVAL_3360 = _EVAL_1885[1:0];
  assign _EVAL_2689 = _EVAL_3360[0];
  assign _EVAL_1174 = _EVAL_3360[1];
  assign _EVAL_469 = _EVAL_1421 ? _EVAL_2689 : _EVAL_1174;
  assign _EVAL_1433 = _EVAL_1174 == _EVAL_2689;
  assign _EVAL_307 = {_EVAL_469,_EVAL_1433};
  assign _EVAL_1570 = _EVAL_517 ? _EVAL_307 : _EVAL_3360;
  assign _EVAL_998 = {_EVAL_1183,_EVAL_2176,_EVAL_2986,_EVAL_1570};
  assign _EVAL_2334 = _EVAL_998[3];
  assign _EVAL_2097 = _EVAL_998[31];
  assign _EVAL_1831 = $signed(_EVAL_2097);
  assign _EVAL_1821 = $unsigned(_EVAL_1831);
  assign _EVAL_2871 = {11{_EVAL_1831}};
  assign _EVAL_1361 = $unsigned(_EVAL_2871);
  assign _EVAL_2597 = _EVAL_998[19:12];
  assign _EVAL_268 = $signed(_EVAL_2597);
  assign _EVAL_3260 = $unsigned(_EVAL_268);
  assign _EVAL_3020 = _EVAL_998[20];
  assign _EVAL_188 = $signed(_EVAL_3020);
  assign _EVAL_332 = $unsigned(_EVAL_188);
  assign _EVAL_1027 = _EVAL_998[30:25];
  assign _EVAL_853 = _EVAL_998[24:21];
  assign _EVAL_3193 = {_EVAL_1821,_EVAL_1361,_EVAL_3260,_EVAL_332,_EVAL_1027,_EVAL_853,1'h0};
  assign _EVAL_1444 = $signed(_EVAL_3193);
  assign _EVAL_2739 = {8{_EVAL_1831}};
  assign _EVAL_1098 = $unsigned(_EVAL_2739);
  assign _EVAL_375 = _EVAL_998[7];
  assign _EVAL_2095 = $signed(_EVAL_375);
  assign _EVAL_2606 = $unsigned(_EVAL_2095);
  assign _EVAL_1220 = _EVAL_998[11:8];
  assign _EVAL_2498 = {_EVAL_1821,_EVAL_1361,_EVAL_1098,_EVAL_2606,_EVAL_1027,_EVAL_1220,1'h0};
  assign _EVAL_3382 = $signed(_EVAL_2498);
  assign _EVAL_1367 = _EVAL_2334 ? $signed(_EVAL_1444) : $signed(_EVAL_3382);
  assign _EVAL_2733 = _EVAL_1657[14];
  assign _EVAL_358 = _EVAL_1657[12];
  assign _EVAL_3130 = _EVAL_358 ? 5'h1f : 5'h0;
  assign _EVAL_554 = _EVAL_1657[6:5];
  assign _EVAL_296 = _EVAL_1657[2];
  assign _EVAL_3263 = _EVAL_1657[11:10];
  assign _EVAL_2344 = _EVAL_1657[4:3];
  assign _EVAL_1200 = {_EVAL_3130,_EVAL_554,_EVAL_296,_EVAL_3263,_EVAL_2344,1'h0};
  assign _EVAL_199 = $signed(_EVAL_1200);
  assign _EVAL_3109 = _EVAL_358 ? 10'h3ff : 10'h0;
  assign _EVAL_1818 = _EVAL_1657[8];
  assign _EVAL_2167 = _EVAL_1657[10:9];
  assign _EVAL_2957 = _EVAL_1657[6];
  assign _EVAL_2244 = _EVAL_1657[7];
  assign _EVAL_2650 = _EVAL_1657[11];
  assign _EVAL_615 = _EVAL_1657[5:3];
  assign _EVAL_749 = {_EVAL_3109,_EVAL_1818,_EVAL_2167,_EVAL_2957,_EVAL_2244,_EVAL_296,_EVAL_2650,_EVAL_615,1'h0};
  assign _EVAL_2328 = $signed(_EVAL_749);
  assign _EVAL_1796 = _EVAL_2733 ? $signed({{8{_EVAL_199[12]}},_EVAL_199}) : $signed(_EVAL_2328);
  assign _EVAL_646 = _EVAL_3316 ? $signed(_EVAL_1367) : $signed({{11{_EVAL_1796[20]}},_EVAL_1796});
  assign _EVAL_859 = $signed(_EVAL_1742) + $signed(_EVAL_646);
  assign _EVAL_2788 = $signed(_EVAL_859);
  assign _EVAL_2605 = $unsigned(_EVAL_2788);
  assign _EVAL_2223 = _EVAL_1336[11:7];
  assign _EVAL_1760 = _EVAL_2223 & 5'h1b;
  assign _EVAL_1596 = 5'h1 == _EVAL_1760;
  assign _EVAL_2061 = _EVAL_1596 ? _EVAL_1163 : _EVAL_1243;
  assign _EVAL_3201 = _EVAL_381 ? _EVAL_2175 : _EVAL_2061;
  assign _EVAL_1780 = _EVAL_3221 ? _EVAL_2605 : _EVAL_3201;
  assign _EVAL_757 = _EVAL_2309 ? _EVAL_233 : _EVAL_1780;
  assign _EVAL_1510 = _EVAL_1257 ? _EVAL_3407 : _EVAL_757;
  assign _EVAL_2136 = _EVAL_1111 ? _EVAL_1602 : _EVAL_1510;
  assign _EVAL_690 = _EVAL_2139 ? _EVAL_1130 : _EVAL_2136;
  assign _EVAL_1260 = _EVAL_2528[1];
  assign _EVAL_820 = _EVAL_3338[15];
  assign _EVAL_997 = _EVAL_1260 & _EVAL_820;
  assign _EVAL_417 = _EVAL_2270[19:5];
  assign _EVAL_647 = _EVAL_2402[15:1];
  assign _EVAL_2894 = _EVAL_417 == _EVAL_647;
  assign _EVAL_572 = _EVAL_997 & _EVAL_2894;
  assign _EVAL_2388 = _EVAL_3338[14];
  assign _EVAL_907 = _EVAL_1260 & _EVAL_2388;
  assign _EVAL_2662 = _EVAL_446[19:5];
  assign _EVAL_889 = _EVAL_2662 == _EVAL_647;
  assign _EVAL_1909 = _EVAL_907 & _EVAL_889;
  assign _EVAL_2424 = _EVAL_3338[13];
  assign _EVAL_3287 = _EVAL_1260 & _EVAL_2424;
  assign _EVAL_341 = _EVAL_3187[19:5];
  assign _EVAL_2898 = _EVAL_341 == _EVAL_647;
  assign _EVAL_335 = _EVAL_3287 & _EVAL_2898;
  assign _EVAL_3153 = _EVAL_3338[12];
  assign _EVAL_2994 = _EVAL_1260 & _EVAL_3153;
  assign _EVAL_2724 = _EVAL_1152[19:5];
  assign _EVAL_243 = _EVAL_2724 == _EVAL_647;
  assign _EVAL_2135 = _EVAL_2994 & _EVAL_243;
  assign _EVAL_3128 = _EVAL_3338[11];
  assign _EVAL_3346 = _EVAL_1260 & _EVAL_3128;
  assign _EVAL_1946 = _EVAL_794[19:5];
  assign _EVAL_1705 = _EVAL_1946 == _EVAL_647;
  assign _EVAL_3048 = _EVAL_3346 & _EVAL_1705;
  assign _EVAL_2370 = _EVAL_3338[10];
  assign _EVAL_1617 = _EVAL_1260 & _EVAL_2370;
  assign _EVAL_2400 = _EVAL_397[19:5];
  assign _EVAL_270 = _EVAL_2400 == _EVAL_647;
  assign _EVAL_1094 = _EVAL_1617 & _EVAL_270;
  assign _EVAL_753 = _EVAL_3338[9];
  assign _EVAL_1218 = _EVAL_1260 & _EVAL_753;
  assign _EVAL_1687 = _EVAL_722[19:5];
  assign _EVAL_1354 = _EVAL_1687 == _EVAL_647;
  assign _EVAL_2405 = _EVAL_1218 & _EVAL_1354;
  assign _EVAL_3373 = _EVAL_3338[8];
  assign _EVAL_815 = _EVAL_1260 & _EVAL_3373;
  assign _EVAL_2757 = _EVAL_2746[19:5];
  assign _EVAL_149 = _EVAL_2757 == _EVAL_647;
  assign _EVAL_1436 = _EVAL_815 & _EVAL_149;
  assign _EVAL_2444 = _EVAL_3338[7];
  assign _EVAL_816 = _EVAL_1260 & _EVAL_2444;
  assign _EVAL_2936 = _EVAL_1352[19:5];
  assign _EVAL_1428 = _EVAL_2936 == _EVAL_647;
  assign _EVAL_3030 = _EVAL_816 & _EVAL_1428;
  assign _EVAL_1974 = _EVAL_3338[6];
  assign _EVAL_2507 = _EVAL_1260 & _EVAL_1974;
  assign _EVAL_1026 = _EVAL_253[19:5];
  assign _EVAL_1524 = _EVAL_1026 == _EVAL_647;
  assign _EVAL_569 = _EVAL_2507 & _EVAL_1524;
  assign _EVAL_1691 = _EVAL_3338[5];
  assign _EVAL_594 = _EVAL_1260 & _EVAL_1691;
  assign _EVAL_977 = _EVAL_2170[19:5];
  assign _EVAL_3218 = _EVAL_977 == _EVAL_647;
  assign _EVAL_2146 = _EVAL_594 & _EVAL_3218;
  assign _EVAL_2297 = _EVAL_3338[4];
  assign _EVAL_2217 = _EVAL_1260 & _EVAL_2297;
  assign _EVAL_221 = _EVAL_1175[19:5];
  assign _EVAL_678 = _EVAL_221 == _EVAL_647;
  assign _EVAL_3275 = _EVAL_2217 & _EVAL_678;
  assign _EVAL_2607 = _EVAL_3338[3];
  assign _EVAL_2839 = _EVAL_1260 & _EVAL_2607;
  assign _EVAL_2277 = _EVAL_3198[19:5];
  assign _EVAL_767 = _EVAL_2277 == _EVAL_647;
  assign _EVAL_2740 = _EVAL_2839 & _EVAL_767;
  assign _EVAL_2111 = _EVAL_3338[2];
  assign _EVAL_2541 = _EVAL_1260 & _EVAL_2111;
  assign _EVAL_1539 = _EVAL_492[19:5];
  assign _EVAL_479 = _EVAL_1539 == _EVAL_647;
  assign _EVAL_420 = _EVAL_2541 & _EVAL_479;
  assign _EVAL_990 = _EVAL_3338[1];
  assign _EVAL_2427 = _EVAL_1260 & _EVAL_990;
  assign _EVAL_1729 = _EVAL_1487[19:5];
  assign _EVAL_2373 = _EVAL_1729 == _EVAL_647;
  assign _EVAL_2495 = _EVAL_2427 & _EVAL_2373;
  assign _EVAL_2261 = _EVAL_3338[0];
  assign _EVAL_1734 = _EVAL_1260 & _EVAL_2261;
  assign _EVAL_2005 = _EVAL_856[19:5];
  assign _EVAL_1808 = _EVAL_2005 == _EVAL_647;
  assign _EVAL_3189 = _EVAL_1734 & _EVAL_1808;
  assign _EVAL_439 = {_EVAL_3030,_EVAL_569,_EVAL_2146,_EVAL_3275,_EVAL_2740,_EVAL_420,_EVAL_2495,_EVAL_3189};
  assign _EVAL_3329 = {_EVAL_572,_EVAL_1909,_EVAL_335,_EVAL_2135,_EVAL_3048,_EVAL_1094,_EVAL_2405,_EVAL_1436,_EVAL_439};
  assign _EVAL_2063 = _EVAL_3329 != 16'h0;
  assign _EVAL_1503 = _EVAL_2063 == 1'h0;
  assign _EVAL_3230 = _EVAL_3189 ? _EVAL_856 : 52'h0;
  assign _EVAL_1363 = _EVAL_2495 ? _EVAL_1487 : 52'h0;
  assign _EVAL_3274 = _EVAL_3230 | _EVAL_1363;
  assign _EVAL_1863 = _EVAL_420 ? _EVAL_492 : 52'h0;
  assign _EVAL_3116 = _EVAL_3274 | _EVAL_1863;
  assign _EVAL_1766 = _EVAL_2740 ? _EVAL_3198 : 52'h0;
  assign _EVAL_2729 = _EVAL_3116 | _EVAL_1766;
  assign _EVAL_2948 = _EVAL_3275 ? _EVAL_1175 : 52'h0;
  assign _EVAL_1599 = _EVAL_2729 | _EVAL_2948;
  assign _EVAL_3245 = _EVAL_2146 ? _EVAL_2170 : 52'h0;
  assign _EVAL_3151 = _EVAL_1599 | _EVAL_3245;
  assign _EVAL_1940 = _EVAL_569 ? _EVAL_253 : 52'h0;
  assign _EVAL_1937 = _EVAL_3151 | _EVAL_1940;
  assign _EVAL_2857 = _EVAL_3030 ? _EVAL_1352 : 52'h0;
  assign _EVAL_552 = _EVAL_1937 | _EVAL_2857;
  assign _EVAL_176 = _EVAL_1436 ? _EVAL_2746 : 52'h0;
  assign _EVAL_1178 = _EVAL_552 | _EVAL_176;
  assign _EVAL_1197 = _EVAL_2405 ? _EVAL_722 : 52'h0;
  assign _EVAL_2162 = _EVAL_1178 | _EVAL_1197;
  assign _EVAL_2343 = _EVAL_1094 ? _EVAL_397 : 52'h0;
  assign _EVAL_1561 = _EVAL_2162 | _EVAL_2343;
  assign _EVAL_654 = _EVAL_3048 ? _EVAL_794 : 52'h0;
  assign _EVAL_936 = _EVAL_1561 | _EVAL_654;
  assign _EVAL_3025 = _EVAL_2135 ? _EVAL_1152 : 52'h0;
  assign _EVAL_2896 = _EVAL_936 | _EVAL_3025;
  assign _EVAL_2253 = _EVAL_335 ? _EVAL_3187 : 52'h0;
  assign _EVAL_1963 = _EVAL_2896 | _EVAL_2253;
  assign _EVAL_389 = _EVAL_1909 ? _EVAL_446 : 52'h0;
  assign _EVAL_941 = _EVAL_1963 | _EVAL_389;
  assign _EVAL_1679 = _EVAL_572 ? _EVAL_2270 : 52'h0;
  assign _EVAL_1540 = _EVAL_941 | _EVAL_1679;
  assign _EVAL_1933 = _EVAL_1540[51:20];
  assign _EVAL_183 = _EVAL_1933[21];
  assign _EVAL_3049 = _EVAL_2402[21];
  assign _EVAL_413 = _EVAL_183 == _EVAL_3049;
  assign _EVAL_1007 = _EVAL_2402[31:21];
  assign _EVAL_1634 = _EVAL_2402[22];
  assign _EVAL_2552 = _EVAL_1634 ^ _EVAL_3049;
  assign _EVAL_2519 = _EVAL_1933[22];
  assign _EVAL_541 = _EVAL_2552 ^ _EVAL_2519;
  assign _EVAL_1289 = _EVAL_1007 - 11'h1;
  assign _EVAL_1396 = _EVAL_1007 + 11'h1;
  assign _EVAL_2403 = _EVAL_541 ? _EVAL_1289 : _EVAL_1396;
  assign _EVAL_2159 = _EVAL_413 ? _EVAL_1007 : _EVAL_2403;
  assign _EVAL_2301 = _EVAL_1503 ? 11'h0 : _EVAL_2159;
  assign _EVAL_241 = _EVAL_1933[20:0];
  assign _EVAL_1432 = {_EVAL_2301,_EVAL_241};
  assign _EVAL_519 = ~ _EVAL_2402;
  assign _EVAL_895 = _EVAL_519 | 32'h7;
  assign _EVAL_617 = ~ _EVAL_895;
  assign _EVAL_811 = _EVAL_617 + 32'h8;
  assign _EVAL_710 = _EVAL_2063 ? 32'h0 : _EVAL_811;
  assign _EVAL_3356 = _EVAL_1432 | _EVAL_710;
  assign _EVAL_1099 = _EVAL_2843 ? _EVAL_2392 : _EVAL_3356;
  assign _EVAL_175 = _EVAL_3296 ? _EVAL_690 : _EVAL_1099;
  assign _EVAL_2690 = _EVAL_175[31:1];
  assign _EVAL_2754 = _EVAL_2690[14:0];
  assign _EVAL_791 = _EVAL_2754[8:0];
  assign _EVAL_3259 = {_EVAL_2172,_EVAL_791};
  assign _EVAL_2131 = _EVAL_3259[8:0];
  assign _EVAL_2660 = _EVAL_2131[3:0];
  assign _EVAL_436 = _EVAL_2131[8:4];
  assign _EVAL_3301 = {_EVAL_2660,_EVAL_436};
  assign _EVAL_770 = _EVAL_3259[17:9];
  assign _EVAL_2704 = _EVAL_770[4:0];
  assign _EVAL_408 = _EVAL_770[8:5];
  assign _EVAL_2985 = {_EVAL_2704,_EVAL_408};
  assign _EVAL_1123 = _EVAL_3301 ^ _EVAL_2985;
  assign _EVAL_2958 = _EVAL_2950[70];
  assign _EVAL_3028 = _EVAL_2950[66];
  assign _EVAL_1536 = _EVAL_2950[63];
  assign _EVAL_1230 = _EVAL_2950[59];
  assign _EVAL_3012 = _EVAL_2950[56];
  assign _EVAL_2166 = _EVAL_2950[52];
  assign _EVAL_1695 = _EVAL_2950[49];
  assign _EVAL_1353 = _EVAL_2950[45];
  assign _EVAL_846 = _EVAL_2950[42];
  assign _EVAL_2612 = _EVAL_2950[38];
  assign _EVAL_1117 = _EVAL_2950[35];
  assign _EVAL_380 = {_EVAL_1695,_EVAL_1353,_EVAL_846,_EVAL_2612,_EVAL_1117};
  assign _EVAL_2907 = _EVAL_2950[31];
  assign _EVAL_1273 = _EVAL_2950[28];
  assign _EVAL_2782 = _EVAL_2950[24];
  assign _EVAL_695 = _EVAL_2950[21];
  assign _EVAL_698 = _EVAL_2950[17];
  assign _EVAL_1087 = _EVAL_2950[14];
  assign _EVAL_2595 = _EVAL_2950[10];
  assign _EVAL_3057 = _EVAL_2950[7];
  assign _EVAL_810 = _EVAL_2950[3];
  assign _EVAL_2657 = _EVAL_2950[0];
  assign _EVAL_1628 = {_EVAL_2907,_EVAL_1273,_EVAL_2782,_EVAL_695,_EVAL_698,_EVAL_1087,_EVAL_2595,_EVAL_3057,_EVAL_810,_EVAL_2657};
  assign _EVAL_878 = _EVAL_2235[14:0];
  assign _EVAL_3026 = {_EVAL_2958,_EVAL_3028,_EVAL_1536,_EVAL_1230,_EVAL_3012,_EVAL_2166,_EVAL_380,_EVAL_1628,_EVAL_878};
  assign _EVAL_484 = _EVAL_3026[8:0];
  assign _EVAL_2107 = _EVAL_484[4:0];
  assign _EVAL_1403 = _EVAL_484[8:5];
  assign _EVAL_1782 = {_EVAL_2107,_EVAL_1403};
  assign _EVAL_2604 = _EVAL_3026[17:9];
  assign _EVAL_1898 = _EVAL_2604[5:0];
  assign _EVAL_157 = _EVAL_2604[8:6];
  assign _EVAL_2641 = {_EVAL_1898,_EVAL_157};
  assign _EVAL_1891 = _EVAL_1782 ^ _EVAL_2641;
  assign _EVAL_2511 = _EVAL_2542__EVAL_2543_data;
  assign _EVAL_2967 = _EVAL_2531[34];
  assign _EVAL_1068 = {MaxPeriodFibonacciLFSR__EVAL_12,MaxPeriodFibonacciLFSR__EVAL_11,MaxPeriodFibonacciLFSR__EVAL_3,MaxPeriodFibonacciLFSR__EVAL_16,MaxPeriodFibonacciLFSR__EVAL_8,MaxPeriodFibonacciLFSR__EVAL_10,MaxPeriodFibonacciLFSR__EVAL_14,MaxPeriodFibonacciLFSR__EVAL_7};
  assign _EVAL_1172 = {MaxPeriodFibonacciLFSR__EVAL_0,MaxPeriodFibonacciLFSR__EVAL_17,MaxPeriodFibonacciLFSR__EVAL_1,MaxPeriodFibonacciLFSR__EVAL,MaxPeriodFibonacciLFSR__EVAL_5,MaxPeriodFibonacciLFSR__EVAL_4,MaxPeriodFibonacciLFSR__EVAL_6,MaxPeriodFibonacciLFSR__EVAL_2,_EVAL_1068};
  assign _EVAL_822 = _EVAL_1172[0];
  assign _EVAL_672 = _EVAL_1172[1];
  assign _EVAL_493 = _EVAL_1172[2];
  assign _EVAL_3272 = _EVAL_1172[3];
  assign _EVAL_3157 = _EVAL_1172[4];
  assign _EVAL_2194 = _EVAL_1172[5];
  assign _EVAL_299 = _EVAL_1172[6];
  assign _EVAL_1489 = _EVAL_1172[7];
  assign _EVAL_686 = _EVAL_1172[8];
  assign _EVAL_2414 = _EVAL_1172[9];
  assign _EVAL_200 = _EVAL_1172[10];
  assign _EVAL_1016 = _EVAL_1172[11];
  assign _EVAL_1089 = _EVAL_1172[12];
  assign _EVAL_2000 = _EVAL_1172[13];
  assign _EVAL_2316 = _EVAL_1172[14];
  assign _EVAL_2779 = _EVAL_1172[15];
  assign _EVAL_2380 = {_EVAL_686,_EVAL_2414,_EVAL_200,_EVAL_1016,_EVAL_1089,_EVAL_2000,_EVAL_2316,_EVAL_2779};
  assign _EVAL_2359 = {_EVAL_822,_EVAL_672,_EVAL_493,_EVAL_3272,_EVAL_3157,_EVAL_2194,_EVAL_299,_EVAL_1489,_EVAL_2380};
  assign _EVAL_1317 = _EVAL_2359[3:0];
  assign _EVAL_616 = 16'h1 << _EVAL_1317;
  assign _EVAL_3188 = _EVAL_2133 & _EVAL_1926;
  assign _EVAL_844 = _EVAL_2293 & _EVAL_3210;
  assign _EVAL_2412 = _EVAL_3188 | _EVAL_844;
  assign _EVAL_996 = _EVAL_2518 & _EVAL_2412;
  assign _EVAL_2039 = _EVAL_204 == 1'h0;
  assign _EVAL_275 = _EVAL_2039 & _EVAL_2384;
  assign _EVAL_1113 = _EVAL_2410 & _EVAL_1528;
  assign _EVAL_522 = _EVAL_1631 & _EVAL_3056;
  assign _EVAL_632 = _EVAL_1113 | _EVAL_522;
  assign _EVAL_1184 = _EVAL_275 & _EVAL_632;
  assign _EVAL_1049 = _EVAL_996 | _EVAL_1184;
  assign _EVAL_1689 = _EVAL_867 == 1'h0;
  assign _EVAL_716 = _EVAL_1689 & _EVAL_2158;
  assign _EVAL_960 = _EVAL_1686 & _EVAL_3208;
  assign _EVAL_437 = _EVAL_1564 & _EVAL_1882;
  assign _EVAL_2995 = _EVAL_960 | _EVAL_437;
  assign _EVAL_805 = _EVAL_716 & _EVAL_2995;
  assign _EVAL_1081 = _EVAL_1049 | _EVAL_805;
  assign _EVAL_715 = _EVAL_2531[66];
  assign _EVAL_2150 = _EVAL_2531[63];
  assign _EVAL_2193 = _EVAL_2531[59];
  assign _EVAL_2824 = _EVAL_2531[56];
  assign _EVAL_2652 = _EVAL_2531[52];
  assign _EVAL_966 = _EVAL_2531[42];
  assign _EVAL_373 = _EVAL_2531[38];
  assign _EVAL_2572 = _EVAL_2531[35];
  assign _EVAL_2345 = {_EVAL_3266,_EVAL_2049,_EVAL_966,_EVAL_373,_EVAL_2572};
  assign _EVAL_3115 = _EVAL_2531[31];
  assign _EVAL_1435 = _EVAL_2531[21];
  assign _EVAL_1044 = _EVAL_2531[17];
  assign _EVAL_2037 = _EVAL_2531[14];
  assign _EVAL_2256 = _EVAL_2531[10];
  assign _EVAL_917 = _EVAL_2531[7];
  assign _EVAL_2239 = _EVAL_2531[3];
  assign _EVAL_1238 = {_EVAL_3115,_EVAL_3139,_EVAL_2387,_EVAL_1435,_EVAL_1044,_EVAL_2037,_EVAL_2256,_EVAL_917,_EVAL_2239,_EVAL_2553};
  assign _EVAL_1864 = {_EVAL_1500,_EVAL_715,_EVAL_2150,_EVAL_2193,_EVAL_2824,_EVAL_2652,_EVAL_2345,_EVAL_1238,_EVAL_2754};
  assign _EVAL_453 = _EVAL_1864[8:0];
  assign _EVAL_3097 = _EVAL_453[4:0];
  assign _EVAL_845 = _EVAL_453[8:5];
  assign _EVAL_2477 = {_EVAL_3097,_EVAL_845};
  assign _EVAL_1075 = _EVAL_1864[17:9];
  assign _EVAL_712 = _EVAL_1075[5:0];
  assign _EVAL_3347 = _EVAL_1075[8:6];
  assign _EVAL_2787 = {_EVAL_712,_EVAL_3347};
  assign _EVAL_288 = _EVAL_2477 ^ _EVAL_2787;
  assign _EVAL_560 = _EVAL_1864[26:18];
  assign _EVAL_2903 = _EVAL_560[6:0];
  assign _EVAL_2161 = _EVAL_560[8:7];
  assign _EVAL_2500 = {_EVAL_2903,_EVAL_2161};
  assign _EVAL_2048 = _EVAL_288 ^ _EVAL_2500;
  assign _EVAL_1131 = _EVAL_1864[35:27];
  assign _EVAL_2125 = _EVAL_1131[7:0];
  assign _EVAL_2186 = _EVAL_1131[8:8];
  assign _EVAL_261 = {_EVAL_2125,_EVAL_2186};
  assign _EVAL_2564 = _EVAL_2048 ^ _EVAL_261;
  assign _EVAL_1213 = predictor_Queue__EVAL_0[2];
  assign _EVAL_1160 = _EVAL_1213 == 1'h0;
  assign _EVAL_2711 = _EVAL_607 == 1'h0;
  assign _EVAL_1763 = _EVAL_2711 & _EVAL_3105;
  assign _EVAL_2949 = _EVAL_972 == 1'h0;
  assign _EVAL_2797 = _EVAL_2168[1];
  assign _EVAL_2993 = _EVAL_2168[0];
  assign _EVAL_165 = _EVAL_2797 == _EVAL_2993;
  assign _EVAL_2559 = _EVAL_306[2];
  assign _EVAL_1822 = _EVAL_2559 == 1'h0;
  assign _EVAL_3236 = _EVAL_947 & _EVAL_1822;
  assign _EVAL_1379 = _EVAL_314[0];
  assign _EVAL_543 = _EVAL_3236 & _EVAL_1379;
  assign _EVAL_2554 = _EVAL_2785[63:48];
  assign _EVAL_368 = _EVAL_2554[15:2];
  assign _EVAL_703 = _EVAL_2554[15:13];
  assign _EVAL_994 = _EVAL_703 == 3'h4;
  assign _EVAL_2147 = _EVAL_2554[6:2];
  assign _EVAL_1800 = _EVAL_2147 == 5'h0;
  assign _EVAL_3239 = _EVAL_2554[1:0];
  assign _EVAL_827 = _EVAL_3239[0];
  assign _EVAL_427 = _EVAL_3239[1];
  assign _EVAL_2706 = _EVAL_1800 ? _EVAL_827 : _EVAL_427;
  assign _EVAL_2616 = _EVAL_427 == _EVAL_827;
  assign _EVAL_1249 = {_EVAL_2706,_EVAL_2616};
  assign _EVAL_3034 = _EVAL_994 ? _EVAL_1249 : _EVAL_3239;
  assign _EVAL_781 = _EVAL_2785[47:32];
  assign _EVAL_237 = _EVAL_781[15:2];
  assign _EVAL_190 = _EVAL_781[15:13];
  assign _EVAL_836 = _EVAL_190 == 3'h4;
  assign _EVAL_2951 = _EVAL_781[6:2];
  assign _EVAL_3244 = _EVAL_2951 == 5'h0;
  assign _EVAL_504 = _EVAL_781[1:0];
  assign _EVAL_1126 = _EVAL_504[0];
  assign _EVAL_1104 = _EVAL_504[1];
  assign _EVAL_3297 = _EVAL_3244 ? _EVAL_1126 : _EVAL_1104;
  assign _EVAL_269 = _EVAL_1104 == _EVAL_1126;
  assign _EVAL_3223 = {_EVAL_3297,_EVAL_269};
  assign _EVAL_265 = _EVAL_836 ? _EVAL_3223 : _EVAL_504;
  assign _EVAL_1431 = _EVAL_2785[31:16];
  assign _EVAL_1598 = _EVAL_1431[15:2];
  assign _EVAL_1063 = _EVAL_1431[15:13];
  assign _EVAL_2687 = _EVAL_1063 == 3'h4;
  assign _EVAL_2418 = _EVAL_1431[6:2];
  assign _EVAL_1294 = _EVAL_2418 == 5'h0;
  assign _EVAL_1658 = _EVAL_1431[1:0];
  assign _EVAL_915 = _EVAL_1658[0];
  assign _EVAL_1383 = _EVAL_1658[1];
  assign _EVAL_929 = _EVAL_1294 ? _EVAL_915 : _EVAL_1383;
  assign _EVAL_2567 = _EVAL_1383 == _EVAL_915;
  assign _EVAL_2254 = {_EVAL_929,_EVAL_2567};
  assign _EVAL_913 = _EVAL_2687 ? _EVAL_2254 : _EVAL_1658;
  assign _EVAL_3197 = _EVAL_2785[15:0];
  assign _EVAL_2237 = _EVAL_3197[15:2];
  assign _EVAL_3369 = _EVAL_3197[15:13];
  assign _EVAL_3242 = _EVAL_3369 == 3'h4;
  assign _EVAL_670 = _EVAL_3197[6:2];
  assign _EVAL_2199 = _EVAL_670 == 5'h0;
  assign _EVAL_3389 = _EVAL_3197[1:0];
  assign _EVAL_2675 = _EVAL_3389[0];
  assign _EVAL_3090 = _EVAL_3389[1];
  assign _EVAL_1669 = _EVAL_2199 ? _EVAL_2675 : _EVAL_3090;
  assign _EVAL_862 = _EVAL_3090 == _EVAL_2675;
  assign _EVAL_472 = {_EVAL_1669,_EVAL_862};
  assign _EVAL_2688 = _EVAL_3242 ? _EVAL_472 : _EVAL_3389;
  assign _EVAL_1641 = {_EVAL_368,_EVAL_3034,_EVAL_237,_EVAL_265,_EVAL_1598,_EVAL_913,_EVAL_2237,_EVAL_2688};
  assign _EVAL_3247 = _EVAL_543 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_2826 = _EVAL_3247[7:0];
  assign _EVAL_2271 = _EVAL_54 | _EVAL_80;
  assign _EVAL_575 = _EVAL_89[2:0];
  assign _EVAL_965 = _EVAL_575 == 3'h0;
  assign _EVAL_2741 = _EVAL_2271 | _EVAL_965;
  assign _EVAL_3381 = _EVAL_2518 & _EVAL_2789;
  assign _EVAL_222 = _EVAL_275 & _EVAL_239;
  assign _EVAL_3021 = _EVAL_3381 | _EVAL_222;
  assign _EVAL_2614 = _EVAL_2950[22];
  assign _EVAL_1645 = _EVAL_2950[20];
  assign _EVAL_3029 = _EVAL_2950[19];
  assign _EVAL_2008 = _EVAL_2950[18];
  assign _EVAL_635 = _EVAL_2950[16];
  assign _EVAL_2829 = _EVAL_2950[15];
  assign _EVAL_2064 = _EVAL_2950[12];
  assign _EVAL_1037 = _EVAL_2950[11];
  assign _EVAL_1794 = _EVAL_2950[9];
  assign _EVAL_219 = _EVAL_2950[6];
  assign _EVAL_487 = _EVAL_2950[5];
  assign _EVAL_2911 = _EVAL_2950[1];
  assign _EVAL_2568 = {_EVAL_2595,_EVAL_1794,_EVAL_3057,_EVAL_219,_EVAL_487,_EVAL_810,_EVAL_3348,_EVAL_2911,_EVAL_2657};
  assign _EVAL_2143 = {_EVAL_2614,_EVAL_1645,_EVAL_3029,_EVAL_2008,_EVAL_635,_EVAL_2829,_EVAL_1087,_EVAL_2064,_EVAL_1037,_EVAL_2568};
  assign _EVAL_1006 = _EVAL_2235[8:0];
  assign _EVAL_326 = {_EVAL_2143,_EVAL_1006};
  assign _EVAL_717 = _EVAL_326[8:0];
  assign _EVAL_1376 = _EVAL_2531[15];
  assign _EVAL_2434 = _EVAL_2531[13];
  assign _EVAL_1931 = _EVAL_2531[11];
  assign _EVAL_843 = {_EVAL_1376,_EVAL_2037,_EVAL_2434,_EVAL_3388,_EVAL_1931};
  assign _EVAL_711 = _EVAL_956 | _EVAL_336;
  assign _EVAL_2508 = _EVAL_1245 & _EVAL_711;
  assign _EVAL_2922 = _EVAL_2950[112];
  assign _EVAL_1616 = _EVAL_2950[105];
  assign _EVAL_2138 = _EVAL_2950[98];
  assign _EVAL_1697 = _EVAL_2950[92];
  assign _EVAL_2279 = _EVAL_2950[85];
  assign _EVAL_441 = _EVAL_2950[79];
  assign _EVAL_2879 = _EVAL_2950[72];
  assign _EVAL_1694 = _EVAL_2950[65];
  assign _EVAL_623 = _EVAL_2950[46];
  assign _EVAL_587 = _EVAL_2950[39];
  assign _EVAL_2211 = _EVAL_2950[32];
  assign _EVAL_153 = _EVAL_2950[26];
  assign _EVAL_3380 = _EVAL_2950[13];
  assign _EVAL_2635 = {_EVAL_2166,_EVAL_623,_EVAL_587,_EVAL_2211,_EVAL_153,_EVAL_3029,_EVAL_3380,_EVAL_219,_EVAL_2657};
  assign _EVAL_676 = {_EVAL_2922,_EVAL_1616,_EVAL_2138,_EVAL_1697,_EVAL_2279,_EVAL_441,_EVAL_2879,_EVAL_1694,_EVAL_1230,_EVAL_2635};
  assign _EVAL_1990 = {_EVAL_676,_EVAL_1006};
  assign _EVAL_1019 = _EVAL_1990[8:0];
  assign _EVAL_590 = _EVAL_1019[5:0];
  assign _EVAL_1739 = _EVAL_1019[8:6];
  assign _EVAL_2496 = {_EVAL_590,_EVAL_1739};
  assign _EVAL_1404 = _EVAL_1990[17:9];
  assign _EVAL_1683 = _EVAL_1404[6:0];
  assign _EVAL_2463 = _EVAL_1404[8:7];
  assign _EVAL_629 = {_EVAL_1683,_EVAL_2463};
  assign _EVAL_729 = _EVAL_2496 ^ _EVAL_629;
  assign _EVAL_1708 = _EVAL_2292 & _EVAL_1176;
  assign _EVAL_976 = _EVAL_3173 == 1'h0;
  assign _EVAL_3004 = _EVAL_1708 & _EVAL_976;
  assign _EVAL_460 = _EVAL_155 & _EVAL_2806;
  assign _EVAL_147 = _EVAL_1199 | _EVAL_460;
  assign _EVAL_2636 = _EVAL_254 == _EVAL_2248;
  assign _EVAL_813 = _EVAL_3054 & _EVAL_2636;
  assign _EVAL_626 = _EVAL_813 ? 3'h4 : 3'h0;
  assign _EVAL_2584 = _EVAL_254 - _EVAL_2248;
  assign _EVAL_1468 = {{1'd0}, _EVAL_2584};
  assign _EVAL_223 = _EVAL_626 | _EVAL_1468;
  assign _EVAL_1778 = _EVAL_223 + 3'h1;
  assign _EVAL_1306 = ~ _EVAL_1778;
  assign _EVAL_350 = _EVAL_2949 == 1'h0;
  assign _EVAL_759 = ~ _EVAL_350;
  assign _EVAL_2747 = {{3'd0}, _EVAL_759};
  assign _EVAL_495 = _EVAL_1306 | _EVAL_2747;
  assign _EVAL_1297 = ~ _EVAL_495;
  assign _EVAL_2743 = _EVAL_1297[2:0];
  assign _EVAL_3302 = _EVAL_2743 == 3'h0;
  assign _EVAL_2071 = _EVAL_2359[15];
  assign _EVAL_1514 = _EVAL_2743 == 3'h1;
  assign _EVAL_851 = _EVAL_2359[14];
  assign _EVAL_444 = _EVAL_2743 == 3'h2;
  assign _EVAL_901 = _EVAL_2359[13];
  assign _EVAL_3066 = _EVAL_444 | _EVAL_901;
  assign _EVAL_665 = _EVAL_851 & _EVAL_3066;
  assign _EVAL_2255 = _EVAL_1514 | _EVAL_665;
  assign _EVAL_2188 = _EVAL_2071 & _EVAL_2255;
  assign _EVAL_945 = _EVAL_3302 | _EVAL_2188;
  assign _EVAL_2360 = _EVAL_147 & _EVAL_945;
  assign _EVAL_2783 = _EVAL_3004 & _EVAL_2360;
  assign _EVAL_693 = _EVAL_3338 | _EVAL_616;
  assign _EVAL_814 = _EVAL_1708 & _EVAL_3173;
  assign _EVAL_1369 = ~ _EVAL_3340;
  assign _EVAL_2804 = {{15'd0}, _EVAL_1369};
  assign _EVAL_606 = _EVAL_3338 & _EVAL_2804;
  assign _EVAL_3146 = _EVAL_43[15:0];
  assign _EVAL_399 = _EVAL_3146[1:0];
  assign _EVAL_1994 = _EVAL_399 != 2'h3;
  assign _EVAL_523 = _EVAL_1886[14:3];
  assign _EVAL_671 = {_EVAL_523, 2'h0};
  assign _EVAL_601 = _EVAL_182 & _EVAL_1412;
  assign _EVAL_1793 = _EVAL_2336 == 1'h0;
  assign _EVAL_2796 = _EVAL_2443 & _EVAL_1793;
  assign _EVAL_248 = _EVAL_1209 == 1'h0;
  assign _EVAL_2407 = _EVAL_713 & _EVAL_248;
  assign _EVAL_2276 = _EVAL_2796 | _EVAL_2407;
  assign _EVAL_2295 = _EVAL_601 & _EVAL_2276;
  assign _EVAL_944 = _EVAL_2518 & _EVAL_2295;
  assign _EVAL_3408 = _EVAL_2621 & _EVAL_248;
  assign _EVAL_2959 = _EVAL_336 == 1'h0;
  assign _EVAL_728 = _EVAL_1245 & _EVAL_2959;
  assign _EVAL_1961 = _EVAL_3408 | _EVAL_728;
  assign _EVAL_2659 = _EVAL_601 & _EVAL_1961;
  assign _EVAL_1384 = _EVAL_275 & _EVAL_2659;
  assign _EVAL_3232 = _EVAL_944 | _EVAL_1384;
  assign _EVAL_2035 = _EVAL_2012 & _EVAL_2959;
  assign _EVAL_2238 = _EVAL_1035 == 1'h0;
  assign _EVAL_2625 = _EVAL_684 & _EVAL_2238;
  assign _EVAL_885 = _EVAL_2035 | _EVAL_2625;
  assign _EVAL_2484 = _EVAL_601 & _EVAL_885;
  assign _EVAL_2385 = _EVAL_716 & _EVAL_2484;
  assign _EVAL_613 = _EVAL_3232 | _EVAL_2385;
  assign _EVAL_3047 = _EVAL_868 == 1'h0;
  assign _EVAL_2719 = _EVAL_3047 & _EVAL_1276;
  assign _EVAL_2241 = _EVAL_902 & _EVAL_2238;
  assign _EVAL_1910 = _EVAL_601 & _EVAL_2241;
  assign _EVAL_2132 = _EVAL_2719 & _EVAL_1910;
  assign _EVAL_3168 = _EVAL_613 | _EVAL_2132;
  assign _EVAL_1749 = _EVAL_3168 == 1'h0;
  assign _EVAL_796 = _EVAL_3050 - 7'h1;
  assign _EVAL_682 = $unsigned(_EVAL_796);
  assign _EVAL_3386 = _EVAL_682[6:0];
  assign _EVAL_1414 = _EVAL_1749 ? _EVAL_3386 : _EVAL_1387;
  assign _EVAL_2988 = _EVAL_1077 ? _EVAL_1414 : _EVAL_1387;
  assign _EVAL_737 = _EVAL_1386 | _EVAL_3261;
  assign _EVAL_2268 = _EVAL_737 == 1'h0;
  assign _EVAL_938 = {{1'd0}, _EVAL_2887};
  assign _EVAL_1825 = _EVAL_1215 ? {{1'd0}, _EVAL_2189} : 2'h2;
  assign _EVAL_3231 = _EVAL_938 <= _EVAL_1825;
  assign _EVAL_2216 = _EVAL_2268 & _EVAL_3231;
  assign _EVAL_3121 = _EVAL_1215 ? 2'h3 : 2'h0;
  assign _EVAL_2767 = _EVAL_2216 ? 2'h2 : _EVAL_3121;
  assign _EVAL_2251 = _EVAL_481 == 3'h1;
  assign _EVAL_2157 = _EVAL_2212 == 2'h1;
  assign _EVAL_1700 = _EVAL_1836 | _EVAL_2447;
  assign _EVAL_3177 = _EVAL_2157 & _EVAL_1700;
  assign _EVAL_2807 = _EVAL_2251 | _EVAL_3177;
  assign _EVAL_1790 = _EVAL_227 == 1'h0;
  assign _EVAL_666 = _EVAL_1790 | _EVAL_900;
  assign _EVAL_804 = _EVAL_2251 & _EVAL_666;
  assign _EVAL_2934 = _EVAL_1677 ? _EVAL_2807 : _EVAL_804;
  assign _EVAL_2821 = _EVAL_3033 & _EVAL_3053;
  assign _EVAL_1390 = _EVAL_1077 & _EVAL_2821;
  assign _EVAL_1535 = _EVAL_113 | _EVAL_1390;
  assign _EVAL_2642 = {_EVAL_2528, 1'h0};
  assign _EVAL_571 = _EVAL_2642 | 3'h1;
  assign _EVAL_1342 = _EVAL_1077 ? _EVAL_571 : {{1'd0}, _EVAL_2528};
  assign _EVAL_1638 = _EVAL_1535 ? 3'h0 : _EVAL_1342;
  assign _EVAL_880 = {predictor_tagged_tables_1__EVAL_8,predictor_tagged_tables_1__EVAL_19,predictor_tagged_tables_1__EVAL_0,predictor_tagged_tables_1__EVAL_13,predictor_tagged_tables_1__EVAL_7,predictor_tagged_tables_1__EVAL_34};
  assign _EVAL_2452 = {predictor_tagged_tables_1__EVAL_25,predictor_tagged_tables_1__EVAL_35,predictor_tagged_tables_1__EVAL_27,predictor_tagged_tables_1__EVAL_18,predictor_tagged_tables_1__EVAL_10,predictor_tagged_tables_1__EVAL_36,_EVAL_880};
  assign _EVAL_2467 = _EVAL_2452[10];
  assign _EVAL_1382 = _EVAL_1886[1:0];
  assign _EVAL_2610 = {{12'd0}, _EVAL_1382};
  assign _EVAL_3172 = _EVAL_671 | _EVAL_2610;
  assign _EVAL_2016 = _EVAL_3172[10:0];
  assign _EVAL_2121 = _EVAL_3172[13:11];
  assign _EVAL_3119 = {{8'd0}, _EVAL_2121};
  assign _EVAL_433 = _EVAL_2016 ^ _EVAL_3119;
  assign _EVAL_1083 = {{128'd0}, _EVAL_433};
  assign _EVAL_2570 = {_EVAL_2928, 11'h0};
  assign _EVAL_797 = _EVAL_1083 ^ _EVAL_2570;
  assign _EVAL_1279 = _EVAL_797[2:0];
  assign _EVAL_2210 = predictor_base_table_0__EVAL_27;
  assign _EVAL_258 = _EVAL_1663 == 1'h0;
  assign _EVAL_1423 = _EVAL_3054 == 1'h0;
  assign _EVAL_750 = _EVAL_2636 & _EVAL_1423;
  assign _EVAL_2468 = _EVAL_750 == 1'h0;
  assign _EVAL_1753 = _EVAL_2081__EVAL_2082_data;
  assign _EVAL_181 = _EVAL_2629 | _EVAL_737;
  assign _EVAL_1188 = _EVAL_1954 | _EVAL_181;
  assign _EVAL_1419 = _EVAL_1188 == 1'h0;
  assign _EVAL_1922 = _EVAL_1673 == 1'h0;
  assign _EVAL_2052 = _EVAL_1419 & _EVAL_1922;
  assign _EVAL_707 = _EVAL_181 == 1'h0;
  assign _EVAL_1062 = _EVAL_700 == 1'h0;
  assign _EVAL_1299 = _EVAL_707 & _EVAL_1062;
  assign _EVAL_2999 = _EVAL_2052 | _EVAL_1299;
  assign _EVAL_3270 = _EVAL_2398 == 1'h0;
  assign _EVAL_366 = _EVAL_2268 & _EVAL_3270;
  assign _EVAL_3154 = _EVAL_2999 | _EVAL_366;
  assign _EVAL_576 = _EVAL_2294 == 1'h0;
  assign _EVAL_513 = _EVAL_1215 & _EVAL_576;
  assign _EVAL_1584 = _EVAL_3154 | _EVAL_513;
  assign _EVAL_1685 = _EVAL_1584 == 1'h0;
  assign _EVAL_2707 = _EVAL_2347 == 1'h0;
  assign _EVAL_1371 = _EVAL_1031 == 1'h0;
  assign _EVAL_274 = _EVAL_3284 == 1'h0;
  assign _EVAL_563 = _EVAL_1954 ? 1'h0 : _EVAL_274;
  assign _EVAL_1145 = _EVAL_1371 ? 1'h1 : _EVAL_563;
  assign _EVAL_1736 = _EVAL_2629 ? 1'h0 : _EVAL_1145;
  assign _EVAL_1889 = _EVAL_258 ? 1'h1 : _EVAL_1736;
  assign _EVAL_1569 = _EVAL_1386 ? 1'h0 : _EVAL_1889;
  assign _EVAL_2446 = _EVAL_2707 ? 1'h1 : _EVAL_1569;
  assign _EVAL_866 = _EVAL_3261 ? 1'h0 : _EVAL_2446;
  assign _EVAL_894 = _EVAL_866 == 1'h0;
  assign _EVAL_2040 = _EVAL_1685 & _EVAL_894;
  assign _EVAL_206 = _EVAL_2040;
  assign _EVAL_883 = _EVAL_2468 ? _EVAL_1753 : _EVAL_206;
  assign _EVAL_2440 = _EVAL_2443 & _EVAL_2336;
  assign _EVAL_466 = _EVAL_713 & _EVAL_1209;
  assign _EVAL_201 = _EVAL_2440 | _EVAL_466;
  assign _EVAL_906 = _EVAL_2742 | _EVAL_3319;
  assign _EVAL_2748 = _EVAL_906 & _EVAL_1887;
  assign _EVAL_1603 = _EVAL_481 == 3'h2;
  assign _EVAL_2001 = _EVAL_1603 == 1'h0;
  assign _EVAL_2299 = _EVAL_2001 & _EVAL_1781;
  assign _EVAL_2054 = _EVAL_2299 ? 9'h0 : 9'h1ff;
  assign _EVAL_3167 = _EVAL_113;
  assign _EVAL_2902 = _EVAL_2550 == 1'h0;
  assign _EVAL_428 = _EVAL_344 + _EVAL_1529;
  assign _EVAL_3200 = {{1'd0}, _EVAL_428};
  assign _EVAL_2851 = _EVAL_2743 + _EVAL_3200;
  assign _EVAL_3110 = _EVAL_2851[2:0];
  assign _EVAL_3044 = _EVAL_3110 < 3'h5;
  assign _EVAL_3327 = _EVAL_2902 & _EVAL_3044;
  assign _EVAL_1255 = _EVAL_2754[2];
  assign _EVAL_1237 = _EVAL_3327 & _EVAL_1255;
  assign _EVAL_2070 = _EVAL_3167 | _EVAL_1237;
  assign _EVAL_1445 = _EVAL_1540[0];
  assign _EVAL_1899 = _EVAL_2402[5:0];
  assign _EVAL_1553 = _EVAL_1899 < 6'h38;
  assign _EVAL_1787 = 32'h1800000 <= tlb__EVAL_37;
  assign _EVAL_2801 = tlb__EVAL_37 <= 32'h1807fff;
  assign _EVAL_2905 = _EVAL_1787 & _EVAL_2801;
  assign _EVAL_1857 = _EVAL_2402[14:0];
  assign _EVAL_1964 = _EVAL_1857 < 15'h7ff8;
  assign _EVAL_3318 = _EVAL_2905 & _EVAL_1964;
  assign _EVAL_1932 = _EVAL_1553 | _EVAL_3318;
  assign _EVAL_3011 = _EVAL_1503 & _EVAL_1932;
  assign _EVAL_1709 = _EVAL_1445 | _EVAL_3011;
  assign _EVAL_1010 = _EVAL_2378 & _EVAL_1709;
  assign _EVAL_834 = _EVAL_2843 ? 1'h0 : _EVAL_1010;
  assign _EVAL_1786 = _EVAL_43[63:48];
  assign _EVAL_1263 = _EVAL_1786[15:13];
  assign _EVAL_1552 = _EVAL_1263 == 3'h4;
  assign _EVAL_3040 = _EVAL_2629 ? _EVAL_700 : _EVAL_1673;
  assign _EVAL_1151 = _EVAL_1386 ? _EVAL_2398 : _EVAL_3040;
  assign _EVAL_2893 = _EVAL_3261 ? _EVAL_2294 : _EVAL_1151;
  assign _EVAL_3183 = _EVAL_2893;
  assign _EVAL_589 = _EVAL_3183;
  assign _EVAL_709 = predictor_base_table_1__EVAL_27;
  assign _EVAL_1340 = _EVAL_1886[2];
  assign _EVAL_855 = _EVAL_1340 == 1'h0;
  assign _EVAL_2087 = _EVAL_393 & _EVAL_956;
  assign _EVAL_2974 = _EVAL_906 | _EVAL_2087;
  assign _EVAL_251 = _EVAL_1276 & _EVAL_2974;
  assign _EVAL_461 = _EVAL_1786[6:2];
  assign _EVAL_2828 = _EVAL_461 == 5'h0;
  assign _EVAL_1639 = _EVAL_1786[1:0];
  assign _EVAL_2282 = _EVAL_1639 >= 2'h2;
  assign _EVAL_3237 = _EVAL_1639 == 2'h0;
  assign _EVAL_1844 = _EVAL_2828 ? _EVAL_2282 : _EVAL_3237;
  assign _EVAL_333 = _EVAL_1993 - 5'h1;
  assign _EVAL_528 = ~ _EVAL_333;
  assign _EVAL_3215 = _EVAL_2828 ? _EVAL_3237 : _EVAL_2282;
  assign _EVAL_2910 = predictor_Queue__EVAL_0[31:3];
  assign _EVAL_2397 = {_EVAL_2910, 2'h0};
  assign _EVAL_841 = predictor_Queue__EVAL_0[1:0];
  assign _EVAL_1186 = {{29'd0}, _EVAL_841};
  assign _EVAL_1915 = _EVAL_2397 | _EVAL_1186;
  assign _EVAL_2015 = _EVAL_1915[13:11];
  assign _EVAL_2633 = {{8'd0}, _EVAL_2015};
  assign _EVAL_2278 = {MaxPeriodFibonacciLFSR_1__EVAL_12,MaxPeriodFibonacciLFSR_1__EVAL_11,MaxPeriodFibonacciLFSR_1__EVAL_3,MaxPeriodFibonacciLFSR_1__EVAL_16,MaxPeriodFibonacciLFSR_1__EVAL_8,MaxPeriodFibonacciLFSR_1__EVAL_10,MaxPeriodFibonacciLFSR_1__EVAL_14,MaxPeriodFibonacciLFSR_1__EVAL_7};
  assign _EVAL_614 = {MaxPeriodFibonacciLFSR_1__EVAL_0,MaxPeriodFibonacciLFSR_1__EVAL_17,MaxPeriodFibonacciLFSR_1__EVAL_1,MaxPeriodFibonacciLFSR_1__EVAL,MaxPeriodFibonacciLFSR_1__EVAL_5,MaxPeriodFibonacciLFSR_1__EVAL_4,MaxPeriodFibonacciLFSR_1__EVAL_6,MaxPeriodFibonacciLFSR_1__EVAL_2,_EVAL_2278};
  assign _EVAL_1138 = _EVAL_614[0];
  assign _EVAL_2615 = _EVAL_614[1];
  assign _EVAL_3070 = _EVAL_614[2];
  assign _EVAL_943 = _EVAL_614[3];
  assign _EVAL_1325 = _EVAL_614[4];
  assign _EVAL_2430 = _EVAL_614[5];
  assign _EVAL_958 = _EVAL_614[6];
  assign _EVAL_1626 = _EVAL_614[7];
  assign _EVAL_583 = _EVAL_614[8];
  assign _EVAL_3317 = _EVAL_614[9];
  assign _EVAL_3219 = _EVAL_614[10];
  assign _EVAL_1167 = _EVAL_614[11];
  assign _EVAL_2768 = _EVAL_614[12];
  assign _EVAL_628 = _EVAL_614[13];
  assign _EVAL_1233 = _EVAL_614[14];
  assign _EVAL_3132 = _EVAL_614[15];
  assign _EVAL_356 = {_EVAL_583,_EVAL_3317,_EVAL_3219,_EVAL_1167,_EVAL_2768,_EVAL_628,_EVAL_1233,_EVAL_3132};
  assign _EVAL_2393 = {_EVAL_1138,_EVAL_2615,_EVAL_3070,_EVAL_943,_EVAL_1325,_EVAL_2430,_EVAL_958,_EVAL_1626,_EVAL_356};
  assign _EVAL_2918 = _EVAL_2393[1:0];
  assign _EVAL_979 = _EVAL_2918 == 2'h1;
  assign _EVAL_708 = _EVAL_2549[11:6];
  assign _EVAL_1880 = {_EVAL_708, 3'h0};
  assign _EVAL_2003 = _EVAL_97[0];
  assign _EVAL_1456 = 23'hff << _EVAL_122;
  assign _EVAL_2537 = _EVAL_1456[7:0];
  assign _EVAL_2267 = ~ _EVAL_2537;
  assign _EVAL_1494 = _EVAL_2267[7:3];
  assign _EVAL_639 = _EVAL_2003 ? _EVAL_1494 : 5'h0;
  assign _EVAL_3144 = _EVAL_639 & _EVAL_528;
  assign _EVAL_2106 = {{4'd0}, _EVAL_3144};
  assign _EVAL_2122 = _EVAL_1880 | _EVAL_2106;
  assign _EVAL_903 = _EVAL_2122[0];
  assign _EVAL_2705 = _EVAL_10 & _EVAL_903;
  assign _EVAL_1357 = {{17'd0}, _EVAL_118};
  assign _EVAL_2437 = _EVAL_94 ^ _EVAL_1357;
  assign _EVAL_1810 = _EVAL_2534[15:0];
  assign _EVAL_1458 = _EVAL_1810[15:13];
  assign _EVAL_1989 = _EVAL_2531[22];
  assign _EVAL_179 = _EVAL_2531[19];
  assign _EVAL_2331 = _EVAL_2531[18];
  assign _EVAL_2626 = _EVAL_2531[9];
  assign _EVAL_2539 = _EVAL_2531[6];
  assign _EVAL_2285 = _EVAL_2531[5];
  assign _EVAL_904 = _EVAL_2531[2];
  assign _EVAL_3332 = _EVAL_2531[1];
  assign _EVAL_1335 = {_EVAL_2626,_EVAL_1711,_EVAL_917,_EVAL_2539,_EVAL_2285,_EVAL_1927,_EVAL_2239,_EVAL_904,_EVAL_3332,_EVAL_2553};
  assign _EVAL_656 = {_EVAL_1989,_EVAL_3264,_EVAL_179,_EVAL_2331,_EVAL_1044,_EVAL_1129,_EVAL_843,_EVAL_1335,_EVAL_2754};
  assign _EVAL_1224 = _EVAL_656[8:0];
  assign _EVAL_1585 = _EVAL_1224[0];
  assign _EVAL_1998 = _EVAL_1224[8:1];
  assign _EVAL_1972 = {_EVAL_1585,_EVAL_1998};
  assign _EVAL_1873 = _EVAL_2251 == 1'h0;
  assign _EVAL_2149 = _EVAL_1873 & _EVAL_1781;
  assign _EVAL_739 = _EVAL_3063 & _EVAL_842;
  assign _EVAL_1750 = _EVAL_3319 & _EVAL_2546;
  assign _EVAL_293 = _EVAL_739 | _EVAL_1750;
  assign _EVAL_2817 = _EVAL_2719 & _EVAL_293;
  assign _EVAL_2944 = _EVAL_3296 ? 1'h0 : _EVAL_834;
  assign _EVAL_3206 = _EVAL_1706[2:1];
  assign _EVAL_850 = _EVAL_3206 == 2'h0;
  assign _EVAL_1071 = _EVAL_2[6:0];
  assign _EVAL_2422 = _EVAL_1071[2];
  assign _EVAL_264 = _EVAL_282 | _EVAL_2133;
  assign _EVAL_2485 = _EVAL_956 | _EVAL_2336;
  assign _EVAL_3401 = _EVAL_2443 & _EVAL_2485;
  assign _EVAL_1001 = _EVAL_264 | _EVAL_3401;
  assign _EVAL_3072 = _EVAL_2518 & _EVAL_1001;
  assign _EVAL_3344 = _EVAL_2330 | _EVAL_2293;
  assign _EVAL_609 = _EVAL_956 | _EVAL_1209;
  assign _EVAL_1727 = _EVAL_713 & _EVAL_609;
  assign _EVAL_3067 = _EVAL_3344 | _EVAL_1727;
  assign _EVAL_3311 = _EVAL_2518 & _EVAL_3067;
  assign _EVAL_2197 = _EVAL_3072 | _EVAL_3311;
  assign _EVAL_1856 = _EVAL_1855 | _EVAL_2410;
  assign _EVAL_1106 = _EVAL_2621 & _EVAL_609;
  assign _EVAL_2119 = _EVAL_1856 | _EVAL_1106;
  assign _EVAL_1939 = _EVAL_2384 & _EVAL_2119;
  assign _EVAL_494 = _EVAL_3106 | _EVAL_1631;
  assign _EVAL_2815 = _EVAL_494 | _EVAL_2508;
  assign _EVAL_1582 = _EVAL_2384 & _EVAL_2815;
  assign _EVAL_1901 = _EVAL_1939 | _EVAL_1582;
  assign _EVAL_3123 = _EVAL_2197 | _EVAL_1901;
  assign _EVAL_1280 = _EVAL_1025 | _EVAL_1686;
  assign _EVAL_1427 = _EVAL_2012 & _EVAL_711;
  assign _EVAL_2777 = _EVAL_1280 | _EVAL_1427;
  assign _EVAL_2677 = _EVAL_2158 & _EVAL_2777;
  assign _EVAL_2013 = _EVAL_970 | _EVAL_1564;
  assign _EVAL_2448 = _EVAL_956 | _EVAL_1035;
  assign _EVAL_2250 = _EVAL_684 & _EVAL_2448;
  assign _EVAL_1947 = _EVAL_2013 | _EVAL_2250;
  assign _EVAL_1332 = _EVAL_2158 & _EVAL_1947;
  assign _EVAL_2303 = _EVAL_2677 | _EVAL_1332;
  assign _EVAL_694 = _EVAL_3123 | _EVAL_2303;
  assign _EVAL_3378 = _EVAL_641 | _EVAL_3063;
  assign _EVAL_2925 = _EVAL_902 & _EVAL_2448;
  assign _EVAL_1676 = _EVAL_3378 | _EVAL_2925;
  assign _EVAL_981 = _EVAL_1276 & _EVAL_1676;
  assign _EVAL_3240 = _EVAL_981 | _EVAL_251;
  assign _EVAL_697 = _EVAL_694 | _EVAL_3240;
  assign _EVAL_2152 = _EVAL_1193 | _EVAL_1537;
  assign _EVAL_1632 = _EVAL_1035 & _EVAL_956;
  assign _EVAL_2676 = _EVAL_2152 | _EVAL_1632;
  assign _EVAL_577 = _EVAL_3105 & _EVAL_2676;
  assign _EVAL_1242 = _EVAL_697 | _EVAL_577;
  assign _EVAL_689 = _EVAL_3064 < 2'h3;
  assign _EVAL_2093 = _EVAL_689 == 1'h0;
  assign _EVAL_832 = _EVAL_3105 & _EVAL_2093;
  assign _EVAL_2202 = _EVAL_3146[15:13];
  assign _EVAL_809 = _EVAL_2202 == 3'h4;
  assign _EVAL_1460 = _EVAL_809 & _EVAL_1994;
  assign _EVAL_2933 = {_EVAL_2829,_EVAL_1087,_EVAL_3380,_EVAL_2064,_EVAL_1037};
  assign _EVAL_3022 = _EVAL_2950[8];
  assign _EVAL_1878 = _EVAL_2950[4];
  assign _EVAL_3055 = {_EVAL_1794,_EVAL_3022,_EVAL_3057,_EVAL_219,_EVAL_487,_EVAL_1878,_EVAL_810,_EVAL_3348,_EVAL_2911,_EVAL_2657};
  assign _EVAL_260 = {_EVAL_2614,_EVAL_1645,_EVAL_3029,_EVAL_2008,_EVAL_698,_EVAL_635,_EVAL_2933,_EVAL_3055,_EVAL_878};
  assign _EVAL_1093 = _EVAL_260[26:18];
  assign _EVAL_3404 = _EVAL_1093[2:0];
  assign _EVAL_2164 = _EVAL_865 & _EVAL_1677;
  assign _EVAL_1170 = _EVAL_2164 == 1'h0;
  assign _EVAL_1359 = _EVAL_374 & _EVAL_1170;
  assign _EVAL_250 = _EVAL_39 & _EVAL_54;
  assign _EVAL_536 = _EVAL_2443 | _EVAL_713;
  assign _EVAL_1328 = _EVAL_536 & _EVAL_542;
  assign _EVAL_1715 = _EVAL_2789 | _EVAL_1328;
  assign _EVAL_2809 = _EVAL_2518 & _EVAL_1715;
  assign _EVAL_1425 = _EVAL_1719 & _EVAL_542;
  assign _EVAL_1370 = _EVAL_239 | _EVAL_1425;
  assign _EVAL_1405 = _EVAL_275 & _EVAL_1370;
  assign _EVAL_3184 = _EVAL_2809 | _EVAL_1405;
  assign _EVAL_1659 = _EVAL_942 & _EVAL_542;
  assign _EVAL_2325 = _EVAL_1688 | _EVAL_1659;
  assign _EVAL_1984 = _EVAL_716 & _EVAL_2325;
  assign _EVAL_3217 = _EVAL_3184 | _EVAL_1984;
  assign _EVAL_3351 = _EVAL_641 | _EVAL_2742;
  assign _EVAL_1803 = _EVAL_740 & _EVAL_542;
  assign _EVAL_226 = _EVAL_3351 | _EVAL_1803;
  assign _EVAL_1533 = _EVAL_2719 & _EVAL_226;
  assign _EVAL_2260 = _EVAL_3217 | _EVAL_1533;
  assign _EVAL_783 = _EVAL_1035 & _EVAL_542;
  assign _EVAL_1977 = _EVAL_1193 | _EVAL_783;
  assign _EVAL_2154 = _EVAL_1763 & _EVAL_1977;
  assign _EVAL_3031 = _EVAL_2260 | _EVAL_2154;
  assign _EVAL_286 = _EVAL_113 ? _EVAL_250 : _EVAL_3031;
  assign _EVAL_2151 = _EVAL_2534[47:32];
  assign _EVAL_649 = _EVAL_2151[6:2];
  assign _EVAL_3058 = _EVAL_649 == 5'h0;
  assign _EVAL_2050 = _EVAL_2950[100];
  assign _EVAL_2275 = _EVAL_51;
  assign _EVAL_1018 = _EVAL_2275;
  assign _EVAL_2790 = _EVAL_1018 ? 1'h1 : _EVAL_2949;
  assign _EVAL_3032 = _EVAL_2790;
  assign _EVAL_916 = _EVAL_139[31:6];
  assign _EVAL_2067 = _EVAL_2531[85];
  assign _EVAL_1479 = _EVAL_2950[43];
  assign _EVAL_1173 = _EVAL_2950[41];
  assign _EVAL_567 = _EVAL_2950[36];
  assign _EVAL_1282 = _EVAL_2950[34];
  assign _EVAL_2916 = _EVAL_2950[29];
  assign _EVAL_1612 = _EVAL_2950[27];
  assign _EVAL_556 = _EVAL_2950[25];
  assign _EVAL_1420 = _EVAL_2950[23];
  assign _EVAL_1783 = {_EVAL_2211,_EVAL_2916,_EVAL_1612,_EVAL_556,_EVAL_1420};
  assign _EVAL_760 = {_EVAL_1645,_EVAL_2008,_EVAL_635,_EVAL_3380,_EVAL_1037,_EVAL_1794,_EVAL_219,_EVAL_1878,_EVAL_3348,_EVAL_2657};
  assign _EVAL_2868 = {_EVAL_623,_EVAL_1479,_EVAL_1173,_EVAL_587,_EVAL_567,_EVAL_1282,_EVAL_1783,_EVAL_760,_EVAL_878};
  assign _EVAL_914 = _EVAL_2531[112];
  assign _EVAL_1430 = _EVAL_2531[106];
  assign _EVAL_2474 = _EVAL_2531[100];
  assign _EVAL_2535 = _EVAL_2531[95];
  assign _EVAL_1437 = _EVAL_2531[89];
  assign _EVAL_3283 = _EVAL_2531[84];
  assign _EVAL_2145 = _EVAL_2531[78];
  assign _EVAL_1712 = _EVAL_2531[72];
  assign _EVAL_3288 = _EVAL_2531[67];
  assign _EVAL_2835 = {_EVAL_2145,_EVAL_1712,_EVAL_3288,_EVAL_667,_EVAL_2824};
  assign _EVAL_1917 = _EVAL_2531[50];
  assign _EVAL_1307 = _EVAL_2531[44];
  assign _EVAL_1042 = _EVAL_2531[39];
  assign _EVAL_2245 = _EVAL_2531[33];
  assign _EVAL_3358 = {_EVAL_1917,_EVAL_1307,_EVAL_1042,_EVAL_2245,_EVAL_3139,_EVAL_1989,_EVAL_1129,_EVAL_1931,_EVAL_2285,_EVAL_2553};
  assign _EVAL_3138 = {_EVAL_914,_EVAL_1430,_EVAL_2474,_EVAL_2535,_EVAL_1437,_EVAL_3283,_EVAL_2835,_EVAL_3358,_EVAL_2754};
  assign _EVAL_2578 = _EVAL_3138[35:27];
  assign _EVAL_1565 = _EVAL_2578[0];
  assign _EVAL_1270 = _EVAL_2578[8:1];
  assign _EVAL_2823 = {_EVAL_1565,_EVAL_1270};
  assign _EVAL_2664 = _EVAL_118[2:1];
  assign _EVAL_730 = _EVAL_548__EVAL_549_data;
  assign _EVAL_1105 = _EVAL_1652__EVAL_1653_data;
  assign _EVAL_790 = _EVAL_481 == 3'h0;
  assign _EVAL_148 = _EVAL_2212 == 2'h0;
  assign _EVAL_2144 = _EVAL_148 & _EVAL_1700;
  assign _EVAL_2760 = _EVAL_790 | _EVAL_2144;
  assign _EVAL_2771 = _EVAL_790 & _EVAL_666;
  assign _EVAL_651 = _EVAL_1677 ? _EVAL_2760 : _EVAL_2771;
  assign _EVAL_3156 = _EVAL_865 & _EVAL_651;
  assign _EVAL_338 = _EVAL_3156 == 1'h0;
  assign _EVAL_470 = _EVAL_338 & _EVAL_3327;
  assign _EVAL_1664 = _EVAL_350 == 1'h0;
  assign _EVAL_2560 = _EVAL_2052 ? 1'h0 : 1'h1;
  assign _EVAL_1956 = _EVAL_2999 ? {{1'd0}, _EVAL_2560} : 2'h2;
  assign _EVAL_1728 = _EVAL_3154 ? _EVAL_1956 : 2'h3;
  assign _EVAL_376 = {{1'd0}, _EVAL_1165};
  assign _EVAL_1331 = {{1'd0}, _EVAL_1748};
  assign _EVAL_266 = _EVAL_2216 ? {{1'd0}, _EVAL_2887} : _EVAL_1825;
  assign _EVAL_580 = _EVAL_1331 <= _EVAL_266;
  assign _EVAL_1824 = _EVAL_707 & _EVAL_580;
  assign _EVAL_2608 = _EVAL_1824 ? {{1'd0}, _EVAL_1748} : _EVAL_266;
  assign _EVAL_1593 = _EVAL_376 <= _EVAL_2608;
  assign _EVAL_2683 = _EVAL_1419 & _EVAL_1593;
  assign _EVAL_1945 = _EVAL_1824 ? 2'h1 : _EVAL_2767;
  assign _EVAL_2221 = _EVAL_2683 ? 2'h0 : _EVAL_1945;
  assign _EVAL_2307 = _EVAL_1584 ? _EVAL_1728 : _EVAL_2221;
  assign _EVAL_636 = _EVAL_2307;
  assign _EVAL_787 = _EVAL_3082__EVAL_3083_data;
  assign _EVAL_561 = _EVAL_1664 ? _EVAL_636 : _EVAL_787;
  assign _EVAL_1511 = _EVAL_1993 == 5'h1;
  assign _EVAL_1157 = _EVAL_639 == 5'h0;
  assign _EVAL_3129 = _EVAL_1511 | _EVAL_1157;
  assign _EVAL_2010 = _EVAL_3129 & _EVAL_10;
  assign _EVAL_146 = _EVAL_10 & _EVAL_2010;
  assign _EVAL_1248 = _EVAL_1848 & _EVAL_1170;
  assign _EVAL_278 = _EVAL_2452[9:1];
  assign _EVAL_2349 = _EVAL_278 == _EVAL_1128;
  assign _EVAL_1410 = _EVAL_1248 & _EVAL_2349;
  assign _EVAL_2080 = {_EVAL_2256,_EVAL_2626,_EVAL_917,_EVAL_2539,_EVAL_2285,_EVAL_2239,_EVAL_904,_EVAL_3332,_EVAL_2553};
  assign _EVAL_1067 = {_EVAL_1989,_EVAL_3264,_EVAL_179,_EVAL_2331,_EVAL_1129,_EVAL_1376,_EVAL_2037,_EVAL_3388,_EVAL_1931,_EVAL_2080};
  assign _EVAL_3387 = {_EVAL_1067,_EVAL_791};
  assign _EVAL_568 = _EVAL_3387[17:9];
  assign _EVAL_946 = _EVAL_568[8:1];
  assign _EVAL_2825 = _EVAL_2151[1:0];
  assign _EVAL_2180 = _EVAL_2825 == 2'h0;
  assign _EVAL_2929 = _EVAL_2825 >= 2'h2;
  assign _EVAL_2931 = _EVAL_3058 ? _EVAL_2180 : _EVAL_2929;
  assign _EVAL_1725 = _EVAL_2531[46];
  assign _EVAL_3043 = _EVAL_2531[43];
  assign _EVAL_785 = _EVAL_2531[36];
  assign _EVAL_854 = _EVAL_2531[29];
  assign _EVAL_1894 = _EVAL_2531[27];
  assign _EVAL_1562 = _EVAL_2531[25];
  assign _EVAL_2492 = _EVAL_2531[23];
  assign _EVAL_1858 = {_EVAL_2521,_EVAL_854,_EVAL_1894,_EVAL_1562,_EVAL_2492};
  assign _EVAL_2002 = {_EVAL_3264,_EVAL_2331,_EVAL_1129,_EVAL_2434,_EVAL_1931,_EVAL_2626,_EVAL_2539,_EVAL_1927,_EVAL_904,_EVAL_2553};
  assign _EVAL_234 = {_EVAL_1725,_EVAL_3043,_EVAL_3299,_EVAL_1042,_EVAL_785,_EVAL_2967,_EVAL_1858,_EVAL_2002,_EVAL_2754};
  assign _EVAL_1936 = _EVAL_234[26:18];
  assign _EVAL_2588 = _EVAL_1936[4:0];
  assign _EVAL_2791 = _EVAL_1387 - 7'h2;
  assign _EVAL_1103 = $unsigned(_EVAL_2791);
  assign _EVAL_1158 = _EVAL_1103[6:0];
  assign _EVAL_1448 = _EVAL_2629 ? _EVAL_1372 : _EVAL_430;
  assign _EVAL_999 = _EVAL_1071[0];
  assign _EVAL_1837 = _EVAL_2518 & _EVAL_201;
  assign _EVAL_2566 = _EVAL_2621 & _EVAL_1209;
  assign _EVAL_2487 = _EVAL_1245 & _EVAL_336;
  assign _EVAL_1806 = _EVAL_2566 | _EVAL_2487;
  assign _EVAL_3307 = _EVAL_275 & _EVAL_1806;
  assign _EVAL_172 = _EVAL_1837 | _EVAL_3307;
  assign _EVAL_1301 = _EVAL_2012 & _EVAL_336;
  assign _EVAL_2609 = _EVAL_684 & _EVAL_1035;
  assign _EVAL_2466 = _EVAL_1301 | _EVAL_2609;
  assign _EVAL_220 = _EVAL_716 & _EVAL_2466;
  assign _EVAL_2805 = _EVAL_172 | _EVAL_220;
  assign _EVAL_2698 = _EVAL_902 & _EVAL_1035;
  assign _EVAL_2891 = _EVAL_2719 & _EVAL_2698;
  assign _EVAL_1908 = _EVAL_2805 | _EVAL_2891;
  assign _EVAL_1350 = _EVAL_719__EVAL_720_data;
  assign _EVAL_2296 = _EVAL_2212 == 2'h3;
  assign _EVAL_2845 = _EVAL_2296 & _EVAL_1700;
  assign _EVAL_456 = _EVAL_1981 | _EVAL_2845;
  assign _EVAL_2886 = _EVAL_314[2];
  assign _EVAL_2482 = _EVAL_3236 & _EVAL_2886;
  assign _EVAL_3304 = _EVAL_43[31:16];
  assign _EVAL_2269 = _EVAL_3304[15:13];
  assign _EVAL_2181 = _EVAL_2269 == 3'h4;
  assign _EVAL_2846 = _EVAL_2534[63:48];
  assign _EVAL_308 = _EVAL_2846[1:0];
  assign _EVAL_1629 = _EVAL_308 == 2'h0;
  assign _EVAL_1459 = {predictor_tagged_tables_2__EVAL_8,predictor_tagged_tables_2__EVAL_19,predictor_tagged_tables_2__EVAL_0,predictor_tagged_tables_2__EVAL_13,predictor_tagged_tables_2__EVAL_7,predictor_tagged_tables_2__EVAL_34};
  assign _EVAL_741 = {predictor_tagged_tables_2__EVAL_25,predictor_tagged_tables_2__EVAL_35,predictor_tagged_tables_2__EVAL_27,predictor_tagged_tables_2__EVAL_18,predictor_tagged_tables_2__EVAL_10,predictor_tagged_tables_2__EVAL_36,_EVAL_1459};
  assign _EVAL_637 = _EVAL_741[9:1];
  assign _EVAL_2601 = _EVAL_3387[8:0];
  assign _EVAL_3213 = _EVAL_568[0];
  assign _EVAL_3088 = {_EVAL_3213,_EVAL_946};
  assign _EVAL_1497 = _EVAL_2601 ^ _EVAL_3088;
  assign _EVAL_1635 = _EVAL_394__EVAL_395_data;
  assign _EVAL_357 = _EVAL_1255 == 1'h0;
  assign _EVAL_1826 = _EVAL_3327 & _EVAL_357;
  assign _EVAL_3069 = _EVAL_3167 | _EVAL_1826;
  assign _EVAL_1110 = _EVAL_3069 == 1'h0;
  assign _EVAL_1543 = _EVAL_1110 & _EVAL_1160;
  assign _EVAL_2200 = predictor_Queue__EVAL_9 != predictor_Queue__EVAL_11;
  assign _EVAL_3233 = predictor_Queue__EVAL_13 | _EVAL_2200;
  assign _EVAL_2182 = _EVAL_3233 == 1'h0;
  assign _EVAL_3013 = _EVAL_1543 ? 1'h1 : _EVAL_2182;
  assign _EVAL_1227 = _EVAL_658__EVAL_659_data;
  assign _EVAL_1973 = _EVAL_2846[15:13];
  assign _EVAL_312 = _EVAL_1973 == 3'h4;
  assign _EVAL_764 = _EVAL_82 - 128'h1;
  assign _EVAL_1854 = $unsigned(_EVAL_764);
  assign _EVAL_298 = _EVAL_2534[31:16];
  assign _EVAL_1185 = _EVAL_298[6:2];
  assign _EVAL_3345 = _EVAL_2291[12];
  assign _EVAL_912 = _EVAL_1102 + 3'h1;
  assign _EVAL_170 = _EVAL_234[17:9];
  assign _EVAL_2778 = _EVAL_170[3:0];
  assign _EVAL_2375 = _EVAL_170[8:4];
  assign _EVAL_2875 = {_EVAL_2778,_EVAL_2375};
  assign _EVAL_655 = _EVAL_1071[1];
  assign _EVAL_1583 = _EVAL_999 ? _EVAL_3155 : _EVAL_837;
  assign _EVAL_1928 = _EVAL_1583[1:0];
  assign _EVAL_465 = _EVAL_1583[127:2];
  assign _EVAL_2432 = {_EVAL_1928,_EVAL_465};
  assign _EVAL_524 = _EVAL_655 ? _EVAL_2432 : _EVAL_1583;
  assign _EVAL_733 = _EVAL_524[127:4];
  assign _EVAL_2716 = _EVAL_2677 | _EVAL_1582;
  assign _EVAL_2090 = _EVAL_2950[61];
  assign _EVAL_1356 = _EVAL_2950[57];
  assign _EVAL_1622 = _EVAL_2950[53];
  assign _EVAL_1581 = _EVAL_2950[37];
  assign _EVAL_236 = {_EVAL_2211,_EVAL_1273,_EVAL_2782,_EVAL_1645,_EVAL_635,_EVAL_2064,_EVAL_3022,_EVAL_1878,_EVAL_2657};
  assign _EVAL_2190 = {_EVAL_2958,_EVAL_1694,_EVAL_2090,_EVAL_1356,_EVAL_1622,_EVAL_1695,_EVAL_1353,_EVAL_1173,_EVAL_1581,_EVAL_236};
  assign _EVAL_1161 = {_EVAL_2190,_EVAL_1006};
  assign _EVAL_429 = _EVAL_1161[17:9];
  assign _EVAL_1095 = _EVAL_429[4:0];
  assign _EVAL_346 = _EVAL_1639 != 2'h3;
  assign _EVAL_1997 = _EVAL_1552 & _EVAL_346;
  assign _EVAL_1278 = {_EVAL_3215,_EVAL_1844};
  assign _EVAL_499 = _EVAL_1997 ? _EVAL_1278 : _EVAL_1639;
  assign _EVAL_2450 = _EVAL_3076;
  assign _EVAL_2617 = _EVAL_2450;
  assign _EVAL_1268 = _EVAL_2640 ? tag_array__EVAL_2 : _EVAL_849;
  assign _EVAL_2420 = _EVAL_1268[20];
  assign _EVAL_1968 = _EVAL_1336 | 16'h3;
  assign _EVAL_3295 = _EVAL_260[17:9];
  assign _EVAL_586 = _EVAL_3295[1:0];
  assign _EVAL_2406 = _EVAL_2402[11:6];
  assign _EVAL_881 = {2'h2,_EVAL_2406};
  assign _EVAL_2602 = _EVAL_1268[19:0];
  assign _EVAL_2892 = _EVAL_3376[12];
  assign _EVAL_475 = _EVAL_2133 & _EVAL_2892;
  assign _EVAL_2114 = _EVAL_2531[105];
  assign _EVAL_2204 = _EVAL_2531[98];
  assign _EVAL_1938 = _EVAL_2531[92];
  assign _EVAL_1418 = _EVAL_2531[79];
  assign _EVAL_303 = _EVAL_2531[26];
  assign _EVAL_2672 = {_EVAL_2652,_EVAL_1725,_EVAL_1042,_EVAL_2521,_EVAL_303,_EVAL_179,_EVAL_2434,_EVAL_2539,_EVAL_2553};
  assign _EVAL_1839 = {_EVAL_914,_EVAL_2114,_EVAL_2204,_EVAL_1938,_EVAL_2067,_EVAL_1418,_EVAL_1712,_EVAL_624,_EVAL_2193,_EVAL_2672};
  assign _EVAL_1057 = {_EVAL_1839,_EVAL_791};
  assign _EVAL_2997 = _EVAL_1057[8:0];
  assign _EVAL_2332 = _EVAL_1365 != _EVAL_1372;
  assign _EVAL_2571 = _EVAL_2332 & _EVAL_1062;
  assign _EVAL_1501 = _EVAL_3063 & _EVAL_3345;
  assign _EVAL_534 = _EVAL_2431 | _EVAL_1501;
  assign _EVAL_808 = _EVAL_139[31:3];
  assign _EVAL_2312 = _EVAL_808[2:0];
  assign _EVAL_1817 = _EVAL_454 >> _EVAL_2312;
  assign _EVAL_644 = _EVAL_1817[0];
  assign _EVAL_2992 = _EVAL_3406 >> _EVAL_2312;
  assign _EVAL_1471 = _EVAL_2992[0];
  assign _EVAL_2442 = _EVAL_644 & _EVAL_1471;
  assign _EVAL_257 = _EVAL_2442 == 1'h0;
  assign _EVAL_2725 = _EVAL_2640 ? tag_array__EVAL_7 : _EVAL_1785;
  assign _EVAL_143 = _EVAL_2725[20];
  assign _EVAL_418 = _EVAL_1859__EVAL_1861_data[7:0];
  assign _EVAL_1515 = _EVAL_2846[6:2];
  assign _EVAL_1698 = _EVAL_1515 == 5'h0;
  assign _EVAL_2224 = _EVAL_308 >= 2'h2;
  assign _EVAL_934 = _EVAL_1698 ? _EVAL_1629 : _EVAL_2224;
  assign _EVAL_1925 = _EVAL_10 == 1'h0;
  assign _EVAL_1526 = _EVAL_1692 | _EVAL_947;
  assign _EVAL_372 = _EVAL_1526 | _EVAL_1953;
  assign _EVAL_1288 = _EVAL_83 | _EVAL_372;
  assign _EVAL_1388 = _EVAL_1288 == 1'h0;
  assign _EVAL_1507 = _EVAL_1925 & _EVAL_1388;
  assign _EVAL_3126 = _EVAL_2902 & _EVAL_3044;
  assign _EVAL_450 = _EVAL_113 | _EVAL_3126;
  assign _EVAL_2700 = _EVAL_1507 & _EVAL_450;
  assign _EVAL_738 = _EVAL_113 ? 1'h0 : _EVAL_2944;
  assign _EVAL_1235 = _EVAL_738 == 1'h0;
  assign _EVAL_2863 = _EVAL_616[0];
  assign _EVAL_2653 = _EVAL_2273[15:1];
  assign _EVAL_831 = _EVAL_3206 - 2'h1;
  assign _EVAL_788 = _EVAL_850 | _EVAL_1957;
  assign _EVAL_1054 = _EVAL_2273 ^ _EVAL_2686;
  assign _EVAL_2941 = _EVAL_1054[20:6];
  assign _EVAL_2935 = _EVAL_2941 == 15'h0;
  assign _EVAL_2377 = {_EVAL_2686,_EVAL_2653,_EVAL_831,_EVAL_788,_EVAL_155,_EVAL_2935};
  assign _EVAL_864 = _EVAL_2950[106];
  assign _EVAL_2038 = _EVAL_2950[95];
  assign _EVAL_3363 = _EVAL_2950[89];
  assign _EVAL_1139 = _EVAL_2950[84];
  assign _EVAL_778 = _EVAL_2950[78];
  assign _EVAL_1682 = _EVAL_2950[67];
  assign _EVAL_3094 = {_EVAL_778,_EVAL_2879,_EVAL_1682,_EVAL_2090,_EVAL_3012};
  assign _EVAL_1879 = _EVAL_2950[50];
  assign _EVAL_621 = _EVAL_2950[44];
  assign _EVAL_879 = _EVAL_2950[33];
  assign _EVAL_2979 = {_EVAL_1879,_EVAL_621,_EVAL_587,_EVAL_879,_EVAL_1273,_EVAL_2614,_EVAL_635,_EVAL_1037,_EVAL_487,_EVAL_2657};
  assign _EVAL_3257 = {_EVAL_2922,_EVAL_864,_EVAL_2050,_EVAL_2038,_EVAL_3363,_EVAL_1139,_EVAL_3094,_EVAL_2979,_EVAL_878};
  assign _EVAL_2831 = _EVAL_3257[17:9];
  assign _EVAL_2717 = _EVAL_2402 ^ _EVAL_2392;
  assign _EVAL_3162 = _EVAL_2717[31:6];
  assign _EVAL_2749 = _EVAL_637 == _EVAL_1755;
  assign _EVAL_467 = _EVAL_2227[6:2];
  assign _EVAL_2056 = _EVAL_467 == 5'h0;
  assign _EVAL_2818 = _EVAL_20;
  assign _EVAL_1222 = _EVAL_3032 & _EVAL_2468;
  assign _EVAL_1696 = _EVAL_2248 + 2'h1;
  assign _EVAL_2981 = _EVAL_1386 ? _EVAL_2882 : _EVAL_1448;
  assign _EVAL_847 = _EVAL_3261 ? _EVAL_2304 : _EVAL_2981;
  assign _EVAL_3325 = _EVAL_2868[8:0];
  assign _EVAL_2184 = _EVAL_3325[8:3];
  assign _EVAL_798 = _EVAL_616[10];
  assign _EVAL_348 = _EVAL_1995 ? 1'h1 : _EVAL_113;
  assign _EVAL_1496 = _EVAL_1077 ? _EVAL_348 : _EVAL_113;
  assign _EVAL_1577 = _EVAL_1496 == 1'h0;
  assign _EVAL_2515 = _EVAL_38 == 1'h0;
  assign _EVAL_792 = _EVAL_1077;
  assign _EVAL_160 = _EVAL_113 ? _EVAL_2515 : _EVAL_792;
  assign _EVAL_2762 = _EVAL_3146[6:2];
  assign _EVAL_2736 = _EVAL_2762 == 5'h0;
  assign _EVAL_705 = _EVAL_399 == 2'h0;
  assign _EVAL_2622 = _EVAL_399 >= 2'h2;
  assign _EVAL_1256 = _EVAL_2736 ? _EVAL_705 : _EVAL_2622;
  assign _EVAL_196 = _EVAL_2736 ? _EVAL_2622 : _EVAL_705;
  assign _EVAL_1137 = {_EVAL_1256,_EVAL_196};
  assign _EVAL_2576 = _EVAL_113 ? _EVAL_89 : _EVAL_175;
  assign _EVAL_3095 = _EVAL_2576[31:1];
  assign _EVAL_1090 = _EVAL_3095[14:0];
  assign _EVAL_1665 = _EVAL_1090[14:3];
  assign _EVAL_3204 = {_EVAL_1665, 2'h0};
  assign _EVAL_1262 = _EVAL_1090[1:0];
  assign _EVAL_620 = {{12'd0}, _EVAL_1262};
  assign _EVAL_1050 = _EVAL_3204 | _EVAL_620;
  assign _EVAL_242 = _EVAL_1810[6:2];
  assign _EVAL_2183 = _EVAL_242 == 5'h0;
  assign _EVAL_496 = _EVAL_1810[1:0];
  assign _EVAL_322 = _EVAL_496 == 2'h0;
  assign _EVAL_2726 = _EVAL_496 >= 2'h2;
  assign _EVAL_2415 = _EVAL_2183 ? _EVAL_322 : _EVAL_2726;
  assign _EVAL_3081 = _EVAL_2183 ? _EVAL_2726 : _EVAL_322;
  assign _EVAL_214 = {_EVAL_2415,_EVAL_3081};
  assign _EVAL_1066 = {predictor_tagged_tables_0__EVAL_8,predictor_tagged_tables_0__EVAL_19,predictor_tagged_tables_0__EVAL_0,predictor_tagged_tables_0__EVAL_13,predictor_tagged_tables_0__EVAL_7,predictor_tagged_tables_0__EVAL_34};
  assign _EVAL_1924 = {predictor_tagged_tables_0__EVAL_25,predictor_tagged_tables_0__EVAL_35,predictor_tagged_tables_0__EVAL_27,predictor_tagged_tables_0__EVAL_18,predictor_tagged_tables_0__EVAL_10,predictor_tagged_tables_0__EVAL_36,_EVAL_1066};
  assign _EVAL_2032 = _EVAL_1924[9:1];
  assign _EVAL_2148 = _EVAL_2032 == _EVAL_1746;
  assign _EVAL_2927 = _EVAL_1359 & _EVAL_2148;
  assign _EVAL_2454 = _EVAL_2950[40];
  assign _EVAL_468 = {_EVAL_695,_EVAL_2008,_EVAL_635,_EVAL_3380,_EVAL_2595,_EVAL_3022,_EVAL_487,_EVAL_3348,_EVAL_2657};
  assign _EVAL_1876 = {_EVAL_623,_EVAL_1479,_EVAL_2454,_EVAL_1581,_EVAL_1117,_EVAL_2211,_EVAL_2916,_EVAL_1612,_EVAL_2782,_EVAL_468};
  assign _EVAL_1684 = {_EVAL_1876,_EVAL_1006};
  assign _EVAL_152 = _EVAL_1684[26:18];
  assign _EVAL_464 = _EVAL_175[31:3];
  assign _EVAL_1203 = _EVAL_464[0];
  assign _EVAL_3191 = _EVAL_1203 == 1'h0;
  assign _EVAL_2441 = _EVAL_2789 | _EVAL_1463;
  assign _EVAL_3192 = _EVAL_2518 & _EVAL_2441;
  assign _EVAL_3079 = _EVAL_44 | _EVAL_113;
  assign _EVAL_1261 = _EVAL_3079;
  assign _EVAL_1578 = _EVAL_616[5];
  assign _EVAL_1774 = _EVAL_43[47:32];
  assign _EVAL_1853 = _EVAL_1774[1:0];
  assign _EVAL_2028 = _EVAL_429[8:5];
  assign _EVAL_1771 = _EVAL_3126 & _EVAL_1203;
  assign _EVAL_2529 = _EVAL_489__EVAL_490_data;
  assign _EVAL_2404 = _EVAL_2580__EVAL_2581_data;
  assign _EVAL_1234 = _EVAL_2468 ? _EVAL_2404 : _EVAL_2450;
  assign _EVAL_2368 = _EVAL_113 | packageanon1_4__EVAL_0;
  assign _EVAL_478 = _EVAL_656[17:9];
  assign _EVAL_2358 = _EVAL_478[1:0];
  assign _EVAL_3313 = _EVAL_478[8:2];
  assign _EVAL_412 = {_EVAL_2358,_EVAL_3313};
  assign _EVAL_2737 = _EVAL_1972 ^ _EVAL_412;
  assign _EVAL_3391 = _EVAL_314[6];
  assign _EVAL_551 = _EVAL_3236 & _EVAL_3391;
  assign _EVAL_1546 = _EVAL_551 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_1513 = _EVAL_2531[40];
  assign _EVAL_2207 = _EVAL_903 == 1'h0;
  assign _EVAL_2319 = _EVAL_10 & _EVAL_2207;
  assign _EVAL_1935 = _EVAL_2918 == 2'h3;
  assign _EVAL_2792 = _EVAL_2319 & _EVAL_1935;
  assign _EVAL_564 = _EVAL_2792 == 1'h0;
  assign _EVAL_1866 = _EVAL_113 | packageanon1_7__EVAL_0;
  assign _EVAL_3268 = _EVAL_2792 | _EVAL_1866;
  assign _EVAL_1108 = _EVAL_564 & _EVAL_3268;
  assign _EVAL_1323 = _EVAL_2868[26:18];
  assign _EVAL_3241 = _EVAL_3058 ? _EVAL_2929 : _EVAL_2180;
  assign _EVAL_177 = _EVAL_1161[8:0];
  assign _EVAL_3051 = _EVAL_177[8:4];
  assign _EVAL_1902 = _EVAL_1303 & _EVAL_1170;
  assign _EVAL_2196 = _EVAL_1323[4:0];
  assign _EVAL_2864 = _EVAL_2274;
  assign _EVAL_2558 = _EVAL_2864 == 1'h0;
  assign _EVAL_1904 = _EVAL_3076 != _EVAL_430;
  assign _EVAL_1022 = _EVAL_1904 & _EVAL_1922;
  assign _EVAL_463 = _EVAL_1954 ? _EVAL_1022 : 1'h0;
  assign _EVAL_2638 = _EVAL_239 | _EVAL_1847;
  assign _EVAL_3120 = _EVAL_2384 & _EVAL_2638;
  assign _EVAL_1462 = _EVAL_1939 | _EVAL_3311;
  assign _EVAL_3343 = _EVAL_1915[10:0];
  assign _EVAL_1474 = _EVAL_3343 ^ _EVAL_2633;
  assign _EVAL_599 = {{128'd0}, _EVAL_1474};
  assign _EVAL_1180 = {predictor_Queue__EVAL_12, 11'h0};
  assign _EVAL_2732 = _EVAL_599 ^ _EVAL_1180;
  assign _EVAL_246 = _EVAL_2732[138:3];
  assign _EVAL_2619 = _EVAL_246[7:0];
  assign _EVAL_1765 = _EVAL_2732[2:0];
  assign _EVAL_2226 = _EVAL_1765 == 3'h6;
  assign _EVAL_1784 = _EVAL_1081 | _EVAL_2817;
  assign _EVAL_3042 = _EVAL_2636 & _EVAL_3054;
  assign _EVAL_2361 = _EVAL_3042 == 1'h0;
  assign _EVAL_1171 = _EVAL_2719 & _EVAL_3351;
  assign _EVAL_1164 = _EVAL_2023__EVAL_2024_data;
  assign _EVAL_3149 = _EVAL_1677 & _EVAL_1790;
  assign _EVAL_2962 = _EVAL_3080 | _EVAL_3149;
  assign _EVAL_2536 = _EVAL_1751 & _EVAL_227;
  assign _EVAL_455 = _EVAL_227 + 1'h1;
  assign _EVAL_367 = _EVAL_2536 ? 1'h1 : _EVAL_455;
  assign _EVAL_277 = _EVAL_2962 ? 1'h0 : _EVAL_367;
  assign _EVAL_2475 = _EVAL_616[11];
  assign _EVAL_3291 = _EVAL_1071[5];
  assign _EVAL_3096 = _EVAL_1071[4];
  assign _EVAL_1499 = _EVAL_1071[3];
  assign _EVAL_1558 = _EVAL_524[3:0];
  assign _EVAL_2547 = {_EVAL_1558,_EVAL_733};
  assign _EVAL_452 = _EVAL_2422 ? _EVAL_2547 : _EVAL_524;
  assign _EVAL_872 = _EVAL_452[7:0];
  assign _EVAL_2417 = _EVAL_452[127:8];
  assign _EVAL_2734 = {_EVAL_872,_EVAL_2417};
  assign _EVAL_2983 = _EVAL_1499 ? _EVAL_2734 : _EVAL_452;
  assign _EVAL_2620 = _EVAL_2983[15:0];
  assign _EVAL_1009 = _EVAL_2983[127:16];
  assign _EVAL_1877 = {_EVAL_2620,_EVAL_1009};
  assign _EVAL_3007 = _EVAL_3096 ? _EVAL_1877 : _EVAL_2983;
  assign _EVAL_2476 = _EVAL_3007[31:0];
  assign _EVAL_2545 = _EVAL_3007[127:32];
  assign _EVAL_2703 = {_EVAL_2476,_EVAL_2545};
  assign _EVAL_2594 = _EVAL_3291 ? _EVAL_2703 : _EVAL_3007;
  assign _EVAL_2813 = _EVAL_2594[63:0];
  assign _EVAL_500 = _EVAL_2594[127:64];
  assign _EVAL_533 = {_EVAL_2813,_EVAL_500};
  assign _EVAL_2109 = _EVAL_2918 == 2'h0;
  assign _EVAL_3227 = _EVAL_2319 & _EVAL_2109;
  assign _EVAL_3315 = _EVAL_494 & _EVAL_2060;
  assign _EVAL_1250 = _EVAL_1993 == 5'h0;
  assign _EVAL_2058 = {predictor_tagged_tables_3__EVAL_8,predictor_tagged_tables_3__EVAL_19,predictor_tagged_tables_3__EVAL_0,predictor_tagged_tables_3__EVAL_13,predictor_tagged_tables_3__EVAL_7,predictor_tagged_tables_3__EVAL_34};
  assign _EVAL_2192 = {predictor_tagged_tables_3__EVAL_25,predictor_tagged_tables_3__EVAL_35,predictor_tagged_tables_3__EVAL_27,predictor_tagged_tables_3__EVAL_18,predictor_tagged_tables_3__EVAL_10,predictor_tagged_tables_3__EVAL_36,_EVAL_2058};
  assign _EVAL_1133 = _EVAL_2192[10];
  assign _EVAL_211 = _EVAL_1688 | _EVAL_3372;
  assign _EVAL_825 = _EVAL_616[7];
  assign _EVAL_826 = _EVAL_1990[26:18];
  assign _EVAL_3062 = _EVAL_826[7:0];
  assign _EVAL_1788 = _EVAL_2482 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_1498 = _EVAL_1788[23:16];
  assign _EVAL_2710 = _EVAL_113 | _EVAL_10;
  assign _EVAL_1754 = _EVAL_2710 ? packageanon1__EVAL : _EVAL_175;
  assign _EVAL_1324 = _EVAL_1754[11:6];
  assign _EVAL_424 = {_EVAL_1324, 3'h0};
  assign _EVAL_2069 = _EVAL_2790 == 1'h0;
  assign _EVAL_2859 = _EVAL_2468 | _EVAL_2069;
  assign _EVAL_1911 = _EVAL_1077 & _EVAL_2859;
  assign _EVAL_2390 = _EVAL_2361 & _EVAL_1911;
  assign _EVAL_2242 = _EVAL_1873 | _EVAL_3149;
  assign _EVAL_1619 = _EVAL_2242 ? 1'h0 : _EVAL_367;
  assign _EVAL_2937 = _EVAL_2212 == 2'h2;
  assign _EVAL_2661 = _EVAL_2937 & _EVAL_1700;
  assign _EVAL_1982 = _EVAL_215__EVAL_216_data;
  assign _EVAL_2042 = _EVAL_3192 | _EVAL_3120;
  assign _EVAL_2491 = _EVAL_2402[31:6];
  assign _EVAL_1024 = _EVAL_995[12];
  assign _EVAL_899 = _EVAL_2825 != 2'h3;
  assign _EVAL_1291 = _EVAL_1050[10:0];
  assign _EVAL_2524 = _EVAL_3257[35:27];
  assign _EVAL_1971 = _EVAL_2524[8:1];
  assign _EVAL_3331 = _EVAL_19 | _EVAL_271;
  assign _EVAL_501 = _EVAL_3331 | _EVAL_344;
  assign _EVAL_2525 = _EVAL_1102 - 3'h1;
  assign _EVAL_449 = $unsigned(_EVAL_2525);
  assign _EVAL_2708 = _EVAL_2158 & _EVAL_3372;
  assign _EVAL_848 = _EVAL_2013 & _EVAL_1310;
  assign _EVAL_3010 = _EVAL_1185 == 5'h0;
  assign _EVAL_1216 = _EVAL_298[1:0];
  assign _EVAL_2259 = _EVAL_1216 >= 2'h2;
  assign _EVAL_1777 = _EVAL_1216 == 2'h0;
  assign _EVAL_2027 = _EVAL_3010 ? _EVAL_2259 : _EVAL_1777;
  assign _EVAL_1391 = _EVAL_326[26:18];
  assign _EVAL_1321 = _EVAL_1391[8:2];
  assign _EVAL_723 = _EVAL_260[35:27];
  assign _EVAL_2065 = _EVAL_723[3:0];
  assign _EVAL_252 = _EVAL_723[8:4];
  assign _EVAL_205 = {_EVAL_2065,_EVAL_252};
  assign _EVAL_2481 = _EVAL_779 == 3'h4;
  assign _EVAL_1398 = _EVAL_995[6:2];
  assign _EVAL_406 = _EVAL_1398 == 5'h0;
  assign _EVAL_1065 = _EVAL_1545[0];
  assign _EVAL_497 = _EVAL_1545[1];
  assign _EVAL_3368 = _EVAL_406 ? _EVAL_1065 : _EVAL_497;
  assign _EVAL_1681 = _EVAL_497 == _EVAL_1065;
  assign _EVAL_2870 = {_EVAL_3368,_EVAL_1681};
  assign _EVAL_2630 = _EVAL_2481 ? _EVAL_2870 : _EVAL_1545;
  assign _EVAL_1741 = _EVAL_113 | packageanon1_1__EVAL_0;
  assign _EVAL_1048 = _EVAL_3304[1:0];
  assign _EVAL_421 = _EVAL_975 & _EVAL_1170;
  assign _EVAL_1486 = _EVAL_2192[9:1];
  assign _EVAL_281 = _EVAL_1486 == _EVAL_954;
  assign _EVAL_1576 = _EVAL_421 & _EVAL_281;
  assign _EVAL_2007 = _EVAL_534 | _EVAL_2748;
  assign _EVAL_1127 = _EVAL_2918 == 2'h2;
  assign _EVAL_3216 = _EVAL_2319 & _EVAL_1127;
  assign _EVAL_602 = _EVAL_3216 == 1'h0;
  assign _EVAL_926 = _EVAL_113 | packageanon1_5__EVAL_0;
  assign _EVAL_162 = _EVAL_3216 | _EVAL_926;
  assign _EVAL_1625 = _EVAL_602 & _EVAL_162;
  assign _EVAL_267 = _EVAL_1686 & _EVAL_1024;
  assign _EVAL_3309 = _EVAL_1343 | _EVAL_267;
  assign _EVAL_289 = _EVAL_3309 | _EVAL_848;
  assign _EVAL_290 = _EVAL_1924[10];
  assign _EVAL_323 = _EVAL_177[3:0];
  assign _EVAL_3214 = {_EVAL_323,_EVAL_3051};
  assign _EVAL_2006 = _EVAL_2518 & _EVAL_1463;
  assign _EVAL_1874 = _EVAL_2384 & _EVAL_1847;
  assign _EVAL_2827 = _EVAL_2006 | _EVAL_1874;
  assign _EVAL_2924 = _EVAL_2827 | _EVAL_2708;
  assign _EVAL_280 = _EVAL_3063 | _EVAL_3319;
  assign _EVAL_1484 = _EVAL_1276 & _EVAL_280;
  assign _EVAL_2694 = _EVAL_2924 | _EVAL_1484;
  assign _EVAL_2989 = _EVAL_3105 & _EVAL_1537;
  assign _EVAL_1667 = _EVAL_2694 | _EVAL_2989;
  assign _EVAL_2364 = _EVAL_2725[19:0];
  assign _EVAL_588 = tlb__EVAL_37[31:12];
  assign _EVAL_3349 = _EVAL_2364 == _EVAL_588;
  assign _EVAL_743 = _EVAL_308 != 2'h3;
  assign _EVAL_1944 = _EVAL_957 == 1'h0;
  assign _EVAL_2932 = _EVAL_2291[6:2];
  assign _EVAL_1905 = _EVAL_2932 == 5'h0;
  assign _EVAL_3205 = _EVAL_1952[0];
  assign _EVAL_2695 = _EVAL_1952[1];
  assign _EVAL_3322 = _EVAL_1905 ? _EVAL_3205 : _EVAL_2695;
  assign _EVAL_1608 = _EVAL_2695 == _EVAL_3205;
  assign _EVAL_1298 = {_EVAL_3322,_EVAL_1608};
  assign _EVAL_2648 = _EVAL_2392[14:0];
  assign _EVAL_1941 = _EVAL_2392;
  assign _EVAL_3164 = _EVAL_2337__EVAL_2338_data;
  assign _EVAL_451 = _EVAL_1664 ? _EVAL_1941 : _EVAL_3164;
  assign _EVAL_2124 = _EVAL_3001__EVAL_3002_data;
  assign _EVAL_2455 = _EVAL_1664 ? _EVAL_2821 : _EVAL_2124;
  assign _EVAL_688 = _EVAL_94[31:3];
  assign _EVAL_869 = {_EVAL_1435,_EVAL_2331,_EVAL_1129,_EVAL_2434,_EVAL_2256,_EVAL_1711,_EVAL_2285,_EVAL_904,_EVAL_2553};
  assign _EVAL_1820 = {_EVAL_1725,_EVAL_3043,_EVAL_1513,_EVAL_1443,_EVAL_2572,_EVAL_2521,_EVAL_854,_EVAL_1894,_EVAL_2387,_EVAL_869};
  assign _EVAL_3353 = {_EVAL_1820,_EVAL_791};
  assign _EVAL_1416 = _EVAL_3353[8:0];
  assign _EVAL_752 = _EVAL_1416[1:0];
  assign _EVAL_1493 = _EVAL_1416[8:2];
  assign _EVAL_1000 = {_EVAL_752,_EVAL_1493};
  assign _EVAL_359 = _EVAL_790 == 1'h0;
  assign _EVAL_2750 = _EVAL_359 | _EVAL_1790;
  assign _EVAL_633 = _EVAL_2750 ? _EVAL_2880 : _EVAL_2413;
  assign _EVAL_986 = _EVAL_359 | _EVAL_3149;
  assign _EVAL_2811 = _EVAL_986 ? 1'h0 : _EVAL_367;
  assign _EVAL_652 = _EVAL_260[8:0];
  assign _EVAL_1422 = _EVAL_652[0];
  assign _EVAL_486 = _EVAL_652[8:1];
  assign _EVAL_1597 = {_EVAL_1422,_EVAL_486};
  assign _EVAL_2195 = _EVAL_3295[8:2];
  assign _EVAL_3150 = {_EVAL_586,_EVAL_2195};
  assign _EVAL_574 = _EVAL_1597 ^ _EVAL_3150;
  assign _EVAL_1015 = _EVAL_1093[8:3];
  assign _EVAL_1166 = {_EVAL_3404,_EVAL_1015};
  assign _EVAL_775 = _EVAL_574 ^ _EVAL_1166;
  assign _EVAL_3366 = _EVAL_775 ^ _EVAL_205;
  assign _EVAL_3397 = {_EVAL_633,_EVAL_2811,_EVAL_3366,_EVAL_1751};
  assign _EVAL_3310 = _EVAL_3138[8:0];
  assign _EVAL_2300 = _EVAL_2227[12];
  assign _EVAL_3375 = _EVAL_2410 & _EVAL_2300;
  assign _EVAL_2639 = _EVAL_858 | _EVAL_3375;
  assign _EVAL_1231 = _EVAL_2639 | _EVAL_3315;
  assign _EVAL_806 = _EVAL_275 & _EVAL_1231;
  assign _EVAL_2565 = _EVAL_3026[35:27];
  assign _EVAL_1179 = _EVAL_2565[8:8];
  assign _EVAL_1393 = _EVAL_1071[6];
  assign _EVAL_1871 = _EVAL_1393 ? _EVAL_533 : _EVAL_2594;
  assign _EVAL_1809 = _EVAL_1871[127:2];
  assign _EVAL_1473 = _EVAL_1873 | _EVAL_1790;
  assign _EVAL_1568 = _EVAL_1473 ? _EVAL_2880 : _EVAL_2413;
  assign _EVAL_2324 = {{1'd0}, _EVAL_1279};
  assign _EVAL_2600 = ~ _EVAL_3406;
  assign _EVAL_2116 = 8'h1 << _EVAL_2312;
  assign _EVAL_3256 = _EVAL_2600 | _EVAL_2116;
  assign _EVAL_3350 = ~ _EVAL_3256;
  assign _EVAL_3091 = _EVAL_1440__EVAL_1441_data;
  assign _EVAL_353 = _EVAL_1336[15:2];
  assign _EVAL_3108 = _EVAL_314[4];
  assign _EVAL_3111 = _EVAL_3236 & _EVAL_3108;
  assign _EVAL_2998 = _EVAL_2864;
  assign _EVAL_2856 = _EVAL_2998;
  assign _EVAL_1347 = _EVAL_314[7];
  assign _EVAL_3371 = _EVAL_3236 & _EVAL_1347;
  assign _EVAL_2506 = _EVAL_3371 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_2912 = _EVAL_1580 == 3'h4;
  assign _EVAL_2628 = _EVAL_1336[6:2];
  assign _EVAL_2632 = _EVAL_2628 == 5'h0;
  assign _EVAL_1464 = _EVAL_3064[0];
  assign _EVAL_978 = _EVAL_3064[1];
  assign _EVAL_1675 = _EVAL_2632 ? _EVAL_1464 : _EVAL_978;
  assign _EVAL_2842 = _EVAL_978 == _EVAL_1464;
  assign _EVAL_2722 = {_EVAL_1675,_EVAL_2842};
  assign _EVAL_886 = _EVAL_2912 ? _EVAL_2722 : _EVAL_3064;
  assign _EVAL_1395 = _EVAL_2291[15:2];
  assign _EVAL_1623 = _EVAL_2755 == 3'h4;
  assign _EVAL_663 = _EVAL_1623 ? _EVAL_1298 : _EVAL_1952;
  assign _EVAL_2371 = {_EVAL_353,_EVAL_886,_EVAL_1395,_EVAL_663};
  assign _EVAL_1587 = _EVAL_995[15:2];
  assign _EVAL_2459 = _EVAL_2227[15:2];
  assign _EVAL_2072 = _EVAL_2068 == 3'h4;
  assign _EVAL_1086 = _EVAL_2056 ? _EVAL_2993 : _EVAL_2797;
  assign _EVAL_714 = {_EVAL_1086,_EVAL_165};
  assign _EVAL_2117 = _EVAL_2072 ? _EVAL_714 : _EVAL_2168;
  assign _EVAL_1013 = {_EVAL_1587,_EVAL_2630,_EVAL_2459,_EVAL_2117};
  assign _EVAL_2011 = {_EVAL_2371,_EVAL_1013};
  assign _EVAL_823 = _EVAL_2468 ? _EVAL_1350 : _EVAL_2011;
  assign _EVAL_1594 = _EVAL_2705 & _EVAL_1127;
  assign _EVAL_2990 = _EVAL_113 | packageanon1_6__EVAL_0;
  assign _EVAL_202 = _EVAL_1594 | _EVAL_2990;
  assign _EVAL_1951 = _EVAL_3026[26:18];
  assign _EVAL_2841 = _EVAL_1951[6:0];
  assign _EVAL_1912 = _EVAL_1951[8:7];
  assign _EVAL_3158 = {_EVAL_2841,_EVAL_1912};
  assign _EVAL_2470 = _EVAL_1891 ^ _EVAL_3158;
  assign _EVAL_2680 = _EVAL_2846[15:2];
  assign _EVAL_2691 = _EVAL_312 & _EVAL_743;
  assign _EVAL_1881 = _EVAL_1698 ? _EVAL_2224 : _EVAL_1629;
  assign _EVAL_1671 = {_EVAL_934,_EVAL_1881};
  assign _EVAL_1101 = _EVAL_2691 ? _EVAL_1671 : _EVAL_308;
  assign _EVAL_1918 = _EVAL_2151[15:2];
  assign _EVAL_1064 = _EVAL_2151[15:13];
  assign _EVAL_1251 = _EVAL_1064 == 3'h4;
  assign _EVAL_2318 = _EVAL_1251 & _EVAL_899;
  assign _EVAL_2469 = {_EVAL_2931,_EVAL_3241};
  assign _EVAL_1451 = _EVAL_2318 ? _EVAL_2469 : _EVAL_2825;
  assign _EVAL_747 = {_EVAL_2680,_EVAL_1101,_EVAL_1918,_EVAL_1451};
  assign _EVAL_3269 = _EVAL_3111 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_2471 = _EVAL_3269[39:32];
  assign _EVAL_1304 = _EVAL_1140__EVAL_1141_data;
  assign _EVAL_1560 = _EVAL_2468 ? _EVAL_1304 : _EVAL_3183;
  assign _EVAL_2670 = _EVAL_3325[2:0];
  assign _EVAL_2169 = {_EVAL_2670,_EVAL_2184};
  assign _EVAL_2735 = _EVAL_2868[17:9];
  assign _EVAL_2812 = _EVAL_2735[3:0];
  assign _EVAL_3199 = _EVAL_2735[8:4];
  assign _EVAL_440 = {_EVAL_2812,_EVAL_3199};
  assign _EVAL_1033 = _EVAL_2169 ^ _EVAL_440;
  assign _EVAL_1884 = _EVAL_1323[8:5];
  assign _EVAL_1723 = {_EVAL_2196,_EVAL_1884};
  assign _EVAL_2838 = _EVAL_1033 ^ _EVAL_1723;
  assign _EVAL_1446 = _EVAL_2868[35:27];
  assign _EVAL_2473 = _EVAL_1446[5:0];
  assign _EVAL_2769 = _EVAL_1446[8:6];
  assign _EVAL_2883 = {_EVAL_2473,_EVAL_2769};
  assign _EVAL_1950 = _EVAL_2838 ^ _EVAL_2883;
  assign _EVAL_802 = _EVAL_3138[26:18];
  assign _EVAL_887 = {1'h0,_EVAL_2406};
  assign _EVAL_1775 = _EVAL_2031 >> _EVAL_887;
  assign _EVAL_2329 = _EVAL_1775[0];
  assign _EVAL_2679 = _EVAL_2602 == _EVAL_588;
  assign _EVAL_1737 = _EVAL_2329 & _EVAL_2679;
  assign _EVAL_225 = _EVAL_1737 & _EVAL_2420;
  assign _EVAL_603 = _EVAL_1336[12];
  assign _EVAL_1872 = _EVAL_1537 & _EVAL_603;
  assign _EVAL_3125 = _EVAL_2396 | _EVAL_1872;
  assign _EVAL_2770 = _EVAL_1763 & _EVAL_3125;
  assign _EVAL_2311 = _EVAL_716 & _EVAL_1688;
  assign _EVAL_2128 = _EVAL_741[11];
  assign _EVAL_457 = _EVAL_1853 == 2'h0;
  assign _EVAL_2715 = _EVAL_449[3];
  assign _EVAL_1875 = _EVAL_449 + 4'h6;
  assign _EVAL_3195 = _EVAL_2715 ? _EVAL_1875 : _EVAL_449;
  assign _EVAL_2920 = {_EVAL_2918,_EVAL_708};
  assign _EVAL_1378 = _EVAL_2031 >> _EVAL_881;
  assign _EVAL_1624 = _EVAL_1378[0];
  assign _EVAL_1958 = _EVAL_656[35:27];
  assign _EVAL_410 = _EVAL_1958[3:0];
  assign _EVAL_661 = _EVAL_1958[8:4];
  assign _EVAL_422 = {_EVAL_410,_EVAL_661};
  assign _EVAL_2094 = _EVAL_2629 ? _EVAL_2721 : _EVAL_1394;
  assign _EVAL_2577 = _EVAL_1386 ? _EVAL_352 : _EVAL_2094;
  assign _EVAL_1392 = _EVAL_1902 & _EVAL_2749;
  assign _EVAL_186 = _EVAL_1392 & _EVAL_2128;
  assign _EVAL_2946 = _EVAL_1529 & _EVAL_145;
  assign _EVAL_1970 = _EVAL_2946 & _EVAL_1944;
  assign _EVAL_3101 = _EVAL_1970 & _EVAL_132;
  assign _EVAL_1707 = {_EVAL_1095,_EVAL_2028};
  assign _EVAL_2780 = _EVAL_656[26:18];
  assign _EVAL_3330 = _EVAL_2780[2:0];
  assign _EVAL_2086 = _EVAL_2780[8:3];
  assign _EVAL_212 = {_EVAL_3330,_EVAL_2086};
  assign _EVAL_742 = _EVAL_234[8:0];
  assign _EVAL_2699 = _EVAL_3304[6:2];
  assign _EVAL_3131 = _EVAL_2699 == 5'h0;
  assign _EVAL_2033 = _EVAL_1048 >= 2'h2;
  assign _EVAL_2869 = _EVAL_1048 == 2'h0;
  assign _EVAL_1409 = _EVAL_3131 ? _EVAL_2033 : _EVAL_2869;
  assign _EVAL_1740 = _EVAL_1765 == 3'h3;
  assign _EVAL_871 = _EVAL_2402[31:3];
  assign _EVAL_2110 = _EVAL_871[2:0];
  assign _EVAL_3074 = _EVAL_454 >> _EVAL_2110;
  assign _EVAL_1296 = _EVAL_1853 != 2'h3;
  assign _EVAL_2497 = _EVAL_2158 & _EVAL_211;
  assign _EVAL_908 = _EVAL_2042 | _EVAL_2497;
  assign _EVAL_510 = _EVAL_3351 | _EVAL_280;
  assign _EVAL_2381 = _EVAL_1276 & _EVAL_510;
  assign _EVAL_1322 = _EVAL_908 | _EVAL_2381;
  assign _EVAL_2752 = _EVAL_3105 & _EVAL_2152;
  assign _EVAL_762 = _EVAL_1322 | _EVAL_2752;
  assign _EVAL_2315 = _EVAL_2629 ? _EVAL_1748 : _EVAL_1165;
  assign _EVAL_2246 = _EVAL_1386 ? _EVAL_2887 : _EVAL_2315;
  assign _EVAL_1196 = _EVAL_3261 ? _EVAL_2189 : _EVAL_2246;
  assign _EVAL_1850 = _EVAL_1970 | _EVAL_271;
  assign _EVAL_2901 = _EVAL_616[14];
  assign _EVAL_596 = _EVAL_3387[26:18];
  assign _EVAL_3037 = _EVAL_1018 & _EVAL_350;
  assign _EVAL_1586 = _EVAL_2524[0];
  assign _EVAL_1302 = {_EVAL_1586,_EVAL_1971};
  assign _EVAL_2089 = _EVAL_46;
  assign _EVAL_3145 = _EVAL_3146[15:2];
  assign _EVAL_897 = _EVAL_981 | _EVAL_1332;
  assign _EVAL_2836 = _EVAL_897 ? 3'h3 : 3'h4;
  assign _EVAL_1744 = _EVAL_2716 ? 3'h2 : _EVAL_2836;
  assign _EVAL_2096 = _EVAL_1462 ? 3'h1 : _EVAL_1744;
  assign _EVAL_1334 = _EVAL_744__EVAL_745_data;
  assign _EVAL_351 = _EVAL_1797 != _EVAL_2304;
  assign _EVAL_789 = _EVAL_351 & _EVAL_576;
  assign _EVAL_969 = _EVAL_1841 != _EVAL_2882;
  assign _EVAL_673 = _EVAL_969 & _EVAL_3270;
  assign _EVAL_807 = _EVAL_2629 ? _EVAL_2571 : _EVAL_463;
  assign _EVAL_967 = _EVAL_1386 ? _EVAL_673 : _EVAL_807;
  assign _EVAL_1314 = _EVAL_3261 ? _EVAL_789 : _EVAL_967;
  assign _EVAL_627 = _EVAL_1314;
  assign _EVAL_1385 = _EVAL_2468 ? _EVAL_1334 : _EVAL_627;
  assign _EVAL_704 = _EVAL_2452[11];
  assign _EVAL_2214 = _EVAL_1410 & _EVAL_704;
  assign _EVAL_2637 = _EVAL_344 | _EVAL_1529;
  assign _EVAL_1043 = _EVAL_372 | _EVAL_2637;
  assign _EVAL_232 = _EVAL_1043 == 1'h0;
  assign _EVAL_2213 = _EVAL_3216 & _EVAL_162;
  assign _EVAL_2763 = _EVAL_1458 == 3'h4;
  assign _EVAL_209 = _EVAL_496 != 2'h3;
  assign _EVAL_1701 = _EVAL_2763 & _EVAL_209;
  assign _EVAL_987 = _EVAL_1701 ? _EVAL_214 : _EVAL_496;
  assign _EVAL_471 = _EVAL_2468 | _EVAL_1077;
  assign _EVAL_2249 = _EVAL_2275 ? 1'h0 : _EVAL_471;
  assign _EVAL_1548 = _EVAL_1664 ? _EVAL_2249 : _EVAL_471;
  assign _EVAL_3229 = _EVAL_2790 & _EVAL_1548;
  assign _EVAL_1842 = _EVAL_3229 != _EVAL_3037;
  assign _EVAL_390 = _EVAL_1774[6:2];
  assign _EVAL_1074 = _EVAL_725__EVAL_726_data;
  assign _EVAL_1795 = ~ _EVAL_2576;
  assign _EVAL_544 = _EVAL_1795 | 32'h1;
  assign _EVAL_1949 = _EVAL_344 == 1'h0;
  assign _EVAL_1381 = {2'h3,_EVAL_2406};
  assign _EVAL_3065 = _EVAL_2031 >> _EVAL_1381;
  assign _EVAL_1764 = _EVAL_3065[0];
  assign _EVAL_2098 = _EVAL_2640 ? tag_array__EVAL_11 : _EVAL_1023;
  assign _EVAL_1865 = _EVAL_2098[19:0];
  assign _EVAL_1417 = _EVAL_1865 == _EVAL_588;
  assign _EVAL_1811 = _EVAL_1764 & _EVAL_1417;
  assign _EVAL_2978 = _EVAL_2098[20];
  assign _EVAL_3280 = _EVAL_1811 & _EVAL_2978;
  assign _EVAL_354 = _EVAL_1624 & _EVAL_3349;
  assign _EVAL_3365 = _EVAL_354 & _EVAL_143;
  assign _EVAL_776 = {1'h1,_EVAL_2406};
  assign _EVAL_921 = _EVAL_2031 >> _EVAL_776;
  assign _EVAL_2243 = _EVAL_921[0];
  assign _EVAL_2939 = _EVAL_2640 ? tag_array__EVAL_1 : _EVAL_3225;
  assign _EVAL_334 = _EVAL_2939[19:0];
  assign _EVAL_3357 = _EVAL_334 == _EVAL_588;
  assign _EVAL_1088 = _EVAL_2243 & _EVAL_3357;
  assign _EVAL_1985 = _EVAL_2939[20];
  assign _EVAL_2505 = _EVAL_1088 & _EVAL_1985;
  assign _EVAL_991 = {1'h0,_EVAL_3280,_EVAL_3365,_EVAL_2505,_EVAL_225};
  assign _EVAL_3140 = _EVAL_742[2:0];
  assign _EVAL_401 = _EVAL_742[8:3];
  assign _EVAL_1722 = {_EVAL_3140,_EVAL_401};
  assign _EVAL_2984 = _EVAL_1722 ^ _EVAL_2875;
  assign _EVAL_3228 = _EVAL_1936[8:5];
  assign _EVAL_1030 = {_EVAL_2588,_EVAL_3228};
  assign _EVAL_2201 = _EVAL_2984 ^ _EVAL_1030;
  assign _EVAL_2926 = _EVAL_1057[26:18];
  assign _EVAL_1999 = _EVAL_2437[3];
  assign _EVAL_1247 = _EVAL_1999 ? 2'h0 : _EVAL_2664;
  assign _EVAL_1555 = {_EVAL_688,_EVAL_1247};
  assign _EVAL_3253 = {{1'd0}, _EVAL_1555};
  assign _EVAL_2555 = _EVAL_3353[17:9];
  assign _EVAL_674 = _EVAL_2555[2:0];
  assign _EVAL_3086 = _EVAL_2555[8:3];
  assign _EVAL_1449 = {_EVAL_674,_EVAL_3086};
  assign _EVAL_1005 = _EVAL_1000 ^ _EVAL_1449;
  assign _EVAL_482 = _EVAL_3353[26:18];
  assign _EVAL_585 = _EVAL_482[3:0];
  assign _EVAL_1316 = _EVAL_482[8:4];
  assign _EVAL_340 = {_EVAL_585,_EVAL_1316};
  assign _EVAL_3354 = _EVAL_1005 ^ _EVAL_340;
  assign _EVAL_1207 = _EVAL_2565[7:0];
  assign _EVAL_294 = {_EVAL_1207,_EVAL_1179};
  assign _EVAL_1757 = _EVAL_2470 ^ _EVAL_294;
  assign _EVAL_669 = _EVAL_1594 == 1'h0;
  assign _EVAL_610 = _EVAL_669 & _EVAL_202;
  assign _EVAL_3046 = _EVAL_2705 & _EVAL_979;
  assign _EVAL_1531 = _EVAL_3046 == 1'h0;
  assign _EVAL_1812 = _EVAL_591 == 1'h0;
  assign _EVAL_2976 = _EVAL_2010 & _EVAL_1812;
  assign _EVAL_488 = 256'h1 << _EVAL_2920;
  assign _EVAL_285 = _EVAL_2031 | _EVAL_488;
  assign _EVAL_1802 = ~ _EVAL_2031;
  assign _EVAL_1406 = _EVAL_1802 | _EVAL_488;
  assign _EVAL_734 = ~ _EVAL_1406;
  assign _EVAL_2889 = _EVAL_1584 & _EVAL_894;
  assign _EVAL_317 = _EVAL_2889;
  assign _EVAL_595 = _EVAL_317;
  assign _EVAL_701 = _EVAL_2011;
  assign _EVAL_985 = _EVAL_1537 & _EVAL_1596;
  assign _EVAL_2457 = _EVAL_1763 & _EVAL_985;
  assign _EVAL_2720 = _EVAL_1784 | _EVAL_2457;
  assign _EVAL_3165 = _EVAL_3394 | _EVAL_2720;
  assign _EVAL_1693 = _EVAL_1119__EVAL_1120_data;
  assign _EVAL_2961 = _EVAL_1664 ? _EVAL_3165 : _EVAL_1693;
  assign _EVAL_3254 = _EVAL_24 == 1'h0;
  assign _EVAL_2057 = _EVAL_206;
  assign _EVAL_3222 = _EVAL_1147__EVAL_1148_data;
  assign _EVAL_1337 = _EVAL_1908;
  assign _EVAL_1704 = _EVAL_2831[7:0];
  assign _EVAL_2265 = _EVAL_826[8:8];
  assign _EVAL_718 = _EVAL_912 >= 4'h6;
  assign _EVAL_3300 = _EVAL_912 - 4'h6;
  assign _EVAL_1606 = _EVAL_718 ? _EVAL_3300 : _EVAL_912;
  assign _EVAL_2987 = _EVAL_616[13];
  assign _EVAL_2669 = predictor_Queue__EVAL_13 & _EVAL_2200;
  assign _EVAL_799 = _EVAL_1924[0];
  assign _EVAL_801 = _EVAL_2001 | _EVAL_1790;
  assign _EVAL_2395 = _EVAL_390 == 5'h0;
  assign _EVAL_2982 = _EVAL_1853 >= 2'h2;
  assign _EVAL_630 = _EVAL_2395 ? _EVAL_457 : _EVAL_2982;
  assign _EVAL_1341 = _EVAL_2395 ? _EVAL_2982 : _EVAL_457;
  assign _EVAL_558 = {_EVAL_630,_EVAL_1341};
  assign _EVAL_1601 = _EVAL_738 & _EVAL_2053;
  assign _EVAL_1265 = _EVAL_1601 & _EVAL_2029;
  assign _EVAL_2322 = _EVAL_1265 ? _EVAL_731 : 1'h1;
  assign _EVAL_980 = _EVAL_450 & _EVAL_2322;
  assign _EVAL_3359 = _EVAL_83 | _EVAL_980;
  assign _EVAL_2203 = _EVAL_1953 | _EVAL_3359;
  assign _EVAL_1194 = _EVAL_1953 & _EVAL_2203;
  assign _EVAL_3362 = predictor_Queue__EVAL_1 & _EVAL_3233;
  assign _EVAL_1339 = _EVAL_3362 & _EVAL_1160;
  assign _EVAL_3190 = _EVAL_1110 & _EVAL_1339;
  assign _EVAL_3298 = _EVAL_1546[55:48];
  assign _EVAL_3374 = _EVAL_1684[17:9];
  assign _EVAL_1703 = _EVAL_3374[2:0];
  assign _EVAL_2772 = _EVAL_2969 | _EVAL_475;
  assign _EVAL_1191 = _EVAL_3344 & _EVAL_3324;
  assign _EVAL_795 = _EVAL_2772 | _EVAL_1191;
  assign _EVAL_2379 = _EVAL_1387 - 7'h1;
  assign _EVAL_507 = $unsigned(_EVAL_2379);
  assign _EVAL_2461 = _EVAL_507[6:0];
  assign _EVAL_2206 = _EVAL_1057[17:9];
  assign _EVAL_2449 = _EVAL_2206[8:7];
  assign _EVAL_1182 = _EVAL_2319 & _EVAL_979;
  assign _EVAL_1319 = _EVAL_1182 == 1'h0;
  assign _EVAL_685 = _EVAL_138;
  assign _EVAL_1776 = _EVAL_3144 > 5'h0;
  assign _EVAL_425 = _EVAL_1776 & _EVAL_2808;
  assign _EVAL_2004 = _EVAL_103 | _EVAL_425;
  assign _EVAL_662 = _EVAL_2149 ? 1'h0 : 1'h1;
  assign _EVAL_2906 = _EVAL_2700 & _EVAL_1235;
  assign _EVAL_2501 = _EVAL_254 + 2'h1;
  assign _EVAL_2017 = _EVAL_319__EVAL_320_data;
  assign _EVAL_1254 = _EVAL_1048 != 2'h3;
  assign _EVAL_1472 = _EVAL_2181 & _EVAL_1254;
  assign _EVAL_345 = _EVAL_3131 ? _EVAL_2869 : _EVAL_2033;
  assign _EVAL_1401 = {_EVAL_345,_EVAL_1409};
  assign _EVAL_1246 = _EVAL_1472 ? _EVAL_1401 : _EVAL_1048;
  assign _EVAL_1849 = _EVAL_2926[7:0];
  assign _EVAL_1055 = _EVAL_596[8:2];
  assign _EVAL_2884 = _EVAL_1774[15:13];
  assign _EVAL_1223 = _EVAL_2884 == 3'h4;
  assign _EVAL_2308 = _EVAL_1223 & _EVAL_1296;
  assign _EVAL_459 = _EVAL_1050[13:11];
  assign _EVAL_940 = {{8'd0}, _EVAL_459};
  assign _EVAL_1034 = _EVAL_1291 ^ _EVAL_940;
  assign _EVAL_2386 = _EVAL_2070 == 1'h0;
  assign _EVAL_592 = _EVAL_2386 & _EVAL_1213;
  assign _EVAL_1747 = _EVAL_3304[15:2];
  assign _EVAL_1710 = _EVAL_1460 ? _EVAL_1137 : _EVAL_399;
  assign _EVAL_1992 = {_EVAL_1747,_EVAL_1246,_EVAL_3145,_EVAL_1710};
  assign _EVAL_337 = _EVAL_865 & _EVAL_2934;
  assign _EVAL_1132 = _EVAL_337 == 1'h0;
  assign _EVAL_1477 = _EVAL_1132 & _EVAL_3327;
  assign _EVAL_905 = _EVAL_3227 == 1'h0;
  assign _EVAL_3273 = _EVAL_1603 | _EVAL_2661;
  assign _EVAL_3174 = _EVAL_1603 & _EVAL_666;
  assign _EVAL_1080 = _EVAL_1677 ? _EVAL_3273 : _EVAL_3174;
  assign _EVAL_173 = _EVAL_865 & _EVAL_1080;
  assign _EVAL_411 = _EVAL_173 == 1'h0;
  assign _EVAL_1485 = _EVAL_3310[6:0];
  assign _EVAL_370 = _EVAL_3310[8:7];
  assign _EVAL_3147 = {_EVAL_1485,_EVAL_370};
  assign _EVAL_2855 = _EVAL_3138[17:9];
  assign _EVAL_1092 = _EVAL_2855[7:0];
  assign _EVAL_1920 = _EVAL_2855[8:8];
  assign _EVAL_2527 = {_EVAL_1092,_EVAL_1920};
  assign _EVAL_1943 = _EVAL_3147 ^ _EVAL_2527;
  assign _EVAL_330 = _EVAL_1943 ^ _EVAL_802;
  assign _EVAL_1293 = _EVAL_330 ^ _EVAL_2823;
  assign _EVAL_2861 = tlb__EVAL_37[31:6];
  assign _EVAL_1942 = {_EVAL_2861, 6'h0};
  assign _EVAL_2586 = _EVAL_2468 ? _EVAL_3091 : _EVAL_2998;
  assign _EVAL_2126 = _EVAL_1475 == 1'h0;
  assign _EVAL_3104 = _EVAL_1970 & _EVAL_2126;
  assign _EVAL_1512 = _EVAL_3104 & _EVAL_1269;
  assign _EVAL_1333 = ~ _EVAL;
  assign _EVAL_2113 = _EVAL_1333 | 32'h1;
  assign _EVAL_1061 = ~ _EVAL_2113;
  assign _EVAL_774 = _EVAL_1664 ? _EVAL_627 : _EVAL_1164;
  assign _EVAL_2280 = _EVAL_2518 & _EVAL_795;
  assign _EVAL_890 = _EVAL_2280 | _EVAL_806;
  assign _EVAL_1509 = _EVAL_716 & _EVAL_289;
  assign _EVAL_1258 = _EVAL_890 | _EVAL_1509;
  assign _EVAL_2489 = _EVAL_234[35:27];
  assign _EVAL_383 = _EVAL_2489[8:6];
  assign _EVAL_392 = _EVAL_2299 ? 1'h0 : 1'h1;
  assign _EVAL_2908 = _EVAL_2001 | _EVAL_1192;
  assign _EVAL_1228 = {_EVAL_392,_EVAL_392,_EVAL_2054,_EVAL_2908};
  assign _EVAL_385 = _EVAL_916[7:0];
  assign _EVAL_2123 = _EVAL_2719 & _EVAL_2007;
  assign _EVAL_1201 = _EVAL_113 | packageanon1_3__EVAL_0;
  assign _EVAL_2858 = _EVAL_1182 | _EVAL_1201;
  assign _EVAL_1615 = _EVAL_83 ? {{7'd0}, _EVAL_121} : _EVAL_2576;
  assign _EVAL_2963 = {{121'd0}, _EVAL_3050};
  assign _EVAL_582 = {{128'd0}, _EVAL_1034};
  assign _EVAL_3182 = {_EVAL_2531, 11'h0};
  assign _EVAL_2409 = _EVAL_582 ^ _EVAL_3182;
  assign _EVAL_171 = _EVAL_2409[138:3];
  assign _EVAL_2526 = _EVAL_171[7:0];
  assign _EVAL_198 = _EVAL_2705 & _EVAL_1935;
  assign _EVAL_1646 = _EVAL_198 == 1'h0;
  assign _EVAL_2429 = _EVAL_113 | packageanon1_8__EVAL_0;
  assign _EVAL_1229 = _EVAL_198 | _EVAL_2429;
  assign _EVAL_3392 = _EVAL_1646 & _EVAL_1229;
  assign _EVAL_600 = _EVAL_1986__EVAL_1987_data;
  assign _EVAL_702 = _EVAL_2489[5:0];
  assign _EVAL_679 = {_EVAL_702,_EVAL_383};
  assign _EVAL_2408 = _EVAL_2201 ^ _EVAL_679;
  assign _EVAL_3383 = _EVAL_871[0];
  assign _EVAL_1900 = _EVAL_3383 == 1'h0;
  assign _EVAL_3052 = _EVAL_132 & _EVAL_1512;
  assign _EVAL_1726 = _EVAL_1161[26:18];
  assign _EVAL_2656 = _EVAL_1726[5:0];
  assign _EVAL_765 = _EVAL_1765 == 3'h1;
  assign _EVAL_448 = _EVAL_2515 & _EVAL_2741;
  assign _EVAL_2026 = _EVAL_1854[6:0];
  assign _EVAL_1135 = _EVAL_448 ? {{121'd0}, _EVAL_2026} : _EVAL_82;
  assign _EVAL_2153 = _EVAL_271 == 1'h0;
  assign _EVAL_2759 = _EVAL_2831[8:8];
  assign _EVAL_283 = _EVAL_1216 != 2'h3;
  assign _EVAL_3170 = _EVAL_3079;
  assign _EVAL_873 = _EVAL_542;
  assign _EVAL_1107 = _EVAL_403__EVAL_404_data;
  assign _EVAL_824 = _EVAL_1664 ? _EVAL_873 : _EVAL_1107;
  assign _EVAL_1264 = _EVAL_2926[8:8];
  assign _EVAL_2647 = {_EVAL_1849,_EVAL_1264};
  assign _EVAL_643 = _EVAL_2549[31:12];
  assign _EVAL_328 = _EVAL_3112__EVAL_3113_data;
  assign _EVAL_1017 = _EVAL_1954 ? 3'h0 : 3'h4;
  assign _EVAL_974 = _EVAL_2629 ? 3'h1 : _EVAL_1017;
  assign _EVAL_3085 = _EVAL_1386 ? 3'h2 : _EVAL_974;
  assign _EVAL_2127 = _EVAL_3261 ? 3'h3 : _EVAL_3085;
  assign _EVAL_1480 = _EVAL_2127;
  assign _EVAL_1713 = _EVAL_2468 ? _EVAL_328 : _EVAL_1480;
  assign _EVAL_1845 = _EVAL_3080 | _EVAL_1790;
  assign _EVAL_910 = _EVAL_1845 ? _EVAL_2880 : _EVAL_2413;
  assign _EVAL_784 = _EVAL_3257[8:0];
  assign _EVAL_2634 = _EVAL_784[6:0];
  assign _EVAL_1505 = _EVAL_784[8:7];
  assign _EVAL_327 = {_EVAL_2634,_EVAL_1505};
  assign _EVAL_2952 = {_EVAL_1704,_EVAL_2759};
  assign _EVAL_2624 = _EVAL_327 ^ _EVAL_2952;
  assign _EVAL_1084 = _EVAL_3257[26:18];
  assign _EVAL_3175 = _EVAL_2624 ^ _EVAL_1084;
  assign _EVAL_1349 = _EVAL_3175 ^ _EVAL_1302;
  assign _EVAL_1253 = {_EVAL_910,_EVAL_277,_EVAL_1349,_EVAL_1751};
  assign _EVAL_1532 = _EVAL_3046 | _EVAL_2368;
  assign _EVAL_382 = _EVAL_1763 & _EVAL_1193;
  assign _EVAL_1320 = _EVAL_501 | _EVAL_2252;
  assign _EVAL_434 = _EVAL_1774[15:2];
  assign _EVAL_2764 = _EVAL_298[15:13];
  assign _EVAL_2305 = _EVAL_1258 | _EVAL_2123;
  assign _EVAL_971 = _EVAL_2305 | _EVAL_2770;
  assign _EVAL_301 = _EVAL_1606[2:0];
  assign _EVAL_426 = _EVAL_3195[2:0];
  assign _EVAL_1738 = _EVAL_1981 & _EVAL_666;
  assign _EVAL_2104 = _EVAL_1677 ? _EVAL_456 : _EVAL_1738;
  assign _EVAL_1789 = _EVAL_865 & _EVAL_2104;
  assign _EVAL_2019 = _EVAL_1789 == 1'h0;
  assign _EVAL_1819 = _EVAL_2019 & _EVAL_3327;
  assign _EVAL_1541 = _EVAL_1102;
  assign _EVAL_1914 = _EVAL_1481__EVAL_1482_data;
  assign _EVAL_2222 = _EVAL_1664 ? _EVAL_1541 : _EVAL_1914;
  assign _EVAL_1450 = _EVAL_359 & _EVAL_1781;
  assign _EVAL_924 = _EVAL_2084 & _EVAL_959;
  assign _EVAL_3118 = _EVAL_2997[5:0];
  assign _EVAL_988 = _EVAL_1077 ? 1'h1 : _EVAL_350;
  assign _EVAL_2850 = _EVAL_2029 & _EVAL_2915;
  assign _EVAL_1656 = _EVAL_2850 ? 1'h1 : _EVAL_957;
  assign _EVAL_3390 = _EVAL_1664 ? _EVAL_1656 : _EVAL_1105;
  assign _EVAL_2914 = _EVAL_386__EVAL_387_data;
  assign _EVAL_2022 = _EVAL_326[17:9];
  assign _EVAL_1840 = _EVAL_2022[0];
  assign _EVAL_1364 = _EVAL_2022[8:1];
  assign _EVAL_2302 = {_EVAL_1840,_EVAL_1364};
  assign _EVAL_2532 = _EVAL_717 ^ _EVAL_2302;
  assign _EVAL_2460 = _EVAL_801 ? _EVAL_2880 : _EVAL_2413;
  assign _EVAL_1267 = _EVAL_3227 | _EVAL_1741;
  assign _EVAL_2654 = _EVAL_3227 & _EVAL_1267;
  assign _EVAL_3355 = _EVAL_36;
  assign _EVAL_151 = _EVAL_2468 ? _EVAL_2914 : _EVAL_1541;
  assign _EVAL_1835 = _EVAL_3362 & _EVAL_1213;
  assign _EVAL_195 = _EVAL_2386 & _EVAL_1835;
  assign _EVAL_2684 = _EVAL_1953 & _EVAL_3254;
  assign _EVAL_2598 = _EVAL_3259[26:18];
  assign _EVAL_640 = _EVAL_2598[5:0];
  assign _EVAL_1438 = _EVAL_3072 ? 3'h0 : _EVAL_2096;
  assign _EVAL_2548 = {_EVAL_1438, 1'h0};
  assign _EVAL_2091 = _EVAL_2548[3];
  assign _EVAL_3148 = _EVAL_2091 ? _EVAL_2175 : _EVAL_3009;
  assign _EVAL_1053 = _EVAL_961__EVAL_962_data;
  assign _EVAL_2800 = _EVAL_3261 ? _EVAL_1259 : _EVAL_2577;
  assign _EVAL_2955 = _EVAL_2800;
  assign _EVAL_692 = _EVAL_2468 ? _EVAL_1053 : _EVAL_2955;
  assign _EVAL_2456 = _EVAL_3214 ^ _EVAL_1707;
  assign _EVAL_435 = _EVAL_1726[8:6];
  assign _EVAL_1906 = {_EVAL_2656,_EVAL_435};
  assign _EVAL_2428 = _EVAL_2456 ^ _EVAL_1906;
  assign _EVAL_1674 = _EVAL_1518__EVAL_1519_data;
  assign _EVAL_2234 = _EVAL_3402 & _EVAL_232;
  assign _EVAL_2494 = _EVAL_2361;
  assign _EVAL_1285 = _EVAL_1684[8:0];
  assign _EVAL_3226 = _EVAL_1285[1:0];
  assign _EVAL_1650 = _EVAL_2177__EVAL_2178_data;
  assign _EVAL_1890 = _EVAL_2468 ? _EVAL_1650 : _EVAL_3165;
  assign _EVAL_2674 = _EVAL_2944 & _EVAL_2053;
  assign _EVAL_2667 = _EVAL_2674 & _EVAL_2029;
  assign _EVAL_1351 = _EVAL_2667 ? _EVAL_1523 : 1'h1;
  assign _EVAL_800 = _EVAL_3021 | _EVAL_2311;
  assign _EVAL_1770 = _EVAL_800 | _EVAL_1171;
  assign _EVAL_263 = _EVAL_1770 | _EVAL_382;
  assign _EVAL_2517 = _EVAL_1667 == 1'h0;
  assign _EVAL_911 = _EVAL_314[1];
  assign _EVAL_677 = _EVAL_3236 & _EVAL_911;
  assign _EVAL_458 = _EVAL_677 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_3271 = _EVAL_458[15:8];
  assign _EVAL_1198 = _EVAL_2229__EVAL_2230_data;
  assign _EVAL_1153 = _EVAL_1664 ? _EVAL_2011 : _EVAL_1198;
  assign _EVAL_1530 = _EVAL_314[5];
  assign _EVAL_398 = _EVAL_3236 & _EVAL_1530;
  assign _EVAL_2784 = _EVAL_398 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_1124 = _EVAL_2784[47:40];
  assign _EVAL_2310 = _EVAL_1873 | _EVAL_1192;
  assign _EVAL_224 = _EVAL_2468 ? _EVAL_1982 : _EVAL_873;
  assign _EVAL_2346 = _EVAL_530__EVAL_531_data;
  assign _EVAL_1590 = _EVAL_411 & _EVAL_3327;
  assign _EVAL_1571 = _EVAL_2548[2:0];
  assign _EVAL_1903 = _EVAL_1664 ? _EVAL_1571 : _EVAL_2346;
  assign _EVAL_2753 = _EVAL_1895__EVAL_1896_data;
  assign _EVAL_3235 = _EVAL_1531 & _EVAL_1532;
  assign _EVAL_1150 = _EVAL_1285[8:2];
  assign _EVAL_891 = {_EVAL_3226,_EVAL_1150};
  assign _EVAL_3073 = _EVAL_3374[8:3];
  assign _EVAL_1012 = {_EVAL_1703,_EVAL_3073};
  assign _EVAL_508 = _EVAL_891 ^ _EVAL_1012;
  assign _EVAL_2953 = _EVAL_152[3:0];
  assign _EVAL_447 = _EVAL_152[8:4];
  assign _EVAL_1225 = {_EVAL_2953,_EVAL_447};
  assign _EVAL_852 = _EVAL_508 ^ _EVAL_1225;
  assign _EVAL_2696 = _EVAL_418 != _EVAL_385;
  assign _EVAL_1286 = _EVAL_1850 == 1'h0;
  assign _EVAL_2665 = _EVAL_931__EVAL_932_data;
  assign _EVAL_1833 = _EVAL_1182 & _EVAL_2858;
  assign _EVAL_1329 = _EVAL_1953 ? {{7'd0}, _EVAL_1846} : _EVAL_1615;
  assign _EVAL_2627 = _EVAL_3074[0];
  assign _EVAL_2372 = _EVAL_1859__EVAL_1860_data[7:0];
  assign _EVAL_2919 = _EVAL_2491[7:0];
  assign _EVAL_2228 = _EVAL_2372 == _EVAL_2919;
  assign _EVAL_3103 = _EVAL_2627 & _EVAL_2228;
  assign _EVAL_2502 = _EVAL_450 == 1'h0;
  assign _EVAL_1212 = _EVAL_2843 & _EVAL_2502;
  assign _EVAL_1360 = _EVAL_982__EVAL_983_data;
  assign _EVAL_483 = _EVAL_1664 ? _EVAL_1480 : _EVAL_1360;
  assign _EVAL_409 = _EVAL_949__EVAL_950_data;
  assign _EVAL_1573 = _EVAL_298[15:2];
  assign _EVAL_668 = _EVAL_1765 == 3'h0;
  assign _EVAL_1156 = _EVAL_273 ? _EVAL_1714 : {{121'd0}, _EVAL_3050};
  assign _EVAL_291 = _EVAL_991 != 5'h0;
  assign _EVAL_1620 = _EVAL_1196;
  assign _EVAL_2247 = _EVAL_2468 ? _EVAL_2665 : _EVAL_1620;
  assign _EVAL_675 = _EVAL_1620;
  assign _EVAL_3176 = _EVAL_3162 != 26'h0;
  assign _EVAL_1852 = _EVAL_924 & _EVAL_3176;
  assign _EVAL_1542 = _EVAL_363__EVAL_364_data;
  assign _EVAL_1020 = _EVAL_2468 ? _EVAL_1542 : _EVAL_1908;
  assign _EVAL_877 = _EVAL_596[1:0];
  assign _EVAL_2786 = {_EVAL_877,_EVAL_1055};
  assign _EVAL_2682 = _EVAL_616[9];
  assign _EVAL_2793 = _EVAL_1716__EVAL_1717_data;
  assign _EVAL_3249 = _EVAL_113 ? _EVAL_2026 : _EVAL_3386;
  assign _EVAL_1730 = 128'h1 << _EVAL_3249;
  assign _EVAL_1046 = _EVAL_2737 ^ _EVAL_212;
  assign _EVAL_2917 = _EVAL_1046 ^ _EVAL_422;
  assign _EVAL_1832 = _EVAL_2506[63:56];
  assign _EVAL_1702 = _EVAL_314[3];
  assign _EVAL_3078 = _EVAL_3236 & _EVAL_1702;
  assign _EVAL_559 = _EVAL_3078 ? _EVAL_2534 : _EVAL_1641;
  assign _EVAL_2209 = _EVAL_559[31:24];
  assign _EVAL_964 = {_EVAL_1832,_EVAL_3298,_EVAL_1124,_EVAL_2471,_EVAL_2209,_EVAL_1498,_EVAL_3271,_EVAL_2826};
  assign _EVAL_1287 = _EVAL_741[10];
  assign _EVAL_2141 = _EVAL_1594 & _EVAL_202;
  assign _EVAL_1389 = _EVAL_1754[5:3];
  assign _EVAL_1040 = _EVAL_1859__EVAL_1860_data[39:8];
  assign _EVAL_2076 = _EVAL_142 == 1'h0;
  assign _EVAL_2438 = {{6'd0}, _EVAL_1389};
  assign _EVAL_1072 = _EVAL_2468 ? _EVAL_600 : _EVAL_2821;
  assign _EVAL_2401 = _EVAL_1765 == 3'h2;
  assign _EVAL_1284 = _EVAL_1391[1:0];
  assign _EVAL_2589 = {_EVAL_1284,_EVAL_1321};
  assign _EVAL_167 = _EVAL_837 | _EVAL_1730;
  assign _EVAL_1666 = ~ _EVAL_1730;
  assign _EVAL_2225 = _EVAL_837 & _EVAL_1666;
  assign _EVAL_1724 = _EVAL_2234 & _EVAL_83;
  assign _EVAL_2215 = _EVAL_1724 ? _EVAL_121 : _EVAL_1846;
  assign _EVAL_1112 = {{7'd0}, _EVAL_2215};
  assign _EVAL_1919 = _EVAL_344 | _EVAL_1692;
  assign _EVAL_2374 = _EVAL_762 == 1'h0;
  assign _EVAL_3305 = _EVAL_3031 & _EVAL_2374;
  assign _EVAL_2942 = _EVAL_2997[8:6];
  assign _EVAL_480 = {_EVAL_3118,_EVAL_2942};
  assign _EVAL_207 = _EVAL_2206[6:0];
  assign _EVAL_498 = {_EVAL_207,_EVAL_2449};
  assign _EVAL_2357 = _EVAL_480 ^ _EVAL_498;
  assign _EVAL_1699 = _EVAL_2357 ^ _EVAL_2647;
  assign _EVAL_2802 = _EVAL_2149 ? 9'h0 : 9'h1ff;
  assign _EVAL_1792 = {_EVAL_662,_EVAL_662,_EVAL_2802,_EVAL_2310};
  assign _EVAL_579 = _EVAL_1664 ? _EVAL_206 : _EVAL_2793;
  assign _EVAL_2483 = _EVAL_2548[2:0];
  assign _EVAL_3202 = _EVAL_2792 & _EVAL_3268;
  assign _EVAL_557 = _EVAL_2852__EVAL_2853_data;
  assign _EVAL_3367 = _EVAL_263 & _EVAL_2517;
  assign _EVAL_608 = _EVAL_89[31:12];
  assign _EVAL_443 = {_EVAL_608,_EVAL_2122,_EVAL_575};
  assign _EVAL_3246 = _EVAL_2010 | _EVAL_113;
  assign _EVAL_1563 = _EVAL_359 | _EVAL_1192;
  assign _EVAL_2820 = _EVAL_1529 & _EVAL_971;
  assign _EVAL_3224 = _EVAL_1664 ? _EVAL_2955 : _EVAL_3222;
  assign _EVAL_3385 = _EVAL_1810[15:2];
  assign _EVAL_539 = itim_array__EVAL_2;
  assign _EVAL_1647 = _EVAL_3165;
  assign _EVAL_1181 = _EVAL_3010 ? _EVAL_1777 : _EVAL_2259;
  assign _EVAL_838 = {_EVAL_1181,_EVAL_2027};
  assign _EVAL_918 = _EVAL_616[3];
  assign _EVAL_2923 = _EVAL_1450 ? 9'h0 : 9'h1ff;
  assign _EVAL_732 = _EVAL_636;
  assign _EVAL_2685 = _EVAL_1450 ? 1'h0 : 1'h1;
  assign _EVAL_379 = {_EVAL_2685,_EVAL_2685,_EVAL_2923,_EVAL_1563};
  assign _EVAL_1338 = _EVAL_616[1];
  assign _EVAL_3045 = _EVAL_616[15];
  assign _EVAL_948 = _EVAL_3335__EVAL_3336_data;
  assign _EVAL_218 = _EVAL_2468 ? _EVAL_948 : 1'h0;
  assign _EVAL_992 = _EVAL_3126 & _EVAL_3191;
  assign _EVAL_1869 = _EVAL_1786[15:2];
  assign _EVAL_1452 = _EVAL_2308 ? _EVAL_558 : _EVAL_1853;
  assign _EVAL_3252 = {_EVAL_1869,_EVAL_499,_EVAL_434,_EVAL_1452};
  assign _EVAL_2340 = {_EVAL_3062,_EVAL_2265};
  assign _EVAL_1326 = _EVAL_616[6];
  assign _EVAL_1447 = _EVAL_198 & _EVAL_1229;
  assign _EVAL_262 = _EVAL_3406 | _EVAL_2116;
  assign _EVAL_923 = _EVAL_2764 == 3'h4;
  assign _EVAL_1609 = _EVAL_923 & _EVAL_283;
  assign _EVAL_292 = _EVAL_1465__EVAL_1466_data;
  assign _EVAL_1380 = _EVAL_1664 ? _EVAL_2963 : _EVAL_292;
  assign _EVAL_154 = _EVAL_454 | _EVAL_2116;
  assign _EVAL_3306 = _EVAL_1541;
  assign _EVAL_2862 = _EVAL_2452[0];
  assign _EVAL_1506 = _EVAL_11;
  assign _EVAL_537 = _EVAL_1664 ? _EVAL_2450 : _EVAL_1635;
  assign _EVAL_840 = _EVAL_1609 ? _EVAL_838 : _EVAL_1216;
  assign _EVAL_780 = {_EVAL_1573,_EVAL_840,_EVAL_3385,_EVAL_987};
  assign _EVAL_3393 = _EVAL_1480;
  assign _EVAL_516 = _EVAL_34;
  assign _EVAL_634 = _EVAL_65;
  assign _EVAL_3036 = _EVAL_2192[0];
  assign _EVAL_593 = _EVAL_1941;
  assign _EVAL_570 = {{29'd0}, _EVAL_2483};
  assign _EVAL_821 = _EVAL_2073__EVAL_2074_data;
  assign _EVAL_1814 = _EVAL_741[0];
  assign _EVAL_1660 = _EVAL_1924[11];
  assign _EVAL_1637 = _EVAL_2927 & _EVAL_1660;
  assign _EVAL_2354 = _EVAL_2667 ? _EVAL_1272 : 1'h1;
  assign _EVAL_1801 = _EVAL_616[4];
  assign _EVAL_2776 = _EVAL_2573__EVAL_2574_data;
  assign _EVAL_545 = _EVAL_2468 ? _EVAL_2776 : _EVAL_2648;
  assign _EVAL_2956 = _EVAL_2591__EVAL_2592_data;
  assign _EVAL_642 = _EVAL_616[2];
  assign _EVAL_1600 = _EVAL_116;
  assign _EVAL_2118 = _EVAL_2963;
  assign _EVAL_2445 = _EVAL_3076 & _EVAL_2558;
  assign _EVAL_1454 = _EVAL_2705 & _EVAL_2109;
  assign _EVAL_2587 = _EVAL_113 | packageanon1_2__EVAL_0;
  assign _EVAL_1429 = _EVAL_1454 | _EVAL_2587;
  assign _EVAL_1348 = _EVAL_1953 == 1'h0;
  assign _EVAL_2416 = _EVAL_1348 & _EVAL_2203;
  assign _EVAL_3194 = _EVAL_2390 != _EVAL_1222;
  assign _EVAL_3134 = _EVAL_257 ? 1'h0 : 1'h1;
  assign _EVAL_2021 = _EVAL_847;
  assign _EVAL_3160 = _EVAL_2021;
  assign _EVAL_3243 = _EVAL_2532 ^ _EVAL_2589;
  assign _EVAL_2513 = _EVAL_1664 ? _EVAL_3183 : _EVAL_2017;
  assign _EVAL_1761 = _EVAL_616[8];
  assign _EVAL_1047 = _EVAL_2468 ? _EVAL_821 : _EVAL_636;
  assign _EVAL_681 = _EVAL_616[12];
  assign _EVAL_3328 = _EVAL_1765 == 3'h7;
  assign _EVAL_772 = _EVAL_627;
  assign _EVAL_2509 = _EVAL_273 ? _EVAL_3329 : {{15'd0}, _EVAL_287};
  assign _EVAL_2522 = _EVAL_729 ^ _EVAL_2340;
  assign _EVAL_1838 = _EVAL_2648;
  assign _EVAL_2348 = _EVAL_2001 | _EVAL_3149;
  assign _EVAL_952 = _EVAL_1664 ? _EVAL_2998 : _EVAL_1227;
  assign _EVAL_909 = _EVAL_1656;
  assign _EVAL_828 = _EVAL_2773__EVAL_2774_data;
  assign _EVAL_2643 = _EVAL_2468 ? _EVAL_828 : _EVAL_317;
  assign _EVAL_2847 = _EVAL_38 | _EVAL_2076;
  assign _EVAL_1003 = _EVAL_1454 == 1'h0;
  assign _EVAL_3124 = _EVAL_1003 & _EVAL_1429;
  assign _EVAL_2651 = _EVAL_2468 ? _EVAL_1674 : _EVAL_1941;
  assign _EVAL_2873 = {_EVAL_1809, 2'h0};
  assign _EVAL_812 = _EVAL_2468 ? _EVAL_557 : _EVAL_1656;
  assign _EVAL_1574 = _EVAL_344 & _EVAL_1286;
  assign _EVAL_438 = _EVAL_1765 == 3'h5;
  assign _EVAL_505 = _EVAL_1664 ? 1'h0 : _EVAL_409;
  assign _EVAL_2034 = _EVAL_873;
  assign _EVAL_1521 = _EVAL_2348 ? 1'h0 : _EVAL_367;
  assign _EVAL_361 = _EVAL_30;
  assign _EVAL_3024 = _EVAL_2468 ? _EVAL_730 : _EVAL_2021;
  assign _EVAL_1843 = _EVAL_2468 ? _EVAL_2529 : _EVAL_2963;
  assign _EVAL_3279 = _EVAL_1377 ? _EVAL_2461 : _EVAL_1387;
  assign _EVAL_415 = _EVAL_316 ? _EVAL_1158 : _EVAL_3279;
  assign _EVAL_2298 = _EVAL_2667 ? _EVAL_2399 : 1'h1;
  assign _EVAL_2562 = _EVAL_113 ? _EVAL_1135 : {{121'd0}, _EVAL_2988};
  assign _EVAL_1745 = _EVAL_424 | _EVAL_2438;
  assign _EVAL_2421 = _EVAL_2712__EVAL_2713_data;
  assign _EVAL_2731 = _EVAL_2598[8:6];
  assign _EVAL_509 = {_EVAL_640,_EVAL_2731};
  assign _EVAL_3339 = _EVAL_2478__EVAL_2479_data;
  assign _EVAL_1457 = _EVAL_1664 ? _EVAL_2648 : _EVAL_3339;
  assign _EVAL_2055 = _EVAL_2821;
  assign _EVAL_3403 = _EVAL_3148 | _EVAL_570;
  assign _EVAL_1408 = _EVAL_3167 | _EVAL_3327;
  assign _EVAL_2945 = _EVAL_2667 ? _EVAL_664 : 1'h1;
  assign _EVAL_2819 = _EVAL_1765 == 3'h4;
  assign _EVAL_2435 = _EVAL_113 == 1'h0;
  assign _EVAL_893 = _EVAL_3046 & _EVAL_1532;
  assign _EVAL_2488 = _EVAL_1320 | _EVAL_1288;
  assign _EVAL_1239 = _EVAL_2192[11];
  assign _EVAL_736 = _EVAL_1576 & _EVAL_1239;
  assign _EVAL_612 = _EVAL_1664 ? _EVAL_2021 : _EVAL_2421;
  assign _EVAL_2611 = _EVAL_1664 ? _EVAL_1620 : _EVAL_1074;
  assign _EVAL_2830 = _EVAL_1664 ? _EVAL_317 : _EVAL_2753;
  assign _EVAL_631 = _EVAL_1123 ^ _EVAL_509;
  assign _EVAL_1690 = _EVAL_1319 & _EVAL_2858;
  assign _EVAL_208 = _EVAL_1454 & _EVAL_1429;
  assign _EVAL_1470 = _EVAL_905 & _EVAL_1267;
  assign _EVAL_2102 = _EVAL_44;
  assign _EVAL_3077 = _EVAL_1497 ^ _EVAL_2786;
  assign _EVAL_526 = _EVAL_2955;
  assign _EVAL_2844 = {_EVAL_1568,_EVAL_1619,_EVAL_1950,_EVAL_1751};
  assign _EVAL_1892 = _EVAL_18;
  assign _EVAL_597 = _EVAL_2468 ? _EVAL_2956 : _EVAL_1571;
  assign _EVAL_2313 = _EVAL_1571;
  assign _EVAL_2362 = {_EVAL_2460,_EVAL_1521,_EVAL_1757,_EVAL_1751};
  assign _EVAL_793 = _EVAL_16;
  assign _EVAL_611 = _EVAL_1664 ? _EVAL_1908 : _EVAL_2511;
  assign predictor_base_table_1__EVAL = _EVAL_2070 | _EVAL_195;
  assign predictor_tagged_tables_2__EVAL_2 = _EVAL_1228[10];
  assign predictor_base_table_0__EVAL_21 = _EVAL_2226 & _EVAL_2669;
  assign predictor_tagged_tables_3__EVAL_3 = _EVAL_1980[1];
  assign predictor_tagged_tables_2__EVAL_4 = _EVAL_228;
  assign predictor_tagged_tables_0__EVAL_20 = _EVAL_379[8];
  assign predictor_base_table_1__EVAL_16 = _EVAL_2819 & _EVAL_2669;
  assign predictor_tagged_tables_1__EVAL_31 = _EVAL_1792[7];
  assign tlb__EVAL_49 = _EVAL_88;
  assign data_arrays_2_1__EVAL = _EVAL_610 | _EVAL_2141;
  assign data_arrays_2_0__EVAL = _EVAL_1625 | _EVAL_2213;
  assign predictor_tagged_tables_1__EVAL_32 = _EVAL_1792[0];
  assign predictor_tagged_tables_1__EVAL_37 = _EVAL_2844[11];
  assign predictor_tagged_tables_2__EVAL_5 = _EVAL_1228[4];
  assign tlb__EVAL_14 = _EVAL_41;
  assign predictor_tagged_tables_1__EVAL_16 = _EVAL_2844[0];
  assign predictor_tagged_tables_1__EVAL_17 = _EVAL_1792[2];
  assign predictor_tagged_tables_0__EVAL_2 = _EVAL_379[10];
  assign predictor_Queue__EVAL_8 = _EVAL_2102;
  assign data_arrays_2_0__EVAL_3 = icache_clock_gate_out;
  assign tlb__EVAL_38 = _EVAL_134;
  assign _EVAL_108 = _EVAL_3104 & _EVAL_1269;
  assign predictor_tagged_tables_0__EVAL_23 = _EVAL_3397[4];
  assign predictor_tagged_tables_1__EVAL_29 = _EVAL_2844[7];
  assign tag_array__EVAL_5 = _EVAL_2918 == 2'h0;
  assign predictor_tagged_tables_0__EVAL_5 = _EVAL_379[4];
  assign predictor_Queue__EVAL = _EVAL_3253;
  assign MaxPeriodFibonacciLFSR_1__EVAL_13 = _EVAL_44;
  assign predictor_tagged_tables_2__EVAL_23 = _EVAL_2362[4];
  assign data_arrays_3_1__EVAL_2 = _EVAL_2705 & _EVAL_1935;
  assign tlb__EVAL_55 = _EVAL_87;
  assign data_arrays_1_0__EVAL_3 = icache_clock_gate_out;
  assign _EVAL_124 = _EVAL_774;
  assign _EVAL_99 = _EVAL_2455;
  assign predictor_tagged_tables_0__EVAL_4 = _EVAL_228;
  assign predictor_base_table_0__EVAL_28 = predictor_Queue__EVAL_9;
  assign data_arrays_2_1__EVAL_1 = _EVAL_1745[8:1];
  assign predictor_tagged_tables_2__EVAL_14 = _EVAL_2362[6];
  assign _EVAL_31 = _EVAL_1903;
  assign packageanon1_6__EVAL = _EVAL_1771 & _EVAL_2298;
  assign _EVAL_26 = _EVAL_2830;
  assign tlb__EVAL_6 = _EVAL_112;
  assign tlb__EVAL_24 = _EVAL_105;
  assign _EVAL_25 = _EVAL_505;
  assign packageanon1_7__EVAL = _EVAL_992 & _EVAL_2945;
  assign predictor_base_table_0__EVAL_25 = _EVAL_2669 == 1'h0;
  assign predictor_tagged_tables_0__EVAL_14 = _EVAL_3397[6];
  assign tlb__EVAL_56 = _EVAL_4;
  assign data_arrays_3_0__EVAL_2 = _EVAL_2319 & _EVAL_1935;
  assign _EVAL_66 = _EVAL_2549;
  assign tlb__EVAL_21 = _EVAL_81;
  assign tag_array__EVAL = _EVAL_1754[11:6];
  assign tlb__EVAL_59 = _EVAL_130;
  assign predictor_tagged_tables_0__EVAL_22 = _EVAL_3397[9];
  assign MaxPeriodFibonacciLFSR__EVAL_15 = icache_clock_gate_out;
  assign tlb__EVAL_16 = _EVAL_3143;
  assign _EVAL_62 = _EVAL_1380;
  assign _EVAL_110 = _EVAL_1953;
  assign tlb__EVAL_40 = _EVAL_50;
  assign predictor_tagged_tables_1__EVAL_26 = _EVAL_2844[3];
  assign tlb__EVAL_8 = _EVAL_74;
  assign data_arrays_0_1__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign predictor_tagged_tables_1__EVAL_11 = _EVAL_865 & _EVAL_2934;
  assign _EVAL_22 = _EVAL_40 & _EVAL_14;
  assign predictor_tagged_tables_2__EVAL_28 = _EVAL_2362[8];
  assign _EVAL_96 = _EVAL_1457;
  assign _EVAL_91 = _EVAL_612;
  assign data_arrays_0_0__EVAL_2 = _EVAL_2319 & _EVAL_2109;
  assign _EVAL_61 = _EVAL_451;
  assign predictor_base_table_0__EVAL_12 = _EVAL_1740 & _EVAL_2669;
  assign predictor_base_table_0__EVAL_18 = _EVAL_668 & _EVAL_2669;
  assign data_arrays_0_1__EVAL_1 = _EVAL_1745[8:1];
  assign predictor_base_table_0__EVAL_20 = _EVAL_2401 & _EVAL_2669;
  assign predictor_tagged_tables_3__EVAL_14 = _EVAL_1253[6];
  assign _EVAL_125 = _EVAL_824;
  assign tlb__EVAL_18 = _EVAL_13;
  assign predictor_tagged_tables_2__EVAL_32 = _EVAL_1228[0];
  assign tlb__EVAL_13 = _EVAL_33;
  assign predictor_base_table_1__EVAL_12 = _EVAL_1740 & _EVAL_2669;
  assign predictor_tagged_tables_1__EVAL_2 = _EVAL_1792[10];
  assign predictor_base_table_0__EVAL_15 = _EVAL_765 & _EVAL_2669;
  assign predictor_tagged_tables_3__EVAL_21 = _EVAL_1253[10];
  assign itim_array__EVAL_1 = _EVAL_1329[14:3];
  assign predictor_tagged_tables_2__EVAL_6 = _EVAL_1228[5];
  assign predictor_base_table_0__EVAL_9 = _EVAL_3069 == 1'h0;
  assign predictor_base_table_1__EVAL_19 = predictor_Queue__EVAL_9;
  assign tag_array__EVAL_13 = icache_clock_gate_out;
  assign data_arrays_3_0__EVAL_3 = icache_clock_gate_out;
  assign predictor_tagged_tables_1__EVAL_24 = _EVAL_2844[1];
  assign predictor_tagged_tables_2__EVAL = _EVAL_1228[11];
  assign predictor_base_table_1__EVAL_4 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_0__EVAL_17 = _EVAL_379[2];
  assign _EVAL_17 = _EVAL_2637 == 1'h0;
  assign predictor_base_table_0__EVAL_14 = predictor_Queue__EVAL_9;
  assign predictor_Queue__EVAL_3 = _EVAL_1506;
  assign tlb__EVAL_30 = _EVAL_70;
  assign data_arrays_2_0__EVAL_2 = _EVAL_2319 & _EVAL_1127;
  assign predictor_tagged_tables_3__EVAL_23 = _EVAL_1253[4];
  assign packageanon1_8__EVAL = _EVAL_1771 & _EVAL_2945;
  assign predictor_tagged_tables_1__EVAL_33 = _EVAL_1792[3];
  assign packageanon1_3__EVAL = _EVAL_992 & _EVAL_2354;
  assign tlb__EVAL_11 = _EVAL_28;
  assign predictor_Queue__EVAL_7 = _EVAL_228;
  assign _EVAL_53 = _EVAL_1153;
  assign tlb__EVAL_50 = _EVAL_93;
  assign predictor_tagged_tables_1__EVAL_30 = _EVAL_1792[6];
  assign predictor_tagged_tables_0__EVAL_6 = _EVAL_379[5];
  assign _EVAL_107 = _EVAL_1522;
  assign predictor_tagged_tables_1__EVAL_4 = _EVAL_228;
  assign tlb__EVAL_62 = _EVAL_58;
  assign predictor_base_table_0__EVAL_23 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_0__EVAL_37 = _EVAL_3397[11];
  assign predictor_tagged_tables_3__EVAL_16 = _EVAL_1253[0];
  assign tlb__EVAL_35 = _EVAL_117;
  assign _EVAL_133 = _EVAL_3402 & _EVAL_232;
  assign tag_array__EVAL_10 = _EVAL_10;
  assign MaxPeriodFibonacciLFSR__EVAL_9 = _EVAL_2292 & _EVAL_1176;
  assign predictor_tagged_tables_0__EVAL_32 = _EVAL_379[0];
  assign predictor_tagged_tables_0__EVAL_28 = _EVAL_3397[8];
  assign predictor_Queue__EVAL_4 = _EVAL_3355;
  assign tlb__EVAL_42 = _EVAL_67;
  assign tlb__EVAL_34 = _EVAL_92;
  assign tlb__EVAL_4 = _EVAL_5;
  assign itim_array__EVAL_3 = _EVAL_2416 | _EVAL_1194;
  assign predictor_base_table_1__EVAL_5 = predictor_Queue__EVAL_9;
  assign predictor_base_table_1__EVAL_15 = _EVAL_765 & _EVAL_2669;
  assign predictor_Queue__EVAL_10 = _EVAL_516;
  assign _EVAL_56 = _EVAL_611;
  assign predictor_tagged_tables_2__EVAL_22 = _EVAL_2362[9];
  assign predictor_tagged_tables_2__EVAL_16 = _EVAL_2362[0];
  assign predictor_base_table_1__EVAL_29 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_2__EVAL_20 = _EVAL_1228[8];
  assign predictor_tagged_tables_3__EVAL_30 = _EVAL_1980[6];
  assign predictor_tagged_tables_1__EVAL = _EVAL_1792[11];
  assign itim_array__EVAL_0 = _EVAL_1953;
  assign itim_array__EVAL = icache_clock_gate_out;
  assign predictor_tagged_tables_0__EVAL_15 = _EVAL_3156 ? _EVAL_3243 : _EVAL_3077;
  assign predictor_tagged_tables_2__EVAL_38 = _EVAL_1228[9];
  assign predictor_tagged_tables_3__EVAL_5 = _EVAL_1980[4];
  assign _EVAL_69 = _EVAL_3292;
  assign packageanon1__EVAL_0 = _EVAL_10 ? _EVAL_443 : _EVAL_89;
  assign predictor_tagged_tables_2__EVAL_30 = _EVAL_1228[6];
  assign data_arrays_0_1__EVAL_3 = icache_clock_gate_out;
  assign predictor_tagged_tables_0__EVAL_29 = _EVAL_3397[7];
  assign tlb__EVAL_41 = _EVAL_27;
  assign tlb__EVAL_20 = _EVAL_44;
  assign tlb__EVAL_19 = _EVAL_6;
  assign predictor_base_table_0__EVAL_5 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_2__EVAL_31 = _EVAL_1228[7];
  assign predictor_tagged_tables_3__EVAL_38 = _EVAL_1980[9];
  assign tlb__EVAL_29 = _EVAL_109;
  assign predictor_tagged_tables_1__EVAL_5 = _EVAL_1792[4];
  assign tlb__EVAL_51 = _EVAL_9;
  assign tlb__EVAL_60 = _EVAL_123;
  assign predictor_tagged_tables_1__EVAL_23 = _EVAL_2844[4];
  assign predictor_tagged_tables_3__EVAL_2 = _EVAL_1980[10];
  assign icache_clock_gate_en = _EVAL_3402 | _EVAL_19;
  assign predictor_tagged_tables_3__EVAL_26 = _EVAL_1253[3];
  assign predictor_tagged_tables_0__EVAL_31 = _EVAL_379[7];
  assign data_arrays_0_0__EVAL_1 = _EVAL_1745[8:1];
  assign data_arrays_3_1__EVAL_1 = _EVAL_1745[8:1];
  assign packageanon1_5__EVAL = _EVAL_992 & _EVAL_2298;
  assign predictor_tagged_tables_3__EVAL_17 = _EVAL_1980[2];
  assign tlb__EVAL_43 = _EVAL_42;
  assign predictor_Queue__EVAL_6 = _EVAL_2873;
  assign predictor_base_table_1__EVAL_23 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_3__EVAL_6 = _EVAL_1980[5];
  assign data_arrays_1_0__EVAL_1 = _EVAL_1745[8:1];
  assign data_arrays_1_0__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign tlb__EVAL_48 = _EVAL_0;
  assign tlb__EVAL_58 = _EVAL_136;
  assign _EVAL_84 = _EVAL_537;
  assign predictor_tagged_tables_3__EVAL_12 = _EVAL_1253[5];
  assign predictor_tagged_tables_1__EVAL_15 = _EVAL_337 ? _EVAL_852 : _EVAL_3354;
  assign predictor_base_table_0__EVAL_19 = predictor_Queue__EVAL_9;
  assign data_arrays_1_1__EVAL = _EVAL_3235 | _EVAL_893;
  assign tlb__EVAL_15 = _EVAL_60;
  assign predictor_tagged_tables_3__EVAL_32 = _EVAL_1980[0];
  assign predictor_tagged_tables_2__EVAL_12 = _EVAL_2362[5];
  assign _EVAL_79 = _EVAL_952;
  assign predictor_tagged_tables_3__EVAL_9 = _EVAL_1819 | _EVAL_1789;
  assign tag_array__EVAL_4 = _EVAL_2906 | _EVAL_146;
  assign _EVAL_76 = _EVAL_1822 ? 3'h0 : 3'h1;
  assign _EVAL_111 = _EVAL_3390;
  assign data_arrays_0_1__EVAL_2 = _EVAL_2705 & _EVAL_2109;
  assign tlb__EVAL_0 = _EVAL_140;
  assign _EVAL_72 = _EVAL_132 & _EVAL_1512;
  assign data_arrays_0_1__EVAL = _EVAL_3124 | _EVAL_208;
  assign data_arrays_0_0__EVAL = _EVAL_1470 | _EVAL_2654;
  assign data_arrays_1_1__EVAL_1 = _EVAL_1745[8:1];
  assign predictor_tagged_tables_1__EVAL_12 = _EVAL_2844[5];
  assign predictor_base_table_0__EVAL_24 = predictor_Queue__EVAL_9 != predictor_Queue__EVAL_11;
  assign data_arrays_2_1__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign predictor_tagged_tables_0__EVAL_21 = _EVAL_3397[10];
  assign predictor_tagged_tables_0__EVAL_3 = _EVAL_379[1];
  assign data_arrays_1_0__EVAL_2 = _EVAL_2319 & _EVAL_979;
  assign predictor_tagged_tables_0__EVAL_12 = _EVAL_3397[5];
  assign tlb__EVAL_57 = _EVAL_2402;
  assign predictor_tagged_tables_3__EVAL_20 = _EVAL_1980[8];
  assign predictor_base_table_0__EVAL_2 = _EVAL_228;
  assign data_arrays_1_0__EVAL = _EVAL_1690 | _EVAL_1833;
  assign packageanon1_1__EVAL = _EVAL_992 & _EVAL_1351;
  assign _EVAL_106 = _EVAL_579;
  assign predictor_tagged_tables_2__EVAL_1 = _EVAL_2362[2];
  assign predictor_tagged_tables_2__EVAL_15 = _EVAL_173 ? _EVAL_2428 : _EVAL_631;
  assign predictor_tagged_tables_3__EVAL_11 = _EVAL_865 & _EVAL_2104;
  assign predictor_base_table_0__EVAL_8 = _EVAL_3190 ? _EVAL_2619 : _EVAL_2526;
  assign tlb__EVAL_28 = _EVAL_7;
  assign predictor_tagged_tables_0__EVAL_33 = _EVAL_379[3];
  assign _EVAL_126 = _EVAL_2513;
  assign predictor_tagged_tables_2__EVAL_11 = _EVAL_865 & _EVAL_1080;
  assign predictor_base_table_1__EVAL_28 = predictor_Queue__EVAL_9;
  assign _EVAL_135 = _EVAL_988;
  assign predictor_tagged_tables_1__EVAL_21 = _EVAL_2844[10];
  assign predictor_tagged_tables_3__EVAL_1 = _EVAL_1253[2];
  assign _EVAL_127 = _EVAL_2961;
  assign data_arrays_1_1__EVAL_2 = _EVAL_2705 & _EVAL_979;
  assign tlb__EVAL_2 = _EVAL_1762;
  assign predictor_base_table_1__EVAL_9 = _EVAL_2070 == 1'h0;
  assign predictor_base_table_1__EVAL_8 = _EVAL_195 ? _EVAL_2619 : _EVAL_2526;
  assign tlb__EVAL_27 = _EVAL_101;
  assign predictor_tagged_tables_1__EVAL_28 = _EVAL_2844[8];
  assign predictor_tagged_tables_1__EVAL_3 = _EVAL_1792[1];
  assign predictor_tagged_tables_3__EVAL = _EVAL_1980[11];
  assign MaxPeriodFibonacciLFSR_1__EVAL_15 = icache_clock_gate_out;
  assign tag_array__EVAL_8 = _EVAL_2918 == 2'h3;
  assign predictor_tagged_tables_2__EVAL_24 = _EVAL_2362[1];
  assign tag_array__EVAL_6 = _EVAL_2918 == 2'h2;
  assign predictor_tagged_tables_2__EVAL_37 = _EVAL_2362[11];
  assign _EVAL_14 = 1'h0;
  assign predictor_base_table_1__EVAL_25 = _EVAL_2669 == 1'h0;
  assign data_arrays_3_0__EVAL = _EVAL_1108 | _EVAL_3202;
  assign tlb__EVAL_33 = _EVAL_119;
  assign data_arrays_2_1__EVAL_2 = _EVAL_2705 & _EVAL_1127;
  assign MaxPeriodFibonacciLFSR_1__EVAL_9 = _EVAL_3129 & _EVAL_10;
  assign predictor_tagged_tables_1__EVAL_14 = _EVAL_2844[6];
  assign data_arrays_2_1__EVAL_3 = icache_clock_gate_out;
  assign predictor_base_table_0__EVAL_11 = _EVAL_438 & _EVAL_2669;
  assign icache_clock_gate_in = _EVAL_57;
  assign predictor_tagged_tables_2__EVAL_3 = _EVAL_1228[1];
  assign predictor_base_table_1__EVAL_3 = _EVAL_3328 & _EVAL_2669;
  assign predictor_base_table_1__EVAL_11 = _EVAL_438 & _EVAL_2669;
  assign predictor_tagged_tables_3__EVAL_31 = _EVAL_1980[7];
  assign predictor_tagged_tables_0__EVAL = _EVAL_379[11];
  assign predictor_tagged_tables_1__EVAL_38 = _EVAL_1792[9];
  assign tlb__EVAL_44 = _EVAL_21;
  assign predictor_tagged_tables_3__EVAL_22 = _EVAL_1253[9];
  assign predictor_base_table_1__EVAL_24 = predictor_Queue__EVAL_9 != predictor_Queue__EVAL_11;
  assign predictor_tagged_tables_2__EVAL_17 = _EVAL_1228[2];
  assign tlb__EVAL_17 = _EVAL_95;
  assign predictor_base_table_1__EVAL_2 = _EVAL_228;
  assign predictor_tagged_tables_0__EVAL_26 = _EVAL_3397[3];
  assign tlb__EVAL = _EVAL_90;
  assign predictor_tagged_tables_3__EVAL_24 = _EVAL_1253[1];
  assign tlb__EVAL_52 = _EVAL_47;
  assign predictor_tagged_tables_2__EVAL_33 = _EVAL_1228[3];
  assign itim_array__EVAL_4 = {_EVAL_747,_EVAL_780};
  assign tlb__EVAL_22 = _EVAL_59;
  assign data_arrays_3_1__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign tlb__EVAL_54 = _EVAL_8;
  assign tag_array__EVAL_12 = {_EVAL_2004,_EVAL_643};
  assign packageanon1_4__EVAL = _EVAL_1771 & _EVAL_2354;
  assign predictor_Queue__EVAL_5 = _EVAL_592 ? 1'h1 : _EVAL_3013;
  assign tlb__EVAL_47 = _EVAL_55;
  assign tlb__EVAL_9 = _EVAL_68;
  assign predictor_tagged_tables_2__EVAL_9 = _EVAL_1590 | _EVAL_173;
  assign data_arrays_2_0__EVAL_1 = _EVAL_1745[8:1];
  assign predictor_base_table_1__EVAL_26 = predictor_Queue__EVAL_9;
  assign predictor_base_table_0__EVAL_4 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_0__EVAL_1 = _EVAL_3397[2];
  assign tlb__EVAL_61 = _EVAL_64;
  assign predictor_tagged_tables_0__EVAL_38 = _EVAL_379[9];
  assign tlb__EVAL_1 = _EVAL_98;
  assign tlb__EVAL_46 = _EVAL_115;
  assign tag_array__EVAL_0 = {_EVAL_2004,_EVAL_643};
  assign data_arrays_0_0__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign predictor_base_table_0__EVAL = _EVAL_3069 | _EVAL_3190;
  assign tag_array__EVAL_14 = {_EVAL_2004,_EVAL_643};
  assign predictor_tagged_tables_3__EVAL_29 = _EVAL_1253[7];
  assign tag_array__EVAL_3 = {_EVAL_2004,_EVAL_643};
  assign MaxPeriodFibonacciLFSR__EVAL_13 = _EVAL_44;
  assign predictor_tagged_tables_0__EVAL_24 = _EVAL_3397[1];
  assign _EVAL_120 = _EVAL_2534;
  assign tlb__EVAL_53 = _EVAL_3;
  assign predictor_base_table_1__EVAL_18 = _EVAL_668 & _EVAL_2669;
  assign predictor_tagged_tables_0__EVAL_9 = _EVAL_470 | _EVAL_3156;
  assign predictor_tagged_tables_0__EVAL_11 = _EVAL_865 & _EVAL_651;
  assign packageanon1_2__EVAL = _EVAL_1771 & _EVAL_1351;
  assign predictor_tagged_tables_3__EVAL_33 = _EVAL_1980[3];
  assign tlb__EVAL_23 = _EVAL_78;
  assign data_arrays_0_0__EVAL_3 = icache_clock_gate_out;
  assign data_arrays_3_1__EVAL_3 = icache_clock_gate_out;
  assign predictor_Queue__EVAL_2 = _EVAL_361;
  assign predictor_base_table_1__EVAL_14 = predictor_Queue__EVAL_9;
  assign predictor_tagged_tables_1__EVAL_9 = _EVAL_1477 | _EVAL_337;
  assign predictor_base_table_1__EVAL_21 = _EVAL_2226 & _EVAL_2669;
  assign tlb__EVAL_32 = _EVAL_52;
  assign tlb__EVAL_31 = _EVAL_100;
  assign predictor_tagged_tables_3__EVAL_4 = _EVAL_228;
  assign predictor_tagged_tables_0__EVAL_16 = _EVAL_3397[0];
  assign tag_array__EVAL_9 = _EVAL_2918 == 2'h1;
  assign tlb__EVAL_5 = _EVAL_73;
  assign tlb__EVAL_45 = _EVAL_57;
  assign predictor_tagged_tables_1__EVAL_1 = _EVAL_2844[2];
  assign data_arrays_3_1__EVAL = _EVAL_3392 | _EVAL_1447;
  assign _EVAL_49 = _EVAL_3224;
  assign tlb__EVAL_36 = _EVAL_35;
  assign data_arrays_3_0__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign predictor_tagged_tables_2__EVAL_29 = _EVAL_2362[7];
  assign _EVAL_86 = _EVAL_483;
  assign predictor_tagged_tables_2__EVAL_26 = _EVAL_2362[3];
  assign tlb__EVAL_12 = _EVAL_71;
  assign tlb__EVAL_7 = _EVAL_114;
  assign predictor_base_table_0__EVAL_29 = predictor_Queue__EVAL_9;
  assign predictor_base_table_1__EVAL_20 = _EVAL_2401 & _EVAL_2669;
  assign tlb__EVAL_3 = _EVAL_23;
  assign predictor_tagged_tables_0__EVAL_30 = _EVAL_379[6];
  assign data_arrays_1_1__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign predictor_tagged_tables_3__EVAL_37 = _EVAL_1253[11];
  assign data_arrays_2_0__EVAL_4 = {_EVAL_3252,_EVAL_1992};
  assign _EVAL_1 = _EVAL_2611;
  assign predictor_tagged_tables_2__EVAL_21 = _EVAL_2362[10];
  assign tlb__EVAL_25 = _EVAL_128;
  assign predictor_tagged_tables_1__EVAL_20 = _EVAL_1792[8];
  assign predictor_tagged_tables_1__EVAL_22 = _EVAL_2844[9];
  assign predictor_tagged_tables_1__EVAL_6 = _EVAL_1792[5];
  assign data_arrays_3_0__EVAL_1 = _EVAL_1745[8:1];
  assign _EVAL_75 = _EVAL_561;
  assign tlb__EVAL_26 = _EVAL_37;
  assign _EVAL_102 = _EVAL_2222;
  assign predictor_tagged_tables_3__EVAL_15 = _EVAL_1789 ? _EVAL_2522 : _EVAL_1699;
  assign predictor_tagged_tables_3__EVAL_28 = _EVAL_1253[8];
  assign data_arrays_1_1__EVAL_3 = icache_clock_gate_out;
  assign predictor_base_table_0__EVAL_3 = _EVAL_3328 & _EVAL_2669;
  assign predictor_base_table_0__EVAL_16 = _EVAL_2819 & _EVAL_2669;
  assign predictor_base_table_0__EVAL_26 = predictor_Queue__EVAL_9;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_215[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_319[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_363[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_386[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_394[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_403[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_489[initvar] = _RAND_6[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_530[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_548[initvar] = _RAND_8[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_658[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_719[initvar] = _RAND_10[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_725[initvar] = _RAND_11[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_744[initvar] = _RAND_12[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_931[initvar] = _RAND_13[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_949[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_961[initvar] = _RAND_15[8:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_982[initvar] = _RAND_16[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1119[initvar] = _RAND_17[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_1140[initvar] = _RAND_18[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1147[initvar] = _RAND_19[8:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_1440[initvar] = _RAND_20[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1465[initvar] = _RAND_21[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1481[initvar] = _RAND_22[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_23 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_1518[initvar] = _RAND_23[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1652[initvar] = _RAND_24[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1716[initvar] = _RAND_25[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_26 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    _EVAL_1767[initvar] = _RAND_26[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_27 = {1{`RANDOM}};
  _RAND_28 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _EVAL_1859[initvar] = _RAND_28[39:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_1895[initvar] = _RAND_29[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_1986[initvar] = _RAND_30[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_31 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_2023[initvar] = _RAND_31[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2073[initvar] = _RAND_32[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2081[initvar] = _RAND_33[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_34 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2177[initvar] = _RAND_34[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_35 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_2229[initvar] = _RAND_35[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_2337[initvar] = _RAND_36[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_2478[initvar] = _RAND_37[14:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_38 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_2542[initvar] = _RAND_38[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_39 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2573[initvar] = _RAND_39[14:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2580[initvar] = _RAND_40[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2591[initvar] = _RAND_41[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_42 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_2712[initvar] = _RAND_42[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_43 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2773[initvar] = _RAND_43[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_44 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_2852[initvar] = _RAND_44[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_3001[initvar] = _RAND_45[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_46 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_3082[initvar] = _RAND_46[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_47 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_3112[initvar] = _RAND_47[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _EVAL_3335[initvar] = _RAND_48[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_155 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_227 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  _EVAL_253 = _RAND_51[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_254 = _RAND_52[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_271 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_287 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_306 = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_314 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_339 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_344 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_352 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_374 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {2{`RANDOM}};
  _EVAL_397 = _RAND_61[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_430 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {2{`RANDOM}};
  _EVAL_446 = _RAND_63[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_454 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_481 = _RAND_65[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  _EVAL_492 = _RAND_66[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_591 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_664 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_700 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {2{`RANDOM}};
  _EVAL_722 = _RAND_70[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_731 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {2{`RANDOM}};
  _EVAL_794 = _RAND_72[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {4{`RANDOM}};
  _EVAL_837 = _RAND_73[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_839 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_849 = _RAND_75[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  _EVAL_856 = _RAND_76[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_865 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_900 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_927 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_928 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_947 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_954 = _RAND_82[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_957 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_959 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_972 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_975 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1004 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1023 = _RAND_88[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1031 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1085 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1102 = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1128 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {2{`RANDOM}};
  _EVAL_1152 = _RAND_93[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1163 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1165 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {2{`RANDOM}};
  _EVAL_1168 = _RAND_96[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{`RANDOM}};
  _EVAL_1175 = _RAND_97[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1176 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1199 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1243 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1244 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1259 = _RAND_102[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1269 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1272 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1303 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1344 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {2{`RANDOM}};
  _EVAL_1352 = _RAND_107[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1372 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_1386 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1387 = _RAND_110[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1394 = _RAND_111[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1412 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1415 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {2{`RANDOM}};
  _EVAL_1434 = _RAND_114[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {2{`RANDOM}};
  _EVAL_1487 = _RAND_115[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1522 = _RAND_116[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1523 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1529 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {2{`RANDOM}};
  _EVAL_1544 = _RAND_119[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1591 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1649 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1663 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1673 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_1692 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_1706 = _RAND_125[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {4{`RANDOM}};
  _EVAL_1714 = _RAND_126[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_1731 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_1746 = _RAND_128[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_1748 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_1755 = _RAND_130[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_1762 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_1785 = _RAND_132[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_1807 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_1836 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_1846 = _RAND_135[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_1848 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_1886 = _RAND_137[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_1953 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_1954 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_1957 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_1993 = _RAND_141[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {8{`RANDOM}};
  _EVAL_2031 = _RAND_142[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2053 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {2{`RANDOM}};
  _EVAL_2062 = _RAND_144[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {2{`RANDOM}};
  _EVAL_2078 = _RAND_145[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2084 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {2{`RANDOM}};
  _EVAL_2170 = _RAND_147[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _EVAL_2189 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _EVAL_2212 = _RAND_149[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _EVAL_2235 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _EVAL_2248 = _RAND_151[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _EVAL_2252 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {2{`RANDOM}};
  _EVAL_2270 = _RAND_153[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _EVAL_2273 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _EVAL_2274 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _EVAL_2292 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _EVAL_2294 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _EVAL_2304 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _EVAL_2347 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _EVAL_2378 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {2{`RANDOM}};
  _EVAL_2383 = _RAND_161[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _EVAL_2392 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _EVAL_2398 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _EVAL_2399 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _EVAL_2402 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _EVAL_2413 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _EVAL_2447 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _EVAL_2518 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _EVAL_2528 = _RAND_169[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {2{`RANDOM}};
  _EVAL_2534 = _RAND_170[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _EVAL_2549 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _EVAL_2550 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _EVAL_2629 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _EVAL_2640 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {2{`RANDOM}};
  _EVAL_2655 = _RAND_175[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _EVAL_2663 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _EVAL_2686 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _EVAL_2721 = _RAND_178[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {2{`RANDOM}};
  _EVAL_2746 = _RAND_179[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {2{`RANDOM}};
  _EVAL_2785 = _RAND_180[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _EVAL_2799 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _EVAL_2806 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _EVAL_2808 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _EVAL_2880 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _EVAL_2882 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _EVAL_2887 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _EVAL_2888 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _EVAL_2915 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {4{`RANDOM}};
  _EVAL_2928 = _RAND_189[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {4{`RANDOM}};
  _EVAL_2950 = _RAND_190[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {2{`RANDOM}};
  _EVAL_2971 = _RAND_191[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _EVAL_3019 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _EVAL_3050 = _RAND_193[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _EVAL_3054 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _EVAL_3089 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _EVAL_3143 = _RAND_196[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _EVAL_3173 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {2{`RANDOM}};
  _EVAL_3187 = _RAND_198[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {2{`RANDOM}};
  _EVAL_3198 = _RAND_199[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _EVAL_3220 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _EVAL_3225 = _RAND_201[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _EVAL_3261 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _EVAL_3284 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _EVAL_3292 = _RAND_204[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _EVAL_3338 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _EVAL_3340 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _EVAL_3370 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _EVAL_3376 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _EVAL_3394 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _EVAL_3402 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _EVAL_3406 = _RAND_211[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_255) begin
    if(_EVAL_215__EVAL_217_en & _EVAL_215__EVAL_217_mask) begin
      _EVAL_215[_EVAL_215__EVAL_217_addr] <= _EVAL_215__EVAL_217_data;
    end
    if(_EVAL_363__EVAL_365_en & _EVAL_363__EVAL_365_mask) begin
      _EVAL_363[_EVAL_363__EVAL_365_addr] <= _EVAL_363__EVAL_365_data;
    end
    if(_EVAL_386__EVAL_388_en & _EVAL_386__EVAL_388_mask) begin
      _EVAL_386[_EVAL_386__EVAL_388_addr] <= _EVAL_386__EVAL_388_data;
    end
    if(_EVAL_489__EVAL_491_en & _EVAL_489__EVAL_491_mask) begin
      _EVAL_489[_EVAL_489__EVAL_491_addr] <= _EVAL_489__EVAL_491_data;
    end
    if(_EVAL_548__EVAL_550_en & _EVAL_548__EVAL_550_mask) begin
      _EVAL_548[_EVAL_548__EVAL_550_addr] <= _EVAL_548__EVAL_550_data;
    end
    if(_EVAL_719__EVAL_721_en & _EVAL_719__EVAL_721_mask) begin
      _EVAL_719[_EVAL_719__EVAL_721_addr] <= _EVAL_719__EVAL_721_data;
    end
    if(_EVAL_744__EVAL_746_en & _EVAL_744__EVAL_746_mask) begin
      _EVAL_744[_EVAL_744__EVAL_746_addr] <= _EVAL_744__EVAL_746_data;
    end
    if(_EVAL_931__EVAL_933_en & _EVAL_931__EVAL_933_mask) begin
      _EVAL_931[_EVAL_931__EVAL_933_addr] <= _EVAL_931__EVAL_933_data;
    end
    if(_EVAL_961__EVAL_963_en & _EVAL_961__EVAL_963_mask) begin
      _EVAL_961[_EVAL_961__EVAL_963_addr] <= _EVAL_961__EVAL_963_data;
    end
    if(_EVAL_1140__EVAL_1142_en & _EVAL_1140__EVAL_1142_mask) begin
      _EVAL_1140[_EVAL_1140__EVAL_1142_addr] <= _EVAL_1140__EVAL_1142_data;
    end
    if(_EVAL_1440__EVAL_1442_en & _EVAL_1440__EVAL_1442_mask) begin
      _EVAL_1440[_EVAL_1440__EVAL_1442_addr] <= _EVAL_1440__EVAL_1442_data;
    end
    if(_EVAL_1518__EVAL_1520_en & _EVAL_1518__EVAL_1520_mask) begin
      _EVAL_1518[_EVAL_1518__EVAL_1520_addr] <= _EVAL_1518__EVAL_1520_data;
    end
    if(_EVAL_1986__EVAL_1988_en & _EVAL_1986__EVAL_1988_mask) begin
      _EVAL_1986[_EVAL_1986__EVAL_1988_addr] <= _EVAL_1986__EVAL_1988_data;
    end
    if(_EVAL_2073__EVAL_2075_en & _EVAL_2073__EVAL_2075_mask) begin
      _EVAL_2073[_EVAL_2073__EVAL_2075_addr] <= _EVAL_2073__EVAL_2075_data;
    end
    if(_EVAL_2081__EVAL_2083_en & _EVAL_2081__EVAL_2083_mask) begin
      _EVAL_2081[_EVAL_2081__EVAL_2083_addr] <= _EVAL_2081__EVAL_2083_data;
    end
    if(_EVAL_2177__EVAL_2179_en & _EVAL_2177__EVAL_2179_mask) begin
      _EVAL_2177[_EVAL_2177__EVAL_2179_addr] <= _EVAL_2177__EVAL_2179_data;
    end
    if(_EVAL_2573__EVAL_2575_en & _EVAL_2573__EVAL_2575_mask) begin
      _EVAL_2573[_EVAL_2573__EVAL_2575_addr] <= _EVAL_2573__EVAL_2575_data;
    end
    if(_EVAL_2580__EVAL_2582_en & _EVAL_2580__EVAL_2582_mask) begin
      _EVAL_2580[_EVAL_2580__EVAL_2582_addr] <= _EVAL_2580__EVAL_2582_data;
    end
    if(_EVAL_2591__EVAL_2593_en & _EVAL_2591__EVAL_2593_mask) begin
      _EVAL_2591[_EVAL_2591__EVAL_2593_addr] <= _EVAL_2591__EVAL_2593_data;
    end
    if(_EVAL_2773__EVAL_2775_en & _EVAL_2773__EVAL_2775_mask) begin
      _EVAL_2773[_EVAL_2773__EVAL_2775_addr] <= _EVAL_2773__EVAL_2775_data;
    end
    if(_EVAL_2852__EVAL_2854_en & _EVAL_2852__EVAL_2854_mask) begin
      _EVAL_2852[_EVAL_2852__EVAL_2854_addr] <= _EVAL_2852__EVAL_2854_data;
    end
    if(_EVAL_3112__EVAL_3114_en & _EVAL_3112__EVAL_3114_mask) begin
      _EVAL_3112[_EVAL_3112__EVAL_3114_addr] <= _EVAL_3112__EVAL_3114_data;
    end
    if(_EVAL_3335__EVAL_3337_en & _EVAL_3335__EVAL_3337_mask) begin
      _EVAL_3335[_EVAL_3335__EVAL_3337_addr] <= _EVAL_3335__EVAL_3337_data;
    end
    if (_EVAL_3170) begin
      _EVAL_254 <= 2'h0;
    end else begin
      if (_EVAL_2390) begin
        _EVAL_254 <= _EVAL_2501;
      end
    end
    if (_EVAL_3170) begin
      _EVAL_2248 <= 2'h0;
    end else begin
      if (_EVAL_1222) begin
        _EVAL_2248 <= _EVAL_1696;
      end
    end
    if (_EVAL_3170) begin
      _EVAL_3054 <= 1'h0;
    end else begin
      if (_EVAL_3194) begin
        _EVAL_3054 <= _EVAL_2390;
      end
    end
  end
  always @(posedge _EVAL_973) begin
    if(_EVAL_319__EVAL_321_en & _EVAL_319__EVAL_321_mask) begin
      _EVAL_319[_EVAL_319__EVAL_321_addr] <= _EVAL_319__EVAL_321_data;
    end
    if(_EVAL_394__EVAL_396_en & _EVAL_394__EVAL_396_mask) begin
      _EVAL_394[_EVAL_394__EVAL_396_addr] <= _EVAL_394__EVAL_396_data;
    end
    if(_EVAL_403__EVAL_405_en & _EVAL_403__EVAL_405_mask) begin
      _EVAL_403[_EVAL_403__EVAL_405_addr] <= _EVAL_403__EVAL_405_data;
    end
    if(_EVAL_530__EVAL_532_en & _EVAL_530__EVAL_532_mask) begin
      _EVAL_530[_EVAL_530__EVAL_532_addr] <= _EVAL_530__EVAL_532_data;
    end
    if(_EVAL_658__EVAL_660_en & _EVAL_658__EVAL_660_mask) begin
      _EVAL_658[_EVAL_658__EVAL_660_addr] <= _EVAL_658__EVAL_660_data;
    end
    if(_EVAL_725__EVAL_727_en & _EVAL_725__EVAL_727_mask) begin
      _EVAL_725[_EVAL_725__EVAL_727_addr] <= _EVAL_725__EVAL_727_data;
    end
    if(_EVAL_949__EVAL_951_en & _EVAL_949__EVAL_951_mask) begin
      _EVAL_949[_EVAL_949__EVAL_951_addr] <= _EVAL_949__EVAL_951_data;
    end
    if(_EVAL_982__EVAL_984_en & _EVAL_982__EVAL_984_mask) begin
      _EVAL_982[_EVAL_982__EVAL_984_addr] <= _EVAL_982__EVAL_984_data;
    end
    if(_EVAL_1119__EVAL_1121_en & _EVAL_1119__EVAL_1121_mask) begin
      _EVAL_1119[_EVAL_1119__EVAL_1121_addr] <= _EVAL_1119__EVAL_1121_data;
    end
    if(_EVAL_1147__EVAL_1149_en & _EVAL_1147__EVAL_1149_mask) begin
      _EVAL_1147[_EVAL_1147__EVAL_1149_addr] <= _EVAL_1147__EVAL_1149_data;
    end
    if(_EVAL_1465__EVAL_1467_en & _EVAL_1465__EVAL_1467_mask) begin
      _EVAL_1465[_EVAL_1465__EVAL_1467_addr] <= _EVAL_1465__EVAL_1467_data;
    end
    if(_EVAL_1481__EVAL_1483_en & _EVAL_1481__EVAL_1483_mask) begin
      _EVAL_1481[_EVAL_1481__EVAL_1483_addr] <= _EVAL_1481__EVAL_1483_data;
    end
    if(_EVAL_1652__EVAL_1654_en & _EVAL_1652__EVAL_1654_mask) begin
      _EVAL_1652[_EVAL_1652__EVAL_1654_addr] <= _EVAL_1652__EVAL_1654_data;
    end
    if(_EVAL_1716__EVAL_1718_en & _EVAL_1716__EVAL_1718_mask) begin
      _EVAL_1716[_EVAL_1716__EVAL_1718_addr] <= _EVAL_1716__EVAL_1718_data;
    end
    if(_EVAL_1895__EVAL_1897_en & _EVAL_1895__EVAL_1897_mask) begin
      _EVAL_1895[_EVAL_1895__EVAL_1897_addr] <= _EVAL_1895__EVAL_1897_data;
    end
    if(_EVAL_2023__EVAL_2025_en & _EVAL_2023__EVAL_2025_mask) begin
      _EVAL_2023[_EVAL_2023__EVAL_2025_addr] <= _EVAL_2023__EVAL_2025_data;
    end
    if(_EVAL_2229__EVAL_2231_en & _EVAL_2229__EVAL_2231_mask) begin
      _EVAL_2229[_EVAL_2229__EVAL_2231_addr] <= _EVAL_2229__EVAL_2231_data;
    end
    if(_EVAL_2337__EVAL_2339_en & _EVAL_2337__EVAL_2339_mask) begin
      _EVAL_2337[_EVAL_2337__EVAL_2339_addr] <= _EVAL_2337__EVAL_2339_data;
    end
    if(_EVAL_2478__EVAL_2480_en & _EVAL_2478__EVAL_2480_mask) begin
      _EVAL_2478[_EVAL_2478__EVAL_2480_addr] <= _EVAL_2478__EVAL_2480_data;
    end
    if(_EVAL_2542__EVAL_2544_en & _EVAL_2542__EVAL_2544_mask) begin
      _EVAL_2542[_EVAL_2542__EVAL_2544_addr] <= _EVAL_2542__EVAL_2544_data;
    end
    if(_EVAL_2712__EVAL_2714_en & _EVAL_2712__EVAL_2714_mask) begin
      _EVAL_2712[_EVAL_2712__EVAL_2714_addr] <= _EVAL_2712__EVAL_2714_data;
    end
    if(_EVAL_3001__EVAL_3003_en & _EVAL_3001__EVAL_3003_mask) begin
      _EVAL_3001[_EVAL_3001__EVAL_3003_addr] <= _EVAL_3001__EVAL_3003_data;
    end
    if(_EVAL_3082__EVAL_3084_en & _EVAL_3082__EVAL_3084_mask) begin
      _EVAL_3082[_EVAL_3082__EVAL_3084_addr] <= _EVAL_3082__EVAL_3084_data;
    end
    if (_EVAL_1261) begin
      _EVAL_972 <= 1'h0;
    end else begin
      if (_EVAL_1842) begin
        _EVAL_972 <= _EVAL_3229;
      end
    end
  end
  always @(posedge icache_clock_gate_out) begin
    if(_EVAL_1767__EVAL_1769_en & _EVAL_1767__EVAL_1769_mask) begin
      _EVAL_1767[_EVAL_1767__EVAL_1769_addr] <= _EVAL_1767__EVAL_1769_data;
    end
    if(_EVAL_1859__EVAL_1862_en & _EVAL_1859__EVAL_1862_mask) begin
      _EVAL_1859[_EVAL_1859__EVAL_1862_addr] <= _EVAL_1859__EVAL_1862_data;
    end
    if (_EVAL_1077) begin
      _EVAL_155 <= _EVAL_3305;
    end
    if (_EVAL_2783) begin
      if (_EVAL_1326) begin
        _EVAL_253 <= _EVAL_2377;
      end
    end
    if (_EVAL_44) begin
      _EVAL_271 <= 1'h0;
    end else begin
      if (_EVAL_2010) begin
        _EVAL_271 <= 1'h0;
      end else begin
        if (_EVAL_3052) begin
          _EVAL_271 <= 1'h1;
        end
      end
    end
    _EVAL_287 <= _EVAL_2509[0];
    if (_EVAL_1724) begin
      _EVAL_306 <= _EVAL_32;
    end
    if (_EVAL_1724) begin
      _EVAL_314 <= _EVAL_85;
    end
    if (_EVAL_273) begin
      if (_EVAL_1577) begin
        if (_EVAL_1949) begin
          _EVAL_344 <= 1'h0;
        end else begin
          _EVAL_344 <= _EVAL_2700;
        end
      end else begin
        _EVAL_344 <= _EVAL_2700;
      end
    end else begin
      _EVAL_344 <= _EVAL_2700;
    end
    if (_EVAL_2783) begin
      if (_EVAL_798) begin
        _EVAL_397 <= _EVAL_2377;
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_2901) begin
        _EVAL_446 <= _EVAL_2377;
      end
    end
    if (_EVAL_77) begin
      if (_EVAL_257) begin
        _EVAL_454 <= _EVAL_154;
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_642) begin
        _EVAL_492 <= _EVAL_2377;
      end
    end
    if (_EVAL_2153) begin
      _EVAL_591 <= 1'h0;
    end else begin
      if (_EVAL_131) begin
        _EVAL_591 <= 1'h1;
      end
    end
    if (_EVAL_344) begin
      _EVAL_664 <= _EVAL_1811;
    end
    if (_EVAL_2783) begin
      if (_EVAL_2682) begin
        _EVAL_722 <= _EVAL_2377;
      end
    end
    if (_EVAL_344) begin
      _EVAL_731 <= _EVAL_2905;
    end
    if (_EVAL_2783) begin
      if (_EVAL_2475) begin
        _EVAL_794 <= _EVAL_2377;
      end
    end
    if (_EVAL_160) begin
      if (_EVAL_286) begin
        _EVAL_837 <= _EVAL_167;
      end else begin
        _EVAL_837 <= _EVAL_2225;
      end
    end
    _EVAL_839 <= _EVAL_3383 & _EVAL_1088;
    if (_EVAL_2640) begin
      _EVAL_849 <= tag_array__EVAL_2;
    end
    if (_EVAL_2783) begin
      if (_EVAL_2863) begin
        _EVAL_856 <= _EVAL_2377;
      end
    end
    _EVAL_927 <= _EVAL_1540[2];
    _EVAL_947 <= _EVAL_1692;
    if (_EVAL_273) begin
      _EVAL_957 <= tlb__EVAL_39;
    end
    _EVAL_959 <= _EVAL_1540[0];
    _EVAL_1004 <= _EVAL_1900 & _EVAL_1737;
    if (_EVAL_2640) begin
      _EVAL_1023 <= tag_array__EVAL_11;
    end
    _EVAL_1085 <= _EVAL_1900 & _EVAL_354;
    if (_EVAL_113) begin
      if (_EVAL_2847) begin
        _EVAL_1102 <= _EVAL_12;
      end else begin
        if (_EVAL_1077) begin
          if (_EVAL_971) begin
            _EVAL_1102 <= _EVAL_301;
          end else begin
            if (_EVAL_2720) begin
              _EVAL_1102 <= _EVAL_426;
            end
          end
        end
      end
    end else begin
      if (_EVAL_1077) begin
        if (_EVAL_971) begin
          _EVAL_1102 <= _EVAL_301;
        end else begin
          if (_EVAL_2720) begin
            _EVAL_1102 <= _EVAL_426;
          end
        end
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_681) begin
        _EVAL_1152 <= _EVAL_2377;
      end
    end
    if (_EVAL_273) begin
      if (_EVAL_2820) begin
        _EVAL_1163 <= _EVAL_3403;
      end else begin
        _EVAL_1163 <= _EVAL_1767__EVAL_1768_data;
      end
    end
    if (_EVAL_1900) begin
      _EVAL_1168 <= data_arrays_1_0__EVAL_0;
    end
    if (_EVAL_2783) begin
      if (_EVAL_1801) begin
        _EVAL_1175 <= _EVAL_2377;
      end
    end
    if (_EVAL_1077) begin
      _EVAL_1176 <= _EVAL_1995;
    end
    if (_EVAL_1077) begin
      _EVAL_1199 <= _EVAL_3367;
    end
    if (_EVAL_273) begin
      _EVAL_1243 <= _EVAL_1040;
    end
    _EVAL_1269 <= _EVAL_1850 == 1'h0;
    if (_EVAL_344) begin
      _EVAL_1272 <= _EVAL_1088;
    end
    _EVAL_1344 <= _EVAL_1900 & _EVAL_1088;
    if (_EVAL_2783) begin
      if (_EVAL_825) begin
        _EVAL_1352 <= _EVAL_2377;
      end
    end
    _EVAL_1387 <= _EVAL_2562[6:0];
    _EVAL_1412 <= _EVAL_1540[1];
    if (_EVAL_3383) begin
      _EVAL_1434 <= data_arrays_1_1__EVAL_0;
    end
    if (_EVAL_2783) begin
      if (_EVAL_1338) begin
        _EVAL_1487 <= _EVAL_2377;
      end
    end
    if (_EVAL_1724) begin
      _EVAL_1522 <= _EVAL_137;
    end
    if (_EVAL_344) begin
      _EVAL_1523 <= _EVAL_1737;
    end
    if (_EVAL_44) begin
      _EVAL_1529 <= 1'h0;
    end else begin
      if (_EVAL_1852) begin
        _EVAL_1529 <= 1'h0;
      end else begin
        if (_EVAL_273) begin
          if (_EVAL_1577) begin
            _EVAL_1529 <= _EVAL_344;
          end else begin
            _EVAL_1529 <= 1'h0;
          end
        end else begin
          _EVAL_1529 <= 1'h0;
        end
      end
    end
    if (_EVAL_1900) begin
      _EVAL_1544 <= data_arrays_0_0__EVAL_0;
    end
    if (_EVAL_44) begin
      _EVAL_1591 <= 1'h0;
    end else begin
      if (_EVAL_273) begin
        _EVAL_1591 <= _EVAL_1649;
      end
    end
    if (_EVAL_113) begin
      _EVAL_1649 <= _EVAL_45;
    end else begin
      if (!(_EVAL_2663)) begin
        _EVAL_1649 <= 1'h1;
      end
    end
    if (_EVAL_44) begin
      _EVAL_1692 <= 1'h0;
    end else begin
      _EVAL_1692 <= _EVAL_1724;
    end
    if (_EVAL_1077) begin
      _EVAL_1706 <= _EVAL_2548;
    end
    if (_EVAL_113) begin
      if (_EVAL_448) begin
        _EVAL_1714 <= {{121'd0}, _EVAL_2026};
      end else begin
        _EVAL_1714 <= _EVAL_82;
      end
    end else begin
      _EVAL_1714 <= {{121'd0}, _EVAL_415};
    end
    if (_EVAL_273) begin
      _EVAL_1731 <= tlb__EVAL_10;
    end
    _EVAL_1762 <= _EVAL_104;
    if (_EVAL_2640) begin
      _EVAL_1785 <= tag_array__EVAL_7;
    end
    _EVAL_1807 <= _EVAL_3383 & _EVAL_1811;
    _EVAL_1846 <= _EVAL_1112[24:0];
    _EVAL_1953 <= _EVAL_947 | _EVAL_2684;
    if (_EVAL_1077) begin
      _EVAL_1957 <= _EVAL_1908;
    end
    if (_EVAL_44) begin
      _EVAL_2031 <= 256'h0;
    end else begin
      if (_EVAL_131) begin
        _EVAL_2031 <= 256'h0;
      end else begin
        if (_EVAL_10) begin
          if (_EVAL_2976) begin
            _EVAL_2031 <= _EVAL_285;
          end else begin
            _EVAL_2031 <= _EVAL_734;
          end
        end
      end
    end
    if (_EVAL_113) begin
      _EVAL_2053 <= 1'h0;
    end else begin
      if (_EVAL_3296) begin
        _EVAL_2053 <= 1'h0;
      end else begin
        if (_EVAL_2843) begin
          _EVAL_2053 <= 1'h0;
        end else begin
          _EVAL_2053 <= _EVAL_1010;
        end
      end
    end
    if (_EVAL_1900) begin
      _EVAL_2062 <= data_arrays_2_0__EVAL_0;
    end
    if (_EVAL_1900) begin
      _EVAL_2078 <= data_arrays_3_0__EVAL_0;
    end
    if (_EVAL_113) begin
      _EVAL_2084 <= 1'h0;
    end else begin
      if (_EVAL_3296) begin
        _EVAL_2084 <= 1'h0;
      end else begin
        if (_EVAL_2843) begin
          _EVAL_2084 <= _EVAL_3173;
        end else begin
          _EVAL_2084 <= _EVAL_2063;
        end
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_1578) begin
        _EVAL_2170 <= _EVAL_2377;
      end
    end
    if (_EVAL_44) begin
      _EVAL_2252 <= 1'h0;
    end else begin
      if (_EVAL_273) begin
        _EVAL_2252 <= _EVAL_1577;
      end else begin
        _EVAL_2252 <= 1'h0;
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_3045) begin
        _EVAL_2270 <= _EVAL_2377;
      end
    end
    if (_EVAL_1077) begin
      _EVAL_2273 <= _EVAL_2392;
    end
    _EVAL_2292 <= _EVAL_1077 & _EVAL_2435;
    if (_EVAL_10) begin
      _EVAL_2378 <= 1'h0;
    end else begin
      if (_EVAL_2700) begin
        _EVAL_2378 <= 1'h1;
      end else begin
        if (_EVAL_1235) begin
          _EVAL_2378 <= 1'h0;
        end
      end
    end
    if (_EVAL_3383) begin
      _EVAL_2383 <= data_arrays_2_1__EVAL_0;
    end
    if (_EVAL_44) begin
      _EVAL_2392 <= _EVAL_1061;
    end else begin
      if (_EVAL_273) begin
        _EVAL_2392 <= _EVAL_2402;
      end
    end
    if (_EVAL_344) begin
      _EVAL_2399 <= _EVAL_354;
    end
    _EVAL_2402 <= ~ _EVAL_544;
    if (_EVAL_44) begin
      _EVAL_2518 <= 1'h0;
    end else begin
      if (_EVAL_113) begin
        _EVAL_2518 <= 1'h0;
      end else begin
        if (_EVAL_1077) begin
          if (_EVAL_1242) begin
            _EVAL_2518 <= 1'h0;
          end else begin
            if (_EVAL_1995) begin
              _EVAL_2518 <= 1'h0;
            end else begin
              _EVAL_2518 <= _EVAL_832;
            end
          end
        end
      end
    end
    _EVAL_2528 <= _EVAL_1638[1:0];
    if (_EVAL_947) begin
      _EVAL_2534 <= _EVAL_964;
    end else begin
      if (_EVAL_1724) begin
        _EVAL_2534 <= _EVAL_63;
      end
    end
    if (_EVAL_1574) begin
      _EVAL_2549 <= _EVAL_1942;
    end
    if (_EVAL_44) begin
      _EVAL_2550 <= 1'h1;
    end else begin
      if (_EVAL_3246) begin
        _EVAL_2550 <= 1'h0;
      end else begin
        if (_EVAL_3101) begin
          _EVAL_2550 <= 1'h1;
        end else begin
          if (_EVAL_2153) begin
            _EVAL_2550 <= 1'h0;
          end
        end
      end
    end
    _EVAL_2640 <= _EVAL_2700 & _EVAL_1235;
    if (_EVAL_3383) begin
      _EVAL_2655 <= data_arrays_3_1__EVAL_0;
    end
    _EVAL_2663 <= _EVAL_113;
    if (_EVAL_1077) begin
      if (_EVAL_2139) begin
        if (_EVAL_474) begin
          _EVAL_2686 <= _EVAL_2257;
        end else begin
          if (_EVAL_2671) begin
            if (_EVAL_919) begin
              _EVAL_2686 <= _EVAL_462;
            end else begin
              _EVAL_2686 <= _EVAL_650;
            end
          end else begin
            if (_EVAL_272) begin
              _EVAL_2686 <= _EVAL_1163;
            end else begin
              _EVAL_2686 <= _EVAL_1243;
            end
          end
        end
      end else begin
        if (_EVAL_1111) begin
          if (_EVAL_1413) begin
            _EVAL_2686 <= _EVAL_391;
          end else begin
            if (_EVAL_955) begin
              if (_EVAL_1029) begin
                _EVAL_2686 <= _EVAL_650;
              end else begin
                _EVAL_2686 <= _EVAL_1205;
              end
            end else begin
              if (_EVAL_2236) begin
                _EVAL_2686 <= _EVAL_1163;
              end else begin
                _EVAL_2686 <= _EVAL_1243;
              end
            end
          end
        end else begin
          if (_EVAL_1257) begin
            if (_EVAL_2623) begin
              _EVAL_2686 <= _EVAL_2490;
            end else begin
              if (_EVAL_431) begin
                if (_EVAL_2938) begin
                  _EVAL_2686 <= _EVAL_1205;
                end else begin
                  _EVAL_2686 <= _EVAL_2232;
                end
              end else begin
                if (_EVAL_3410) begin
                  _EVAL_2686 <= _EVAL_1163;
                end else begin
                  _EVAL_2686 <= _EVAL_1243;
                end
              end
            end
          end else begin
            if (_EVAL_2309) begin
              if (_EVAL_1315) begin
                _EVAL_2686 <= _EVAL_2079;
              end else begin
                if (_EVAL_3209) begin
                  if (_EVAL_2866) begin
                    _EVAL_2686 <= _EVAL_2232;
                  end else begin
                    _EVAL_2686 <= _EVAL_2175;
                  end
                end else begin
                  if (_EVAL_1644) begin
                    _EVAL_2686 <= _EVAL_1163;
                  end else begin
                    _EVAL_2686 <= _EVAL_1243;
                  end
                end
              end
            end else begin
              if (_EVAL_3221) begin
                _EVAL_2686 <= _EVAL_2605;
              end else begin
                if (_EVAL_381) begin
                  _EVAL_2686 <= _EVAL_2175;
                end else begin
                  if (_EVAL_1596) begin
                    _EVAL_2686 <= _EVAL_1163;
                  end else begin
                    _EVAL_2686 <= _EVAL_1243;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_1761) begin
        _EVAL_2746 <= _EVAL_2377;
      end
    end
    if (_EVAL_1919) begin
      _EVAL_2785 <= _EVAL_539;
    end
    _EVAL_2799 <= _EVAL_3383 & _EVAL_1737;
    if (_EVAL_1077) begin
      _EVAL_2806 <= _EVAL_2445;
    end
    if (_EVAL_10) begin
      _EVAL_2808 <= _EVAL_2004;
    end
    _EVAL_2888 <= _EVAL_3383 & _EVAL_354;
    if (_EVAL_344) begin
      _EVAL_2915 <= _EVAL_291;
    end
    if (_EVAL_3383) begin
      _EVAL_2971 <= data_arrays_0_1__EVAL_0;
    end
    _EVAL_3050 <= _EVAL_1156[6:0];
    _EVAL_3143 <= _EVAL_29;
    if (_EVAL_273) begin
      _EVAL_3173 <= _EVAL_2084;
    end
    if (_EVAL_2783) begin
      if (_EVAL_2987) begin
        _EVAL_3187 <= _EVAL_2377;
      end
    end
    if (_EVAL_2783) begin
      if (_EVAL_918) begin
        _EVAL_3198 <= _EVAL_2377;
      end
    end
    _EVAL_3220 <= _EVAL_1900 & _EVAL_1811;
    if (_EVAL_2640) begin
      _EVAL_3225 <= tag_array__EVAL_1;
    end
    if (_EVAL_1724) begin
      _EVAL_3292 <= _EVAL_15;
    end
    if (_EVAL_273) begin
      _EVAL_3340 <= _EVAL_287;
    end
    if (_EVAL_44) begin
      _EVAL_3370 <= 1'h1;
    end else begin
      _EVAL_3370 <= _EVAL_1212;
    end
    if (_EVAL_1077) begin
      if (_EVAL_832) begin
        _EVAL_3376 <= _EVAL_1968;
      end
    end
    if (_EVAL_273) begin
      _EVAL_3394 <= _EVAL_3103;
    end
    if (_EVAL_77) begin
      if (_EVAL_257) begin
        _EVAL_3406 <= _EVAL_262;
      end else begin
        if (_EVAL_2696) begin
          _EVAL_3406 <= _EVAL_3350;
        end
      end
    end
  end
  always @(posedge _EVAL_228) begin
    if (_EVAL_361) begin
      _EVAL_227 <= _EVAL_685;
    end
    if (_EVAL_2102) begin
      _EVAL_339 <= 1'h0;
    end else begin
      _EVAL_339 <= _EVAL_1408;
    end
    if (_EVAL_339) begin
      _EVAL_352 <= _EVAL_637;
    end
    _EVAL_374 <= _EVAL_338 & _EVAL_3327;
    if (_EVAL_339) begin
      _EVAL_430 <= _EVAL_1660;
    end
    if (_EVAL_361) begin
      _EVAL_481 <= _EVAL_2818;
    end
    if (_EVAL_339) begin
      _EVAL_700 <= _EVAL_2862;
    end
    _EVAL_865 <= _EVAL_361;
    if (_EVAL_361) begin
      _EVAL_900 <= _EVAL_793;
    end
    if (_EVAL_339) begin
      _EVAL_928 <= _EVAL_186;
    end
    if (_EVAL_3327) begin
      _EVAL_954 <= _EVAL_1293;
    end
    _EVAL_975 <= _EVAL_2019 & _EVAL_3327;
    if (_EVAL_339) begin
      _EVAL_1031 <= _EVAL_1248;
    end
    if (_EVAL_3327) begin
      _EVAL_1128 <= _EVAL_2408;
    end
    if (_EVAL_339) begin
      _EVAL_1165 <= _EVAL_290;
    end
    if (_EVAL_339) begin
      _EVAL_1244 <= _EVAL_2214;
    end
    if (_EVAL_339) begin
      _EVAL_1259 <= _EVAL_1486;
    end
    _EVAL_1303 <= _EVAL_411 & _EVAL_3327;
    if (_EVAL_339) begin
      _EVAL_1372 <= _EVAL_704;
    end
    if (_EVAL_339) begin
      _EVAL_1386 <= _EVAL_1392;
    end
    if (_EVAL_339) begin
      _EVAL_1394 <= _EVAL_2032;
    end
    if (_EVAL_339) begin
      _EVAL_1415 <= _EVAL_736;
    end
    if (_EVAL_339) begin
      _EVAL_1663 <= _EVAL_1902;
    end
    if (_EVAL_339) begin
      _EVAL_1673 <= _EVAL_799;
    end
    if (_EVAL_3327) begin
      _EVAL_1746 <= _EVAL_2917;
    end
    if (_EVAL_339) begin
      _EVAL_1748 <= _EVAL_2467;
    end
    if (_EVAL_3327) begin
      _EVAL_1755 <= _EVAL_2564;
    end
    if (_EVAL_361) begin
      _EVAL_1836 <= _EVAL_634;
    end
    _EVAL_1848 <= _EVAL_1132 & _EVAL_3327;
    if (_EVAL_1408) begin
      _EVAL_1886 <= _EVAL_1090;
    end
    if (_EVAL_339) begin
      _EVAL_1954 <= _EVAL_2927;
    end
    if (_EVAL_339) begin
      _EVAL_2189 <= _EVAL_1133;
    end
    if (_EVAL_361) begin
      _EVAL_2212 <= _EVAL_1600;
    end
    if (_EVAL_361) begin
      _EVAL_2235 <= _EVAL_3253;
    end
    if (_EVAL_339) begin
      if (_EVAL_1340) begin
        _EVAL_2274 <= predictor_base_table_1__EVAL_13;
      end else begin
        if (_EVAL_855) begin
          _EVAL_2274 <= predictor_base_table_0__EVAL_13;
        end else begin
          _EVAL_2274 <= 1'h0;
        end
      end
    end
    if (_EVAL_339) begin
      _EVAL_2294 <= _EVAL_3036;
    end
    if (_EVAL_339) begin
      _EVAL_2304 <= _EVAL_1239;
    end
    if (_EVAL_339) begin
      _EVAL_2347 <= _EVAL_421;
    end
    if (_EVAL_339) begin
      _EVAL_2398 <= _EVAL_1814;
    end
    if (_EVAL_361) begin
      _EVAL_2413 <= _EVAL_2089;
    end
    if (_EVAL_361) begin
      _EVAL_2447 <= _EVAL_1892;
    end
    if (_EVAL_339) begin
      _EVAL_2629 <= _EVAL_1410;
    end
    if (_EVAL_339) begin
      _EVAL_2721 <= _EVAL_278;
    end
    if (_EVAL_361) begin
      _EVAL_2880 <= _EVAL_1506;
    end
    if (_EVAL_339) begin
      _EVAL_2882 <= _EVAL_2128;
    end
    if (_EVAL_339) begin
      _EVAL_2887 <= _EVAL_1287;
    end
    if (_EVAL_1408) begin
      _EVAL_2928 <= _EVAL_2531;
    end
    if (_EVAL_361) begin
      _EVAL_2950 <= _EVAL_2873;
    end
    if (_EVAL_339) begin
      _EVAL_3019 <= _EVAL_1637;
    end
    if (_EVAL_339) begin
      if (_EVAL_1340) begin
        if (4'h8 == _EVAL_2324) begin
          _EVAL_3089 <= predictor_base_table_1__EVAL_13;
        end else begin
          if (3'h7 == _EVAL_1279) begin
            _EVAL_3089 <= predictor_base_table_1__EVAL_10;
          end else begin
            if (3'h6 == _EVAL_1279) begin
              _EVAL_3089 <= predictor_base_table_1__EVAL_22;
            end else begin
              if (3'h5 == _EVAL_1279) begin
                _EVAL_3089 <= predictor_base_table_1__EVAL_6;
              end else begin
                if (3'h4 == _EVAL_1279) begin
                  _EVAL_3089 <= predictor_base_table_1__EVAL_0;
                end else begin
                  if (3'h3 == _EVAL_1279) begin
                    _EVAL_3089 <= predictor_base_table_1__EVAL_17;
                  end else begin
                    if (3'h2 == _EVAL_1279) begin
                      _EVAL_3089 <= predictor_base_table_1__EVAL_7;
                    end else begin
                      if (3'h1 == _EVAL_1279) begin
                        _EVAL_3089 <= predictor_base_table_1__EVAL_1;
                      end else begin
                        _EVAL_3089 <= _EVAL_709;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_EVAL_855) begin
          if (4'h8 == _EVAL_2324) begin
            _EVAL_3089 <= predictor_base_table_0__EVAL_13;
          end else begin
            if (3'h7 == _EVAL_1279) begin
              _EVAL_3089 <= predictor_base_table_0__EVAL_10;
            end else begin
              if (3'h6 == _EVAL_1279) begin
                _EVAL_3089 <= predictor_base_table_0__EVAL_22;
              end else begin
                if (3'h5 == _EVAL_1279) begin
                  _EVAL_3089 <= predictor_base_table_0__EVAL_6;
                end else begin
                  if (3'h4 == _EVAL_1279) begin
                    _EVAL_3089 <= predictor_base_table_0__EVAL_0;
                  end else begin
                    if (3'h3 == _EVAL_1279) begin
                      _EVAL_3089 <= predictor_base_table_0__EVAL_17;
                    end else begin
                      if (3'h2 == _EVAL_1279) begin
                        _EVAL_3089 <= predictor_base_table_0__EVAL_7;
                      end else begin
                        if (3'h1 == _EVAL_1279) begin
                          _EVAL_3089 <= predictor_base_table_0__EVAL_1;
                        end else begin
                          _EVAL_3089 <= _EVAL_2210;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          _EVAL_3089 <= 1'h0;
        end
      end
    end
    if (_EVAL_339) begin
      _EVAL_3261 <= _EVAL_1576;
    end
    if (_EVAL_339) begin
      _EVAL_3284 <= _EVAL_1359;
    end
  end
  always @(posedge _EVAL_57) begin
    if (_EVAL_44) begin
      _EVAL_1993 <= 5'h0;
    end else begin
      if (_EVAL_10) begin
        if (_EVAL_1250) begin
          if (_EVAL_2003) begin
            _EVAL_1993 <= _EVAL_1494;
          end else begin
            _EVAL_1993 <= 5'h0;
          end
        end else begin
          _EVAL_1993 <= _EVAL_333;
        end
      end
    end
    if (_EVAL_48) begin
      _EVAL_3338 <= 16'h0;
    end else begin
      if (_EVAL_2783) begin
        _EVAL_3338 <= _EVAL_693;
      end else begin
        if (_EVAL_814) begin
          _EVAL_3338 <= _EVAL_606;
        end
      end
    end
    _EVAL_3402 <= _EVAL_2488 | _EVAL_2494;
  end
endmodule
