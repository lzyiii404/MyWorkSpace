//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_2_assert(
  input         _EVAL_1,
  input  [2:0]  _EVAL_3,
  input         _EVAL_9,
  input  [31:0] _EVAL_13,
  input         _EVAL_15,
  input  [1:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input         _EVAL_36,
  input         _EVAL_38,
  input  [3:0]  _EVAL_40,
  input         _EVAL_42,
  input  [2:0]  _EVAL_45,
  input         _EVAL_51,
  input         _EVAL_54,
  input  [3:0]  _EVAL_56,
  input         _EVAL_60,
  input  [2:0]  _EVAL_61,
  input  [2:0]  _EVAL_62,
  input  [7:0]  _EVAL_67,
  input  [31:0] _EVAL_69,
  input  [3:0]  _EVAL_71,
  input  [3:0]  _EVAL_77,
  input         _EVAL_82,
  input         _EVAL_84,
  input  [2:0]  _EVAL_90,
  input         _EVAL_101,
  input         _EVAL_103,
  input         _EVAL_113,
  input  [31:0] _EVAL_114,
  input  [3:0]  _EVAL_117,
  input  [7:0]  _EVAL_121,
  input         _EVAL_122,
  input  [5:0]  _EVAL_127,
  input         _EVAL_366,
  input  [2:0]  _EVAL_261,
  input  [1:0]  _EVAL_441,
  input         _EVAL_178,
  input  [1:0]  _EVAL_229,
  input         _EVAL_435,
  input         _EVAL_520,
  input         _EVAL_460,
  input         _EVAL_297,
  input  [1:0]  _EVAL_140,
  input         _EVAL_479,
  input         _EVAL_341,
  input         _EVAL_166,
  input         _EVAL_215,
  input         _EVAL_290,
  input         _EVAL_591,
  input         _EVAL_199,
  input         _EVAL_158,
  input         _EVAL_327,
  input         _EVAL_539,
  input  [2:0]  _EVAL_620,
  input         _EVAL_563,
  input         _EVAL_523,
  input         _EVAL_422,
  input  [82:0] _EVAL_396,
  input         _EVAL_187,
  input         _EVAL_139,
  input         _EVAL_311,
  input  [6:0]  _EVAL_235,
  input         _EVAL_569,
  input  [82:0] _EVAL_614,
  input         _EVAL_378,
  input         _EVAL_243,
  input  [6:0]  _EVAL_170
);
  wire [5:0] TLMonitor_1__EVAL;
  wire  TLMonitor_1__EVAL_0;
  wire [2:0] TLMonitor_1__EVAL_1;
  wire [5:0] TLMonitor_1__EVAL_2;
  wire [2:0] TLMonitor_1__EVAL_3;
  wire  TLMonitor_1__EVAL_4;
  wire  TLMonitor_1__EVAL_5;
  wire  TLMonitor_1__EVAL_6;
  wire [3:0] TLMonitor_1__EVAL_7;
  wire  TLMonitor_1__EVAL_8;
  wire  TLMonitor_1__EVAL_9;
  wire  TLMonitor_1__EVAL_10;
  wire  TLMonitor_1__EVAL_11;
  wire  TLMonitor_1__EVAL_12;
  wire [7:0] TLMonitor_1__EVAL_13;
  wire  TLMonitor_1__EVAL_14;
  wire [2:0] TLMonitor_1__EVAL_15;
  wire [1:0] TLMonitor_1__EVAL_16;
  wire [31:0] TLMonitor_1__EVAL_17;
  wire [3:0] TLMonitor_1__EVAL_18;
  wire [3:0] TLMonitor__EVAL;
  wire [31:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire [3:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [2:0] TLMonitor__EVAL_7;
  wire [31:0] TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire [3:0] TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire [1:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [1:0] TLMonitor__EVAL_14;
  wire [3:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire [2:0] TLMonitor__EVAL_17;
  wire  TLMonitor__EVAL_18;
  wire  TLMonitor__EVAL_19;
  wire [7:0] TLMonitor__EVAL_20;
  wire [3:0] TLMonitor__EVAL_21;
  wire [2:0] TLMonitor__EVAL_22;
  wire  TLMonitor__EVAL_23;
  wire [31:0] TLMonitor__EVAL_24;
  wire  TLMonitor__EVAL_25;
  wire  TLMonitor__EVAL_26;
  wire  TLMonitor__EVAL_27;
  wire  TLMonitor__EVAL_28;
  wire  TLMonitor__EVAL_29;
  wire [3:0] TLMonitor__EVAL_30;
  wire [2:0] TLMonitor__EVAL_31;
  wire  TLMonitor__EVAL_32;
  wire  _EVAL_155;
  wire  _EVAL_197;
  wire  _EVAL_152;
  wire  _EVAL_544;
  wire  _EVAL_147;
  wire  _EVAL_489;
  wire  _EVAL_252;
  wire  _EVAL_527;
  wire  _EVAL_482;
  wire  _EVAL_530;
  wire  _EVAL_212;
  wire  _EVAL_535;
  wire  _EVAL_583;
  wire  _EVAL_542;
  wire  _EVAL_551;
  wire  _EVAL_165;
  wire  _EVAL_303;
  wire  _EVAL_560;
  wire  _EVAL_617;
  wire  _EVAL_465;
  wire  _EVAL_352;
  wire  _EVAL_440;
  wire  _EVAL_411;
  wire  _EVAL_493;
  wire  _EVAL_616;
  wire  _EVAL_305;
  wire  _EVAL_599;
  wire  _EVAL_301;
  wire  _EVAL_444;
  wire  _EVAL_534;
  wire  _EVAL_232;
  wire  _EVAL_285;
  wire  _EVAL_304;
  wire  _EVAL_218;
  wire  _EVAL_367;
  wire  _EVAL_291;
  wire  _EVAL_552;
  wire  _EVAL_470;
  wire  _EVAL_295;
  wire  _EVAL_413;
  wire  _EVAL_494;
  wire  _EVAL_448;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_543;
  wire  _EVAL_363;
  wire  _EVAL_156;
  wire  _EVAL_286;
  wire  _EVAL_462;
  wire  _EVAL_438;
  wire  _EVAL_258;
  wire  _EVAL_167;
  wire  _EVAL_259;
  wire  _EVAL_168;
  wire  _EVAL_611;
  wire  _EVAL_375;
  wire  _EVAL_556;
  wire  _EVAL_579;
  wire  _EVAL_141;
  wire  _EVAL_238;
  wire  _EVAL_143;
  wire  _EVAL_393;
  wire  _EVAL_195;
  wire  _EVAL_528;
  wire  _EVAL_279;
  wire  _EVAL_260;
  wire  _EVAL_510;
  wire  _EVAL_423;
  wire  _EVAL_237;
  wire  _EVAL_205;
  wire  _EVAL_233;
  wire  _EVAL_292;
  wire  _EVAL_317;
  wire  _EVAL_264;
  wire  _EVAL_606;
  SiFive__EVAL_1_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14),
    ._EVAL_15(TLMonitor_1__EVAL_15),
    ._EVAL_16(TLMonitor_1__EVAL_16),
    ._EVAL_17(TLMonitor_1__EVAL_17),
    ._EVAL_18(TLMonitor_1__EVAL_18)
  );
  SiFive__EVAL_0_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18),
    ._EVAL_19(TLMonitor__EVAL_19),
    ._EVAL_20(TLMonitor__EVAL_20),
    ._EVAL_21(TLMonitor__EVAL_21),
    ._EVAL_22(TLMonitor__EVAL_22),
    ._EVAL_23(TLMonitor__EVAL_23),
    ._EVAL_24(TLMonitor__EVAL_24),
    ._EVAL_25(TLMonitor__EVAL_25),
    ._EVAL_26(TLMonitor__EVAL_26),
    ._EVAL_27(TLMonitor__EVAL_27),
    ._EVAL_28(TLMonitor__EVAL_28),
    ._EVAL_29(TLMonitor__EVAL_29),
    ._EVAL_30(TLMonitor__EVAL_30),
    ._EVAL_31(TLMonitor__EVAL_31),
    ._EVAL_32(TLMonitor__EVAL_32)
  );
  assign _EVAL_155 = _EVAL_178 == 1'h0;
  assign _EVAL_197 = _EVAL_435 == 1'h0;
  assign _EVAL_152 = _EVAL_520 == 1'h0;
  assign _EVAL_544 = _EVAL_197 | _EVAL_152;
  assign _EVAL_147 = _EVAL_435 | _EVAL_520;
  assign _EVAL_489 = _EVAL_147 == 1'h0;
  assign _EVAL_252 = _EVAL_460 == 1'h0;
  assign _EVAL_527 = _EVAL_489 | _EVAL_252;
  assign _EVAL_482 = _EVAL_544 & _EVAL_527;
  assign _EVAL_530 = _EVAL_482 | _EVAL_51;
  assign _EVAL_212 = _EVAL_530 == 1'h0;
  assign _EVAL_535 = _EVAL_441 == _EVAL_441;
  assign _EVAL_583 = _EVAL_229 == _EVAL_229;
  assign _EVAL_542 = _EVAL_583 | _EVAL_51;
  assign _EVAL_551 = _EVAL_542 == 1'h0;
  assign _EVAL_165 = _EVAL_535 | _EVAL_51;
  assign _EVAL_303 = _EVAL_158 == 1'h0;
  assign _EVAL_560 = _EVAL_341 | _EVAL_166;
  assign _EVAL_617 = _EVAL_303 | _EVAL_560;
  assign _EVAL_465 = _EVAL_617 | _EVAL_51;
  assign _EVAL_352 = _EVAL_341 == 1'h0;
  assign _EVAL_440 = _EVAL_166 == 1'h0;
  assign _EVAL_411 = _EVAL_352 | _EVAL_440;
  assign _EVAL_493 = _EVAL_165 == 1'h0;
  assign _EVAL_616 = _EVAL_563 | _EVAL_139;
  assign _EVAL_305 = _EVAL_616 | _EVAL_187;
  assign _EVAL_599 = _EVAL_523 | _EVAL_422;
  assign _EVAL_301 = _EVAL_155 | _EVAL_599;
  assign _EVAL_444 = _EVAL_301 | _EVAL_51;
  assign _EVAL_534 = _EVAL_444 == 1'h0;
  assign _EVAL_232 = _EVAL_591 == 1'h0;
  assign _EVAL_285 = _EVAL_147 | _EVAL_460;
  assign _EVAL_304 = _EVAL_232 | _EVAL_285;
  assign _EVAL_218 = _EVAL_304 | _EVAL_51;
  assign _EVAL_367 = _EVAL_539 == 1'h0;
  assign _EVAL_291 = _EVAL_367 | _EVAL_305;
  assign _EVAL_552 = _EVAL_465 == 1'h0;
  assign _EVAL_470 = _EVAL_616 == 1'h0;
  assign _EVAL_295 = _EVAL_140 == _EVAL_140;
  assign _EVAL_413 = _EVAL_295 | _EVAL_51;
  assign _EVAL_494 = _EVAL_413 == 1'h0;
  assign _EVAL_448 = _EVAL_261 == _EVAL_261;
  assign _EVAL_328 = _EVAL_297 == 1'h0;
  assign _EVAL_329 = _EVAL_479 == 1'h0;
  assign _EVAL_543 = _EVAL_328 | _EVAL_329;
  assign _EVAL_363 = _EVAL_139 == 1'h0;
  assign _EVAL_156 = _EVAL_523 == 1'h0;
  assign _EVAL_286 = _EVAL_422 == 1'h0;
  assign _EVAL_462 = _EVAL_156 | _EVAL_286;
  assign _EVAL_438 = _EVAL_462 | _EVAL_51;
  assign _EVAL_258 = _EVAL_438 == 1'h0;
  assign _EVAL_167 = _EVAL_218 == 1'h0;
  assign _EVAL_259 = _EVAL_543 | _EVAL_51;
  assign _EVAL_168 = _EVAL_297 | _EVAL_479;
  assign _EVAL_611 = _EVAL_563 == 1'h0;
  assign _EVAL_375 = _EVAL_611 | _EVAL_363;
  assign _EVAL_556 = _EVAL_366 == 1'h0;
  assign _EVAL_579 = _EVAL_187 == 1'h0;
  assign _EVAL_141 = _EVAL_448 | _EVAL_51;
  assign _EVAL_238 = _EVAL_141 == 1'h0;
  assign _EVAL_143 = _EVAL_620 == _EVAL_620;
  assign _EVAL_393 = _EVAL_143 | _EVAL_51;
  assign _EVAL_195 = _EVAL_411 | _EVAL_51;
  assign _EVAL_528 = _EVAL_259 == 1'h0;
  assign _EVAL_279 = _EVAL_291 | _EVAL_51;
  assign _EVAL_260 = _EVAL_556 | _EVAL_168;
  assign _EVAL_510 = _EVAL_260 | _EVAL_51;
  assign _EVAL_423 = _EVAL_393 == 1'h0;
  assign _EVAL_237 = _EVAL_279 == 1'h0;
  assign _EVAL_205 = _EVAL_470 | _EVAL_579;
  assign _EVAL_233 = _EVAL_375 & _EVAL_205;
  assign _EVAL_292 = _EVAL_195 == 1'h0;
  assign _EVAL_317 = _EVAL_233 | _EVAL_51;
  assign _EVAL_264 = _EVAL_317 == 1'h0;
  assign _EVAL_606 = _EVAL_510 == 1'h0;
  assign TLMonitor__EVAL_26 = _EVAL_42;
  assign TLMonitor_1__EVAL_1 = _EVAL_45;
  assign TLMonitor__EVAL_17 = _EVAL_90;
  assign TLMonitor_1__EVAL = _EVAL_127;
  assign TLMonitor__EVAL_22 = _EVAL_396[82:80];
  assign TLMonitor__EVAL_12 = _EVAL_31;
  assign TLMonitor__EVAL_0 = _EVAL_33;
  assign TLMonitor__EVAL_25 = _EVAL_569 | _EVAL_378;
  assign TLMonitor__EVAL_11 = _EVAL_61;
  assign TLMonitor_1__EVAL_13 = _EVAL_121;
  assign TLMonitor__EVAL_13 = _EVAL_113;
  assign TLMonitor_1__EVAL_14 = _EVAL_84;
  assign TLMonitor__EVAL_4 = _EVAL_71;
  assign TLMonitor_1__EVAL_10 = _EVAL_101;
  assign TLMonitor__EVAL_30 = _EVAL_40;
  assign TLMonitor__EVAL_32 = _EVAL_36;
  assign TLMonitor__EVAL_8 = _EVAL_69;
  assign TLMonitor__EVAL_5 = _EVAL_396[65];
  assign TLMonitor_1__EVAL_5 = _EVAL_60;
  assign TLMonitor_1__EVAL_18 = _EVAL_614[77:74];
  assign TLMonitor__EVAL_3 = _EVAL_396[66];
  assign TLMonitor_1__EVAL_6 = _EVAL_614[65];
  assign TLMonitor_1__EVAL_7 = _EVAL_117;
  assign TLMonitor_1__EVAL_2 = _EVAL_170[5:0];
  assign TLMonitor__EVAL_16 = _EVAL_54;
  assign TLMonitor__EVAL = _EVAL_396[77:74];
  assign TLMonitor__EVAL_14 = _EVAL_396[79:78];
  assign TLMonitor__EVAL_29 = _EVAL_396[0];
  assign TLMonitor__EVAL_18 = _EVAL_101;
  assign TLMonitor__EVAL_1 = _EVAL_9;
  assign TLMonitor__EVAL_24 = _EVAL_114;
  assign TLMonitor_1__EVAL_3 = _EVAL_614[82:80];
  assign TLMonitor_1__EVAL_16 = _EVAL_614[79:78];
  assign TLMonitor__EVAL_10 = _EVAL_235[3:0];
  assign TLMonitor__EVAL_31 = _EVAL_62;
  assign TLMonitor_1__EVAL_0 = _EVAL_327 ? _EVAL_539 : _EVAL_215;
  assign TLMonitor_1__EVAL_8 = _EVAL_15;
  assign TLMonitor__EVAL_27 = _EVAL_103;
  assign TLMonitor_1__EVAL_9 = _EVAL_614[66];
  assign TLMonitor__EVAL_19 = _EVAL_1;
  assign TLMonitor_1__EVAL_12 = _EVAL_311 | _EVAL_243;
  assign TLMonitor__EVAL_20 = _EVAL_67;
  assign TLMonitor_1__EVAL_11 = _EVAL_614[0];
  assign TLMonitor_1__EVAL_15 = _EVAL_3;
  assign TLMonitor__EVAL_9 = _EVAL_290 ? _EVAL_591 : _EVAL_199;
  assign TLMonitor__EVAL_6 = _EVAL_82;
  assign TLMonitor_1__EVAL_17 = _EVAL_13;
  assign TLMonitor_1__EVAL_4 = _EVAL_51;
  assign TLMonitor__EVAL_2 = _EVAL_122;
  assign TLMonitor__EVAL_7 = _EVAL_32;
  assign TLMonitor__EVAL_15 = _EVAL_56;
  assign TLMonitor__EVAL_23 = _EVAL_38;
  assign TLMonitor__EVAL_28 = _EVAL_51;
  assign TLMonitor__EVAL_21 = _EVAL_77;
  always @(posedge _EVAL_101) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_493) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a924c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_493) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_494) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_528) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_423) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_551) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a924c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a924c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_528) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_552) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a924c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_551) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_534) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_552) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_606) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a924c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_606) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
