//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_53_assert(
  input  [2:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [31:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [5:0] _EVAL_36;
  reg [31:0] _RAND_0;
  reg [5:0] _EVAL_59;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_64;
  reg [31:0] _RAND_2;
  reg  _EVAL_105;
  reg [31:0] _RAND_3;
  reg  _EVAL_152;
  reg [31:0] _RAND_4;
  reg  _EVAL_157;
  reg [31:0] _RAND_5;
  reg [31:0] _EVAL_163;
  reg [31:0] _RAND_6;
  reg [5:0] _EVAL_221;
  reg [31:0] _RAND_7;
  reg [5:0] _EVAL_233;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_241;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_246;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_249;
  reg [31:0] _RAND_11;
  reg [2:0] _EVAL_256;
  reg [31:0] _RAND_12;
  reg [31:0] _EVAL_269;
  reg [31:0] _RAND_13;
  wire  _EVAL_141;
  wire  _EVAL_276;
  wire [5:0] _EVAL_177;
  wire  _EVAL_186;
  wire [1:0] _EVAL_296;
  wire [1:0] _EVAL_127;
  wire  _EVAL_206;
  wire [31:0] _EVAL_220;
  wire [32:0] _EVAL_65;
  wire [32:0] _EVAL_95;
  wire  _EVAL_33;
  wire  _EVAL_275;
  wire  _EVAL_245;
  wire  _EVAL_281;
  wire  _EVAL_280;
  wire  _EVAL_26;
  wire [31:0] _EVAL_271;
  wire [32:0] _EVAL_175;
  wire  _EVAL_219;
  wire  _EVAL_184;
  wire  _EVAL_261;
  wire  _EVAL_97;
  wire  _EVAL_117;
  wire  _EVAL_79;
  wire  _EVAL_201;
  wire  _EVAL_22;
  wire  _EVAL_240;
  wire  _EVAL_260;
  wire  _EVAL_124;
  wire  _EVAL_212;
  wire  _EVAL_143;
  wire [31:0] _EVAL_42;
  wire [32:0] _EVAL_90;
  wire [32:0] _EVAL_46;
  wire [32:0] _EVAL_160;
  wire [22:0] _EVAL_287;
  wire [7:0] _EVAL_48;
  wire [7:0] _EVAL_100;
  wire [31:0] _EVAL_165;
  wire [31:0] _EVAL_62;
  wire  _EVAL_192;
  wire  _EVAL_198;
  wire [31:0] _EVAL_31;
  wire [32:0] _EVAL_199;
  wire [32:0] _EVAL_252;
  wire [32:0] _EVAL_34;
  wire  _EVAL_224;
  wire  _EVAL_102;
  wire [5:0] _EVAL_209;
  wire [5:0] _EVAL_255;
  wire  _EVAL_151;
  wire [31:0] _EVAL_270;
  wire [32:0] _EVAL_204;
  wire [32:0] _EVAL_291;
  wire [32:0] _EVAL_251;
  wire  _EVAL_24;
  wire [31:0] _EVAL_264;
  wire [32:0] _EVAL_15;
  wire [32:0] _EVAL_267;
  wire [32:0] _EVAL_229;
  wire  _EVAL_72;
  wire  _EVAL_180;
  wire [32:0] _EVAL_215;
  wire [32:0] _EVAL_99;
  wire  _EVAL_166;
  wire  _EVAL_294;
  wire  _EVAL_91;
  wire  _EVAL_257;
  wire [32:0] _EVAL_41;
  wire [32:0] _EVAL_149;
  wire [32:0] _EVAL_277;
  wire  _EVAL_128;
  wire  _EVAL_30;
  wire [31:0] _EVAL_21;
  wire [32:0] _EVAL_55;
  wire [32:0] _EVAL_32;
  wire [32:0] _EVAL_195;
  wire  _EVAL_182;
  wire  _EVAL_286;
  wire [32:0] _EVAL_53;
  wire  _EVAL_216;
  wire  _EVAL_106;
  wire [31:0] _EVAL_173;
  wire [32:0] _EVAL_136;
  wire [32:0] _EVAL_56;
  wire [32:0] _EVAL_129;
  wire  _EVAL_236;
  wire  _EVAL_148;
  wire  _EVAL_292;
  wire  _EVAL_285;
  wire  _EVAL_248;
  wire  _EVAL_19;
  wire  _EVAL_44;
  wire  _EVAL_109;
  wire  _EVAL_227;
  wire  _EVAL_290;
  wire  _EVAL_47;
  wire  _EVAL_189;
  wire [3:0] _EVAL_161;
  wire  _EVAL_176;
  wire  _EVAL_89;
  wire  _EVAL_168;
  wire  _EVAL_54;
  wire  _EVAL_153;
  wire  _EVAL_145;
  wire  _EVAL_107;
  wire  _EVAL_123;
  wire  _EVAL_172;
  wire  _EVAL_84;
  wire  _EVAL_162;
  wire  _EVAL_27;
  wire  _EVAL_235;
  wire  _EVAL_74;
  wire [1:0] _EVAL_170;
  wire  _EVAL_197;
  wire  _EVAL_283;
  wire  _EVAL_92;
  wire  _EVAL_67;
  wire  _EVAL_211;
  wire  _EVAL_49;
  wire  _EVAL_25;
  wire [1:0] _EVAL_265;
  wire  _EVAL_16;
  wire  _EVAL_96;
  wire  _EVAL_222;
  wire  _EVAL_98;
  wire  _EVAL_58;
  wire  _EVAL_103;
  wire  _EVAL_188;
  wire  _EVAL_23;
  wire  _EVAL_78;
  wire  _EVAL_125;
  wire  _EVAL_119;
  wire [22:0] _EVAL_258;
  wire [7:0] _EVAL_147;
  wire [7:0] _EVAL_203;
  wire [5:0] _EVAL_88;
  wire [5:0] _EVAL_156;
  wire  _EVAL_137;
  wire  _EVAL_230;
  wire  _EVAL_200;
  wire  _EVAL_181;
  wire  _EVAL_218;
  wire  _EVAL_150;
  wire  _EVAL_239;
  wire  _EVAL_131;
  wire  _EVAL_185;
  wire  _EVAL_234;
  wire  _EVAL_146;
  wire  _EVAL_142;
  wire  _EVAL_40;
  wire  _EVAL_112;
  wire  _EVAL_50;
  wire [3:0] _EVAL_60;
  wire [3:0] _EVAL_37;
  wire [3:0] _EVAL_43;
  wire  _EVAL_279;
  wire  _EVAL_52;
  wire  _EVAL_158;
  wire  _EVAL_214;
  wire  _EVAL_244;
  wire [31:0] _EVAL_45;
  wire  _EVAL_225;
  wire  _EVAL_101;
  wire  _EVAL_57;
  wire  _EVAL_295;
  wire  _EVAL_144;
  wire  _EVAL_268;
  wire  _EVAL_116;
  wire  _EVAL_110;
  wire  _EVAL_61;
  wire  _EVAL_190;
  wire  _EVAL_135;
  wire  _EVAL_159;
  wire  _EVAL_83;
  wire  _EVAL_169;
  wire  _EVAL_254;
  wire  _EVAL_263;
  wire  _EVAL_28;
  wire  _EVAL_250;
  wire  _EVAL_242;
  wire  _EVAL_118;
  wire  _EVAL_272;
  wire  _EVAL_75;
  wire  _EVAL_66;
  wire  _EVAL_213;
  wire  _EVAL_126;
  wire  _EVAL_293;
  wire  _EVAL_237;
  wire  _EVAL_17;
  wire  _EVAL_134;
  wire  _EVAL_69;
  wire  _EVAL_282;
  wire  _EVAL_87;
  wire  _EVAL_217;
  wire  _EVAL_104;
  wire  _EVAL_183;
  wire  _EVAL_29;
  wire  _EVAL_18;
  wire  _EVAL_278;
  wire  _EVAL_63;
  wire  _EVAL_179;
  wire  _EVAL_266;
  wire  _EVAL_68;
  wire  _EVAL_133;
  wire  _EVAL_194;
  wire  _EVAL_114;
  wire  _EVAL_130;
  wire  _EVAL_139;
  wire  _EVAL_93;
  wire  _EVAL_85;
  wire  _EVAL_140;
  wire [5:0] _EVAL_210;
  wire  _EVAL_35;
  wire  _EVAL_187;
  wire  _EVAL_289;
  wire  _EVAL_138;
  wire  _EVAL_274;
  wire  _EVAL_253;
  wire  _EVAL_120;
  wire  _EVAL_164;
  wire  _EVAL_228;
  wire  _EVAL_82;
  wire  _EVAL_171;
  wire  _EVAL_238;
  wire  _EVAL_77;
  wire  _EVAL_247;
  wire  _EVAL_121;
  wire  _EVAL_262;
  wire  _EVAL_111;
  wire  _EVAL_232;
  wire  _EVAL_167;
  wire  _EVAL_70;
  wire  _EVAL_297;
  wire  _EVAL_202;
  wire  _EVAL_73;
  wire  _EVAL_154;
  wire  _EVAL_81;
  wire  _EVAL_207;
  wire  _EVAL_20;
  wire  _EVAL_259;
  wire  _EVAL_288;
  wire  _EVAL_284;
  wire  _EVAL_205;
  wire  _EVAL_39;
  wire  _EVAL_76;
  wire  _EVAL_51;
  wire  _EVAL_178;
  wire  _EVAL_71;
  wire  _EVAL_94;
  wire  _EVAL_122;
  wire  _EVAL_273;
  wire  _EVAL_196;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_141 = _EVAL_12 == 1'h0;
  assign _EVAL_276 = _EVAL_141 | _EVAL_1;
  assign _EVAL_177 = _EVAL_59 - 6'h1;
  assign _EVAL_186 = _EVAL_13[0];
  assign _EVAL_296 = 2'h1 << _EVAL_186;
  assign _EVAL_127 = _EVAL_296 | 2'h1;
  assign _EVAL_206 = _EVAL_127[0];
  assign _EVAL_220 = _EVAL_4 ^ 32'h1900000;
  assign _EVAL_65 = {1'b0,$signed(_EVAL_220)};
  assign _EVAL_95 = $signed(_EVAL_65) & $signed(-33'sh2000);
  assign _EVAL_33 = _EVAL_233 == 6'h0;
  assign _EVAL_275 = _EVAL_33 == 1'h0;
  assign _EVAL_245 = _EVAL_11 & _EVAL_275;
  assign _EVAL_281 = _EVAL_10 == 3'h0;
  assign _EVAL_280 = _EVAL == 3'h6;
  assign _EVAL_26 = _EVAL_11 & _EVAL_280;
  assign _EVAL_271 = _EVAL_4 ^ 32'hc000000;
  assign _EVAL_175 = {1'b0,$signed(_EVAL_271)};
  assign _EVAL_219 = _EVAL_13 >= 4'h2;
  assign _EVAL_184 = _EVAL_127[1];
  assign _EVAL_261 = _EVAL_4[1];
  assign _EVAL_97 = _EVAL_184 & _EVAL_261;
  assign _EVAL_117 = _EVAL_219 | _EVAL_97;
  assign _EVAL_79 = _EVAL_219 | _EVAL_1;
  assign _EVAL_201 = _EVAL_4 == _EVAL_163;
  assign _EVAL_22 = _EVAL_201 | _EVAL_1;
  assign _EVAL_240 = _EVAL_22 == 1'h0;
  assign _EVAL_260 = _EVAL[2];
  assign _EVAL_124 = _EVAL_2 == 1'h0;
  assign _EVAL_212 = _EVAL_124 | _EVAL_1;
  assign _EVAL_143 = _EVAL_212 == 1'h0;
  assign _EVAL_42 = _EVAL_4 ^ 32'h2000000;
  assign _EVAL_90 = {1'b0,$signed(_EVAL_42)};
  assign _EVAL_46 = $signed(_EVAL_90) & $signed(-33'sh10000);
  assign _EVAL_160 = $signed(_EVAL_46);
  assign _EVAL_287 = 23'hff << _EVAL_13;
  assign _EVAL_48 = _EVAL_287[7:0];
  assign _EVAL_100 = ~ _EVAL_48;
  assign _EVAL_165 = {{24'd0}, _EVAL_100};
  assign _EVAL_62 = _EVAL_4 & _EVAL_165;
  assign _EVAL_192 = _EVAL_62 == 32'h0;
  assign _EVAL_198 = _EVAL_192 | _EVAL_1;
  assign _EVAL_31 = _EVAL_4 ^ 32'h3000;
  assign _EVAL_199 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_252 = $signed(_EVAL_199) & $signed(-33'sh1000);
  assign _EVAL_34 = $signed(_EVAL_252);
  assign _EVAL_224 = $signed(_EVAL_34) == $signed(33'sh0);
  assign _EVAL_102 = _EVAL_260 == 1'h0;
  assign _EVAL_209 = _EVAL_100[7:2];
  assign _EVAL_255 = _EVAL_233 - 6'h1;
  assign _EVAL_151 = _EVAL_13 <= 4'h6;
  assign _EVAL_270 = _EVAL_4 ^ 32'h40000000;
  assign _EVAL_204 = {1'b0,$signed(_EVAL_270)};
  assign _EVAL_291 = $signed(_EVAL_204) & $signed(-33'sh2000);
  assign _EVAL_251 = $signed(_EVAL_291);
  assign _EVAL_24 = $signed(_EVAL_251) == $signed(33'sh0);
  assign _EVAL_264 = _EVAL_4 ^ 32'h80000000;
  assign _EVAL_15 = {1'b0,$signed(_EVAL_264)};
  assign _EVAL_267 = $signed(_EVAL_15) & $signed(-33'sh20000);
  assign _EVAL_229 = $signed(_EVAL_267);
  assign _EVAL_72 = $signed(_EVAL_229) == $signed(33'sh0);
  assign _EVAL_180 = _EVAL_24 | _EVAL_72;
  assign _EVAL_215 = $signed(_EVAL_175) & $signed(-33'sh4000000);
  assign _EVAL_99 = $signed(_EVAL_215);
  assign _EVAL_166 = $signed(_EVAL_99) == $signed(33'sh0);
  assign _EVAL_294 = _EVAL_180 | _EVAL_166;
  assign _EVAL_91 = $signed(_EVAL_160) == $signed(33'sh0);
  assign _EVAL_257 = _EVAL_294 | _EVAL_91;
  assign _EVAL_41 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_149 = $signed(_EVAL_41) & $signed(-33'sh5000);
  assign _EVAL_277 = $signed(_EVAL_149);
  assign _EVAL_128 = $signed(_EVAL_277) == $signed(33'sh0);
  assign _EVAL_30 = _EVAL_257 | _EVAL_128;
  assign _EVAL_21 = _EVAL_4 ^ 32'h1800000;
  assign _EVAL_55 = {1'b0,$signed(_EVAL_21)};
  assign _EVAL_32 = $signed(_EVAL_55) & $signed(-33'sh8000);
  assign _EVAL_195 = $signed(_EVAL_32);
  assign _EVAL_182 = $signed(_EVAL_195) == $signed(33'sh0);
  assign _EVAL_286 = _EVAL_30 | _EVAL_182;
  assign _EVAL_53 = $signed(_EVAL_95);
  assign _EVAL_216 = $signed(_EVAL_53) == $signed(33'sh0);
  assign _EVAL_106 = _EVAL_286 | _EVAL_216;
  assign _EVAL_173 = _EVAL_4 ^ 32'h20000000;
  assign _EVAL_136 = {1'b0,$signed(_EVAL_173)};
  assign _EVAL_56 = $signed(_EVAL_136) & $signed(-33'sh2000);
  assign _EVAL_129 = $signed(_EVAL_56);
  assign _EVAL_236 = $signed(_EVAL_129) == $signed(33'sh0);
  assign _EVAL_148 = _EVAL_106 | _EVAL_236;
  assign _EVAL_292 = _EVAL_151 & _EVAL_148;
  assign _EVAL_285 = _EVAL_13 <= 4'h8;
  assign _EVAL_248 = _EVAL_285 & _EVAL_224;
  assign _EVAL_19 = _EVAL_292 | _EVAL_248;
  assign _EVAL_44 = _EVAL_19 | _EVAL_1;
  assign _EVAL_109 = _EVAL_44 == 1'h0;
  assign _EVAL_227 = _EVAL_261 == 1'h0;
  assign _EVAL_290 = _EVAL_4[0];
  assign _EVAL_47 = _EVAL_227 & _EVAL_290;
  assign _EVAL_189 = _EVAL_206 & _EVAL_47;
  assign _EVAL_161 = ~ _EVAL_9;
  assign _EVAL_176 = _EVAL_161 == 4'h0;
  assign _EVAL_89 = _EVAL_176 | _EVAL_1;
  assign _EVAL_168 = _EVAL_89 == 1'h0;
  assign _EVAL_54 = _EVAL_59 == 6'h0;
  assign _EVAL_153 = _EVAL_54 == 1'h0;
  assign _EVAL_145 = _EVAL_14 & _EVAL_153;
  assign _EVAL_107 = _EVAL_10 == _EVAL_249;
  assign _EVAL_123 = _EVAL_107 | _EVAL_1;
  assign _EVAL_172 = _EVAL_224 | _EVAL_166;
  assign _EVAL_84 = _EVAL_172 | _EVAL_91;
  assign _EVAL_162 = _EVAL_84 | _EVAL_128;
  assign _EVAL_27 = _EVAL_8 & _EVAL_11;
  assign _EVAL_235 = _EVAL_36 == 6'h0;
  assign _EVAL_74 = _EVAL_27 & _EVAL_235;
  assign _EVAL_170 = _EVAL_74 ? 2'h1 : 2'h0;
  assign _EVAL_197 = _EVAL_170[0];
  assign _EVAL_283 = _EVAL_6 & _EVAL_14;
  assign _EVAL_92 = _EVAL_221 == 6'h0;
  assign _EVAL_67 = _EVAL_283 & _EVAL_92;
  assign _EVAL_211 = _EVAL_10 == 3'h6;
  assign _EVAL_49 = _EVAL_211 == 1'h0;
  assign _EVAL_25 = _EVAL_67 & _EVAL_49;
  assign _EVAL_265 = _EVAL_25 ? 2'h1 : 2'h0;
  assign _EVAL_16 = _EVAL_265[0];
  assign _EVAL_96 = _EVAL_197 != _EVAL_16;
  assign _EVAL_222 = _EVAL_197 == 1'h0;
  assign _EVAL_98 = _EVAL_96 | _EVAL_222;
  assign _EVAL_58 = _EVAL_7 == _EVAL_246;
  assign _EVAL_103 = _EVAL_248 | _EVAL_1;
  assign _EVAL_188 = _EVAL_103 == 1'h0;
  assign _EVAL_23 = _EVAL_3 == _EVAL_157;
  assign _EVAL_78 = _EVAL_23 | _EVAL_1;
  assign _EVAL_125 = _EVAL_78 == 1'h0;
  assign _EVAL_119 = _EVAL_10[0];
  assign _EVAL_258 = 23'hff << _EVAL_0;
  assign _EVAL_147 = _EVAL_258[7:0];
  assign _EVAL_203 = ~ _EVAL_147;
  assign _EVAL_88 = _EVAL_203[7:2];
  assign _EVAL_156 = _EVAL_221 - 6'h1;
  assign _EVAL_137 = _EVAL == _EVAL_256;
  assign _EVAL_230 = _EVAL_290 == 1'h0;
  assign _EVAL_200 = _EVAL_261 & _EVAL_230;
  assign _EVAL_181 = _EVAL_206 & _EVAL_200;
  assign _EVAL_218 = _EVAL_151 & _EVAL_72;
  assign _EVAL_150 = _EVAL_261 & _EVAL_290;
  assign _EVAL_239 = _EVAL_206 & _EVAL_150;
  assign _EVAL_131 = _EVAL_117 | _EVAL_239;
  assign _EVAL_185 = _EVAL_117 | _EVAL_181;
  assign _EVAL_234 = _EVAL_184 & _EVAL_227;
  assign _EVAL_146 = _EVAL_219 | _EVAL_234;
  assign _EVAL_142 = _EVAL_146 | _EVAL_189;
  assign _EVAL_40 = _EVAL_227 & _EVAL_230;
  assign _EVAL_112 = _EVAL_206 & _EVAL_40;
  assign _EVAL_50 = _EVAL_146 | _EVAL_112;
  assign _EVAL_60 = {_EVAL_131,_EVAL_185,_EVAL_142,_EVAL_50};
  assign _EVAL_37 = ~ _EVAL_60;
  assign _EVAL_43 = _EVAL_9 & _EVAL_37;
  assign _EVAL_279 = _EVAL_43 == 4'h0;
  assign _EVAL_52 = _EVAL_197 | _EVAL_105;
  assign _EVAL_158 = _EVAL_52 | _EVAL_1;
  assign _EVAL_214 = _EVAL_79 == 1'h0;
  assign _EVAL_244 = _EVAL_27 | _EVAL_283;
  assign _EVAL_45 = _EVAL_269 + 32'h1;
  assign _EVAL_225 = _EVAL_7 == 2'h0;
  assign _EVAL_101 = _EVAL_225 | _EVAL_1;
  assign _EVAL_57 = _EVAL_101 == 1'h0;
  assign _EVAL_295 = _EVAL == 3'h5;
  assign _EVAL_144 = _EVAL_11 & _EVAL_295;
  assign _EVAL_268 = _EVAL_13 <= 4'h2;
  assign _EVAL_116 = _EVAL_162 | _EVAL_182;
  assign _EVAL_110 = _EVAL_116 | _EVAL_216;
  assign _EVAL_61 = _EVAL_110 | _EVAL_236;
  assign _EVAL_190 = _EVAL_268 & _EVAL_61;
  assign _EVAL_135 = _EVAL_190 | _EVAL_1;
  assign _EVAL_159 = _EVAL_124 | _EVAL_12;
  assign _EVAL_83 = _EVAL_159 | _EVAL_1;
  assign _EVAL_169 = _EVAL_83 == 1'h0;
  assign _EVAL_254 = _EVAL_10 == 3'h4;
  assign _EVAL_263 = _EVAL == 3'h3;
  assign _EVAL_28 = _EVAL == 3'h4;
  assign _EVAL_250 = _EVAL_11 & _EVAL_28;
  assign _EVAL_242 = _EVAL_13 == _EVAL_241;
  assign _EVAL_118 = _EVAL_123 == 1'h0;
  assign _EVAL_272 = _EVAL_10 == 3'h2;
  assign _EVAL_75 = _EVAL_198 == 1'h0;
  assign _EVAL_66 = _EVAL == 3'h0;
  assign _EVAL_213 = _EVAL_135 == 1'h0;
  assign _EVAL_126 = _EVAL_7 != 2'h2;
  assign _EVAL_293 = _EVAL_126 | _EVAL_1;
  assign _EVAL_237 = _EVAL_293 == 1'h0;
  assign _EVAL_17 = _EVAL_137 | _EVAL_1;
  assign _EVAL_134 = _EVAL_17 == 1'h0;
  assign _EVAL_69 = _EVAL == 3'h1;
  assign _EVAL_282 = _EVAL_279 | _EVAL_1;
  assign _EVAL_87 = _EVAL_242 | _EVAL_1;
  assign _EVAL_217 = _EVAL_10 == 3'h5;
  assign _EVAL_104 = _EVAL_14 & _EVAL_217;
  assign _EVAL_183 = _EVAL_10 == 3'h1;
  assign _EVAL_29 = _EVAL_105 == 1'h0;
  assign _EVAL_18 = plusarg_reader_out == 32'h0;
  assign _EVAL_278 = _EVAL_29 | _EVAL_18;
  assign _EVAL_63 = _EVAL_269 < plusarg_reader_out;
  assign _EVAL_179 = _EVAL_278 | _EVAL_63;
  assign _EVAL_266 = _EVAL_179 | _EVAL_1;
  assign _EVAL_68 = _EVAL_266 == 1'h0;
  assign _EVAL_133 = _EVAL_0 >= 4'h2;
  assign _EVAL_194 = _EVAL_0 == _EVAL_64;
  assign _EVAL_114 = _EVAL_194 | _EVAL_1;
  assign _EVAL_130 = _EVAL_98 | _EVAL_1;
  assign _EVAL_139 = _EVAL_283 & _EVAL_54;
  assign _EVAL_93 = _EVAL_105 | _EVAL_197;
  assign _EVAL_85 = ~ _EVAL_16;
  assign _EVAL_140 = _EVAL_93 & _EVAL_85;
  assign _EVAL_210 = _EVAL_36 - 6'h1;
  assign _EVAL_35 = _EVAL_218 | _EVAL_1;
  assign _EVAL_187 = _EVAL_35 == 1'h0;
  assign _EVAL_289 = _EVAL_58 | _EVAL_1;
  assign _EVAL_138 = _EVAL_10 <= 3'h6;
  assign _EVAL_274 = _EVAL_138 | _EVAL_1;
  assign _EVAL_253 = _EVAL_274 == 1'h0;
  assign _EVAL_120 = _EVAL_11 & _EVAL_66;
  assign _EVAL_164 = _EVAL_9 == _EVAL_60;
  assign _EVAL_228 = _EVAL_164 | _EVAL_1;
  assign _EVAL_82 = _EVAL_2 == _EVAL_152;
  assign _EVAL_171 = _EVAL_82 | _EVAL_1;
  assign _EVAL_238 = _EVAL_171 == 1'h0;
  assign _EVAL_77 = _EVAL_289 == 1'h0;
  assign _EVAL_247 = _EVAL_29 | _EVAL_1;
  assign _EVAL_121 = _EVAL == 3'h7;
  assign _EVAL_262 = _EVAL_276 == 1'h0;
  assign _EVAL_111 = _EVAL_14 & _EVAL_183;
  assign _EVAL_232 = _EVAL_7 <= 2'h2;
  assign _EVAL_167 = _EVAL_232 | _EVAL_1;
  assign _EVAL_70 = _EVAL_167 == 1'h0;
  assign _EVAL_297 = _EVAL_133 | _EVAL_1;
  assign _EVAL_202 = _EVAL_297 == 1'h0;
  assign _EVAL_73 = _EVAL_27 & _EVAL_33;
  assign _EVAL_154 = _EVAL == 3'h2;
  assign _EVAL_81 = _EVAL_11 & _EVAL_263;
  assign _EVAL_207 = _EVAL_14 & _EVAL_272;
  assign _EVAL_20 = _EVAL_14 & _EVAL_254;
  assign _EVAL_259 = _EVAL_247 == 1'h0;
  assign _EVAL_288 = _EVAL_14 & _EVAL_211;
  assign _EVAL_284 = _EVAL_87 == 1'h0;
  assign _EVAL_205 = _EVAL_14 & _EVAL_281;
  assign _EVAL_39 = _EVAL_1 == 1'h0;
  assign _EVAL_76 = _EVAL_158 == 1'h0;
  assign _EVAL_51 = _EVAL_228 == 1'h0;
  assign _EVAL_178 = _EVAL_11 & _EVAL_154;
  assign _EVAL_71 = _EVAL_130 == 1'h0;
  assign _EVAL_94 = _EVAL_114 == 1'h0;
  assign _EVAL_122 = _EVAL_11 & _EVAL_121;
  assign _EVAL_273 = _EVAL_11 & _EVAL_69;
  assign _EVAL_196 = _EVAL_282 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_36 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_59 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_105 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_152 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_157 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_163 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_221 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_233 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_241 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_246 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_249 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_256 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_269 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_5) begin
    if (_EVAL_1) begin
      _EVAL_36 <= 6'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_235) begin
          if (_EVAL_102) begin
            _EVAL_36 <= _EVAL_209;
          end else begin
            _EVAL_36 <= 6'h0;
          end
        end else begin
          _EVAL_36 <= _EVAL_210;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_59 <= 6'h0;
    end else begin
      if (_EVAL_283) begin
        if (_EVAL_54) begin
          if (_EVAL_119) begin
            _EVAL_59 <= _EVAL_88;
          end else begin
            _EVAL_59 <= 6'h0;
          end
        end else begin
          _EVAL_59 <= _EVAL_177;
        end
      end
    end
    if (_EVAL_139) begin
      _EVAL_64 <= _EVAL_0;
    end
    if (_EVAL_1) begin
      _EVAL_105 <= 1'h0;
    end else begin
      _EVAL_105 <= _EVAL_140;
    end
    if (_EVAL_139) begin
      _EVAL_152 <= _EVAL_2;
    end
    if (_EVAL_139) begin
      _EVAL_157 <= _EVAL_3;
    end
    if (_EVAL_73) begin
      _EVAL_163 <= _EVAL_4;
    end
    if (_EVAL_1) begin
      _EVAL_221 <= 6'h0;
    end else begin
      if (_EVAL_283) begin
        if (_EVAL_92) begin
          if (_EVAL_119) begin
            _EVAL_221 <= _EVAL_88;
          end else begin
            _EVAL_221 <= 6'h0;
          end
        end else begin
          _EVAL_221 <= _EVAL_156;
        end
      end
    end
    if (_EVAL_1) begin
      _EVAL_233 <= 6'h0;
    end else begin
      if (_EVAL_27) begin
        if (_EVAL_33) begin
          if (_EVAL_102) begin
            _EVAL_233 <= _EVAL_209;
          end else begin
            _EVAL_233 <= 6'h0;
          end
        end else begin
          _EVAL_233 <= _EVAL_255;
        end
      end
    end
    if (_EVAL_73) begin
      _EVAL_241 <= _EVAL_13;
    end
    if (_EVAL_139) begin
      _EVAL_246 <= _EVAL_7;
    end
    if (_EVAL_139) begin
      _EVAL_249 <= _EVAL_10;
    end
    if (_EVAL_73) begin
      _EVAL_256 <= _EVAL;
    end
    if (_EVAL_1) begin
      _EVAL_269 <= 32'h0;
    end else begin
      if (_EVAL_244) begin
        _EVAL_269 <= 32'h0;
      end else begin
        _EVAL_269 <= _EVAL_45;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b954c816)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(116506c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac26eb40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45f2f3ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbb81728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b19fcb6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba28fd9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2297f7cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e7b0b67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66b5f7d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51b238c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1661524)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c5ec967)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f6bd04b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3d52980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1adfe509)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d318f3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(241c2ce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9514fca7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d16d8d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b47e6d97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68b774dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42cb08da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fd8715c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b22b3fc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(746a35ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4e61cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e912bffd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82c5765c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d4e414)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f94657a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d968708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1b7e973)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ccf762f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5267dbf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f78b77c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6caaf1cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b59705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(315a61e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7109585b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d081859)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec4250d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bd8322c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f053bb09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b24b78e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(259a954)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe0b24b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a13bc1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ce0b4d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(511c5d11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e99c765)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adfed718)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3db2455)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c117fbfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d52abedd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5273662)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a1a1ce8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d89ae924)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33aa10ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(266385e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
