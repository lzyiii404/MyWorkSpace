//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_112(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [31:0] _EVAL_6,
  output [29:0] _EVAL_7,
  output [31:0] _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  output [2:0]  _EVAL_13,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  input  [29:0] _EVAL_16,
  output [6:0]  _EVAL_17,
  output [3:0]  _EVAL_18,
  output [2:0]  _EVAL_19,
  output        _EVAL_20,
  input  [6:0]  _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output [31:0] _EVAL_25,
  output [3:0]  _EVAL_26,
  output        _EVAL_27,
  output [3:0]  _EVAL_28,
  input  [31:0] _EVAL_29,
  output [6:0]  _EVAL_30,
  input  [3:0]  _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input  [6:0]  _EVAL_34,
  output [1:0]  _EVAL_35,
  output        _EVAL_36,
  output [2:0]  _EVAL_37,
  output        _EVAL_38,
  input         _EVAL_39,
  input  [3:0]  _EVAL_40
);
  reg  _EVAL_43;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_49;
  reg [31:0] _RAND_1;
  reg  _EVAL_90;
  reg [31:0] _RAND_2;
  reg  _EVAL_99;
  reg [31:0] _RAND_3;
  reg  _EVAL_141;
  reg [31:0] _RAND_4;
  reg  _EVAL_143;
  reg [31:0] _RAND_5;
  reg  _EVAL_160;
  reg [31:0] _RAND_6;
  reg  _EVAL_170;
  reg [31:0] _RAND_7;
  reg  _EVAL_173;
  reg [31:0] _RAND_8;
  reg  _EVAL_204;
  reg [31:0] _RAND_9;
  reg  _EVAL_212;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_216;
  reg [31:0] _RAND_11;
  reg  _EVAL_219;
  reg [31:0] _RAND_12;
  reg [5:0] _EVAL_244;
  reg [31:0] _RAND_13;
  reg  _EVAL_273;
  reg [31:0] _RAND_14;
  reg  _EVAL_293;
  reg [31:0] _RAND_15;
  reg  _EVAL_296;
  reg [31:0] _RAND_16;
  reg  _EVAL_302;
  reg [31:0] _RAND_17;
  reg  _EVAL_326;
  reg [31:0] _RAND_18;
  reg [3:0] _EVAL_334;
  reg [31:0] _RAND_19;
  reg  _EVAL_336;
  reg [31:0] _RAND_20;
  reg  _EVAL_338;
  reg [31:0] _RAND_21;
  reg  _EVAL_344;
  reg [31:0] _RAND_22;
  reg  _EVAL_357;
  reg [31:0] _RAND_23;
  reg  _EVAL_358;
  reg [31:0] _RAND_24;
  reg [3:0] _EVAL_359;
  reg [31:0] _RAND_25;
  reg  _EVAL_370;
  reg [31:0] _RAND_26;
  reg  _EVAL_401;
  reg [31:0] _RAND_27;
  reg  _EVAL_410;
  reg [31:0] _RAND_28;
  reg  _EVAL_413;
  reg [31:0] _RAND_29;
  reg [5:0] _EVAL_474;
  reg [31:0] _RAND_30;
  reg  _EVAL_476;
  reg [31:0] _RAND_31;
  reg  _EVAL_490;
  reg [31:0] _RAND_32;
  reg  _EVAL_491;
  reg [31:0] _RAND_33;
  reg  _EVAL_501;
  reg [31:0] _RAND_34;
  reg [3:0] _EVAL_503;
  reg [31:0] _RAND_35;
  reg  _EVAL_511;
  reg [31:0] _RAND_36;
  reg  _EVAL_553;
  reg [31:0] _RAND_37;
  reg  _EVAL_556;
  reg [31:0] _RAND_38;
  reg  _EVAL_569;
  reg [31:0] _RAND_39;
  reg  _EVAL_598;
  reg [31:0] _RAND_40;
  reg  _EVAL_603;
  reg [31:0] _RAND_41;
  reg  _EVAL_623;
  reg [31:0] _RAND_42;
  reg  _EVAL_630;
  reg [31:0] _RAND_43;
  reg  _EVAL_634;
  reg [31:0] _RAND_44;
  reg  _EVAL_640;
  reg [31:0] _RAND_45;
  wire  _EVAL_346;
  wire [3:0] _EVAL_291;
  wire  _EVAL_282;
  wire [2:0] _EVAL_387;
  wire  _EVAL_199;
  wire  _EVAL_178;
  wire  _EVAL_87;
  wire  _EVAL_211;
  wire  _EVAL_595;
  wire  _EVAL_619;
  wire  _EVAL_521;
  wire  _EVAL_218;
  wire  _EVAL_455;
  wire  _EVAL_464;
  wire [29:0] _EVAL_260;
  wire [30:0] _EVAL_202;
  wire [30:0] _EVAL_116;
  wire [30:0] _EVAL_295;
  wire  _EVAL_487;
  wire [1:0] _EVAL_187;
  wire [29:0] _EVAL_284;
  wire [30:0] _EVAL_84;
  wire [30:0] _EVAL_55;
  wire [30:0] _EVAL_451;
  wire  _EVAL_51;
  wire [1:0] _EVAL_197;
  wire [1:0] _EVAL_612;
  wire [2:0] _EVAL_75;
  wire [29:0] _EVAL_201;
  wire [30:0] _EVAL_520;
  wire [30:0] _EVAL_261;
  wire [30:0] _EVAL_243;
  wire  _EVAL_74;
  wire [2:0] _EVAL_222;
  wire [2:0] _EVAL_114;
  wire [30:0] _EVAL_149;
  wire [30:0] _EVAL_183;
  wire [30:0] _EVAL_163;
  wire  _EVAL_380;
  wire [2:0] _EVAL_460;
  wire [2:0] _EVAL_221;
  wire [3:0] _EVAL_303;
  wire [29:0] _EVAL_298;
  wire [30:0] _EVAL_593;
  wire [30:0] _EVAL_544;
  wire [30:0] _EVAL_418;
  wire  _EVAL_446;
  wire [3:0] _EVAL_79;
  wire [3:0] _EVAL_400;
  wire [29:0] _EVAL_409;
  wire [30:0] _EVAL_288;
  wire [30:0] _EVAL_399;
  wire [30:0] _EVAL_59;
  wire  _EVAL_226;
  wire [1:0] _EVAL_481;
  wire [3:0] _EVAL_255;
  wire [3:0] _EVAL_287;
  wire [29:0] _EVAL_354;
  wire [30:0] _EVAL_405;
  wire [30:0] _EVAL_541;
  wire [30:0] _EVAL_41;
  wire  _EVAL_180;
  wire [2:0] _EVAL_574;
  wire [3:0] _EVAL_292;
  wire [3:0] _EVAL_104;
  wire [29:0] _EVAL_624;
  wire [30:0] _EVAL_352;
  wire [30:0] _EVAL_353;
  wire [30:0] _EVAL_238;
  wire  _EVAL_552;
  wire [2:0] _EVAL_614;
  wire [3:0] _EVAL_305;
  wire [3:0] _EVAL_513;
  wire  _EVAL_534;
  wire  _EVAL_286;
  wire  _EVAL_373;
  wire  _EVAL_144;
  wire  _EVAL_531;
  wire  _EVAL_453;
  wire  _EVAL_497;
  wire  _EVAL_158;
  wire  _EVAL_421;
  wire  _EVAL_91;
  wire  _EVAL_396;
  wire  _EVAL_347;
  wire  _EVAL_97;
  wire  _EVAL_181;
  wire  _EVAL_443;
  wire  _EVAL_319;
  wire  _EVAL_546;
  wire  _EVAL_45;
  wire  _EVAL_361;
  wire  _EVAL_190;
  wire  _EVAL_109;
  wire  _EVAL_414;
  wire  _EVAL_83;
  wire  _EVAL_482;
  wire  _EVAL_262;
  wire  _EVAL_191;
  wire  _EVAL_375;
  wire  _EVAL_335;
  wire  _EVAL_322;
  wire  _EVAL_206;
  wire  _EVAL_472;
  wire  _EVAL_281;
  wire  _EVAL_454;
  wire  _EVAL_571;
  wire  _EVAL_516;
  wire  _EVAL_120;
  wire  _EVAL_54;
  wire  _EVAL_313;
  wire  _EVAL_189;
  wire  _EVAL_263;
  wire  _EVAL_139;
  wire  _EVAL_417;
  wire  _EVAL_235;
  wire  _EVAL_389;
  wire  _EVAL_393;
  wire  _EVAL_580;
  wire  _EVAL_617;
  wire  _EVAL_404;
  wire  _EVAL_386;
  wire  _EVAL_80;
  wire  _EVAL_426;
  wire  _EVAL_150;
  wire  _EVAL_473;
  wire  _EVAL_465;
  wire  _EVAL_374;
  wire  _EVAL_304;
  wire  _EVAL_558;
  wire  _EVAL_323;
  wire  _EVAL_533;
  wire  _EVAL_557;
  wire  _EVAL_266;
  wire  _EVAL_441;
  wire  _EVAL_394;
  wire  _EVAL_562;
  wire  _EVAL_331;
  wire  _EVAL_519;
  wire  _EVAL_483;
  wire  _EVAL_493;
  wire  _EVAL_589;
  wire [22:0] _EVAL_363;
  wire  _EVAL_532;
  wire  _EVAL_103;
  wire [7:0] _EVAL_411;
  wire [7:0] _EVAL_175;
  wire [5:0] _EVAL_110;
  wire [5:0] _EVAL_567;
  wire [5:0] _EVAL_655;
  wire  _EVAL_650;
  wire [22:0] _EVAL_161;
  wire [7:0] _EVAL_184;
  wire  _EVAL_648;
  wire  _EVAL_642;
  wire  _EVAL_535;
  wire [7:0] _EVAL_164;
  wire [5:0] _EVAL_343;
  wire  _EVAL_341;
  wire  _EVAL_438;
  assign _EVAL_346 = _EVAL_244 == 6'h0;
  assign _EVAL_291 = _EVAL_34[6:3];
  assign _EVAL_282 = _EVAL_291 == 4'h8;
  assign _EVAL_387 = _EVAL_34[2:0];
  assign _EVAL_199 = 3'h1 <= _EVAL_387;
  assign _EVAL_178 = _EVAL_282 & _EVAL_199;
  assign _EVAL_87 = _EVAL_178 & _EVAL_346;
  assign _EVAL_211 = _EVAL_370 | _EVAL_501;
  assign _EVAL_595 = _EVAL_211 | _EVAL_630;
  assign _EVAL_619 = _EVAL_595 | _EVAL_344;
  assign _EVAL_521 = _EVAL_619 | _EVAL_476;
  assign _EVAL_218 = _EVAL_521 | _EVAL_43;
  assign _EVAL_455 = _EVAL_218 | _EVAL_273;
  assign _EVAL_464 = _EVAL_87 & _EVAL_455;
  assign _EVAL_260 = _EVAL_16 ^ 30'h1000;
  assign _EVAL_202 = {1'b0,$signed(_EVAL_260)};
  assign _EVAL_116 = $signed(_EVAL_202) & $signed(31'sh2b105000);
  assign _EVAL_295 = $signed(_EVAL_116);
  assign _EVAL_487 = $signed(_EVAL_295) == $signed(31'sh0);
  assign _EVAL_187 = {{1'd0}, _EVAL_487};
  assign _EVAL_284 = _EVAL_16 ^ 30'h8000000;
  assign _EVAL_84 = {1'b0,$signed(_EVAL_284)};
  assign _EVAL_55 = $signed(_EVAL_84) & $signed(31'sh28000000);
  assign _EVAL_451 = $signed(_EVAL_55);
  assign _EVAL_51 = $signed(_EVAL_451) == $signed(31'sh0);
  assign _EVAL_197 = _EVAL_51 ? 2'h3 : 2'h0;
  assign _EVAL_612 = _EVAL_187 | _EVAL_197;
  assign _EVAL_75 = {{1'd0}, _EVAL_612};
  assign _EVAL_201 = _EVAL_16 ^ 30'h2000000;
  assign _EVAL_520 = {1'b0,$signed(_EVAL_201)};
  assign _EVAL_261 = $signed(_EVAL_520) & $signed(31'sh2b100000);
  assign _EVAL_243 = $signed(_EVAL_261);
  assign _EVAL_74 = $signed(_EVAL_243) == $signed(31'sh0);
  assign _EVAL_222 = _EVAL_74 ? 3'h5 : 3'h0;
  assign _EVAL_114 = _EVAL_75 | _EVAL_222;
  assign _EVAL_149 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_183 = $signed(_EVAL_149) & $signed(31'sh2b105000);
  assign _EVAL_163 = $signed(_EVAL_183);
  assign _EVAL_380 = $signed(_EVAL_163) == $signed(31'sh0);
  assign _EVAL_460 = _EVAL_380 ? 3'h7 : 3'h0;
  assign _EVAL_221 = _EVAL_114 | _EVAL_460;
  assign _EVAL_303 = {{1'd0}, _EVAL_221};
  assign _EVAL_298 = _EVAL_16 ^ 30'h1000000;
  assign _EVAL_593 = {1'b0,$signed(_EVAL_298)};
  assign _EVAL_544 = $signed(_EVAL_593) & $signed(31'sh2b100000);
  assign _EVAL_418 = $signed(_EVAL_544);
  assign _EVAL_446 = $signed(_EVAL_418) == $signed(31'sh0);
  assign _EVAL_79 = _EVAL_446 ? 4'h8 : 4'h0;
  assign _EVAL_400 = _EVAL_303 | _EVAL_79;
  assign _EVAL_409 = _EVAL_16 ^ 30'h1100000;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_409)};
  assign _EVAL_399 = $signed(_EVAL_288) & $signed(31'sh2b104000);
  assign _EVAL_59 = $signed(_EVAL_399);
  assign _EVAL_226 = $signed(_EVAL_59) == $signed(31'sh0);
  assign _EVAL_481 = _EVAL_226 ? 2'h2 : 2'h0;
  assign _EVAL_255 = {{2'd0}, _EVAL_481};
  assign _EVAL_287 = _EVAL_400 | _EVAL_255;
  assign _EVAL_354 = _EVAL_16 ^ 30'h4000;
  assign _EVAL_405 = {1'b0,$signed(_EVAL_354)};
  assign _EVAL_541 = $signed(_EVAL_405) & $signed(31'sh2b105000);
  assign _EVAL_41 = $signed(_EVAL_541);
  assign _EVAL_180 = $signed(_EVAL_41) == $signed(31'sh0);
  assign _EVAL_574 = _EVAL_180 ? 3'h4 : 3'h0;
  assign _EVAL_292 = {{1'd0}, _EVAL_574};
  assign _EVAL_104 = _EVAL_287 | _EVAL_292;
  assign _EVAL_624 = _EVAL_16 ^ 30'h20000000;
  assign _EVAL_352 = {1'b0,$signed(_EVAL_624)};
  assign _EVAL_353 = $signed(_EVAL_352) & $signed(31'sh2b104000);
  assign _EVAL_238 = $signed(_EVAL_353);
  assign _EVAL_552 = $signed(_EVAL_238) == $signed(31'sh0);
  assign _EVAL_614 = _EVAL_552 ? 3'h6 : 3'h0;
  assign _EVAL_305 = {{1'd0}, _EVAL_614};
  assign _EVAL_513 = _EVAL_104 | _EVAL_305;
  assign _EVAL_534 = _EVAL_513 == 4'h0;
  assign _EVAL_286 = _EVAL_503 != _EVAL_513;
  assign _EVAL_373 = _EVAL_534 | _EVAL_286;
  assign _EVAL_144 = _EVAL_464 & _EVAL_373;
  assign _EVAL_531 = _EVAL_291 == 4'h0;
  assign _EVAL_453 = _EVAL_531 & _EVAL_346;
  assign _EVAL_497 = _EVAL_326 | _EVAL_160;
  assign _EVAL_158 = _EVAL_497 | _EVAL_569;
  assign _EVAL_421 = _EVAL_158 | _EVAL_302;
  assign _EVAL_91 = _EVAL_421 | _EVAL_143;
  assign _EVAL_396 = _EVAL_91 | _EVAL_553;
  assign _EVAL_347 = _EVAL_396 | _EVAL_336;
  assign _EVAL_97 = _EVAL_347 | _EVAL_338;
  assign _EVAL_181 = _EVAL_453 & _EVAL_97;
  assign _EVAL_443 = _EVAL_359 != _EVAL_513;
  assign _EVAL_319 = _EVAL_534 | _EVAL_443;
  assign _EVAL_546 = _EVAL_181 & _EVAL_319;
  assign _EVAL_45 = _EVAL_144 | _EVAL_546;
  assign _EVAL_361 = _EVAL_291 == 4'h1;
  assign _EVAL_190 = _EVAL_361 & _EVAL_346;
  assign _EVAL_109 = _EVAL_634 | _EVAL_141;
  assign _EVAL_414 = _EVAL_109 | _EVAL_598;
  assign _EVAL_83 = _EVAL_414 | _EVAL_293;
  assign _EVAL_482 = _EVAL_83 | _EVAL_170;
  assign _EVAL_262 = _EVAL_482 | _EVAL_603;
  assign _EVAL_191 = _EVAL_262 | _EVAL_410;
  assign _EVAL_375 = _EVAL_191 | _EVAL_173;
  assign _EVAL_335 = _EVAL_190 & _EVAL_375;
  assign _EVAL_322 = _EVAL_216 != _EVAL_513;
  assign _EVAL_206 = _EVAL_534 | _EVAL_322;
  assign _EVAL_472 = _EVAL_335 & _EVAL_206;
  assign _EVAL_281 = _EVAL_45 | _EVAL_472;
  assign _EVAL_454 = _EVAL_291 == 4'h2;
  assign _EVAL_571 = _EVAL_454 & _EVAL_346;
  assign _EVAL_516 = _EVAL_556 | _EVAL_99;
  assign _EVAL_120 = _EVAL_516 | _EVAL_296;
  assign _EVAL_54 = _EVAL_120 | _EVAL_490;
  assign _EVAL_313 = _EVAL_54 | _EVAL_511;
  assign _EVAL_189 = _EVAL_313 | _EVAL_623;
  assign _EVAL_263 = _EVAL_189 | _EVAL_204;
  assign _EVAL_139 = _EVAL_263 | _EVAL_90;
  assign _EVAL_417 = _EVAL_571 & _EVAL_139;
  assign _EVAL_235 = _EVAL_49 != _EVAL_513;
  assign _EVAL_389 = _EVAL_534 | _EVAL_235;
  assign _EVAL_393 = _EVAL_417 & _EVAL_389;
  assign _EVAL_580 = _EVAL_281 | _EVAL_393;
  assign _EVAL_617 = _EVAL_291 == 4'h3;
  assign _EVAL_404 = _EVAL_617 & _EVAL_346;
  assign _EVAL_386 = _EVAL_219 | _EVAL_413;
  assign _EVAL_80 = _EVAL_386 | _EVAL_640;
  assign _EVAL_426 = _EVAL_80 | _EVAL_357;
  assign _EVAL_150 = _EVAL_426 | _EVAL_212;
  assign _EVAL_473 = _EVAL_150 | _EVAL_491;
  assign _EVAL_465 = _EVAL_473 | _EVAL_358;
  assign _EVAL_374 = _EVAL_465 | _EVAL_401;
  assign _EVAL_304 = _EVAL_404 & _EVAL_374;
  assign _EVAL_558 = _EVAL_334 != _EVAL_513;
  assign _EVAL_323 = _EVAL_534 | _EVAL_558;
  assign _EVAL_533 = _EVAL_304 & _EVAL_323;
  assign _EVAL_557 = _EVAL_580 | _EVAL_533;
  assign _EVAL_266 = _EVAL_557 == 1'h0;
  assign _EVAL_441 = _EVAL_24 & _EVAL_266;
  assign _EVAL_394 = _EVAL_441 & _EVAL_9;
  assign _EVAL_562 = _EVAL_346 & _EVAL_394;
  assign _EVAL_331 = _EVAL_474 == 6'h0;
  assign _EVAL_519 = _EVAL_2 != 3'h6;
  assign _EVAL_483 = _EVAL_331 & _EVAL_519;
  assign _EVAL_493 = _EVAL_4 & _EVAL_5;
  assign _EVAL_589 = _EVAL_483 & _EVAL_493;
  assign _EVAL_363 = 23'hff << _EVAL_31;
  assign _EVAL_532 = _EVAL[2];
  assign _EVAL_103 = _EVAL_532 == 1'h0;
  assign _EVAL_411 = _EVAL_363[7:0];
  assign _EVAL_175 = ~ _EVAL_411;
  assign _EVAL_110 = _EVAL_175[7:2];
  assign _EVAL_567 = _EVAL_244 - 6'h1;
  assign _EVAL_655 = _EVAL_474 - 6'h1;
  assign _EVAL_650 = _EVAL_394 & _EVAL_454;
  assign _EVAL_161 = 23'hff << _EVAL_40;
  assign _EVAL_184 = _EVAL_161[7:0];
  assign _EVAL_648 = _EVAL_394 & _EVAL_361;
  assign _EVAL_642 = _EVAL_394 & _EVAL_617;
  assign _EVAL_535 = _EVAL_2[0];
  assign _EVAL_164 = ~ _EVAL_184;
  assign _EVAL_343 = _EVAL_164[7:2];
  assign _EVAL_341 = _EVAL_394 & _EVAL_178;
  assign _EVAL_438 = _EVAL_394 & _EVAL_531;
  assign _EVAL_37 = _EVAL_2;
  assign _EVAL_33 = _EVAL_23;
  assign _EVAL_8 = _EVAL_6;
  assign _EVAL_36 = _EVAL_5;
  assign _EVAL_35 = _EVAL_15;
  assign _EVAL_7 = _EVAL_16;
  assign _EVAL_10 = _EVAL_4;
  assign _EVAL_19 = _EVAL;
  assign _EVAL_32 = _EVAL_9 & _EVAL_266;
  assign _EVAL_12 = _EVAL_24 & _EVAL_266;
  assign _EVAL_17 = _EVAL_34;
  assign _EVAL_20 = _EVAL_14;
  assign _EVAL_18 = _EVAL_40;
  assign _EVAL_13 = _EVAL_22;
  assign _EVAL_26 = _EVAL_31;
  assign _EVAL_27 = _EVAL_1;
  assign _EVAL_38 = _EVAL_39;
  assign _EVAL_25 = _EVAL_29;
  assign _EVAL_28 = _EVAL_3;
  assign _EVAL_30 = _EVAL_21;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_43 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_49 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_90 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_99 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_141 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_143 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_160 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_170 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_173 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_204 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_212 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_216 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_219 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_244 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_273 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_293 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_296 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_302 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_326 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_334 = _RAND_19[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_336 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_338 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_344 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_357 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_358 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_359 = _RAND_25[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_370 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_401 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_410 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_413 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_474 = _RAND_30[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_476 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_490 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_491 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_501 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_503 = _RAND_35[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_511 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_553 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_556 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_569 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_598 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_603 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_623 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_630 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_634 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_640 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL_11) begin
      _EVAL_43 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h46 == _EVAL_21) begin
          _EVAL_43 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h46 == _EVAL_34) begin
              _EVAL_43 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h46 == _EVAL_34) begin
            _EVAL_43 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_650) begin
      _EVAL_49 <= _EVAL_513;
    end
    if (_EVAL_11) begin
      _EVAL_90 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h17 == _EVAL_21) begin
          _EVAL_90 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h17 == _EVAL_34) begin
              _EVAL_90 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h17 == _EVAL_34) begin
            _EVAL_90 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_99 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h11 == _EVAL_21) begin
          _EVAL_99 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h11 == _EVAL_34) begin
              _EVAL_99 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h11 == _EVAL_34) begin
            _EVAL_99 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_141 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h9 == _EVAL_21) begin
          _EVAL_141 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h9 == _EVAL_34) begin
              _EVAL_141 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h9 == _EVAL_34) begin
            _EVAL_141 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_143 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h4 == _EVAL_21) begin
          _EVAL_143 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h4 == _EVAL_34) begin
              _EVAL_143 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h4 == _EVAL_34) begin
            _EVAL_143 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_160 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1 == _EVAL_21) begin
          _EVAL_160 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1 == _EVAL_34) begin
              _EVAL_160 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1 == _EVAL_34) begin
            _EVAL_160 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_170 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'hc == _EVAL_21) begin
          _EVAL_170 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'hc == _EVAL_34) begin
              _EVAL_170 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'hc == _EVAL_34) begin
            _EVAL_170 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_173 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'hf == _EVAL_21) begin
          _EVAL_173 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'hf == _EVAL_34) begin
              _EVAL_173 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'hf == _EVAL_34) begin
            _EVAL_173 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_204 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h16 == _EVAL_21) begin
          _EVAL_204 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h16 == _EVAL_34) begin
              _EVAL_204 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h16 == _EVAL_34) begin
            _EVAL_204 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_212 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1c == _EVAL_21) begin
          _EVAL_212 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1c == _EVAL_34) begin
              _EVAL_212 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1c == _EVAL_34) begin
            _EVAL_212 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_648) begin
      _EVAL_216 <= _EVAL_513;
    end
    if (_EVAL_11) begin
      _EVAL_219 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h18 == _EVAL_21) begin
          _EVAL_219 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h18 == _EVAL_34) begin
              _EVAL_219 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h18 == _EVAL_34) begin
            _EVAL_219 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_244 <= 6'h0;
    end else begin
      if (_EVAL_394) begin
        if (_EVAL_346) begin
          if (_EVAL_103) begin
            _EVAL_244 <= _EVAL_110;
          end else begin
            _EVAL_244 <= 6'h0;
          end
        end else begin
          _EVAL_244 <= _EVAL_567;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_273 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h47 == _EVAL_21) begin
          _EVAL_273 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h47 == _EVAL_34) begin
              _EVAL_273 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h47 == _EVAL_34) begin
            _EVAL_273 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_293 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'hb == _EVAL_21) begin
          _EVAL_293 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'hb == _EVAL_34) begin
              _EVAL_293 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'hb == _EVAL_34) begin
            _EVAL_293 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_296 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h12 == _EVAL_21) begin
          _EVAL_296 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h12 == _EVAL_34) begin
              _EVAL_296 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h12 == _EVAL_34) begin
            _EVAL_296 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_302 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h3 == _EVAL_21) begin
          _EVAL_302 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h3 == _EVAL_34) begin
              _EVAL_302 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h3 == _EVAL_34) begin
            _EVAL_302 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_326 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h0 == _EVAL_21) begin
          _EVAL_326 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h0 == _EVAL_34) begin
              _EVAL_326 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h0 == _EVAL_34) begin
            _EVAL_326 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_642) begin
      _EVAL_334 <= _EVAL_513;
    end
    if (_EVAL_11) begin
      _EVAL_336 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h6 == _EVAL_21) begin
          _EVAL_336 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h6 == _EVAL_34) begin
              _EVAL_336 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h6 == _EVAL_34) begin
            _EVAL_336 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_338 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h7 == _EVAL_21) begin
          _EVAL_338 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h7 == _EVAL_34) begin
              _EVAL_338 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h7 == _EVAL_34) begin
            _EVAL_338 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_344 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h44 == _EVAL_21) begin
          _EVAL_344 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h44 == _EVAL_34) begin
              _EVAL_344 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h44 == _EVAL_34) begin
            _EVAL_344 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_357 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1b == _EVAL_21) begin
          _EVAL_357 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1b == _EVAL_34) begin
              _EVAL_357 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1b == _EVAL_34) begin
            _EVAL_357 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_358 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1e == _EVAL_21) begin
          _EVAL_358 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1e == _EVAL_34) begin
              _EVAL_358 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1e == _EVAL_34) begin
            _EVAL_358 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_438) begin
      _EVAL_359 <= _EVAL_513;
    end
    if (_EVAL_11) begin
      _EVAL_370 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h41 == _EVAL_21) begin
          _EVAL_370 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h41 == _EVAL_34) begin
              _EVAL_370 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h41 == _EVAL_34) begin
            _EVAL_370 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_401 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1f == _EVAL_21) begin
          _EVAL_401 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1f == _EVAL_34) begin
              _EVAL_401 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1f == _EVAL_34) begin
            _EVAL_401 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_410 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'he == _EVAL_21) begin
          _EVAL_410 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'he == _EVAL_34) begin
              _EVAL_410 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'he == _EVAL_34) begin
            _EVAL_410 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_413 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h19 == _EVAL_21) begin
          _EVAL_413 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h19 == _EVAL_34) begin
              _EVAL_413 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h19 == _EVAL_34) begin
            _EVAL_413 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_474 <= 6'h0;
    end else begin
      if (_EVAL_493) begin
        if (_EVAL_331) begin
          if (_EVAL_535) begin
            _EVAL_474 <= _EVAL_343;
          end else begin
            _EVAL_474 <= 6'h0;
          end
        end else begin
          _EVAL_474 <= _EVAL_655;
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_476 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h45 == _EVAL_21) begin
          _EVAL_476 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h45 == _EVAL_34) begin
              _EVAL_476 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h45 == _EVAL_34) begin
            _EVAL_476 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_490 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h13 == _EVAL_21) begin
          _EVAL_490 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h13 == _EVAL_34) begin
              _EVAL_490 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h13 == _EVAL_34) begin
            _EVAL_490 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_491 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1d == _EVAL_21) begin
          _EVAL_491 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1d == _EVAL_34) begin
              _EVAL_491 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1d == _EVAL_34) begin
            _EVAL_491 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_501 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h42 == _EVAL_21) begin
          _EVAL_501 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h42 == _EVAL_34) begin
              _EVAL_501 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h42 == _EVAL_34) begin
            _EVAL_501 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_341) begin
      _EVAL_503 <= _EVAL_513;
    end
    if (_EVAL_11) begin
      _EVAL_511 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h14 == _EVAL_21) begin
          _EVAL_511 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h14 == _EVAL_34) begin
              _EVAL_511 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h14 == _EVAL_34) begin
            _EVAL_511 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_553 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h5 == _EVAL_21) begin
          _EVAL_553 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h5 == _EVAL_34) begin
              _EVAL_553 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h5 == _EVAL_34) begin
            _EVAL_553 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_556 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h10 == _EVAL_21) begin
          _EVAL_556 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h10 == _EVAL_34) begin
              _EVAL_556 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h10 == _EVAL_34) begin
            _EVAL_556 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_569 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h2 == _EVAL_21) begin
          _EVAL_569 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h2 == _EVAL_34) begin
              _EVAL_569 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h2 == _EVAL_34) begin
            _EVAL_569 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_598 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'ha == _EVAL_21) begin
          _EVAL_598 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'ha == _EVAL_34) begin
              _EVAL_598 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'ha == _EVAL_34) begin
            _EVAL_598 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_603 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'hd == _EVAL_21) begin
          _EVAL_603 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'hd == _EVAL_34) begin
              _EVAL_603 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'hd == _EVAL_34) begin
            _EVAL_603 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_623 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h15 == _EVAL_21) begin
          _EVAL_623 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h15 == _EVAL_34) begin
              _EVAL_623 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h15 == _EVAL_34) begin
            _EVAL_623 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_630 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h43 == _EVAL_21) begin
          _EVAL_630 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h43 == _EVAL_34) begin
              _EVAL_630 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h43 == _EVAL_34) begin
            _EVAL_630 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_634 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h8 == _EVAL_21) begin
          _EVAL_634 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h8 == _EVAL_34) begin
              _EVAL_634 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h8 == _EVAL_34) begin
            _EVAL_634 <= 1'h1;
          end
        end
      end
    end
    if (_EVAL_11) begin
      _EVAL_640 <= 1'h0;
    end else begin
      if (_EVAL_589) begin
        if (7'h1a == _EVAL_21) begin
          _EVAL_640 <= 1'h0;
        end else begin
          if (_EVAL_562) begin
            if (7'h1a == _EVAL_34) begin
              _EVAL_640 <= 1'h1;
            end
          end
        end
      end else begin
        if (_EVAL_562) begin
          if (7'h1a == _EVAL_34) begin
            _EVAL_640 <= 1'h1;
          end
        end
      end
    end
  end
endmodule
