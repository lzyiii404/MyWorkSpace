//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_142_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [6:0]  _EVAL_2,
  input         _EVAL_3,
  input  [6:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input  [24:0] _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [1:0]  _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_22;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_1;
  reg  _EVAL_39;
  reg [31:0] _RAND_2;
  reg [6:0] _EVAL_70;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_81;
  reg [31:0] _RAND_4;
  reg [72:0] _EVAL_102;
  reg [95:0] _RAND_5;
  reg [6:0] _EVAL_103;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_120;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_155;
  reg [31:0] _RAND_8;
  reg [24:0] _EVAL_179;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_194;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_238;
  reg [31:0] _RAND_11;
  reg  _EVAL_247;
  reg [31:0] _RAND_12;
  reg [2:0] _EVAL_281;
  reg [31:0] _RAND_13;
  reg [2:0] _EVAL_305;
  reg [31:0] _RAND_14;
  reg [3:0] _EVAL_311;
  reg [31:0] _RAND_15;
  reg [31:0] _EVAL_316;
  reg [31:0] _RAND_16;
  wire  _EVAL_329;
  wire  _EVAL_234;
  wire  _EVAL_64;
  wire [1:0] _EVAL_38;
  wire [1:0] _EVAL_63;
  wire  _EVAL_26;
  wire  _EVAL_303;
  wire  _EVAL_324;
  wire  _EVAL_211;
  wire  _EVAL_304;
  wire  _EVAL_322;
  wire  _EVAL_173;
  wire  _EVAL_306;
  wire  _EVAL_223;
  wire  _EVAL_167;
  wire  _EVAL_145;
  wire  _EVAL_197;
  wire  _EVAL_65;
  wire  _EVAL_54;
  wire  _EVAL_108;
  wire  _EVAL_37;
  wire  _EVAL_239;
  wire  _EVAL_127;
  wire  _EVAL_98;
  wire  _EVAL_86;
  wire  _EVAL_168;
  wire  _EVAL_228;
  wire [3:0] _EVAL_106;
  wire [3:0] _EVAL_283;
  wire [3:0] _EVAL_34;
  wire  _EVAL_93;
  wire [12:0] _EVAL_48;
  wire [5:0] _EVAL_330;
  wire [5:0] _EVAL_299;
  wire [24:0] _EVAL_166;
  wire [24:0] _EVAL_66;
  wire  _EVAL_140;
  wire  _EVAL_58;
  wire  _EVAL_163;
  wire  _EVAL_72;
  wire  _EVAL_325;
  wire  _EVAL_112;
  wire  _EVAL_31;
  wire  _EVAL_73;
  wire  _EVAL_24;
  wire  _EVAL_236;
  wire  _EVAL_191;
  wire  _EVAL_208;
  wire  _EVAL_180;
  wire  _EVAL_71;
  wire  _EVAL_35;
  wire [3:0] _EVAL_159;
  wire  _EVAL_258;
  wire [2:0] _EVAL_138;
  wire  _EVAL_130;
  wire  _EVAL_94;
  wire  _EVAL_121;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_294;
  wire  _EVAL_69;
  wire [12:0] _EVAL_288;
  wire [5:0] _EVAL_40;
  wire [5:0] _EVAL_263;
  wire  _EVAL_276;
  wire  _EVAL_185;
  wire  _EVAL_286;
  wire [24:0] _EVAL_251;
  wire [25:0] _EVAL_217;
  wire [25:0] _EVAL_91;
  wire [25:0] _EVAL_90;
  wire  _EVAL_111;
  wire  _EVAL_273;
  wire  _EVAL_218;
  wire  _EVAL_147;
  wire [24:0] _EVAL_157;
  wire [25:0] _EVAL_23;
  wire [25:0] _EVAL_55;
  wire [25:0] _EVAL_242;
  wire  _EVAL_321;
  wire  _EVAL_207;
  wire  _EVAL_181;
  wire  _EVAL_57;
  wire  _EVAL_323;
  wire  _EVAL_328;
  wire  _EVAL_119;
  wire  _EVAL_265;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_74;
  wire  _EVAL_332;
  wire  _EVAL_293;
  wire  _EVAL_78;
  wire [127:0] _EVAL_314;
  wire [127:0] _EVAL_287;
  wire [72:0] _EVAL_60;
  wire  _EVAL_25;
  wire  _EVAL_53;
  wire  _EVAL_320;
  wire  _EVAL_260;
  wire  _EVAL_213;
  wire  _EVAL_227;
  wire  _EVAL_115;
  wire  _EVAL_96;
  wire  _EVAL_221;
  wire  _EVAL_266;
  wire  _EVAL_315;
  wire [127:0] _EVAL_136;
  wire [127:0] _EVAL_156;
  wire [72:0] _EVAL_170;
  wire  _EVAL_250;
  wire  _EVAL_224;
  wire  _EVAL_129;
  wire  _EVAL_19;
  wire  _EVAL_301;
  wire  _EVAL_30;
  wire  _EVAL_201;
  wire  _EVAL_319;
  wire [3:0] _EVAL_226;
  wire  _EVAL_20;
  wire  _EVAL_302;
  wire  _EVAL_62;
  wire  _EVAL_79;
  wire  _EVAL_285;
  wire  _EVAL_212;
  wire  _EVAL_203;
  wire  _EVAL_259;
  wire  _EVAL_313;
  wire  _EVAL_152;
  wire  _EVAL_45;
  wire  _EVAL_125;
  wire  _EVAL_134;
  wire  _EVAL_249;
  wire  _EVAL_82;
  wire  _EVAL_177;
  wire  _EVAL_36;
  wire  _EVAL_97;
  wire  _EVAL_171;
  wire  _EVAL_244;
  wire  _EVAL_327;
  wire  _EVAL_296;
  wire [3:0] _EVAL_278;
  wire  _EVAL_76;
  wire  _EVAL_289;
  wire  _EVAL_231;
  wire  _EVAL_75;
  wire  _EVAL_150;
  wire  _EVAL_205;
  wire  _EVAL_220;
  wire [72:0] _EVAL_252;
  wire [72:0] _EVAL_33;
  wire  _EVAL_295;
  wire  _EVAL_80;
  wire  _EVAL_279;
  wire  _EVAL_270;
  wire [3:0] _EVAL_269;
  wire [3:0] _EVAL_149;
  wire [3:0] _EVAL_246;
  wire  _EVAL_162;
  wire  _EVAL_50;
  wire  _EVAL_307;
  wire  _EVAL_196;
  wire [2:0] _EVAL_165;
  wire  _EVAL_104;
  wire  _EVAL_214;
  wire  _EVAL_160;
  wire  _EVAL_215;
  wire [3:0] _EVAL_114;
  wire  _EVAL_189;
  wire  _EVAL_186;
  wire  _EVAL_209;
  wire  _EVAL_183;
  wire  _EVAL_318;
  wire  _EVAL_92;
  wire  _EVAL_326;
  wire  _EVAL_154;
  wire  _EVAL_241;
  wire  _EVAL_174;
  wire  _EVAL_216;
  wire  _EVAL_240;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_176;
  wire  _EVAL_255;
  wire  _EVAL_253;
  wire  _EVAL_200;
  wire  _EVAL_46;
  wire [3:0] _EVAL_133;
  wire  _EVAL_158;
  wire  _EVAL_188;
  wire  _EVAL_184;
  wire  _EVAL_195;
  wire  _EVAL_146;
  wire  _EVAL_67;
  wire  _EVAL_256;
  wire  _EVAL_131;
  wire  _EVAL_232;
  wire  _EVAL_190;
  wire  _EVAL_153;
  wire  _EVAL_132;
  wire  _EVAL_110;
  wire  _EVAL_109;
  wire  _EVAL_172;
  wire  _EVAL_187;
  wire [3:0] _EVAL_116;
  wire  _EVAL_47;
  wire  _EVAL_300;
  wire  _EVAL_135;
  wire  _EVAL_123;
  wire  _EVAL_267;
  wire  _EVAL_128;
  wire  _EVAL_137;
  wire  _EVAL_245;
  wire  _EVAL_192;
  wire  _EVAL_59;
  wire  _EVAL_113;
  wire [31:0] _EVAL_141;
  wire  _EVAL_284;
  wire  _EVAL_169;
  wire  _EVAL_237;
  wire  _EVAL_88;
  wire  _EVAL_41;
  wire  _EVAL_83;
  wire  _EVAL_124;
  wire  _EVAL_117;
  wire  _EVAL_175;
  wire  _EVAL_277;
  wire  _EVAL_87;
  wire  _EVAL_233;
  wire  _EVAL_42;
  wire  _EVAL_222;
  wire  _EVAL_243;
  wire  _EVAL_290;
  wire [72:0] _EVAL_95;
  wire  _EVAL_317;
  wire  _EVAL_84;
  wire  _EVAL_254;
  wire  _EVAL_105;
  wire [72:0] _EVAL_99;
  wire  _EVAL_275;
  wire  _EVAL_101;
  wire  _EVAL_248;
  wire  _EVAL_139;
  wire  _EVAL_122;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_49;
  wire  _EVAL_268;
  wire  _EVAL_219;
  wire  _EVAL_182;
  wire  _EVAL_100;
  wire  _EVAL_202;
  wire [72:0] _EVAL_225;
  wire  _EVAL_229;
  wire  _EVAL_126;
  wire  _EVAL_21;
  wire  _EVAL_144;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_291;
  wire [72:0] _EVAL_68;
  wire  _EVAL_77;
  wire  _EVAL_143;
  wire  _EVAL_309;
  wire  _EVAL_235;
  wire  _EVAL_331;
  wire  _EVAL_148;
  wire  _EVAL_178;
  wire  _EVAL_308;
  wire  _EVAL_151;
  wire  _EVAL_193;
  wire  _EVAL_161;
  wire  _EVAL_27;
  wire  _EVAL_264;
  wire  _EVAL_257;
  wire  _EVAL_230;
  wire  _EVAL_29;
  wire  _EVAL_292;
  wire  _EVAL_280;
  wire  _EVAL_61;
  wire  _EVAL_118;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_329 = _EVAL_6 == _EVAL_32;
  assign _EVAL_234 = _EVAL_15 >= 3'h2;
  assign _EVAL_64 = _EVAL_15[0];
  assign _EVAL_38 = 2'h1 << _EVAL_64;
  assign _EVAL_63 = _EVAL_38 | 2'h1;
  assign _EVAL_26 = _EVAL_63[1];
  assign _EVAL_303 = _EVAL_11[1];
  assign _EVAL_324 = _EVAL_26 & _EVAL_303;
  assign _EVAL_211 = _EVAL_234 | _EVAL_324;
  assign _EVAL_304 = _EVAL_63[0];
  assign _EVAL_322 = _EVAL_11[0];
  assign _EVAL_173 = _EVAL_303 & _EVAL_322;
  assign _EVAL_306 = _EVAL_304 & _EVAL_173;
  assign _EVAL_223 = _EVAL_211 | _EVAL_306;
  assign _EVAL_167 = _EVAL_322 == 1'h0;
  assign _EVAL_145 = _EVAL_303 & _EVAL_167;
  assign _EVAL_197 = _EVAL_304 & _EVAL_145;
  assign _EVAL_65 = _EVAL_211 | _EVAL_197;
  assign _EVAL_54 = _EVAL_303 == 1'h0;
  assign _EVAL_108 = _EVAL_26 & _EVAL_54;
  assign _EVAL_37 = _EVAL_234 | _EVAL_108;
  assign _EVAL_239 = _EVAL_54 & _EVAL_322;
  assign _EVAL_127 = _EVAL_304 & _EVAL_239;
  assign _EVAL_98 = _EVAL_37 | _EVAL_127;
  assign _EVAL_86 = _EVAL_54 & _EVAL_167;
  assign _EVAL_168 = _EVAL_304 & _EVAL_86;
  assign _EVAL_228 = _EVAL_37 | _EVAL_168;
  assign _EVAL_106 = {_EVAL_223,_EVAL_65,_EVAL_98,_EVAL_228};
  assign _EVAL_283 = ~ _EVAL_106;
  assign _EVAL_34 = _EVAL_9 & _EVAL_283;
  assign _EVAL_93 = _EVAL_34 == 4'h0;
  assign _EVAL_48 = 13'h3f << _EVAL_15;
  assign _EVAL_330 = _EVAL_48[5:0];
  assign _EVAL_299 = ~ _EVAL_330;
  assign _EVAL_166 = {{19'd0}, _EVAL_299};
  assign _EVAL_66 = _EVAL_11 & _EVAL_166;
  assign _EVAL_140 = _EVAL_66 == 25'h0;
  assign _EVAL_58 = _EVAL_140 | _EVAL_18;
  assign _EVAL_163 = _EVAL_3 == 1'h0;
  assign _EVAL_72 = _EVAL_163 | _EVAL_7;
  assign _EVAL_325 = _EVAL_72 | _EVAL_18;
  assign _EVAL_112 = _EVAL_325 == 1'h0;
  assign _EVAL_31 = _EVAL_15 == _EVAL_22;
  assign _EVAL_73 = _EVAL_31 | _EVAL_18;
  assign _EVAL_24 = _EVAL != 3'h0;
  assign _EVAL_236 = _EVAL_194 == 4'h0;
  assign _EVAL_191 = _EVAL_236 == 1'h0;
  assign _EVAL_208 = _EVAL_5 & _EVAL_191;
  assign _EVAL_180 = _EVAL_2 == 7'h48;
  assign _EVAL_71 = _EVAL_2 == 7'h40;
  assign _EVAL_35 = _EVAL_180 | _EVAL_71;
  assign _EVAL_159 = _EVAL_2[6:3];
  assign _EVAL_258 = _EVAL_159 == 4'h8;
  assign _EVAL_138 = _EVAL_2[2:0];
  assign _EVAL_130 = 3'h1 <= _EVAL_138;
  assign _EVAL_94 = _EVAL_258 & _EVAL_130;
  assign _EVAL_121 = _EVAL_35 | _EVAL_94;
  assign _EVAL_271 = _EVAL_2 == 7'h20;
  assign _EVAL_272 = _EVAL_121 | _EVAL_271;
  assign _EVAL_294 = _EVAL_159 == 4'h0;
  assign _EVAL_69 = _EVAL_272 | _EVAL_294;
  assign _EVAL_288 = 13'h3f << _EVAL_6;
  assign _EVAL_40 = _EVAL_288[5:0];
  assign _EVAL_263 = ~ _EVAL_40;
  assign _EVAL_276 = _EVAL_311 == 4'h0;
  assign _EVAL_185 = _EVAL_276 == 1'h0;
  assign _EVAL_286 = _EVAL_12 & _EVAL_185;
  assign _EVAL_251 = _EVAL_11 ^ 25'h1800000;
  assign _EVAL_217 = {1'b0,$signed(_EVAL_251)};
  assign _EVAL_91 = $signed(_EVAL_217) & $signed(-26'sh8000);
  assign _EVAL_90 = $signed(_EVAL_91);
  assign _EVAL_111 = $signed(_EVAL_90) == $signed(26'sh0);
  assign _EVAL_273 = _EVAL_1 <= 3'h6;
  assign _EVAL_218 = _EVAL_273 | _EVAL_18;
  assign _EVAL_147 = _EVAL_15 <= 3'h6;
  assign _EVAL_157 = _EVAL_11 ^ 25'h1900000;
  assign _EVAL_23 = {1'b0,$signed(_EVAL_157)};
  assign _EVAL_55 = $signed(_EVAL_23) & $signed(-26'sh2000);
  assign _EVAL_242 = $signed(_EVAL_55);
  assign _EVAL_321 = $signed(_EVAL_242) == $signed(26'sh0);
  assign _EVAL_207 = _EVAL_111 | _EVAL_321;
  assign _EVAL_181 = _EVAL_147 & _EVAL_207;
  assign _EVAL_57 = _EVAL_181 | _EVAL_18;
  assign _EVAL_323 = _EVAL_57 == 1'h0;
  assign _EVAL_328 = _EVAL_93 | _EVAL_18;
  assign _EVAL_119 = _EVAL_16 == 2'h0;
  assign _EVAL_265 = _EVAL_119 | _EVAL_18;
  assign _EVAL_261 = plusarg_reader_out == 32'h0;
  assign _EVAL_262 = _EVAL <= 3'h4;
  assign _EVAL_74 = _EVAL_262 | _EVAL_18;
  assign _EVAL_332 = _EVAL_10 & _EVAL_5;
  assign _EVAL_293 = _EVAL_155 == 4'h0;
  assign _EVAL_78 = _EVAL_332 & _EVAL_293;
  assign _EVAL_314 = 128'h1 << _EVAL_2;
  assign _EVAL_287 = _EVAL_78 ? _EVAL_314 : 128'h0;
  assign _EVAL_60 = _EVAL_287[72:0];
  assign _EVAL_25 = _EVAL_329 | _EVAL_18;
  assign _EVAL_53 = _EVAL_25 == 1'h0;
  assign _EVAL_320 = _EVAL_13 == 3'h2;
  assign _EVAL_260 = _EVAL_5 & _EVAL_320;
  assign _EVAL_213 = _EVAL_4 == 7'h20;
  assign _EVAL_227 = _EVAL_17 & _EVAL_12;
  assign _EVAL_115 = _EVAL_120 == 4'h0;
  assign _EVAL_96 = _EVAL_227 & _EVAL_115;
  assign _EVAL_221 = _EVAL_1 == 3'h6;
  assign _EVAL_266 = _EVAL_221 == 1'h0;
  assign _EVAL_315 = _EVAL_96 & _EVAL_266;
  assign _EVAL_136 = 128'h1 << _EVAL_4;
  assign _EVAL_156 = _EVAL_315 ? _EVAL_136 : 128'h0;
  assign _EVAL_170 = _EVAL_156[72:0];
  assign _EVAL_250 = _EVAL_60 != _EVAL_170;
  assign _EVAL_224 = _EVAL_60 != 73'h0;
  assign _EVAL_129 = _EVAL_224 == 1'h0;
  assign _EVAL_19 = _EVAL_250 | _EVAL_129;
  assign _EVAL_301 = _EVAL_19 | _EVAL_18;
  assign _EVAL_30 = _EVAL_1 == _EVAL_281;
  assign _EVAL_201 = _EVAL_30 | _EVAL_18;
  assign _EVAL_319 = _EVAL_4 == 7'h48;
  assign _EVAL_226 = _EVAL_311 - 4'h1;
  assign _EVAL_20 = _EVAL_13[2];
  assign _EVAL_302 = _EVAL_3 == _EVAL_39;
  assign _EVAL_62 = _EVAL_302 | _EVAL_18;
  assign _EVAL_79 = _EVAL == 3'h0;
  assign _EVAL_285 = _EVAL_79 | _EVAL_18;
  assign _EVAL_212 = _EVAL_285 == 1'h0;
  assign _EVAL_203 = _EVAL_11 == _EVAL_179;
  assign _EVAL_259 = _EVAL_203 | _EVAL_18;
  assign _EVAL_313 = _EVAL_62 == 1'h0;
  assign _EVAL_152 = _EVAL_0 == _EVAL_247;
  assign _EVAL_45 = _EVAL_152 | _EVAL_18;
  assign _EVAL_125 = _EVAL_45 == 1'h0;
  assign _EVAL_134 = _EVAL_159 == 4'h1;
  assign _EVAL_249 = _EVAL_69 | _EVAL_134;
  assign _EVAL_82 = _EVAL_159 == 4'h2;
  assign _EVAL_177 = _EVAL_249 | _EVAL_82;
  assign _EVAL_36 = _EVAL_159 == 4'h3;
  assign _EVAL_97 = _EVAL_177 | _EVAL_36;
  assign _EVAL_171 = _EVAL_97 | _EVAL_18;
  assign _EVAL_244 = _EVAL_4 == _EVAL_70;
  assign _EVAL_327 = _EVAL_244 | _EVAL_18;
  assign _EVAL_296 = _EVAL_1[0];
  assign _EVAL_278 = _EVAL_263[5:2];
  assign _EVAL_76 = _EVAL_13 == _EVAL_305;
  assign _EVAL_289 = _EVAL_76 | _EVAL_18;
  assign _EVAL_231 = _EVAL_8 == 1'h0;
  assign _EVAL_75 = _EVAL_231 | _EVAL_18;
  assign _EVAL_150 = _EVAL_75 == 1'h0;
  assign _EVAL_205 = _EVAL_7 == 1'h0;
  assign _EVAL_220 = _EVAL_205 | _EVAL_18;
  assign _EVAL_252 = _EVAL_60 | _EVAL_102;
  assign _EVAL_33 = _EVAL_252 >> _EVAL_4;
  assign _EVAL_295 = _EVAL_33[0];
  assign _EVAL_80 = _EVAL_1 == 3'h2;
  assign _EVAL_279 = _EVAL_316 < plusarg_reader_out;
  assign _EVAL_270 = _EVAL_20 == 1'h0;
  assign _EVAL_269 = _EVAL_299[5:2];
  assign _EVAL_149 = _EVAL_194 - 4'h1;
  assign _EVAL_246 = _EVAL_4[6:3];
  assign _EVAL_162 = _EVAL_246 == 4'h8;
  assign _EVAL_50 = _EVAL_6 >= 3'h2;
  assign _EVAL_307 = _EVAL_4 == 7'h40;
  assign _EVAL_196 = _EVAL_319 | _EVAL_307;
  assign _EVAL_165 = _EVAL_4[2:0];
  assign _EVAL_104 = 3'h1 <= _EVAL_165;
  assign _EVAL_214 = _EVAL_162 & _EVAL_104;
  assign _EVAL_160 = _EVAL_196 | _EVAL_214;
  assign _EVAL_215 = _EVAL_160 | _EVAL_213;
  assign _EVAL_114 = _EVAL_120 - 4'h1;
  assign _EVAL_189 = _EVAL_301 == 1'h0;
  assign _EVAL_186 = _EVAL_246 == 4'h0;
  assign _EVAL_209 = _EVAL_215 | _EVAL_186;
  assign _EVAL_183 = _EVAL_246 == 4'h1;
  assign _EVAL_318 = _EVAL_209 | _EVAL_183;
  assign _EVAL_92 = _EVAL_246 == 4'h2;
  assign _EVAL_326 = _EVAL_318 | _EVAL_92;
  assign _EVAL_154 = _EVAL_246 == 4'h3;
  assign _EVAL_241 = _EVAL_326 | _EVAL_154;
  assign _EVAL_174 = _EVAL_241 | _EVAL_18;
  assign _EVAL_216 = _EVAL_174 == 1'h0;
  assign _EVAL_240 = _EVAL_102 != 73'h0;
  assign _EVAL_198 = _EVAL_240 == 1'h0;
  assign _EVAL_199 = _EVAL_198 | _EVAL_261;
  assign _EVAL_176 = _EVAL_199 | _EVAL_279;
  assign _EVAL_255 = _EVAL_176 | _EVAL_18;
  assign _EVAL_253 = _EVAL_220 == 1'h0;
  assign _EVAL_200 = _EVAL_13 == 3'h6;
  assign _EVAL_46 = _EVAL_1 == 3'h5;
  assign _EVAL_133 = ~ _EVAL_9;
  assign _EVAL_158 = _EVAL_133 == 4'h0;
  assign _EVAL_188 = _EVAL_158 | _EVAL_18;
  assign _EVAL_184 = _EVAL_188 == 1'h0;
  assign _EVAL_195 = _EVAL <= 3'h3;
  assign _EVAL_146 = _EVAL_195 | _EVAL_18;
  assign _EVAL_67 = _EVAL_16 == _EVAL_238;
  assign _EVAL_256 = _EVAL_67 | _EVAL_18;
  assign _EVAL_131 = _EVAL_256 == 1'h0;
  assign _EVAL_232 = 3'h6 == _EVAL_15;
  assign _EVAL_190 = _EVAL_71 ? _EVAL_232 : 1'h0;
  assign _EVAL_153 = _EVAL_190 | _EVAL_18;
  assign _EVAL_132 = _EVAL_153 == 1'h0;
  assign _EVAL_110 = _EVAL_15 <= 3'h2;
  assign _EVAL_109 = _EVAL_110 & _EVAL_321;
  assign _EVAL_172 = _EVAL_109 | _EVAL_18;
  assign _EVAL_187 = _EVAL_58 == 1'h0;
  assign _EVAL_116 = _EVAL_155 - 4'h1;
  assign _EVAL_47 = _EVAL_1 == 3'h0;
  assign _EVAL_300 = _EVAL_1 == 3'h4;
  assign _EVAL_135 = _EVAL_13 == 3'h3;
  assign _EVAL_123 = _EVAL == _EVAL_81;
  assign _EVAL_267 = _EVAL_1 == 3'h1;
  assign _EVAL_128 = _EVAL_12 & _EVAL_267;
  assign _EVAL_137 = _EVAL_5 & _EVAL_200;
  assign _EVAL_245 = _EVAL_13 == 3'h7;
  assign _EVAL_192 = _EVAL_13 == 3'h0;
  assign _EVAL_59 = _EVAL_12 & _EVAL_47;
  assign _EVAL_113 = _EVAL_16 != 2'h2;
  assign _EVAL_141 = _EVAL_316 + 32'h1;
  assign _EVAL_284 = _EVAL_163 | _EVAL_18;
  assign _EVAL_169 = _EVAL_18 == 1'h0;
  assign _EVAL_237 = _EVAL_13 == 3'h1;
  assign _EVAL_88 = _EVAL_234 | _EVAL_18;
  assign _EVAL_41 = _EVAL_123 | _EVAL_18;
  assign _EVAL_83 = _EVAL_41 == 1'h0;
  assign _EVAL_124 = _EVAL <= 3'h2;
  assign _EVAL_117 = _EVAL_124 | _EVAL_18;
  assign _EVAL_175 = _EVAL_117 == 1'h0;
  assign _EVAL_277 = _EVAL_12 & _EVAL_300;
  assign _EVAL_87 = _EVAL_9 == _EVAL_106;
  assign _EVAL_233 = _EVAL_87 | _EVAL_18;
  assign _EVAL_42 = _EVAL_233 == 1'h0;
  assign _EVAL_222 = _EVAL_50 | _EVAL_18;
  assign _EVAL_243 = _EVAL_73 == 1'h0;
  assign _EVAL_290 = _EVAL_24 | _EVAL_18;
  assign _EVAL_95 = _EVAL_102 >> _EVAL_2;
  assign _EVAL_317 = _EVAL_95[0];
  assign _EVAL_84 = _EVAL_317 == 1'h0;
  assign _EVAL_254 = _EVAL_5 & _EVAL_245;
  assign _EVAL_105 = _EVAL_327 == 1'h0;
  assign _EVAL_99 = _EVAL_102 | _EVAL_60;
  assign _EVAL_275 = _EVAL_16 <= 2'h2;
  assign _EVAL_101 = _EVAL_259 == 1'h0;
  assign _EVAL_248 = _EVAL_113 | _EVAL_18;
  assign _EVAL_139 = _EVAL_5 & _EVAL_135;
  assign _EVAL_122 = _EVAL_2 == _EVAL_103;
  assign _EVAL_43 = _EVAL_122 | _EVAL_18;
  assign _EVAL_44 = _EVAL_43 == 1'h0;
  assign _EVAL_49 = _EVAL_5 & _EVAL_237;
  assign _EVAL_268 = _EVAL_255 == 1'h0;
  assign _EVAL_219 = _EVAL_171 == 1'h0;
  assign _EVAL_182 = _EVAL_146 == 1'h0;
  assign _EVAL_100 = _EVAL_218 == 1'h0;
  assign _EVAL_202 = _EVAL_84 | _EVAL_18;
  assign _EVAL_225 = ~ _EVAL_170;
  assign _EVAL_229 = _EVAL_295 | _EVAL_18;
  assign _EVAL_126 = _EVAL_229 == 1'h0;
  assign _EVAL_21 = _EVAL_202 == 1'h0;
  assign _EVAL_144 = _EVAL_328 == 1'h0;
  assign _EVAL_297 = _EVAL_201 == 1'h0;
  assign _EVAL_298 = _EVAL_5 & _EVAL_192;
  assign _EVAL_291 = _EVAL_332 | _EVAL_227;
  assign _EVAL_68 = _EVAL_99 & _EVAL_225;
  assign _EVAL_77 = _EVAL_275 | _EVAL_18;
  assign _EVAL_143 = _EVAL_265 == 1'h0;
  assign _EVAL_309 = _EVAL_74 == 1'h0;
  assign _EVAL_235 = _EVAL_227 & _EVAL_276;
  assign _EVAL_331 = _EVAL_172 == 1'h0;
  assign _EVAL_148 = _EVAL_12 & _EVAL_221;
  assign _EVAL_178 = _EVAL_332 & _EVAL_236;
  assign _EVAL_308 = _EVAL_13 == 3'h5;
  assign _EVAL_151 = _EVAL_290 == 1'h0;
  assign _EVAL_193 = _EVAL_5 & _EVAL_308;
  assign _EVAL_161 = _EVAL_222 == 1'h0;
  assign _EVAL_27 = _EVAL_13 == 3'h4;
  assign _EVAL_264 = _EVAL_289 == 1'h0;
  assign _EVAL_257 = _EVAL_77 == 1'h0;
  assign _EVAL_230 = _EVAL_88 == 1'h0;
  assign _EVAL_29 = _EVAL_12 & _EVAL_80;
  assign _EVAL_292 = _EVAL_248 == 1'h0;
  assign _EVAL_280 = _EVAL_284 == 1'h0;
  assign _EVAL_61 = _EVAL_5 & _EVAL_27;
  assign _EVAL_118 = _EVAL_12 & _EVAL_46;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_32 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_70 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_81 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  _EVAL_102 = _RAND_5[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_103 = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_120 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_155 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_179 = _RAND_9[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_194 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_238 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_247 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_281 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_305 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_311 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_316 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL_178) begin
      _EVAL_22 <= _EVAL_15;
    end
    if (_EVAL_235) begin
      _EVAL_32 <= _EVAL_6;
    end
    if (_EVAL_235) begin
      _EVAL_39 <= _EVAL_3;
    end
    if (_EVAL_235) begin
      _EVAL_70 <= _EVAL_4;
    end
    if (_EVAL_178) begin
      _EVAL_81 <= _EVAL;
    end
    if (_EVAL_18) begin
      _EVAL_102 <= 73'h0;
    end else begin
      _EVAL_102 <= _EVAL_68;
    end
    if (_EVAL_178) begin
      _EVAL_103 <= _EVAL_2;
    end
    if (_EVAL_18) begin
      _EVAL_120 <= 4'h0;
    end else begin
      if (_EVAL_227) begin
        if (_EVAL_115) begin
          if (_EVAL_296) begin
            _EVAL_120 <= _EVAL_278;
          end else begin
            _EVAL_120 <= 4'h0;
          end
        end else begin
          _EVAL_120 <= _EVAL_114;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_155 <= 4'h0;
    end else begin
      if (_EVAL_332) begin
        if (_EVAL_293) begin
          if (_EVAL_270) begin
            _EVAL_155 <= _EVAL_269;
          end else begin
            _EVAL_155 <= 4'h0;
          end
        end else begin
          _EVAL_155 <= _EVAL_116;
        end
      end
    end
    if (_EVAL_178) begin
      _EVAL_179 <= _EVAL_11;
    end
    if (_EVAL_18) begin
      _EVAL_194 <= 4'h0;
    end else begin
      if (_EVAL_332) begin
        if (_EVAL_236) begin
          if (_EVAL_270) begin
            _EVAL_194 <= _EVAL_269;
          end else begin
            _EVAL_194 <= 4'h0;
          end
        end else begin
          _EVAL_194 <= _EVAL_149;
        end
      end
    end
    if (_EVAL_235) begin
      _EVAL_238 <= _EVAL_16;
    end
    if (_EVAL_235) begin
      _EVAL_247 <= _EVAL_0;
    end
    if (_EVAL_235) begin
      _EVAL_281 <= _EVAL_1;
    end
    if (_EVAL_178) begin
      _EVAL_305 <= _EVAL_13;
    end
    if (_EVAL_18) begin
      _EVAL_311 <= 4'h0;
    end else begin
      if (_EVAL_227) begin
        if (_EVAL_276) begin
          if (_EVAL_296) begin
            _EVAL_311 <= _EVAL_278;
          end else begin
            _EVAL_311 <= 4'h0;
          end
        end else begin
          _EVAL_311 <= _EVAL_226;
        end
      end
    end
    if (_EVAL_18) begin
      _EVAL_316 <= 32'h0;
    end else begin
      if (_EVAL_291) begin
        _EVAL_316 <= 32'h0;
      end else begin
        _EVAL_316 <= _EVAL_141;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5abcc2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1b7c7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(267fcd32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d00a0395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58c24c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59e8f6fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4ebd854)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1d0a2a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb42fc84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccc55f4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97fe61d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35ce1840)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccfa8fef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e91edbfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2ad3224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(993f0c13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f4a7358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1668dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348db9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50419eed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a013e7df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c18c4bcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77a284d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1e8ff24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef7b9854)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(305d6e18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e0566ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3199ff1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1540c7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7958049d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4af4dc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(739bd5f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a340a62b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7a9639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a578362a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(529c4971)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b372fd4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7fd8230)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49dfc7d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6736a5c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c4788a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5cf91c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50d53d99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4240400)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f83f7421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92f8741e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4df9a90c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(676c0f75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(982367c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2adb4555)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91572910)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b22c503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae2e2697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(280bff8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4df0be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5ee0245)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77618a7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce586b64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c11333a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9e3d679)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daab676a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5cd8124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f431d29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eefb4a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7d23788)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c2cd585)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_331) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b6cf57c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5151ffc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(febfa2dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ea74a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c00d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81ad4dea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b07184b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de8e85eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93801e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79d0c18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c9fac93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb58fff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(940f913a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a48bd5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903d4557)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(774c7bc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(732cd825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f67241b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(980863e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cead48d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e87633)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea5f76d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab5b64b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f55b33df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c4b3860)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87199c6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72329dbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4015c7cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba19b907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
