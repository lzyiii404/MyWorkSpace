//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_111_assert(
  input  [2:0]  _EVAL,
  input  [6:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [6:0]  _EVAL_14,
  input  [1:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [29:0] _EVAL_18
);
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_20;
  reg [31:0] _RAND_0;
  reg [72:0] _EVAL_26;
  reg [95:0] _RAND_1;
  reg [5:0] _EVAL_59;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_112;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_167;
  reg [31:0] _RAND_4;
  reg [1:0] _EVAL_187;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_189;
  reg [31:0] _RAND_6;
  reg  _EVAL_207;
  reg [31:0] _RAND_7;
  reg [6:0] _EVAL_241;
  reg [31:0] _RAND_8;
  reg [6:0] _EVAL_242;
  reg [31:0] _RAND_9;
  reg  _EVAL_271;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_273;
  reg [31:0] _RAND_11;
  reg [5:0] _EVAL_278;
  reg [31:0] _RAND_12;
  reg [29:0] _EVAL_284;
  reg [31:0] _RAND_13;
  reg [5:0] _EVAL_304;
  reg [31:0] _RAND_14;
  reg [3:0] _EVAL_331;
  reg [31:0] _RAND_15;
  reg [5:0] _EVAL_339;
  reg [31:0] _RAND_16;
  wire  _EVAL_357;
  wire  _EVAL_309;
  wire  _EVAL_51;
  wire  _EVAL_154;
  wire  _EVAL_58;
  wire  _EVAL_288;
  wire  _EVAL_160;
  wire [72:0] _EVAL_292;
  wire  _EVAL_316;
  wire  _EVAL_127;
  wire  _EVAL_260;
  wire  _EVAL_78;
  wire  _EVAL_206;
  wire  _EVAL_291;
  wire [29:0] _EVAL_194;
  wire [30:0] _EVAL_131;
  wire [30:0] _EVAL_140;
  wire [30:0] _EVAL_86;
  wire  _EVAL_252;
  wire  _EVAL_62;
  wire  _EVAL_145;
  wire  _EVAL_36;
  wire  _EVAL_176;
  wire  _EVAL_30;
  wire  _EVAL_214;
  wire  _EVAL_138;
  wire  _EVAL_74;
  wire  _EVAL_352;
  wire  _EVAL_57;
  wire [22:0] _EVAL_31;
  wire [7:0] _EVAL_226;
  wire [7:0] _EVAL_94;
  wire [5:0] _EVAL_38;
  wire  _EVAL_298;
  wire  _EVAL_239;
  wire  _EVAL_110;
  wire  _EVAL_56;
  wire  _EVAL_329;
  wire  _EVAL_179;
  wire [127:0] _EVAL_186;
  wire [127:0] _EVAL_87;
  wire [72:0] _EVAL_70;
  wire [72:0] _EVAL_113;
  wire  _EVAL_326;
  wire  _EVAL_21;
  wire  _EVAL_193;
  wire [3:0] _EVAL_208;
  wire  _EVAL_143;
  wire  _EVAL_47;
  wire [22:0] _EVAL_268;
  wire  _EVAL_297;
  wire [1:0] _EVAL_308;
  wire [1:0] _EVAL_166;
  wire  _EVAL_46;
  wire  _EVAL_243;
  wire  _EVAL_65;
  wire  _EVAL_96;
  wire  _EVAL_332;
  wire  _EVAL_294;
  wire  _EVAL_60;
  wire  _EVAL_99;
  wire [3:0] _EVAL_324;
  wire  _EVAL_348;
  wire  _EVAL_318;
  wire  _EVAL_121;
  wire  _EVAL_205;
  wire  _EVAL_24;
  wire [3:0] _EVAL_275;
  wire  _EVAL_199;
  wire [2:0] _EVAL_266;
  wire  _EVAL_192;
  wire  _EVAL_203;
  wire  _EVAL_334;
  wire  _EVAL_55;
  wire  _EVAL_184;
  wire  _EVAL_163;
  wire  _EVAL_233;
  wire [2:0] _EVAL_89;
  wire  _EVAL_296;
  wire  _EVAL_264;
  wire [29:0] _EVAL_134;
  wire [29:0] _EVAL_123;
  wire [30:0] _EVAL_210;
  wire [30:0] _EVAL_54;
  wire [30:0] _EVAL_253;
  wire  _EVAL_235;
  wire  _EVAL_133;
  wire  _EVAL_311;
  wire  _EVAL_152;
  wire  _EVAL_258;
  wire  _EVAL_67;
  wire  _EVAL_340;
  wire  _EVAL_282;
  wire  _EVAL_172;
  wire  _EVAL_128;
  wire  _EVAL_114;
  wire  _EVAL_333;
  wire  _EVAL_283;
  wire [7:0] _EVAL_146;
  wire [7:0] _EVAL_93;
  wire [5:0] _EVAL_290;
  wire [5:0] _EVAL_336;
  wire  _EVAL_90;
  wire [29:0] _EVAL_88;
  wire [30:0] _EVAL_25;
  wire [30:0] _EVAL_202;
  wire [30:0] _EVAL_219;
  wire  _EVAL_306;
  wire  _EVAL_42;
  wire  _EVAL_244;
  wire  _EVAL_168;
  wire [5:0] _EVAL_287;
  wire  _EVAL_66;
  wire  _EVAL_129;
  wire  _EVAL_347;
  wire  _EVAL_213;
  wire  _EVAL_136;
  wire  _EVAL_119;
  wire  _EVAL_234;
  wire  _EVAL_248;
  wire  _EVAL_141;
  wire  _EVAL_338;
  wire  _EVAL_267;
  wire  _EVAL_73;
  wire  _EVAL_76;
  wire  _EVAL_276;
  wire [29:0] _EVAL_171;
  wire [30:0] _EVAL_217;
  wire  _EVAL_27;
  wire  _EVAL_102;
  wire [29:0] _EVAL_126;
  wire  _EVAL_200;
  wire  _EVAL_173;
  wire  _EVAL_107;
  wire  _EVAL_295;
  wire  _EVAL_274;
  wire  _EVAL_72;
  wire  _EVAL_153;
  wire  _EVAL_277;
  wire  _EVAL_44;
  wire  _EVAL_169;
  wire  _EVAL_84;
  wire [29:0] _EVAL_191;
  wire [30:0] _EVAL_351;
  wire [30:0] _EVAL_178;
  wire [30:0] _EVAL_197;
  wire  _EVAL_103;
  wire [29:0] _EVAL_180;
  wire [30:0] _EVAL_43;
  wire [30:0] _EVAL_321;
  wire [30:0] _EVAL_325;
  wire  _EVAL_101;
  wire  _EVAL_245;
  wire [30:0] _EVAL_343;
  wire [30:0] _EVAL_29;
  wire [30:0] _EVAL_261;
  wire  _EVAL_317;
  wire  _EVAL_307;
  wire [30:0] _EVAL_105;
  wire [30:0] _EVAL_40;
  wire  _EVAL_64;
  wire  _EVAL_204;
  wire  _EVAL_358;
  wire  _EVAL_125;
  wire  _EVAL_116;
  wire [5:0] _EVAL_122;
  wire  _EVAL_354;
  wire  _EVAL_83;
  wire  _EVAL_300;
  wire  _EVAL_224;
  wire  _EVAL_230;
  wire  _EVAL_158;
  wire  _EVAL_302;
  wire  _EVAL_137;
  wire  _EVAL_320;
  wire  _EVAL_45;
  wire  _EVAL_195;
  wire  _EVAL_270;
  wire  _EVAL_289;
  wire  _EVAL_212;
  wire  _EVAL_161;
  wire  _EVAL_118;
  wire  _EVAL_183;
  wire  _EVAL_188;
  wire  _EVAL_218;
  wire  _EVAL_344;
  wire  _EVAL_319;
  wire  _EVAL_50;
  wire  _EVAL_34;
  wire  _EVAL_259;
  wire  _EVAL_77;
  wire  _EVAL_359;
  wire  _EVAL_211;
  wire  _EVAL_28;
  wire  _EVAL_164;
  wire  _EVAL_305;
  wire  _EVAL_281;
  wire  _EVAL_303;
  wire  _EVAL_91;
  wire  _EVAL_132;
  wire  _EVAL_39;
  wire  _EVAL_198;
  wire  _EVAL_41;
  wire  _EVAL_360;
  wire  _EVAL_97;
  wire  _EVAL_115;
  wire  _EVAL_215;
  wire  _EVAL_106;
  wire  _EVAL_85;
  wire  _EVAL_269;
  wire  _EVAL_256;
  wire  _EVAL_190;
  wire [3:0] _EVAL_254;
  wire  _EVAL_155;
  wire  _EVAL_149;
  wire  _EVAL_301;
  wire  _EVAL_63;
  wire [127:0] _EVAL_139;
  wire [127:0] _EVAL_130;
  wire  _EVAL_310;
  wire [31:0] _EVAL_355;
  wire  _EVAL_313;
  wire  _EVAL_251;
  wire  _EVAL_156;
  wire  _EVAL_237;
  wire  _EVAL_81;
  wire  _EVAL_222;
  wire  _EVAL_328;
  wire  _EVAL_71;
  wire  _EVAL_162;
  wire  _EVAL_151;
  wire  _EVAL_120;
  wire [3:0] _EVAL_246;
  wire [3:0] _EVAL_80;
  wire  _EVAL_147;
  wire  _EVAL_236;
  wire  _EVAL_111;
  wire  _EVAL_356;
  wire  _EVAL_263;
  wire  _EVAL_53;
  wire  _EVAL_157;
  wire  _EVAL_257;
  wire  _EVAL_209;
  wire  _EVAL_35;
  wire  _EVAL_221;
  wire  _EVAL_346;
  wire  _EVAL_142;
  wire  _EVAL_181;
  wire  _EVAL_150;
  wire  _EVAL_79;
  wire  _EVAL_223;
  wire  _EVAL_49;
  wire  _EVAL_108;
  wire  _EVAL_238;
  wire  _EVAL_220;
  wire [72:0] _EVAL_315;
  wire [72:0] _EVAL_52;
  wire  _EVAL_185;
  wire  _EVAL_337;
  wire  _EVAL_159;
  wire  _EVAL_196;
  wire  _EVAL_109;
  wire  _EVAL_124;
  wire  _EVAL_293;
  wire  _EVAL_32;
  wire  _EVAL_19;
  wire  _EVAL_23;
  wire  _EVAL_353;
  wire  _EVAL_249;
  wire [72:0] _EVAL_341;
  wire  _EVAL_165;
  wire  _EVAL_22;
  wire  _EVAL_100;
  wire  _EVAL_327;
  wire  _EVAL_144;
  wire [72:0] _EVAL_286;
  wire  _EVAL_227;
  wire  _EVAL_135;
  wire [5:0] _EVAL_232;
  wire  _EVAL_345;
  wire  _EVAL_349;
  wire  _EVAL_342;
  wire [72:0] _EVAL_98;
  wire  _EVAL_61;
  wire  _EVAL_265;
  wire  _EVAL_225;
  wire  _EVAL_272;
  wire  _EVAL_216;
  wire  _EVAL_250;
  wire  _EVAL_92;
  wire  _EVAL_82;
  wire  _EVAL_148;
  wire  _EVAL_262;
  wire  _EVAL_75;
  wire  _EVAL_312;
  wire  _EVAL_279;
  wire  _EVAL_322;
  wire  _EVAL_335;
  wire  _EVAL_201;
  wire  _EVAL_280;
  wire  _EVAL_240;
  wire  _EVAL_231;
  wire  _EVAL_170;
  wire  _EVAL_228;
  wire  _EVAL_48;
  wire  _EVAL_314;
  wire  _EVAL_247;
  wire  _EVAL_174;
  wire  _EVAL_229;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_357 = _EVAL <= 3'h3;
  assign _EVAL_309 = _EVAL_357 | _EVAL_12;
  assign _EVAL_51 = _EVAL_11 == 1'h0;
  assign _EVAL_154 = _EVAL_51 | _EVAL_12;
  assign _EVAL_58 = _EVAL <= 3'h4;
  assign _EVAL_288 = _EVAL_58 | _EVAL_12;
  assign _EVAL_160 = _EVAL_288 == 1'h0;
  assign _EVAL_292 = _EVAL_26 >> _EVAL_14;
  assign _EVAL_316 = _EVAL_292[0];
  assign _EVAL_127 = _EVAL_316 == 1'h0;
  assign _EVAL_260 = _EVAL_15 == 2'h0;
  assign _EVAL_78 = _EVAL_260 | _EVAL_12;
  assign _EVAL_206 = _EVAL_304 == 6'h0;
  assign _EVAL_291 = _EVAL_206 == 1'h0;
  assign _EVAL_194 = _EVAL_18 ^ 30'h3000;
  assign _EVAL_131 = {1'b0,$signed(_EVAL_194)};
  assign _EVAL_140 = $signed(_EVAL_131) & $signed(-31'sh1000);
  assign _EVAL_86 = $signed(_EVAL_140);
  assign _EVAL_252 = $signed(_EVAL_86) == $signed(31'sh0);
  assign _EVAL_62 = _EVAL_9 == 3'h0;
  assign _EVAL_145 = _EVAL_17 == 3'h0;
  assign _EVAL_36 = _EVAL_10 & _EVAL_145;
  assign _EVAL_176 = _EVAL_14 == _EVAL_242;
  assign _EVAL_30 = _EVAL_176 | _EVAL_12;
  assign _EVAL_214 = _EVAL_2 == 1'h0;
  assign _EVAL_138 = _EVAL_214 | _EVAL_12;
  assign _EVAL_74 = _EVAL_138 == 1'h0;
  assign _EVAL_352 = _EVAL_9[2];
  assign _EVAL_57 = _EVAL_352 == 1'h0;
  assign _EVAL_31 = 23'hff << _EVAL_8;
  assign _EVAL_226 = _EVAL_31[7:0];
  assign _EVAL_94 = ~ _EVAL_226;
  assign _EVAL_38 = _EVAL_94[7:2];
  assign _EVAL_298 = _EVAL_13 & _EVAL_10;
  assign _EVAL_239 = _EVAL_278 == 6'h0;
  assign _EVAL_110 = _EVAL_298 & _EVAL_239;
  assign _EVAL_56 = _EVAL_17 == 3'h6;
  assign _EVAL_329 = _EVAL_56 == 1'h0;
  assign _EVAL_179 = _EVAL_110 & _EVAL_329;
  assign _EVAL_186 = 128'h1 << _EVAL_0;
  assign _EVAL_87 = _EVAL_179 ? _EVAL_186 : 128'h0;
  assign _EVAL_70 = _EVAL_87[72:0];
  assign _EVAL_113 = ~ _EVAL_70;
  assign _EVAL_326 = _EVAL_18 == _EVAL_284;
  assign _EVAL_21 = _EVAL_326 | _EVAL_12;
  assign _EVAL_193 = _EVAL_21 == 1'h0;
  assign _EVAL_208 = ~ _EVAL_4;
  assign _EVAL_143 = _EVAL_208 == 4'h0;
  assign _EVAL_47 = _EVAL_143 | _EVAL_12;
  assign _EVAL_268 = 23'hff << _EVAL_6;
  assign _EVAL_297 = _EVAL_8[0];
  assign _EVAL_308 = 2'h1 << _EVAL_297;
  assign _EVAL_166 = _EVAL_308 | 2'h1;
  assign _EVAL_46 = _EVAL_166[1];
  assign _EVAL_243 = _EVAL_9 == 3'h7;
  assign _EVAL_65 = _EVAL_16 & _EVAL_243;
  assign _EVAL_96 = _EVAL_9 == 3'h3;
  assign _EVAL_332 = _EVAL == 3'h0;
  assign _EVAL_294 = _EVAL_9 == 3'h4;
  assign _EVAL_60 = _EVAL_16 & _EVAL_294;
  assign _EVAL_99 = _EVAL_339 == 6'h0;
  assign _EVAL_324 = _EVAL_14[6:3];
  assign _EVAL_348 = _EVAL_324 == 4'h2;
  assign _EVAL_318 = _EVAL_9 == _EVAL_167;
  assign _EVAL_121 = _EVAL_0 == 7'h48;
  assign _EVAL_205 = _EVAL_0 == 7'h40;
  assign _EVAL_24 = _EVAL_121 | _EVAL_205;
  assign _EVAL_275 = _EVAL_0[6:3];
  assign _EVAL_199 = _EVAL_275 == 4'h8;
  assign _EVAL_266 = _EVAL_0[2:0];
  assign _EVAL_192 = 3'h1 <= _EVAL_266;
  assign _EVAL_203 = _EVAL_199 & _EVAL_192;
  assign _EVAL_334 = _EVAL_24 | _EVAL_203;
  assign _EVAL_55 = _EVAL_0 == 7'h20;
  assign _EVAL_184 = _EVAL_334 | _EVAL_55;
  assign _EVAL_163 = _EVAL_275 == 4'h0;
  assign _EVAL_233 = _EVAL_184 | _EVAL_163;
  assign _EVAL_89 = _EVAL_14[2:0];
  assign _EVAL_296 = 3'h1 <= _EVAL_89;
  assign _EVAL_264 = _EVAL_332 | _EVAL_12;
  assign _EVAL_134 = {{22'd0}, _EVAL_94};
  assign _EVAL_123 = _EVAL_18 ^ 30'h20000000;
  assign _EVAL_210 = {1'b0,$signed(_EVAL_123)};
  assign _EVAL_54 = $signed(_EVAL_210) & $signed(-31'sh2000);
  assign _EVAL_253 = $signed(_EVAL_54);
  assign _EVAL_235 = $signed(_EVAL_253) == $signed(31'sh0);
  assign _EVAL_133 = _EVAL_9 == 3'h6;
  assign _EVAL_311 = _EVAL_16 & _EVAL_133;
  assign _EVAL_152 = _EVAL_17[0];
  assign _EVAL_258 = _EVAL_17 == _EVAL_189;
  assign _EVAL_67 = _EVAL_258 | _EVAL_12;
  assign _EVAL_340 = _EVAL_67 == 1'h0;
  assign _EVAL_282 = _EVAL_26 != 73'h0;
  assign _EVAL_172 = _EVAL_282 == 1'h0;
  assign _EVAL_128 = _EVAL_8 <= 4'h8;
  assign _EVAL_114 = _EVAL_128 & _EVAL_252;
  assign _EVAL_333 = _EVAL_114 | _EVAL_12;
  assign _EVAL_283 = _EVAL_59 == 6'h0;
  assign _EVAL_146 = _EVAL_268[7:0];
  assign _EVAL_93 = ~ _EVAL_146;
  assign _EVAL_290 = _EVAL_93[7:2];
  assign _EVAL_336 = _EVAL_59 - 6'h1;
  assign _EVAL_90 = _EVAL_8 <= 4'h2;
  assign _EVAL_88 = _EVAL_18 ^ 30'h1900000;
  assign _EVAL_25 = {1'b0,$signed(_EVAL_88)};
  assign _EVAL_202 = $signed(_EVAL_25) & $signed(-31'sh2000);
  assign _EVAL_219 = $signed(_EVAL_202);
  assign _EVAL_306 = $signed(_EVAL_219) == $signed(31'sh0);
  assign _EVAL_42 = _EVAL_252 | _EVAL_306;
  assign _EVAL_244 = _EVAL_90 & _EVAL_42;
  assign _EVAL_168 = _EVAL_244 | _EVAL_12;
  assign _EVAL_287 = _EVAL_278 - 6'h1;
  assign _EVAL_66 = plusarg_reader_out == 32'h0;
  assign _EVAL_129 = _EVAL_17 <= 3'h6;
  assign _EVAL_347 = _EVAL_129 | _EVAL_12;
  assign _EVAL_213 = _EVAL_347 == 1'h0;
  assign _EVAL_136 = _EVAL != 3'h0;
  assign _EVAL_119 = _EVAL_8 >= 4'h2;
  assign _EVAL_234 = _EVAL_18[1];
  assign _EVAL_248 = _EVAL_46 & _EVAL_234;
  assign _EVAL_141 = _EVAL_119 | _EVAL_248;
  assign _EVAL_338 = _EVAL_309 == 1'h0;
  assign _EVAL_267 = _EVAL_324 == 4'h0;
  assign _EVAL_73 = _EVAL_1 == 1'h0;
  assign _EVAL_76 = _EVAL_324 == 4'h3;
  assign _EVAL_276 = _EVAL_7 == _EVAL_207;
  assign _EVAL_171 = _EVAL_18 ^ 30'h1800000;
  assign _EVAL_217 = {1'b0,$signed(_EVAL_171)};
  assign _EVAL_27 = _EVAL_9 == 3'h2;
  assign _EVAL_102 = _EVAL <= 3'h2;
  assign _EVAL_126 = _EVAL_18 & _EVAL_134;
  assign _EVAL_200 = _EVAL_126 == 30'h0;
  assign _EVAL_173 = _EVAL_200 | _EVAL_12;
  assign _EVAL_107 = _EVAL_173 == 1'h0;
  assign _EVAL_295 = _EVAL_14 == 7'h40;
  assign _EVAL_274 = 4'h6 == _EVAL_8;
  assign _EVAL_72 = _EVAL_295 ? _EVAL_274 : 1'h0;
  assign _EVAL_153 = _EVAL_72 | _EVAL_12;
  assign _EVAL_277 = _EVAL_153 == 1'h0;
  assign _EVAL_44 = _EVAL_6 >= 4'h2;
  assign _EVAL_169 = _EVAL_44 | _EVAL_12;
  assign _EVAL_84 = _EVAL_169 == 1'h0;
  assign _EVAL_191 = _EVAL_18 ^ 30'hc000000;
  assign _EVAL_351 = {1'b0,$signed(_EVAL_191)};
  assign _EVAL_178 = $signed(_EVAL_351) & $signed(-31'sh4000000);
  assign _EVAL_197 = $signed(_EVAL_178);
  assign _EVAL_103 = $signed(_EVAL_197) == $signed(31'sh0);
  assign _EVAL_180 = _EVAL_18 ^ 30'h2000000;
  assign _EVAL_43 = {1'b0,$signed(_EVAL_180)};
  assign _EVAL_321 = $signed(_EVAL_43) & $signed(-31'sh10000);
  assign _EVAL_325 = $signed(_EVAL_321);
  assign _EVAL_101 = $signed(_EVAL_325) == $signed(31'sh0);
  assign _EVAL_245 = _EVAL_103 | _EVAL_101;
  assign _EVAL_343 = {1'b0,$signed(_EVAL_18)};
  assign _EVAL_29 = $signed(_EVAL_343) & $signed(-31'sh5000);
  assign _EVAL_261 = $signed(_EVAL_29);
  assign _EVAL_317 = $signed(_EVAL_261) == $signed(31'sh0);
  assign _EVAL_307 = _EVAL_245 | _EVAL_317;
  assign _EVAL_105 = $signed(_EVAL_217) & $signed(-31'sh8000);
  assign _EVAL_40 = $signed(_EVAL_105);
  assign _EVAL_64 = $signed(_EVAL_40) == $signed(31'sh0);
  assign _EVAL_204 = _EVAL_307 | _EVAL_64;
  assign _EVAL_358 = _EVAL_204 | _EVAL_306;
  assign _EVAL_125 = _EVAL_358 | _EVAL_235;
  assign _EVAL_116 = _EVAL_5 & _EVAL_16;
  assign _EVAL_122 = _EVAL_304 - 6'h1;
  assign _EVAL_354 = _EVAL_14 == 7'h48;
  assign _EVAL_83 = _EVAL_354 | _EVAL_295;
  assign _EVAL_300 = _EVAL_324 == 4'h8;
  assign _EVAL_224 = _EVAL_300 & _EVAL_296;
  assign _EVAL_230 = _EVAL_83 | _EVAL_224;
  assign _EVAL_158 = _EVAL_14 == 7'h20;
  assign _EVAL_302 = _EVAL_230 | _EVAL_158;
  assign _EVAL_137 = _EVAL_302 | _EVAL_267;
  assign _EVAL_320 = _EVAL_324 == 4'h1;
  assign _EVAL_45 = _EVAL_137 | _EVAL_320;
  assign _EVAL_195 = _EVAL_45 | _EVAL_348;
  assign _EVAL_270 = _EVAL_195 | _EVAL_76;
  assign _EVAL_289 = _EVAL_270 | _EVAL_12;
  assign _EVAL_212 = _EVAL_289 == 1'h0;
  assign _EVAL_161 = _EVAL_78 == 1'h0;
  assign _EVAL_118 = _EVAL_6 == _EVAL_331;
  assign _EVAL_183 = _EVAL_172 | _EVAL_66;
  assign _EVAL_188 = _EVAL_112 < plusarg_reader_out;
  assign _EVAL_218 = _EVAL_183 | _EVAL_188;
  assign _EVAL_344 = _EVAL_8 <= 4'h6;
  assign _EVAL_319 = _EVAL_118 | _EVAL_12;
  assign _EVAL_50 = _EVAL_275 == 4'h2;
  assign _EVAL_34 = _EVAL_116 & _EVAL_206;
  assign _EVAL_259 = _EVAL_344 & _EVAL_125;
  assign _EVAL_77 = _EVAL_114 | _EVAL_259;
  assign _EVAL_359 = _EVAL_77 | _EVAL_12;
  assign _EVAL_211 = _EVAL_166[0];
  assign _EVAL_28 = _EVAL_18[0];
  assign _EVAL_164 = _EVAL_234 & _EVAL_28;
  assign _EVAL_305 = _EVAL_211 & _EVAL_164;
  assign _EVAL_281 = _EVAL_141 | _EVAL_305;
  assign _EVAL_303 = _EVAL_73 | _EVAL_12;
  assign _EVAL_91 = _EVAL_303 == 1'h0;
  assign _EVAL_132 = _EVAL_28 == 1'h0;
  assign _EVAL_39 = _EVAL_234 & _EVAL_132;
  assign _EVAL_198 = _EVAL_211 & _EVAL_39;
  assign _EVAL_41 = _EVAL_141 | _EVAL_198;
  assign _EVAL_360 = _EVAL_234 == 1'h0;
  assign _EVAL_97 = _EVAL_46 & _EVAL_360;
  assign _EVAL_115 = _EVAL_119 | _EVAL_97;
  assign _EVAL_215 = _EVAL_360 & _EVAL_28;
  assign _EVAL_106 = _EVAL_211 & _EVAL_215;
  assign _EVAL_85 = _EVAL_115 | _EVAL_106;
  assign _EVAL_269 = _EVAL_360 & _EVAL_132;
  assign _EVAL_256 = _EVAL_211 & _EVAL_269;
  assign _EVAL_190 = _EVAL_115 | _EVAL_256;
  assign _EVAL_254 = {_EVAL_281,_EVAL_41,_EVAL_85,_EVAL_190};
  assign _EVAL_155 = _EVAL_4 == _EVAL_254;
  assign _EVAL_149 = _EVAL_155 | _EVAL_12;
  assign _EVAL_301 = _EVAL_149 == 1'h0;
  assign _EVAL_63 = _EVAL_116 & _EVAL_99;
  assign _EVAL_139 = 128'h1 << _EVAL_14;
  assign _EVAL_130 = _EVAL_63 ? _EVAL_139 : 128'h0;
  assign _EVAL_310 = _EVAL_116 | _EVAL_298;
  assign _EVAL_355 = _EVAL_112 + 32'h1;
  assign _EVAL_313 = _EVAL_8 == _EVAL_20;
  assign _EVAL_251 = _EVAL_313 | _EVAL_12;
  assign _EVAL_156 = _EVAL_283 == 1'h0;
  assign _EVAL_237 = _EVAL_102 | _EVAL_12;
  assign _EVAL_81 = _EVAL_319 == 1'h0;
  assign _EVAL_222 = _EVAL_0 == _EVAL_241;
  assign _EVAL_328 = _EVAL_222 | _EVAL_12;
  assign _EVAL_71 = _EVAL_328 == 1'h0;
  assign _EVAL_162 = _EVAL == _EVAL_273;
  assign _EVAL_151 = _EVAL_162 | _EVAL_12;
  assign _EVAL_120 = _EVAL_151 == 1'h0;
  assign _EVAL_246 = ~ _EVAL_254;
  assign _EVAL_80 = _EVAL_4 & _EVAL_246;
  assign _EVAL_147 = _EVAL_80 == 4'h0;
  assign _EVAL_236 = _EVAL_147 | _EVAL_12;
  assign _EVAL_111 = _EVAL_236 == 1'h0;
  assign _EVAL_356 = _EVAL_127 | _EVAL_12;
  assign _EVAL_263 = _EVAL_275 == 4'h1;
  assign _EVAL_53 = _EVAL_233 | _EVAL_263;
  assign _EVAL_157 = _EVAL_53 | _EVAL_50;
  assign _EVAL_257 = _EVAL_275 == 4'h3;
  assign _EVAL_209 = _EVAL_157 | _EVAL_257;
  assign _EVAL_35 = _EVAL_119 | _EVAL_12;
  assign _EVAL_221 = _EVAL_15 == _EVAL_187;
  assign _EVAL_346 = _EVAL_221 | _EVAL_12;
  assign _EVAL_142 = _EVAL_9 == 3'h5;
  assign _EVAL_181 = _EVAL_16 & _EVAL_142;
  assign _EVAL_150 = _EVAL_15 != 2'h2;
  assign _EVAL_79 = _EVAL_150 | _EVAL_12;
  assign _EVAL_223 = _EVAL_79 == 1'h0;
  assign _EVAL_49 = _EVAL_17 == 3'h4;
  assign _EVAL_108 = _EVAL_16 & _EVAL_62;
  assign _EVAL_238 = _EVAL_276 | _EVAL_12;
  assign _EVAL_220 = _EVAL_238 == 1'h0;
  assign _EVAL_315 = _EVAL_130[72:0];
  assign _EVAL_52 = _EVAL_26 | _EVAL_315;
  assign _EVAL_185 = _EVAL_16 & _EVAL_291;
  assign _EVAL_337 = _EVAL_154 == 1'h0;
  assign _EVAL_159 = _EVAL_73 | _EVAL_11;
  assign _EVAL_196 = _EVAL_159 | _EVAL_12;
  assign _EVAL_109 = _EVAL_196 == 1'h0;
  assign _EVAL_124 = _EVAL_298 & _EVAL_283;
  assign _EVAL_293 = _EVAL_209 | _EVAL_12;
  assign _EVAL_32 = _EVAL_293 == 1'h0;
  assign _EVAL_19 = _EVAL_16 & _EVAL_96;
  assign _EVAL_23 = _EVAL_9 == 3'h1;
  assign _EVAL_353 = _EVAL_12 == 1'h0;
  assign _EVAL_249 = _EVAL_168 == 1'h0;
  assign _EVAL_341 = _EVAL_315 | _EVAL_26;
  assign _EVAL_165 = _EVAL_318 | _EVAL_12;
  assign _EVAL_22 = _EVAL_165 == 1'h0;
  assign _EVAL_100 = _EVAL_218 | _EVAL_12;
  assign _EVAL_327 = _EVAL_17 == 3'h2;
  assign _EVAL_144 = _EVAL_136 | _EVAL_12;
  assign _EVAL_286 = _EVAL_52 & _EVAL_113;
  assign _EVAL_227 = _EVAL_16 & _EVAL_27;
  assign _EVAL_135 = _EVAL_10 & _EVAL_49;
  assign _EVAL_232 = _EVAL_339 - 6'h1;
  assign _EVAL_345 = _EVAL_15 <= 2'h2;
  assign _EVAL_349 = _EVAL_345 | _EVAL_12;
  assign _EVAL_342 = _EVAL_349 == 1'h0;
  assign _EVAL_98 = _EVAL_341 >> _EVAL_0;
  assign _EVAL_61 = _EVAL_1 == _EVAL_271;
  assign _EVAL_265 = _EVAL_61 | _EVAL_12;
  assign _EVAL_225 = _EVAL_265 == 1'h0;
  assign _EVAL_272 = _EVAL_346 == 1'h0;
  assign _EVAL_216 = _EVAL_98[0];
  assign _EVAL_250 = _EVAL_216 | _EVAL_12;
  assign _EVAL_92 = _EVAL_47 == 1'h0;
  assign _EVAL_82 = _EVAL_333 == 1'h0;
  assign _EVAL_148 = _EVAL_17 == 3'h1;
  assign _EVAL_262 = _EVAL_17 == 3'h5;
  assign _EVAL_75 = _EVAL_10 & _EVAL_262;
  assign _EVAL_312 = _EVAL_100 == 1'h0;
  assign _EVAL_279 = _EVAL_30 == 1'h0;
  assign _EVAL_322 = _EVAL_16 & _EVAL_23;
  assign _EVAL_335 = _EVAL_251 == 1'h0;
  assign _EVAL_201 = _EVAL_35 == 1'h0;
  assign _EVAL_280 = _EVAL_10 & _EVAL_156;
  assign _EVAL_240 = _EVAL_10 & _EVAL_148;
  assign _EVAL_231 = _EVAL_359 == 1'h0;
  assign _EVAL_170 = _EVAL_264 == 1'h0;
  assign _EVAL_228 = _EVAL_356 == 1'h0;
  assign _EVAL_48 = _EVAL_250 == 1'h0;
  assign _EVAL_314 = _EVAL_144 == 1'h0;
  assign _EVAL_247 = _EVAL_237 == 1'h0;
  assign _EVAL_174 = _EVAL_10 & _EVAL_56;
  assign _EVAL_229 = _EVAL_10 & _EVAL_327;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _EVAL_26 = _RAND_1[72:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_59 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_112 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_167 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_187 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_189 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_207 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_241 = _RAND_8[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_242 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_271 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_273 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_278 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_284 = _RAND_13[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_304 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_331 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_339 = _RAND_16[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_3) begin
    if (_EVAL_34) begin
      _EVAL_20 <= _EVAL_8;
    end
    if (_EVAL_12) begin
      _EVAL_26 <= 73'h0;
    end else begin
      _EVAL_26 <= _EVAL_286;
    end
    if (_EVAL_12) begin
      _EVAL_59 <= 6'h0;
    end else begin
      if (_EVAL_298) begin
        if (_EVAL_283) begin
          if (_EVAL_152) begin
            _EVAL_59 <= _EVAL_290;
          end else begin
            _EVAL_59 <= 6'h0;
          end
        end else begin
          _EVAL_59 <= _EVAL_336;
        end
      end
    end
    if (_EVAL_12) begin
      _EVAL_112 <= 32'h0;
    end else begin
      if (_EVAL_310) begin
        _EVAL_112 <= 32'h0;
      end else begin
        _EVAL_112 <= _EVAL_355;
      end
    end
    if (_EVAL_34) begin
      _EVAL_167 <= _EVAL_9;
    end
    if (_EVAL_124) begin
      _EVAL_187 <= _EVAL_15;
    end
    if (_EVAL_124) begin
      _EVAL_189 <= _EVAL_17;
    end
    if (_EVAL_124) begin
      _EVAL_207 <= _EVAL_7;
    end
    if (_EVAL_124) begin
      _EVAL_241 <= _EVAL_0;
    end
    if (_EVAL_34) begin
      _EVAL_242 <= _EVAL_14;
    end
    if (_EVAL_124) begin
      _EVAL_271 <= _EVAL_1;
    end
    if (_EVAL_34) begin
      _EVAL_273 <= _EVAL;
    end
    if (_EVAL_12) begin
      _EVAL_278 <= 6'h0;
    end else begin
      if (_EVAL_298) begin
        if (_EVAL_239) begin
          if (_EVAL_152) begin
            _EVAL_278 <= _EVAL_290;
          end else begin
            _EVAL_278 <= 6'h0;
          end
        end else begin
          _EVAL_278 <= _EVAL_287;
        end
      end
    end
    if (_EVAL_34) begin
      _EVAL_284 <= _EVAL_18;
    end
    if (_EVAL_12) begin
      _EVAL_304 <= 6'h0;
    end else begin
      if (_EVAL_116) begin
        if (_EVAL_206) begin
          if (_EVAL_57) begin
            _EVAL_304 <= _EVAL_38;
          end else begin
            _EVAL_304 <= 6'h0;
          end
        end else begin
          _EVAL_304 <= _EVAL_122;
        end
      end
    end
    if (_EVAL_124) begin
      _EVAL_331 <= _EVAL_6;
    end
    if (_EVAL_12) begin
      _EVAL_339 <= 6'h0;
    end else begin
      if (_EVAL_116) begin
        if (_EVAL_99) begin
          if (_EVAL_57) begin
            _EVAL_339 <= _EVAL_38;
          end else begin
            _EVAL_339 <= 6'h0;
          end
        end else begin
          _EVAL_339 <= _EVAL_232;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df6bddda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a818495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90746b0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30f8028a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7d1e217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c370f6a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0e70e88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd7e2a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93f5d4d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(280239bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e3749c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5488cd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d829688a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(511712e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfde321)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5d09779)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f5713b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_337) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff6c8c12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f66139ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0925afc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(282352cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7328be1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eec1b8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2871df9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e980a4df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(485dcabd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(682edd7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_335) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_340) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4516cc9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66af9345)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f94376b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7664386a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa86548)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(707beff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27487583)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f46c3ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44871a8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cda20ae3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2035895d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed40b550)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6be95a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1fcdbe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34a403ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_337) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d619868c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_335) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99f819d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b48ea2f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_337) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(353ac12e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e71d68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(522ae2b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f13a073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d94296a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(605e05da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca519a2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6bcfd4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a57c8fd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba53ee37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff9b5726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(136d20a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_340) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8da39979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_337) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88642cba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3904b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afe063b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca8b9cad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47777fb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a21bbd74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a9d892)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcc7cee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c59a1c9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4153c56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e49ac531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffccf4de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca514aa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eca431f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adeb79ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c739570b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d1ee487)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bae2429)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b1dae0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854e2ca9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e59c314)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b80148)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e8757a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d25ac706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61d5ffa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b39b9699)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4657a292)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f8981f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd0f38c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b91dde1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c0c2874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
