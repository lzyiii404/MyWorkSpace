//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_213_assert(
  input          _EVAL,
  input  [3:0]   _EVAL_1,
  input          _EVAL_2,
  input  [2:0]   _EVAL_3,
  input          _EVAL_4,
  input  [1:0]   _EVAL_6,
  input  [2:0]   _EVAL_9,
  input          _EVAL_11,
  input  [1:0]   _EVAL_12,
  input          _EVAL_13,
  input  [3:0]   _EVAL_14,
  input  [2:0]   _EVAL_15,
  input          _EVAL_18,
  input  [2:0]   _EVAL_21,
  input  [11:0]  _EVAL_23,
  input          _EVAL_28,
  input          _EVAL_30,
  input  [8:0]   _EVAL_32,
  input          _EVAL_41,
  input          _EVAL_48,
  input  [11:0]  _EVAL_51,
  input          _EVAL_616,
  input          _EVAL_734,
  input  [1:0]   _EVAL_838,
  input          _EVAL_1829,
  input  [2:0]   _EVAL_2167,
  input  [31:0]  _EVAL_1582,
  input          _EVAL_1048,
  input          _EVAL_644,
  input  [511:0] _EVAL_631,
  input          _EVAL_502,
  input          _EVAL_1760,
  input  [31:0]  _EVAL_332,
  input  [7:0]   _EVAL_1017,
  input          _EVAL_1486,
  input          _EVAL_681,
  input          _EVAL_2076,
  input  [63:0]  _EVAL_1421,
  input          _EVAL_680,
  input          _EVAL_139,
  input          _EVAL_1971,
  input          _EVAL_749,
  input  [7:0]   _EVAL_573,
  input          _EVAL_1387,
  input          _EVAL_1145,
  input  [7:0]   _EVAL_1563,
  input          _EVAL_758,
  input          _EVAL_886,
  input          _EVAL_57,
  input  [7:0]   _EVAL_1753,
  input          _EVAL_1638,
  input          _EVAL_857,
  input          _EVAL_1093,
  input          _EVAL_568,
  input          _EVAL_214,
  input          _EVAL_1732,
  input          _EVAL_1303,
  input          _EVAL_2178,
  input          _EVAL_1311,
  input          _EVAL_1501,
  input          _EVAL_1709,
  input          _EVAL_614,
  input          _EVAL_129,
  input          _EVAL_1286,
  input          _EVAL_299,
  input          _EVAL_637,
  input          _EVAL_1608,
  input          _EVAL_994,
  input          _EVAL_328,
  input          _EVAL_2095,
  input          _EVAL_986,
  input          _EVAL_1845,
  input  [9:0]   _EVAL_190,
  input          _EVAL_1188,
  input          _EVAL_1831,
  input          _EVAL_556,
  input          _EVAL_1558,
  input          _EVAL_1654,
  input          _EVAL_1680,
  input          _EVAL_2102,
  input          _EVAL_1570,
  input          _EVAL_233,
  input          _EVAL_418,
  input          _EVAL_1532,
  input          _EVAL_2088,
  input          _EVAL_1551,
  input          _EVAL_166,
  input          _EVAL_1163,
  input          _EVAL_1317,
  input          _EVAL_1192,
  input          _EVAL_1296,
  input          _EVAL_1133,
  input          _EVAL_958,
  input          _EVAL_1171,
  input          _EVAL_1490,
  input          _EVAL_884,
  input          _EVAL_408,
  input          _EVAL_483,
  input          _EVAL_620,
  input          _EVAL_559,
  input          _EVAL_1708,
  input          _EVAL_1752,
  input          _EVAL_2195,
  input          _EVAL_669,
  input          _EVAL_1237,
  input          _EVAL_1242,
  input          _EVAL_686,
  input          _EVAL_191,
  input          _EVAL_221,
  input          _EVAL_1003,
  input          _EVAL_957,
  input          _EVAL_2068,
  input          _EVAL_469,
  input          _EVAL_361,
  input          _EVAL_164,
  input          _EVAL_1838,
  input          _EVAL_1885,
  input          _EVAL_1592,
  input          _EVAL_435,
  input          _EVAL_2192,
  input          _EVAL_590,
  input          _EVAL_1535,
  input          _EVAL_1103,
  input          _EVAL_1750,
  input          _EVAL_1071,
  input          _EVAL_1773,
  input          _EVAL_1998,
  input          _EVAL_517,
  input          _EVAL_833,
  input          _EVAL_320,
  input          _EVAL_1677,
  input          _EVAL_1598,
  input          _EVAL_1820,
  input          _EVAL_319,
  input          _EVAL_1480,
  input          _EVAL_728,
  input          _EVAL_1225,
  input          _EVAL_1889,
  input          _EVAL_141,
  input          _EVAL_175,
  input          _EVAL_1222,
  input          _EVAL_1847,
  input          _EVAL_1391,
  input          _EVAL_953,
  input          _EVAL_1959,
  input          _EVAL_256,
  input          _EVAL_172,
  input          _EVAL_2011,
  input          _EVAL_989,
  input          _EVAL_979,
  input          _EVAL_349,
  input          _EVAL_1153,
  input          _EVAL_1988,
  input          _EVAL_1429,
  input          _EVAL_1703,
  input          _EVAL_2224,
  input          _EVAL_311,
  input          _EVAL_766,
  input          _EVAL_1766,
  input          _EVAL_1997,
  input          _EVAL_1813,
  input          _EVAL_1987,
  input          _EVAL_1534,
  input          _EVAL_1435,
  input          _EVAL_1147,
  input          _EVAL_2079,
  input          _EVAL_1890,
  input          _EVAL_589,
  input          _EVAL_1973,
  input          _EVAL_1711,
  input          _EVAL_598,
  input          _EVAL_260,
  input          _EVAL_487,
  input          _EVAL_685,
  input          _EVAL_1671,
  input          _EVAL_60,
  input          _EVAL_1542,
  input          _EVAL_322,
  input          _EVAL_1441,
  input          _EVAL_1047,
  input          _EVAL_783,
  input          _EVAL_1627,
  input          _EVAL_840,
  input          _EVAL_1210,
  input          _EVAL_1864,
  input  [2:0]   _EVAL_1511,
  input          _EVAL_841,
  input          _EVAL_155,
  input          _EVAL_1082,
  input          _EVAL_923,
  input          _EVAL_1589,
  input          _EVAL_135,
  input          _EVAL_1357,
  input          _EVAL_88,
  input          _EVAL_555,
  input          _EVAL_2222,
  input          _EVAL_371,
  input          _EVAL_1430,
  input          _EVAL_1066,
  input          _EVAL_1806,
  input          _EVAL_1316,
  input          _EVAL_2109,
  input  [15:0]  _EVAL_744,
  input          _EVAL_1465,
  input          _EVAL_1977,
  input          _EVAL_1101,
  input          _EVAL_1428,
  input          _EVAL_1822,
  input          _EVAL_1902,
  input          _EVAL_1789,
  input          _EVAL_2194,
  input          _EVAL_444,
  input          _EVAL_1413,
  input          _EVAL_822,
  input          _EVAL_611,
  input          _EVAL_208,
  input          _EVAL_2152,
  input          _EVAL_777,
  input          _EVAL_2230,
  input          _EVAL_666,
  input          _EVAL_1022,
  input          _EVAL_1337,
  input          _EVAL_1310,
  input          _EVAL_2218,
  input          _EVAL_2020,
  input          _EVAL_1401,
  input          _EVAL_577,
  input          _EVAL_622,
  input          _EVAL_1230,
  input          _EVAL_1821,
  input          _EVAL_1111,
  input          _EVAL_2108,
  input          _EVAL_1271,
  input          _EVAL_312,
  input          _EVAL_872,
  input          _EVAL_2191,
  input          _EVAL_1906,
  input          _EVAL_866,
  input          _EVAL_1049,
  input          _EVAL_1425,
  input          _EVAL_1197,
  input          _EVAL_1105,
  input          _EVAL_503,
  input          _EVAL_69,
  input          _EVAL_1095,
  input          _EVAL_1326,
  input          _EVAL_207,
  input          _EVAL_383,
  input          _EVAL_2200,
  input          _EVAL_1976,
  input          _EVAL_472,
  input          _EVAL_887,
  input          _EVAL_785,
  input  [2:0]   _EVAL_1892,
  input          _EVAL_1517,
  input          _EVAL_1371,
  input          _EVAL_567,
  input          _EVAL_498,
  input          _EVAL_929,
  input          _EVAL_1092,
  input          _EVAL_1113,
  input          _EVAL_179,
  input          _EVAL_1406,
  input  [2:0]   _EVAL_431,
  input          _EVAL_511,
  input          _EVAL_1717,
  input          _EVAL_1936,
  input          _EVAL_2038,
  input          _EVAL_2014,
  input          _EVAL_1622,
  input          _EVAL_1870,
  input          _EVAL_2032,
  input          _EVAL_108,
  input          _EVAL_1612,
  input          _EVAL_981,
  input          _EVAL_786,
  input          _EVAL_1541,
  input          _EVAL_670,
  input          _EVAL_706,
  input          _EVAL_1191,
  input          _EVAL_1460,
  input          _EVAL_712,
  input          _EVAL_718,
  input          _EVAL_521,
  input          _EVAL_1873,
  input          _EVAL_404,
  input          _EVAL_1918,
  input          _EVAL_933,
  input          _EVAL_80,
  input          _EVAL_588,
  input          _EVAL_969,
  input          _EVAL_2134,
  input          _EVAL_875,
  input          _EVAL_2170,
  input          _EVAL_805,
  input          _EVAL_1218,
  input          _EVAL_1688,
  input  [13:0]  _EVAL_156,
  input          _EVAL_1115,
  input          _EVAL_1158,
  input          _EVAL_279,
  input          _EVAL_2048,
  input          _EVAL_703,
  input          _EVAL_1353,
  input          _EVAL_103,
  input          _EVAL_784,
  input          _EVAL_671,
  input          _EVAL_1787,
  input          _EVAL_149,
  input          _EVAL_543,
  input          _EVAL_2034,
  input          _EVAL_1797,
  input          _EVAL_2144,
  input          _EVAL_1433,
  input          _EVAL_112,
  input          _EVAL_1522,
  input          _EVAL_362,
  input          _EVAL_912,
  input  [2:0]   _EVAL_867,
  input          _EVAL_1938,
  input          _EVAL_678,
  input          _EVAL_1643,
  input          _EVAL_2139,
  input          _EVAL_694,
  input          _EVAL_1939,
  input          _EVAL_449,
  input          sb2tlOpt__EVAL_11,
  input          sb2tlOpt__EVAL_25
);
  wire  TLMonitor__EVAL;
  wire [2:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [2:0] TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire [3:0] TLMonitor__EVAL_9;
  wire [1:0] TLMonitor__EVAL_10;
  wire [8:0] TLMonitor__EVAL_11;
  wire [1:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire  TLMonitor_1__EVAL;
  wire [11:0] TLMonitor_1__EVAL_0;
  wire [11:0] TLMonitor_1__EVAL_1;
  wire [1:0] TLMonitor_1__EVAL_2;
  wire  TLMonitor_1__EVAL_3;
  wire  TLMonitor_1__EVAL_4;
  wire [2:0] TLMonitor_1__EVAL_5;
  wire [3:0] TLMonitor_1__EVAL_6;
  wire [1:0] TLMonitor_1__EVAL_7;
  wire [2:0] TLMonitor_1__EVAL_8;
  wire  TLMonitor_1__EVAL_9;
  wire [2:0] TLMonitor_1__EVAL_10;
  wire  TLMonitor_1__EVAL_11;
  wire  TLMonitor_1__EVAL_12;
  wire  TLMonitor_1__EVAL_13;
  wire [11:0] TLMonitor_1__EVAL_14;
  wire [5:0] _EVAL_1267;
  wire  _EVAL_927;
  wire  _EVAL_1151;
  wire  _EVAL_1497;
  wire  _EVAL_967;
  wire  _EVAL_978;
  wire  _EVAL_2123;
  wire  _EVAL_592;
  wire  _EVAL_2022;
  wire  _EVAL_1102;
  wire  _EVAL_338;
  wire  _EVAL_280;
  wire  _EVAL_294;
  wire  _EVAL_1124;
  wire  _EVAL_316;
  wire  _EVAL_1073;
  wire  _EVAL_1444;
  wire  _EVAL_1467;
  wire  _EVAL_1013;
  wire  _EVAL_1178;
  wire [2:0] _EVAL_1978;
  wire  _EVAL_1220;
  wire  _EVAL_2107;
  wire  _EVAL_269;
  wire  _EVAL_1521;
  wire  _EVAL_494;
  wire  _EVAL_973;
  wire  _EVAL_250;
  wire  _EVAL_850;
  wire  _EVAL_1723;
  wire  _EVAL_1336;
  wire  _EVAL_689;
  wire  _EVAL_951;
  wire  _EVAL_564;
  wire  _EVAL_102;
  wire  _EVAL_1792;
  wire  _EVAL_525;
  wire  _EVAL_1676;
  wire  _EVAL_2124;
  wire  _EVAL_1143;
  wire  _EVAL_402;
  wire  _EVAL_456;
  wire  _EVAL_1027;
  wire [3:0] _EVAL_1539;
  wire  _EVAL_2064;
  wire  _EVAL_546;
  wire  _EVAL_2065;
  wire  _EVAL_1149;
  wire  _EVAL_154;
  wire  _EVAL_939;
  wire  _EVAL_798;
  wire  _EVAL_844;
  wire  _EVAL_578;
  wire  _EVAL_1030;
  wire  _EVAL_946;
  wire  _EVAL_1705;
  wire  _EVAL_2132;
  wire  _EVAL_1645;
  wire  _EVAL_922;
  wire [14:0] _EVAL_1748;
  wire  _EVAL_1142;
  wire  _EVAL_275;
  wire  _EVAL_1109;
  wire  _EVAL_2213;
  wire  _EVAL_2176;
  wire  _EVAL_926;
  wire  _EVAL_1784;
  wire  _EVAL_1106;
  wire  _EVAL_1172;
  wire  _EVAL_1689;
  wire [3:0] _EVAL_599;
  wire  _EVAL_58;
  wire  _EVAL_510;
  wire [4:0] _EVAL_1168;
  wire  _EVAL_1278;
  wire  _EVAL_1552;
  wire  _EVAL_499;
  wire  _EVAL_134;
  wire  _EVAL_1369;
  wire  _EVAL_2168;
  wire  _EVAL_1601;
  wire  _EVAL_2231;
  wire  _EVAL_1867;
  wire  _EVAL_762;
  wire  _EVAL_1647;
  wire  _EVAL_2005;
  wire  _EVAL_526;
  wire  _EVAL_1035;
  wire  _EVAL_1075;
  wire  _EVAL_477;
  wire  _EVAL_1388;
  wire  _EVAL_997;
  wire  _EVAL_2193;
  wire [1:0] _EVAL_1208;
  wire  _EVAL_286;
  wire  _EVAL_1659;
  wire  _EVAL_807;
  wire  _EVAL_1355;
  wire  _EVAL_911;
  wire  _EVAL_1203;
  wire  _EVAL_1527;
  wire  _EVAL_2209;
  wire  _EVAL_972;
  wire  _EVAL_2143;
  wire  _EVAL_1559;
  wire  _EVAL_337;
  wire  _EVAL_2151;
  wire  _EVAL_1032;
  wire  _EVAL_1228;
  wire  _EVAL_365;
  wire  _EVAL_674;
  wire  _EVAL_842;
  wire  _EVAL_314;
  wire  _EVAL_1937;
  wire  _EVAL_1779;
  wire  _EVAL_1363;
  wire  _EVAL_1557;
  wire  _EVAL_1289;
  wire  _EVAL_150;
  wire  _EVAL_585;
  wire  _EVAL_396;
  wire  _EVAL_369;
  wire  _EVAL_379;
  wire [6:0] _EVAL_913;
  wire  _EVAL_580;
  wire  _EVAL_1442;
  wire [1:0] _EVAL_249;
  wire  _EVAL_1553;
  wire  _EVAL_1894;
  wire  _EVAL_1288;
  wire  _EVAL_2188;
  wire  _EVAL_1202;
  wire  _EVAL_949;
  wire  _EVAL_1802;
  wire  _EVAL_1426;
  wire  _EVAL_1684;
  wire  _EVAL_2180;
  wire  _EVAL_595;
  wire  _EVAL_2083;
  wire [3:0] _EVAL_1913;
  wire  _EVAL_2033;
  wire  _EVAL_931;
  wire  _EVAL_1625;
  wire  _EVAL_1519;
  wire  _EVAL_992;
  wire  _EVAL_1281;
  wire  _EVAL_1675;
  wire  _EVAL_1257;
  wire  _EVAL_1526;
  wire  _EVAL_2089;
  wire  _EVAL_1097;
  wire  _EVAL_664;
  wire  _EVAL_1828;
  wire  _EVAL_2112;
  wire  _EVAL_1248;
  wire  _EVAL_746;
  wire  _EVAL_2024;
  wire  _EVAL_1882;
  wire  _EVAL_1897;
  wire  _EVAL_1835;
  wire  _EVAL_1262;
  wire  _EVAL_1718;
  wire  _EVAL_2009;
  wire  _EVAL_282;
  wire  _EVAL_1655;
  wire  _EVAL_1214;
  wire  _EVAL_1945;
  wire  _EVAL_938;
  wire  _EVAL_2042;
  wire  _EVAL_2052;
  wire  _EVAL_1445;
  wire  _EVAL_684;
  wire  _EVAL_829;
  wire  _EVAL_2120;
  wire  _EVAL_425;
  wire  _EVAL_754;
  wire  _EVAL_1809;
  wire  _EVAL_1529;
  wire  _EVAL_493;
  wire  _EVAL_1734;
  wire  _EVAL_977;
  wire  _EVAL_974;
  wire  _EVAL_1575;
  wire  _EVAL_802;
  wire  _EVAL_601;
  wire  _EVAL_479;
  wire  _EVAL_1016;
  wire  _EVAL_890;
  wire  _EVAL_1236;
  wire  _EVAL_1468;
  wire  _EVAL_430;
  wire  _EVAL_893;
  wire  _EVAL_235;
  wire  _EVAL_748;
  wire  _EVAL_178;
  wire  _EVAL_1619;
  wire  _EVAL_821;
  wire  _EVAL_730;
  wire  _EVAL_424;
  wire  _EVAL_163;
  wire  _EVAL_2135;
  wire  _EVAL_1623;
  wire  _EVAL_1181;
  wire  _EVAL_1170;
  wire  _EVAL_1868;
  wire  _EVAL_1816;
  wire  _EVAL_288;
  wire  _EVAL_343;
  wire  _EVAL_1287;
  wire  _EVAL_582;
  wire  _EVAL_2043;
  wire  _EVAL_775;
  wire  _EVAL_2171;
  wire  _EVAL_1967;
  wire  _EVAL_1321;
  wire  _EVAL_624;
  wire  _EVAL_572;
  wire  _EVAL_1907;
  wire  _EVAL_2007;
  wire  _EVAL_1514;
  wire  _EVAL_791;
  wire  _EVAL_1679;
  wire  _EVAL_996;
  wire  _EVAL_497;
  wire  _EVAL_765;
  wire  _EVAL_1431;
  wire  _EVAL_947;
  wire  _EVAL_1513;
  wire  _EVAL_2189;
  wire  _EVAL_146;
  wire  _EVAL_1620;
  wire  _EVAL_226;
  wire  _EVAL_1666;
  wire  _EVAL_184;
  wire  _EVAL_1778;
  wire  _EVAL_661;
  wire  _EVAL_1165;
  wire  _EVAL_2196;
  wire  _EVAL_1999;
  wire  _EVAL_604;
  wire  _EVAL_132;
  wire  _EVAL_1332;
  wire  _EVAL_1586;
  wire  _EVAL_1525;
  wire  _EVAL_1849;
  wire  _EVAL_1033;
  wire  _EVAL_717;
  wire  _EVAL_176;
  wire  _EVAL_397;
  wire  _EVAL_1333;
  wire  _EVAL_1576;
  wire  _EVAL_1661;
  wire  _EVAL_640;
  wire  _EVAL_960;
  wire  _EVAL_937;
  wire  _EVAL_549;
  wire  _EVAL_832;
  wire  _EVAL_1507;
  wire  _EVAL_243;
  wire  _EVAL_308;
  wire  _EVAL_2207;
  wire  _EVAL_1150;
  wire  _EVAL_725;
  wire  _EVAL_711;
  wire  _EVAL_231;
  wire  _EVAL_1568;
  wire  _EVAL_427;
  wire  _EVAL_675;
  wire  _EVAL_1759;
  wire  _EVAL_1624;
  wire  _EVAL_426;
  wire  _EVAL_97;
  wire  _EVAL_1255;
  wire  _EVAL_991;
  wire  _EVAL_1373;
  wire  _EVAL_1875;
  wire  _EVAL_584;
  wire  _EVAL_676;
  wire  _EVAL_161;
  wire  _EVAL_1031;
  wire  _EVAL_1272;
  wire  _EVAL_93;
  wire [10:0] _EVAL_1440;
  wire  _EVAL_238;
  wire  _EVAL_1338;
  wire  _EVAL_429;
  wire  _EVAL_1886;
  wire  _EVAL_982;
  wire  _EVAL_2131;
  wire  _EVAL_1144;
  wire  _EVAL_1453;
  wire  _EVAL_1488;
  wire  _EVAL_2203;
  wire  _EVAL_679;
  wire  _EVAL_2100;
  wire  _EVAL_629;
  wire  _EVAL_1757;
  wire  _EVAL_983;
  wire  _EVAL_242;
  wire  _EVAL_1613;
  wire  _EVAL_1924;
  wire  _EVAL_267;
  wire  _EVAL_1364;
  wire  _EVAL_956;
  wire  _EVAL_999;
  wire  _EVAL_419;
  wire  _EVAL_119;
  wire  _EVAL_99;
  wire  _EVAL_1410;
  wire  _EVAL_1259;
  wire  _EVAL_1358;
  wire  _EVAL_944;
  wire  _EVAL_1084;
  wire  _EVAL_1099;
  wire  _EVAL_1342;
  wire  _EVAL_89;
  wire  _EVAL_1217;
  wire  _EVAL_1280;
  wire  _EVAL_1837;
  wire  _EVAL_1110;
  wire  _EVAL_1510;
  wire  _EVAL_812;
  wire  _EVAL_966;
  wire  _EVAL_768;
  wire  _EVAL_448;
  wire  _EVAL_2035;
  wire  _EVAL_1621;
  wire  _EVAL_551;
  wire  _EVAL_1434;
  wire  _EVAL_2061;
  wire  _EVAL_302;
  wire  _EVAL_1063;
  wire  _EVAL_1670;
  wire  _EVAL_1825;
  wire  _EVAL_1481;
  wire  _EVAL_1530;
  wire  _EVAL_2037;
  wire  _EVAL_2053;
  wire  _EVAL_797;
  wire  _EVAL_2008;
  wire  _EVAL_1399;
  wire  _EVAL_271;
  wire  _EVAL_708;
  wire  _EVAL_87;
  wire  _EVAL_759;
  wire  _EVAL_1941;
  wire  _EVAL_917;
  wire  _EVAL_202;
  wire  _EVAL_1817;
  wire  _EVAL_1128;
  wire  _EVAL_932;
  wire  _EVAL_815;
  wire  _EVAL_71;
  wire  _EVAL_995;
  wire  _EVAL_1162;
  wire  _EVAL_1077;
  wire  _EVAL_876;
  wire  _EVAL_2237;
  wire  _EVAL_853;
  wire  _EVAL_1626;
  wire  _EVAL_2049;
  wire  _EVAL_2016;
  wire  _EVAL_2002;
  wire  _EVAL_1574;
  wire  _EVAL_1629;
  wire  _EVAL_304;
  wire  _EVAL_1963;
  wire [11:0] _EVAL_1087;
  wire  _EVAL_998;
  wire  _EVAL_2066;
  wire  _EVAL_2198;
  wire [3:0] _EVAL_2039;
  wire  _EVAL_1899;
  wire  _EVAL_1061;
  wire  _EVAL_1340;
  wire  _EVAL_1673;
  wire  _EVAL_128;
  wire  _EVAL_602;
  wire  _EVAL_1211;
  wire  _EVAL_223;
  wire  _EVAL_2221;
  wire  _EVAL_198;
  wire  _EVAL_412;
  wire  _EVAL_615;
  wire  _EVAL_707;
  wire  _EVAL_851;
  wire  _EVAL_1018;
  wire  _EVAL_1786;
  wire  _EVAL_2119;
  wire  _EVAL_780;
  wire  _EVAL_617;
  wire  _EVAL_1823;
  wire  _EVAL_1761;
  wire  _EVAL_1126;
  wire  _EVAL_1682;
  wire  _EVAL_111;
  wire  _EVAL_1957;
  wire  _EVAL_1660;
  wire  _EVAL_1117;
  wire  _EVAL_2145;
  wire  _EVAL_1026;
  wire  _EVAL_84;
  wire  _EVAL_1846;
  wire  _EVAL_1347;
  wire  _EVAL_2091;
  wire  _EVAL_1378;
  wire  _EVAL_1617;
  wire  _EVAL_1385;
  wire  _EVAL_1348;
  wire  _EVAL_1981;
  wire  _EVAL_1727;
  wire  _EVAL_1974;
  wire  _EVAL_2122;
  wire  _EVAL_1693;
  wire  _EVAL_2063;
  wire  _EVAL_550;
  wire  _EVAL_414;
  wire  _EVAL_1268;
  wire  _EVAL_537;
  wire  _EVAL_340;
  wire  _EVAL_138;
  wire  _EVAL_536;
  wire  _EVAL_963;
  wire  _EVAL_837;
  wire  _EVAL_1382;
  wire  _EVAL_609;
  wire  _EVAL_733;
  wire  _EVAL_1418;
  wire  _EVAL_816;
  wire  _EVAL_400;
  wire  _EVAL_910;
  wire  _EVAL_788;
  wire  _EVAL_1389;
  wire  _EVAL_755;
  wire  _EVAL_1024;
  wire  _EVAL_466;
  wire  _EVAL_1025;
  wire  _EVAL_1651;
  wire  _EVAL_849;
  wire  _EVAL_1650;
  wire  _EVAL_283;
  wire  _EVAL_1290;
  wire  _EVAL_800;
  wire  _EVAL_1235;
  wire  _EVAL_432;
  wire  _EVAL_919;
  wire  _EVAL_2055;
  wire  _EVAL_1585;
  wire  _EVAL_1450;
  wire  _EVAL_2099;
  wire  _EVAL_1118;
  wire  _EVAL_1058;
  wire  _EVAL_1489;
  wire  _EVAL_1983;
  wire  _EVAL_587;
  wire  _EVAL_405;
  wire  _EVAL_698;
  wire  _EVAL_1341;
  wire  _EVAL_586;
  wire  _EVAL_1423;
  wire  _EVAL_265;
  wire  _EVAL_852;
  wire  _EVAL_2121;
  wire  _EVAL_2173;
  wire  _EVAL_1043;
  wire  _EVAL_641;
  wire  _EVAL_1788;
  wire  _EVAL_147;
  wire  _EVAL_1956;
  wire  _EVAL_1550;
  wire  _EVAL_2023;
  wire  _EVAL_1764;
  wire  _EVAL_1876;
  wire  _EVAL_2010;
  wire  _EVAL_1015;
  wire  _EVAL_1663;
  wire  _EVAL_289;
  wire  _EVAL_378;
  wire  _EVAL_563;
  wire  _EVAL_1852;
  wire  _EVAL_1865;
  wire  _EVAL_1712;
  wire  _EVAL_976;
  wire  _EVAL_700;
  wire  _EVAL_683;
  wire  _EVAL_1699;
  wire  _EVAL_1735;
  wire  _EVAL_1763;
  wire  _EVAL_1496;
  wire  _EVAL_1330;
  wire  _EVAL_216;
  wire  _EVAL_1164;
  wire  _EVAL_2183;
  wire  _EVAL_1972;
  wire  _EVAL_183;
  wire  _EVAL_1839;
  wire  _EVAL_984;
  wire  _EVAL_645;
  wire  _EVAL_952;
  wire  _EVAL_1884;
  wire  _EVAL_723;
  wire  _EVAL_2003;
  wire  _EVAL_81;
  wire  _EVAL_1746;
  wire  _EVAL_870;
  wire  _EVAL_2186;
  wire  _EVAL_2072;
  wire  _EVAL_764;
  wire  _EVAL_197;
  wire  _EVAL_421;
  wire  _EVAL_524;
  wire  _EVAL_1395;
  wire  _EVAL_83;
  wire  _EVAL_903;
  wire  _EVAL_2141;
  wire  _EVAL_2074;
  wire  _EVAL_2105;
  wire  _EVAL_1505;
  wire  _EVAL_2142;
  wire  _EVAL_1002;
  wire  _EVAL_1901;
  wire  _EVAL_1728;
  wire  _EVAL_1683;
  wire  _EVAL_474;
  wire  _EVAL_346;
  wire  _EVAL_86;
  wire  _EVAL_394;
  wire  _EVAL_834;
  wire  _EVAL_1713;
  wire  _EVAL_1681;
  wire  _EVAL_1767;
  wire  _EVAL_2223;
  wire  _EVAL_830;
  wire  _EVAL_389;
  wire  _EVAL_258;
  wire  _EVAL_1231;
  wire  _EVAL_239;
  wire  _EVAL_1611;
  wire  _EVAL_638;
  wire  _EVAL_888;
  wire  _EVAL_542;
  wire  _EVAL_1896;
  wire  _EVAL_1891;
  wire  _EVAL_1692;
  wire  _EVAL_1506;
  wire  _EVAL_1848;
  wire  _EVAL_1738;
  wire  _EVAL_605;
  wire  _EVAL_534;
  wire  _EVAL_341;
  wire  _EVAL_413;
  wire  _EVAL_1375;
  wire  _EVAL_1614;
  wire  _EVAL_2040;
  wire  _EVAL_597;
  wire  _EVAL_1351;
  wire  _EVAL_167;
  wire  _EVAL_2078;
  wire  _EVAL_541;
  wire  _EVAL_825;
  wire  _EVAL_2084;
  wire  _EVAL_1437;
  wire  _EVAL_187;
  wire  _EVAL_2098;
  wire  _EVAL_1028;
  wire  _EVAL_2085;
  wire  _EVAL_2149;
  wire  _EVAL_2140;
  wire  _EVAL_1328;
  wire  _EVAL_2028;
  wire  _EVAL_687;
  wire  _EVAL_1895;
  wire  _EVAL_1714;
  wire  _EVAL_1477;
  wire  _EVAL_2050;
  wire  _EVAL_571;
  wire  _EVAL_1498;
  wire  _EVAL_227;
  wire  _EVAL_1223;
  wire  _EVAL_484;
  wire  _EVAL_993;
  wire  _EVAL_1566;
  wire  _EVAL_1600;
  wire  _EVAL_297;
  wire  _EVAL_367;
  wire  _EVAL_1080;
  wire  _EVAL_902;
  wire  _EVAL_1775;
  wire  _EVAL_1871;
  wire  _EVAL_793;
  wire  _EVAL_863;
  wire  _EVAL_158;
  wire  _EVAL_1950;
  wire  _EVAL_252;
  wire  _EVAL_1039;
  wire  _EVAL_535;
  wire  _EVAL_1412;
  wire  _EVAL_626;
  wire  _EVAL_878;
  wire  _EVAL_745;
  wire  _EVAL_1634;
  wire  _EVAL_1934;
  wire  _EVAL_1783;
  wire  _EVAL_2062;
  wire  _EVAL_1186;
  wire  _EVAL_1804;
  wire  _EVAL_2227;
  wire  _EVAL_1365;
  wire  _EVAL_607;
  wire  _EVAL_489;
  wire  _EVAL_1949;
  wire  _EVAL_1224;
  wire  _EVAL_1390;
  wire  _EVAL_78;
  wire  _EVAL_1130;
  wire  _EVAL_1457;
  wire  _EVAL_292;
  wire  _EVAL_1922;
  wire  _EVAL_1587;
  wire  _EVAL_91;
  wire  _EVAL_828;
  wire  _EVAL_206;
  wire  _EVAL_735;
  wire  _EVAL_1733;
  wire  _EVAL_1438;
  wire  _EVAL_691;
  wire  _EVAL_2206;
  wire  _EVAL_891;
  wire  _EVAL_954;
  wire  _EVAL_1515;
  wire  _EVAL_509;
  wire  _EVAL_2175;
  wire  _EVAL_1955;
  wire  _EVAL_1159;
  wire  _EVAL_1674;
  wire  _EVAL_1300;
  wire  _EVAL_1730;
  wire  _EVAL_1883;
  wire  _EVAL_677;
  wire  _EVAL_1910;
  wire  _EVAL_1258;
  wire  _EVAL_520;
  wire  _EVAL_1455;
  wire  _EVAL_1801;
  wire  _EVAL_215;
  wire  _EVAL_1343;
  wire  _EVAL_476;
  wire  _EVAL_1544;
  wire  _EVAL_1408;
  wire  _EVAL_1122;
  wire  _EVAL_720;
  wire  _EVAL_2128;
  wire  _EVAL_76;
  SiFive__EVAL_211_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  SiFive__EVAL_212_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14)
  );
  assign _EVAL_1267 = _EVAL_1582[28:23];
  assign _EVAL_927 = _EVAL_1048 & _EVAL_644;
  assign _EVAL_1151 = _EVAL_631[267];
  assign _EVAL_1497 = _EVAL_927 & _EVAL_1151;
  assign _EVAL_967 = _EVAL_1497 & _EVAL_502;
  assign _EVAL_978 = _EVAL_927 & _EVAL_1760;
  assign _EVAL_2123 = _EVAL_978 & _EVAL_502;
  assign _EVAL_592 = _EVAL_1017 != 8'h0;
  assign _EVAL_2022 = _EVAL_2123 & _EVAL_592;
  assign _EVAL_1102 = _EVAL_927 & _EVAL_1486;
  assign _EVAL_338 = _EVAL_631[271];
  assign _EVAL_280 = _EVAL_749 & _EVAL_338;
  assign _EVAL_294 = _EVAL_280 & _EVAL_502;
  assign _EVAL_1124 = _EVAL_294 & _EVAL_1387;
  assign _EVAL_316 = _EVAL_631[266];
  assign _EVAL_1073 = _EVAL_927 & _EVAL_316;
  assign _EVAL_1444 = _EVAL_1073 & _EVAL_502;
  assign _EVAL_1467 = _EVAL_631[260];
  assign _EVAL_1013 = _EVAL_749 & _EVAL_1467;
  assign _EVAL_1178 = _EVAL_1013 & _EVAL_502;
  assign _EVAL_1978 = _EVAL_1582[31:29];
  assign _EVAL_1220 = _EVAL_1978 != 3'h0;
  assign _EVAL_2107 = _EVAL_749 & _EVAL_1151;
  assign _EVAL_269 = _EVAL_2107 & _EVAL_502;
  assign _EVAL_1521 = _EVAL_269 & _EVAL_758;
  assign _EVAL_494 = _EVAL_927 & _EVAL_886;
  assign _EVAL_973 = _EVAL_494 & _EVAL_502;
  assign _EVAL_250 = _EVAL_1563 != 8'h0;
  assign _EVAL_850 = _EVAL_973 & _EVAL_250;
  assign _EVAL_1723 = _EVAL_631[259];
  assign _EVAL_1336 = _EVAL_749 & _EVAL_1723;
  assign _EVAL_689 = _EVAL_1336 & _EVAL_502;
  assign _EVAL_951 = _EVAL_689 & _EVAL_1638;
  assign _EVAL_564 = _EVAL_631[270];
  assign _EVAL_102 = _EVAL_927 & _EVAL_564;
  assign _EVAL_1792 = _EVAL_102 & _EVAL_502;
  assign _EVAL_525 = _EVAL_1421[17];
  assign _EVAL_1676 = _EVAL_1303 & _EVAL_525;
  assign _EVAL_2124 = _EVAL_1676 & _EVAL_680;
  assign _EVAL_1143 = _EVAL_1582[6];
  assign _EVAL_402 = _EVAL_2124 & _EVAL_1143;
  assign _EVAL_456 = _EVAL_1303 & _EVAL_299;
  assign _EVAL_1027 = _EVAL_456 & _EVAL_680;
  assign _EVAL_1539 = _EVAL_1582[3:0];
  assign _EVAL_2064 = _EVAL_1539 != 4'h0;
  assign _EVAL_546 = _EVAL_1027 & _EVAL_2064;
  assign _EVAL_2065 = _EVAL_927 & _EVAL_637;
  assign _EVAL_1149 = _EVAL_2065 & _EVAL_502;
  assign _EVAL_154 = _EVAL_1149 & _EVAL_592;
  assign _EVAL_939 = _EVAL_1582[11];
  assign _EVAL_798 = _EVAL_328 & _EVAL_939;
  assign _EVAL_844 = _EVAL_927 & _EVAL_1845;
  assign _EVAL_578 = _EVAL_844 & _EVAL_502;
  assign _EVAL_1030 = _EVAL_190 != 10'h0;
  assign _EVAL_946 = _EVAL_578 & _EVAL_1030;
  assign _EVAL_1705 = _EVAL_927 & _EVAL_1188;
  assign _EVAL_2132 = _EVAL_927 & _EVAL_469;
  assign _EVAL_1645 = _EVAL_2132 & _EVAL_502;
  assign _EVAL_922 = _EVAL_1645 & _EVAL_592;
  assign _EVAL_1748 = _EVAL_1582[15:1];
  assign _EVAL_1142 = _EVAL_1748 == 15'h7fff;
  assign _EVAL_275 = _EVAL_631[262];
  assign _EVAL_1109 = _EVAL_749 & _EVAL_275;
  assign _EVAL_2213 = _EVAL_1109 & _EVAL_502;
  assign _EVAL_2176 = _EVAL_2213 & _EVAL_175;
  assign _EVAL_926 = _EVAL_927 & _EVAL_1391;
  assign _EVAL_1784 = _EVAL_927 & _EVAL_129;
  assign _EVAL_1106 = _EVAL_1421[18];
  assign _EVAL_1172 = _EVAL_1303 & _EVAL_1106;
  assign _EVAL_1689 = _EVAL_1172 & _EVAL_680;
  assign _EVAL_599 = _EVAL_1582[15:12];
  assign _EVAL_58 = _EVAL_599 != 4'h0;
  assign _EVAL_510 = _EVAL_1689 & _EVAL_58;
  assign _EVAL_1168 = _EVAL_1582[28:24];
  assign _EVAL_1278 = _EVAL_1168 == 5'h1f;
  assign _EVAL_1552 = _EVAL_328 & _EVAL_1278;
  assign _EVAL_499 = _EVAL_631[264];
  assign _EVAL_134 = _EVAL_749 & _EVAL_499;
  assign _EVAL_1369 = _EVAL_134 & _EVAL_502;
  assign _EVAL_2168 = _EVAL_1369 & _EVAL_175;
  assign _EVAL_1601 = _EVAL_631[257];
  assign _EVAL_2231 = _EVAL_749 & _EVAL_1601;
  assign _EVAL_1867 = _EVAL_2231 & _EVAL_502;
  assign _EVAL_762 = _EVAL_1867 & _EVAL_1387;
  assign _EVAL_1647 = _EVAL_927 & _EVAL_172;
  assign _EVAL_2005 = _EVAL_1647 & _EVAL_502;
  assign _EVAL_526 = _EVAL_573 != 8'h0;
  assign _EVAL_1035 = _EVAL_2005 & _EVAL_526;
  assign _EVAL_1075 = _EVAL_1784 & _EVAL_502;
  assign _EVAL_477 = _EVAL_1753 != 8'h0;
  assign _EVAL_1388 = _EVAL_2123 & _EVAL_477;
  assign _EVAL_997 = _EVAL_2224 == 1'h0;
  assign _EVAL_2193 = _EVAL_599 == 4'hf;
  assign _EVAL_1208 = {{1'd0}, _EVAL_616};
  assign _EVAL_286 = _EVAL_1582[12];
  assign _EVAL_1659 = _EVAL_927 & _EVAL_275;
  assign _EVAL_807 = _EVAL_1659 & _EVAL_502;
  assign _EVAL_1355 = _EVAL_807 & _EVAL_250;
  assign _EVAL_911 = _EVAL_1421[0];
  assign _EVAL_1203 = _EVAL_2076 & _EVAL_911;
  assign _EVAL_1527 = _EVAL_1203 & _EVAL_311;
  assign _EVAL_2209 = _EVAL_631[256];
  assign _EVAL_972 = _EVAL_749 & _EVAL_2209;
  assign _EVAL_2143 = _EVAL_972 & _EVAL_502;
  assign _EVAL_1559 = _EVAL_927 & _EVAL_1987;
  assign _EVAL_337 = _EVAL_1559 & _EVAL_502;
  assign _EVAL_2151 = _EVAL_337 & _EVAL_250;
  assign _EVAL_1032 = _EVAL_927 & _EVAL_2079;
  assign _EVAL_1228 = _EVAL_631[269];
  assign _EVAL_365 = _EVAL_927 & _EVAL_1228;
  assign _EVAL_674 = _EVAL_365 & _EVAL_502;
  assign _EVAL_842 = _EVAL_674 & _EVAL_592;
  assign _EVAL_314 = _EVAL_631[263];
  assign _EVAL_1937 = _EVAL_631[0];
  assign _EVAL_1779 = _EVAL_749 & _EVAL_1937;
  assign _EVAL_1363 = _EVAL_1779 & _EVAL_1441;
  assign _EVAL_1557 = _EVAL_1363 & _EVAL_758;
  assign _EVAL_1289 = _EVAL_926 & _EVAL_502;
  assign _EVAL_150 = _EVAL_1027 & _EVAL_286;
  assign _EVAL_585 = _EVAL_1705 & _EVAL_502;
  assign _EVAL_396 = _EVAL_585 & _EVAL_477;
  assign _EVAL_369 = _EVAL_1303 & _EVAL_989;
  assign _EVAL_379 = _EVAL_369 & _EVAL_680;
  assign _EVAL_913 = _EVAL_1582[11:5];
  assign _EVAL_580 = _EVAL_913 != 7'h0;
  assign _EVAL_1442 = _EVAL_379 & _EVAL_580;
  assign _EVAL_249 = _EVAL_1582[21:20];
  assign _EVAL_1553 = _EVAL_249 == 2'h3;
  assign _EVAL_1894 = _EVAL_749 & _EVAL_316;
  assign _EVAL_1288 = _EVAL_1894 & _EVAL_502;
  assign _EVAL_2188 = _EVAL_1303 & _EVAL_911;
  assign _EVAL_1202 = _EVAL_2188 & _EVAL_311;
  assign _EVAL_949 = _EVAL_631[268];
  assign _EVAL_1802 = _EVAL_927 & _EVAL_949;
  assign _EVAL_1426 = _EVAL_1802 & _EVAL_502;
  assign _EVAL_1684 = _EVAL_1426 & _EVAL_477;
  assign _EVAL_2180 = _EVAL_631[258];
  assign _EVAL_595 = _EVAL_927 & _EVAL_2180;
  assign _EVAL_2083 = _EVAL_631[265];
  assign _EVAL_1913 = _EVAL_1582[7:4];
  assign _EVAL_2033 = _EVAL_1913 != 4'h0;
  assign _EVAL_931 = _EVAL_1027 & _EVAL_2033;
  assign _EVAL_1625 = _EVAL_749 & _EVAL_2180;
  assign _EVAL_1519 = _EVAL_1625 & _EVAL_502;
  assign _EVAL_992 = _EVAL_1519 & _EVAL_1387;
  assign _EVAL_1281 = _EVAL_927 & _EVAL_2083;
  assign _EVAL_1675 = _EVAL_1281 & _EVAL_502;
  assign _EVAL_1257 = _EVAL_927 & _EVAL_499;
  assign _EVAL_1526 = _EVAL_1257 & _EVAL_502;
  assign _EVAL_2089 = _EVAL_1526 & _EVAL_526;
  assign _EVAL_1097 = _EVAL_927 & _EVAL_1534;
  assign _EVAL_664 = _EVAL_1097 & _EVAL_502;
  assign _EVAL_1828 = _EVAL_664 & _EVAL_526;
  assign _EVAL_2112 = _EVAL_1913 == 4'hf;
  assign _EVAL_1248 = _EVAL_328 & _EVAL_2112;
  assign _EVAL_746 = _EVAL_631[275];
  assign _EVAL_2024 = _EVAL_749 & _EVAL_746;
  assign _EVAL_1882 = _EVAL_2024 & _EVAL_502;
  assign _EVAL_1897 = _EVAL_1882 & _EVAL_175;
  assign _EVAL_1835 = _EVAL_1971 == 1'h0;
  assign _EVAL_1262 = _EVAL_1835 & _EVAL_997;
  assign _EVAL_1718 = _EVAL_1262 & _EVAL_555;
  assign _EVAL_2009 = _EVAL_1718 & _EVAL_2222;
  assign _EVAL_282 = _EVAL_2143 & _EVAL_1387;
  assign _EVAL_1655 = _EVAL_927 & _EVAL_338;
  assign _EVAL_1214 = _EVAL_1655 & _EVAL_502;
  assign _EVAL_1945 = _EVAL_1214 & _EVAL_526;
  assign _EVAL_938 = _EVAL_749 & _EVAL_2083;
  assign _EVAL_2042 = _EVAL_749 & _EVAL_314;
  assign _EVAL_2052 = _EVAL_2042 & _EVAL_502;
  assign _EVAL_1445 = _EVAL_2052 & _EVAL_1638;
  assign _EVAL_684 = _EVAL_749 & _EVAL_1228;
  assign _EVAL_829 = _EVAL_684 & _EVAL_502;
  assign _EVAL_2120 = _EVAL_829 & _EVAL_1638;
  assign _EVAL_425 = sb2tlOpt__EVAL_11 | sb2tlOpt__EVAL_25;
  assign _EVAL_754 = _EVAL_425 & _EVAL_1997;
  assign _EVAL_1809 = _EVAL_754 & _EVAL_1806;
  assign _EVAL_1529 = _EVAL_425 & _EVAL_1147;
  assign _EVAL_493 = _EVAL_1529 & _EVAL_1806;
  assign _EVAL_1734 = _EVAL_631[274];
  assign _EVAL_977 = _EVAL_927 & _EVAL_1734;
  assign _EVAL_974 = _EVAL_977 & _EVAL_502;
  assign _EVAL_1575 = _EVAL_974 & _EVAL_592;
  assign _EVAL_802 = _EVAL_11 == 1'h0;
  assign _EVAL_601 = _EVAL_2222 == 1'h0;
  assign _EVAL_479 = _EVAL_802 | _EVAL_601;
  assign _EVAL_1016 = _EVAL_744 != 16'h0;
  assign _EVAL_890 = _EVAL_927 & _EVAL_1429;
  assign _EVAL_1236 = _EVAL_890 & _EVAL_502;
  assign _EVAL_1468 = _EVAL_1236 & _EVAL_526;
  assign _EVAL_430 = _EVAL_631[207];
  assign _EVAL_893 = _EVAL_749 & _EVAL_430;
  assign _EVAL_235 = _EVAL_927 & _EVAL_1937;
  assign _EVAL_748 = _EVAL_927 & _EVAL_1210;
  assign _EVAL_178 = _EVAL_748 & _EVAL_502;
  assign _EVAL_1619 = _EVAL_1582[4];
  assign _EVAL_821 = _EVAL_379 & _EVAL_1619;
  assign _EVAL_730 = _EVAL_967 & _EVAL_477;
  assign _EVAL_424 = _EVAL_1303 & _EVAL_1902;
  assign _EVAL_163 = _EVAL_424 & _EVAL_680;
  assign _EVAL_2135 = _EVAL_1748 != 15'h0;
  assign _EVAL_1623 = _EVAL_163 & _EVAL_2135;
  assign _EVAL_1181 = _EVAL_2052 & _EVAL_1387;
  assign _EVAL_1170 = _EVAL_595 & _EVAL_502;
  assign _EVAL_1868 = _EVAL_1170 & _EVAL_526;
  assign _EVAL_1816 = _EVAL_1149 & _EVAL_477;
  assign _EVAL_288 = _EVAL_631[272];
  assign _EVAL_343 = _EVAL_749 & _EVAL_288;
  assign _EVAL_1287 = _EVAL_343 & _EVAL_502;
  assign _EVAL_582 = _EVAL_1287 & _EVAL_1387;
  assign _EVAL_2043 = _EVAL_822 & _EVAL_1142;
  assign _EVAL_775 = _EVAL_1582[5];
  assign _EVAL_2171 = _EVAL_2124 & _EVAL_775;
  assign _EVAL_1967 = _EVAL_2143 & _EVAL_175;
  assign _EVAL_1321 = _EVAL_2124 & _EVAL_349;
  assign _EVAL_624 = _EVAL_749 & _EVAL_949;
  assign _EVAL_572 = _EVAL_927 & _EVAL_288;
  assign _EVAL_1907 = _EVAL_572 & _EVAL_502;
  assign _EVAL_2007 = _EVAL_1907 & _EVAL_592;
  assign _EVAL_1514 = _EVAL_664 & _EVAL_477;
  assign _EVAL_791 = _EVAL_379 & _EVAL_1517;
  assign _EVAL_1679 = _EVAL_2123 & _EVAL_250;
  assign _EVAL_996 = _EVAL_1645 & _EVAL_477;
  assign _EVAL_497 = _EVAL_1214 & _EVAL_250;
  assign _EVAL_765 = _EVAL_927 & _EVAL_2209;
  assign _EVAL_1431 = _EVAL_765 & _EVAL_502;
  assign _EVAL_947 = _EVAL_1431 & _EVAL_250;
  assign _EVAL_1513 = _EVAL_1075 & _EVAL_1030;
  assign _EVAL_2189 = _EVAL_749 & _EVAL_564;
  assign _EVAL_146 = _EVAL_2189 & _EVAL_502;
  assign _EVAL_1620 = _EVAL_146 & _EVAL_1387;
  assign _EVAL_226 = _EVAL_749 & _EVAL_1734;
  assign _EVAL_1666 = _EVAL_226 & _EVAL_502;
  assign _EVAL_184 = _EVAL_1666 & _EVAL_175;
  assign _EVAL_1778 = _EVAL_631[276];
  assign _EVAL_661 = _EVAL_927 & _EVAL_1778;
  assign _EVAL_1165 = _EVAL_661 & _EVAL_502;
  assign _EVAL_2196 = _EVAL_1165 & _EVAL_526;
  assign _EVAL_1999 = _EVAL_829 & _EVAL_1387;
  assign _EVAL_604 = _EVAL_631[273];
  assign _EVAL_132 = _EVAL_927 & _EVAL_604;
  assign _EVAL_1332 = _EVAL_132 & _EVAL_502;
  assign _EVAL_1586 = _EVAL_1332 & _EVAL_592;
  assign _EVAL_1525 = _EVAL_425 & _EVAL_2011;
  assign _EVAL_1849 = _EVAL_249 != 2'h0;
  assign _EVAL_1033 = _EVAL_2124 & _EVAL_1849;
  assign _EVAL_717 = _EVAL_1421[19];
  assign _EVAL_176 = _EVAL_1303 & _EVAL_717;
  assign _EVAL_397 = _EVAL_1645 & _EVAL_526;
  assign _EVAL_1333 = _EVAL_1289 & _EVAL_526;
  assign _EVAL_1576 = _EVAL_2076 & _EVAL_525;
  assign _EVAL_1661 = _EVAL_1576 & _EVAL_680;
  assign _EVAL_640 = _EVAL_1582[18];
  assign _EVAL_960 = _EVAL_1661 & _EVAL_640;
  assign _EVAL_937 = _EVAL_927 & _EVAL_1601;
  assign _EVAL_549 = _EVAL_937 & _EVAL_502;
  assign _EVAL_832 = _EVAL_1582[19];
  assign _EVAL_1507 = _EVAL_2124 & _EVAL_832;
  assign _EVAL_243 = _EVAL_425 & _EVAL_1113;
  assign _EVAL_308 = _EVAL_243 & _EVAL_1806;
  assign _EVAL_2207 = _EVAL_308 & _EVAL_179;
  assign _EVAL_1150 = _EVAL_1178 & _EVAL_175;
  assign _EVAL_725 = _EVAL_973 & _EVAL_477;
  assign _EVAL_711 = _EVAL_1582[7];
  assign _EVAL_231 = _EVAL_2124 & _EVAL_711;
  assign _EVAL_1568 = _EVAL_1675 & _EVAL_526;
  assign _EVAL_427 = _EVAL_1426 & _EVAL_526;
  assign _EVAL_675 = _EVAL_589 | _EVAL_30;
  assign _EVAL_1759 = _EVAL_675 == 1'h0;
  assign _EVAL_1624 = _EVAL_1582[8];
  assign _EVAL_426 = _EVAL_1661 & _EVAL_1624;
  assign _EVAL_97 = _EVAL_1214 & _EVAL_477;
  assign _EVAL_1255 = _EVAL_1288 & _EVAL_175;
  assign _EVAL_991 = _EVAL_2005 & _EVAL_592;
  assign _EVAL_1373 = _EVAL_631[206];
  assign _EVAL_1875 = _EVAL_749 & _EVAL_1373;
  assign _EVAL_584 = _EVAL_1875 & _EVAL_502;
  assign _EVAL_676 = _EVAL_2123 & _EVAL_526;
  assign _EVAL_161 = _EVAL_1426 & _EVAL_592;
  assign _EVAL_1031 = _EVAL_927 & _EVAL_1723;
  assign _EVAL_1272 = _EVAL_1031 & _EVAL_502;
  assign _EVAL_93 = _EVAL_1272 & _EVAL_250;
  assign _EVAL_1440 = _EVAL_1582[23:13];
  assign _EVAL_238 = _EVAL_1440 == 11'h7ff;
  assign _EVAL_1338 = _EVAL_328 & _EVAL_238;
  assign _EVAL_429 = _EVAL_1661 & _EVAL_349;
  assign _EVAL_1886 = _EVAL_927 & _EVAL_1789;
  assign _EVAL_982 = _EVAL_1886 & _EVAL_502;
  assign _EVAL_2131 = _EVAL_982 & _EVAL_250;
  assign _EVAL_1144 = _EVAL_585 & _EVAL_250;
  assign _EVAL_1453 = _EVAL_749 & _EVAL_1778;
  assign _EVAL_1488 = _EVAL_1453 & _EVAL_502;
  assign _EVAL_2203 = _EVAL_1582[9];
  assign _EVAL_679 = _EVAL_2124 & _EVAL_2203;
  assign _EVAL_2100 = _EVAL_2143 & _EVAL_1638;
  assign _EVAL_629 = _EVAL_938 & _EVAL_502;
  assign _EVAL_1757 = _EVAL_629 & _EVAL_1387;
  assign _EVAL_983 = _EVAL_1582[13];
  assign _EVAL_242 = _EVAL_1661 & _EVAL_983;
  assign _EVAL_1613 = _EVAL_979 & _EVAL_1870;
  assign _EVAL_1924 = _EVAL_927 & _EVAL_1467;
  assign _EVAL_267 = _EVAL_1924 & _EVAL_502;
  assign _EVAL_1364 = _EVAL_379 & _EVAL_1220;
  assign _EVAL_956 = _EVAL_1666 & _EVAL_1638;
  assign _EVAL_999 = _EVAL_674 & _EVAL_250;
  assign _EVAL_419 = _EVAL_1170 & _EVAL_477;
  assign _EVAL_119 = _EVAL_1526 & _EVAL_477;
  assign _EVAL_99 = _EVAL_2076 & _EVAL_717;
  assign _EVAL_1410 = _EVAL_1440 != 11'h0;
  assign _EVAL_1259 = _EVAL_893 & _EVAL_502;
  assign _EVAL_1358 = _EVAL_624 & _EVAL_502;
  assign _EVAL_944 = _EVAL_1358 & _EVAL_1638;
  assign _EVAL_1084 = _EVAL_927 & _EVAL_498;
  assign _EVAL_1099 = _EVAL_1084 & _EVAL_502;
  assign _EVAL_1342 = _EVAL_178 & _EVAL_477;
  assign _EVAL_89 = _EVAL_1202 & _EVAL_2178;
  assign _EVAL_1217 = _EVAL_163 & _EVAL_1016;
  assign _EVAL_1280 = _EVAL_629 & _EVAL_1638;
  assign _EVAL_1837 = _EVAL_1829 == 1'h0;
  assign _EVAL_1110 = _EVAL_1303 & _EVAL_568;
  assign _EVAL_1510 = _EVAL_1110 & _EVAL_680;
  assign _EVAL_812 = _EVAL_267 & _EVAL_250;
  assign _EVAL_966 = _EVAL_1236 & _EVAL_250;
  assign _EVAL_768 = _EVAL_1582[10];
  assign _EVAL_448 = _EVAL_1289 & _EVAL_250;
  assign _EVAL_2035 = _EVAL_927 & _EVAL_746;
  assign _EVAL_1621 = _EVAL_332 != 32'h0;
  assign _EVAL_551 = _EVAL_1527 & _EVAL_214;
  assign _EVAL_1434 = _EVAL_927 & _EVAL_1373;
  assign _EVAL_2061 = _EVAL_1434 & _EVAL_502;
  assign _EVAL_302 = _EVAL_2061 & _EVAL_1621;
  assign _EVAL_1063 = _EVAL_1358 & _EVAL_175;
  assign _EVAL_1670 = _EVAL_1661 & _EVAL_939;
  assign _EVAL_1825 = _EVAL_1102 & _EVAL_502;
  assign _EVAL_1481 = _EVAL_1825 & _EVAL_250;
  assign _EVAL_1530 = _EVAL_749 & _EVAL_604;
  assign _EVAL_2037 = _EVAL_1530 & _EVAL_502;
  assign _EVAL_2053 = _EVAL_2037 & _EVAL_1387;
  assign _EVAL_797 = _EVAL_549 & _EVAL_526;
  assign _EVAL_2008 = _EVAL_629 & _EVAL_758;
  assign _EVAL_1399 = _EVAL_1661 & _EVAL_1517;
  assign _EVAL_271 = _EVAL_967 & _EVAL_250;
  assign _EVAL_708 = _EVAL_267 & _EVAL_526;
  assign _EVAL_87 = _EVAL_332 == 32'hffffffff;
  assign _EVAL_759 = _EVAL_2143 & _EVAL_758;
  assign _EVAL_1941 = _EVAL_99 & _EVAL_680;
  assign _EVAL_917 = _EVAL_2035 & _EVAL_502;
  assign _EVAL_202 = _EVAL_917 & _EVAL_592;
  assign _EVAL_1817 = _EVAL_1892 != 3'h0;
  assign _EVAL_1128 = _EVAL_1027 & _EVAL_1817;
  assign _EVAL_932 = _EVAL_927 & _EVAL_2095;
  assign _EVAL_815 = _EVAL_1867 & _EVAL_758;
  assign _EVAL_71 = _EVAL_2124 & _EVAL_2064;
  assign _EVAL_995 = _EVAL_932 & _EVAL_502;
  assign _EVAL_1162 = _EVAL_927 & _EVAL_57;
  assign _EVAL_1077 = _EVAL_176 & _EVAL_680;
  assign _EVAL_876 = _EVAL_1077 & _EVAL_2178;
  assign _EVAL_2237 = _EVAL_967 & _EVAL_526;
  assign _EVAL_853 = _EVAL_917 & _EVAL_250;
  assign _EVAL_1626 = _EVAL_631[261];
  assign _EVAL_2049 = _EVAL_749 & _EVAL_1626;
  assign _EVAL_2016 = _EVAL_2049 & _EVAL_502;
  assign _EVAL_2002 = _EVAL_2016 & _EVAL_175;
  assign _EVAL_1574 = _EVAL_927 & _EVAL_2200;
  assign _EVAL_1629 = _EVAL_1574 & _EVAL_502;
  assign _EVAL_304 = _EVAL_1629 & _EVAL_1030;
  assign _EVAL_1963 = _EVAL_337 & _EVAL_526;
  assign _EVAL_1087 = _EVAL_1582[11:0];
  assign _EVAL_998 = _EVAL_1488 & _EVAL_175;
  assign _EVAL_2066 = _EVAL_1582[3];
  assign _EVAL_2198 = _EVAL_979 & _EVAL_2066;
  assign _EVAL_2039 = _EVAL_1582[23:20];
  assign _EVAL_1899 = _EVAL_2039 != 4'h0;
  assign _EVAL_1061 = _EVAL_1689 & _EVAL_1899;
  assign _EVAL_1340 = _EVAL_1267 == 6'h3f;
  assign _EVAL_1673 = _EVAL_979 & _EVAL_1340;
  assign _EVAL_128 = _EVAL_927 & _EVAL_1082;
  assign _EVAL_602 = _EVAL_128 & _EVAL_502;
  assign _EVAL_1211 = _EVAL_602 & _EVAL_477;
  assign _EVAL_223 = _EVAL_629 & _EVAL_175;
  assign _EVAL_2221 = _EVAL_674 & _EVAL_526;
  assign _EVAL_198 = _EVAL_1792 & _EVAL_250;
  assign _EVAL_412 = _EVAL_1829 & _EVAL_616;
  assign _EVAL_615 = _EVAL_1162 & _EVAL_502;
  assign _EVAL_707 = _EVAL_615 & _EVAL_477;
  assign _EVAL_851 = _EVAL_1689 & _EVAL_588;
  assign _EVAL_1018 = _EVAL_1661 & _EVAL_768;
  assign _EVAL_1786 = _EVAL_995 & _EVAL_250;
  assign _EVAL_2119 = _EVAL_1363 & _EVAL_1638;
  assign _EVAL_780 = _EVAL_927 & _EVAL_430;
  assign _EVAL_617 = _EVAL_780 & _EVAL_502;
  assign _EVAL_1823 = _EVAL_617 & _EVAL_1621;
  assign _EVAL_1761 = _EVAL_631[192];
  assign _EVAL_1126 = _EVAL_1661 & _EVAL_775;
  assign _EVAL_1682 = _EVAL_1165 & _EVAL_477;
  assign _EVAL_111 = _EVAL_1444 & _EVAL_592;
  assign _EVAL_1957 = _EVAL_1582[14];
  assign _EVAL_1660 = _EVAL_1661 & _EVAL_1957;
  assign _EVAL_1117 = _EVAL_549 & _EVAL_250;
  assign _EVAL_2145 = _EVAL_2016 & _EVAL_758;
  assign _EVAL_1026 = _EVAL_927 & _EVAL_314;
  assign _EVAL_84 = _EVAL_1026 & _EVAL_502;
  assign _EVAL_1846 = _EVAL_84 & _EVAL_250;
  assign _EVAL_1347 = _EVAL_1907 & _EVAL_250;
  assign _EVAL_2091 = _EVAL_1369 & _EVAL_1638;
  assign _EVAL_1378 = _EVAL_749 & _EVAL_1761;
  assign _EVAL_1617 = _EVAL_1378 & _EVAL_502;
  assign _EVAL_1385 = _EVAL_1907 & _EVAL_526;
  assign _EVAL_1348 = _EVAL_1236 & _EVAL_592;
  assign _EVAL_1981 = _EVAL_1978 == 3'h7;
  assign _EVAL_1727 = _EVAL_1519 & _EVAL_1638;
  assign _EVAL_1974 = _EVAL_927 & _EVAL_1761;
  assign _EVAL_2122 = _EVAL_328 & _EVAL_286;
  assign _EVAL_1693 = _EVAL_1582[1];
  assign _EVAL_2063 = _EVAL_979 & _EVAL_1693;
  assign _EVAL_550 = _EVAL_2076 & _EVAL_1106;
  assign _EVAL_414 = _EVAL_550 & _EVAL_680;
  assign _EVAL_1268 = _EVAL_927 & _EVAL_1626;
  assign _EVAL_537 = _EVAL_664 & _EVAL_592;
  assign _EVAL_340 = _EVAL_1431 & _EVAL_592;
  assign _EVAL_138 = _EVAL_1617 & _EVAL_87;
  assign _EVAL_536 = _EVAL_1267 != 6'h0;
  assign _EVAL_963 = _EVAL_2016 & _EVAL_1638;
  assign _EVAL_837 = _EVAL_1027 & _EVAL_939;
  assign _EVAL_1382 = _EVAL_1099 & _EVAL_592;
  assign _EVAL_609 = _EVAL_1303 & _EVAL_361;
  assign _EVAL_733 = _EVAL_84 & _EVAL_526;
  assign _EVAL_1418 = _EVAL_1168 != 5'h0;
  assign _EVAL_816 = _EVAL_664 & _EVAL_250;
  assign _EVAL_400 = _EVAL_2037 & _EVAL_1638;
  assign _EVAL_910 = _EVAL_178 & _EVAL_250;
  assign _EVAL_788 = _EVAL_414 & _EVAL_2193;
  assign _EVAL_1389 = _EVAL_146 & _EVAL_1638;
  assign _EVAL_755 = _EVAL_1525 & _EVAL_1806;
  assign _EVAL_1024 = _EVAL_1526 & _EVAL_250;
  assign _EVAL_466 = _EVAL_674 & _EVAL_477;
  assign _EVAL_1025 = _EVAL_1666 & _EVAL_758;
  assign _EVAL_1651 = _EVAL_1661 & _EVAL_1143;
  assign _EVAL_849 = _EVAL_163 & _EVAL_1870;
  assign _EVAL_1650 = _EVAL_609 & _EVAL_680;
  assign _EVAL_283 = _EVAL_1650 & _EVAL_2178;
  assign _EVAL_1290 = _EVAL_294 & _EVAL_758;
  assign _EVAL_800 = _EVAL_1526 & _EVAL_592;
  assign _EVAL_1235 = _EVAL_973 & _EVAL_592;
  assign _EVAL_432 = _EVAL_2124 & _EVAL_1957;
  assign _EVAL_919 = _EVAL_1444 & _EVAL_477;
  assign _EVAL_2055 = _EVAL_1867 & _EVAL_175;
  assign _EVAL_1585 = _EVAL_269 & _EVAL_175;
  assign _EVAL_1450 = _EVAL_1882 & _EVAL_758;
  assign _EVAL_2099 = _EVAL_1661 & _EVAL_1553;
  assign _EVAL_1118 = _EVAL_1236 & _EVAL_477;
  assign _EVAL_1058 = _EVAL_1792 & _EVAL_592;
  assign _EVAL_1489 = _EVAL_1032 & _EVAL_502;
  assign _EVAL_1983 = _EVAL_1268 & _EVAL_502;
  assign _EVAL_587 = _EVAL_1983 & _EVAL_477;
  assign _EVAL_405 = _EVAL_479 | _EVAL_555;
  assign _EVAL_698 = _EVAL_405 | _EVAL_30;
  assign _EVAL_1341 = _EVAL_698 == 1'h0;
  assign _EVAL_586 = _EVAL_1867 & _EVAL_1638;
  assign _EVAL_1423 = _EVAL_979 & _EVAL_1981;
  assign _EVAL_265 = _EVAL_379 & _EVAL_1693;
  assign _EVAL_852 = _EVAL_1178 & _EVAL_1638;
  assign _EVAL_2121 = _EVAL_703 == 1'h0;
  assign _EVAL_2173 = _EVAL_178 & _EVAL_526;
  assign _EVAL_1043 = _EVAL_2124 & _EVAL_286;
  assign _EVAL_641 = _EVAL_1272 & _EVAL_477;
  assign _EVAL_1788 = _EVAL_1332 & _EVAL_526;
  assign _EVAL_147 = _EVAL_2052 & _EVAL_175;
  assign _EVAL_1956 = _EVAL_2052 & _EVAL_758;
  assign _EVAL_1550 = _EVAL_1027 & _EVAL_1418;
  assign _EVAL_2023 = _EVAL_1358 & _EVAL_758;
  assign _EVAL_1764 = _EVAL_1170 & _EVAL_250;
  assign _EVAL_1876 = _EVAL_1178 & _EVAL_758;
  assign _EVAL_2010 = _EVAL_2213 & _EVAL_1387;
  assign _EVAL_1015 = _EVAL_1582[21];
  assign _EVAL_1663 = _EVAL_1488 & _EVAL_758;
  assign _EVAL_289 = _EVAL_555 == 1'h0;
  assign _EVAL_378 = _EVAL_689 & _EVAL_175;
  assign _EVAL_563 = _EVAL_1511 != 3'h0;
  assign _EVAL_1852 = _EVAL_1787 == 1'h0;
  assign _EVAL_1865 = _EVAL_2121 & _EVAL_1852;
  assign _EVAL_1712 = _EVAL_1865 & _EVAL_875;
  assign _EVAL_976 = _EVAL_1882 & _EVAL_1387;
  assign _EVAL_700 = _EVAL_2167 == 3'h0;
  assign _EVAL_683 = _EVAL_425 & _EVAL_700;
  assign _EVAL_1699 = _EVAL_979 & _EVAL_1619;
  assign _EVAL_1735 = _EVAL_1792 & _EVAL_526;
  assign _EVAL_1763 = _EVAL_829 & _EVAL_175;
  assign _EVAL_1496 = _EVAL_2039 == 4'hf;
  assign _EVAL_1330 = _EVAL_1825 & _EVAL_526;
  assign _EVAL_216 = _EVAL_267 & _EVAL_592;
  assign _EVAL_1164 = _EVAL_1178 & _EVAL_1387;
  assign _EVAL_2183 = _EVAL_1332 & _EVAL_250;
  assign _EVAL_1972 = _EVAL_431 != 3'h0;
  assign _EVAL_183 = _EVAL_379 & _EVAL_1972;
  assign _EVAL_1839 = _EVAL_1289 & _EVAL_592;
  assign _EVAL_984 = _EVAL_838 == 2'h3;
  assign _EVAL_645 = _EVAL_917 & _EVAL_526;
  assign _EVAL_952 = _EVAL_1087 == 12'hfff;
  assign _EVAL_1884 = _EVAL_414 & _EVAL_952;
  assign _EVAL_723 = _EVAL_414 & _EVAL_588;
  assign _EVAL_2003 = _EVAL_1907 & _EVAL_477;
  assign _EVAL_81 = _EVAL_974 & _EVAL_526;
  assign _EVAL_1746 = _EVAL_2213 & _EVAL_1638;
  assign _EVAL_870 = _EVAL_615 & _EVAL_592;
  assign _EVAL_2186 = _EVAL_1539 == 4'hf;
  assign _EVAL_2072 = _EVAL_328 & _EVAL_2186;
  assign _EVAL_764 = _EVAL_1519 & _EVAL_175;
  assign _EVAL_197 = _EVAL_1666 & _EVAL_1387;
  assign _EVAL_421 = _EVAL_1661 & _EVAL_711;
  assign _EVAL_524 = _EVAL_379 & _EVAL_536;
  assign _EVAL_1395 = _EVAL_982 & _EVAL_592;
  assign _EVAL_83 = _EVAL_1444 & _EVAL_526;
  assign _EVAL_903 = _EVAL_1941 & _EVAL_214;
  assign _EVAL_2141 = _EVAL_829 & _EVAL_758;
  assign _EVAL_2074 = _EVAL_967 & _EVAL_592;
  assign _EVAL_2105 = _EVAL_1289 & _EVAL_477;
  assign _EVAL_1505 = _EVAL_178 & _EVAL_592;
  assign _EVAL_2142 = _EVAL_995 & _EVAL_526;
  assign _EVAL_1002 = _EVAL_1582[17];
  assign _EVAL_1901 = _EVAL_1661 & _EVAL_1002;
  assign _EVAL_1728 = _EVAL_1272 & _EVAL_526;
  assign _EVAL_1683 = _EVAL_1426 & _EVAL_250;
  assign _EVAL_474 = _EVAL_1675 & _EVAL_477;
  assign _EVAL_346 = _EVAL_1262 & _EVAL_289;
  assign _EVAL_86 = _EVAL_379 & _EVAL_349;
  assign _EVAL_394 = _EVAL_379 & _EVAL_1015;
  assign _EVAL_834 = _EVAL_1087 != 12'h0;
  assign _EVAL_1713 = _EVAL_1689 & _EVAL_834;
  assign _EVAL_1681 = _EVAL_1983 & _EVAL_526;
  assign _EVAL_1767 = _EVAL_2037 & _EVAL_175;
  assign _EVAL_2223 = _EVAL_1809 & _EVAL_179;
  assign _EVAL_830 = _EVAL_1661 & _EVAL_1619;
  assign _EVAL_389 = _EVAL_1149 & _EVAL_250;
  assign _EVAL_258 = _EVAL_689 & _EVAL_758;
  assign _EVAL_1231 = _EVAL_1825 & _EVAL_592;
  assign _EVAL_239 = _EVAL_1431 & _EVAL_526;
  assign _EVAL_1611 = _EVAL_1332 & _EVAL_477;
  assign _EVAL_638 = _EVAL_269 & _EVAL_1638;
  assign _EVAL_888 = _EVAL_1974 & _EVAL_502;
  assign _EVAL_542 = _EVAL_888 & _EVAL_1621;
  assign _EVAL_1896 = _EVAL_2016 & _EVAL_1387;
  assign _EVAL_1891 = _EVAL_1661 & _EVAL_286;
  assign _EVAL_1692 = _EVAL_1792 & _EVAL_477;
  assign _EVAL_1506 = _EVAL_269 & _EVAL_1387;
  assign _EVAL_1848 = _EVAL_1287 & _EVAL_175;
  assign _EVAL_1738 = _EVAL_84 & _EVAL_592;
  assign _EVAL_605 = _EVAL_493 & _EVAL_179;
  assign _EVAL_534 = _EVAL_807 & _EVAL_592;
  assign _EVAL_341 = _EVAL_337 & _EVAL_477;
  assign _EVAL_413 = _EVAL_1661 & _EVAL_588;
  assign _EVAL_1375 = _EVAL_1825 & _EVAL_477;
  assign _EVAL_1614 = _EVAL_1488 & _EVAL_1387;
  assign _EVAL_2040 = _EVAL_1027 & _EVAL_1410;
  assign _EVAL_597 = _EVAL_974 & _EVAL_477;
  assign _EVAL_1351 = _EVAL_425 & _EVAL_1813;
  assign _EVAL_167 = _EVAL_1214 & _EVAL_592;
  assign _EVAL_2078 = _EVAL_1358 & _EVAL_1387;
  assign _EVAL_541 = _EVAL_1582[2];
  assign _EVAL_825 = _EVAL_979 & _EVAL_541;
  assign _EVAL_2084 = _EVAL_1837 & _EVAL_616;
  assign _EVAL_1437 = _EVAL_379 & _EVAL_2066;
  assign _EVAL_187 = _EVAL_2005 & _EVAL_477;
  assign _EVAL_2098 = _EVAL_1645 & _EVAL_250;
  assign _EVAL_1028 = _EVAL_1661 & _EVAL_2186;
  assign _EVAL_2085 = _EVAL_689 & _EVAL_1387;
  assign _EVAL_2149 = _EVAL_1170 & _EVAL_592;
  assign _EVAL_2140 = _EVAL_30 == 1'h0;
  assign _EVAL_1328 = _EVAL_1288 & _EVAL_1638;
  assign _EVAL_2028 = _EVAL_615 & _EVAL_250;
  assign _EVAL_687 = _EVAL_379 & _EVAL_1709;
  assign _EVAL_1895 = _EVAL_602 & _EVAL_592;
  assign _EVAL_1714 = _EVAL_995 & _EVAL_477;
  assign _EVAL_1477 = _EVAL_379 & _EVAL_563;
  assign _EVAL_2050 = _EVAL_549 & _EVAL_477;
  assign _EVAL_571 = _EVAL_584 & _EVAL_87;
  assign _EVAL_1498 = _EVAL_979 & _EVAL_1015;
  assign _EVAL_227 = _EVAL_1149 & _EVAL_526;
  assign _EVAL_1223 = _EVAL_913 == 7'h7f;
  assign _EVAL_484 = _EVAL_294 & _EVAL_175;
  assign _EVAL_993 = _EVAL_414 & _EVAL_1496;
  assign _EVAL_1566 = _EVAL_235 & _EVAL_1441;
  assign _EVAL_1600 = _EVAL_1510 & _EVAL_2178;
  assign _EVAL_297 = _EVAL_2124 & _EVAL_768;
  assign _EVAL_367 = _EVAL_2037 & _EVAL_758;
  assign _EVAL_1080 = _EVAL_1288 & _EVAL_1387;
  assign _EVAL_902 = _EVAL_146 & _EVAL_758;
  assign _EVAL_1775 = _EVAL_346 & _EVAL_984;
  assign _EVAL_1871 = _EVAL_2005 & _EVAL_250;
  assign _EVAL_793 = _EVAL_1165 & _EVAL_250;
  assign _EVAL_863 = _EVAL_1259 & _EVAL_87;
  assign _EVAL_158 = _EVAL_2124 & _EVAL_1517;
  assign _EVAL_1950 = _EVAL_1287 & _EVAL_758;
  assign _EVAL_252 = _EVAL_2124 & _EVAL_1624;
  assign _EVAL_1039 = _EVAL_146 & _EVAL_175;
  assign _EVAL_535 = _EVAL_1369 & _EVAL_758;
  assign _EVAL_1412 = _EVAL_337 & _EVAL_592;
  assign _EVAL_626 = _EVAL_379 & _EVAL_541;
  assign _EVAL_878 = _EVAL_585 & _EVAL_526;
  assign _EVAL_745 = _EVAL_683 & _EVAL_1806;
  assign _EVAL_1634 = _EVAL_745 & _EVAL_179;
  assign _EVAL_1934 = _EVAL_267 & _EVAL_477;
  assign _EVAL_1783 = _EVAL_1208 == 2'h3;
  assign _EVAL_2062 = _EVAL_1099 & _EVAL_477;
  assign _EVAL_1186 = _EVAL_2124 & _EVAL_1619;
  assign _EVAL_1804 = _EVAL_807 & _EVAL_477;
  assign _EVAL_2227 = _EVAL_1519 & _EVAL_758;
  assign _EVAL_1365 = _EVAL_84 & _EVAL_477;
  assign _EVAL_607 = _EVAL_1675 & _EVAL_250;
  assign _EVAL_489 = _EVAL_2124 & _EVAL_588;
  assign _EVAL_1949 = _EVAL_1661 & _EVAL_2203;
  assign _EVAL_1224 = _EVAL_2124 & _EVAL_983;
  assign _EVAL_1390 = _EVAL_602 & _EVAL_250;
  assign _EVAL_78 = _EVAL_1689 & _EVAL_563;
  assign _EVAL_1130 = _EVAL_1489 & _EVAL_1030;
  assign _EVAL_1457 = _EVAL_995 & _EVAL_592;
  assign _EVAL_292 = _EVAL_1099 & _EVAL_250;
  assign _EVAL_1922 = _EVAL_982 & _EVAL_526;
  assign _EVAL_1587 = _EVAL_1566 & _EVAL_477;
  assign _EVAL_91 = _EVAL_979 & _EVAL_1223;
  assign _EVAL_828 = _EVAL_2124 & _EVAL_939;
  assign _EVAL_206 = _EVAL_379 & _EVAL_1870;
  assign _EVAL_735 = _EVAL_1675 & _EVAL_592;
  assign _EVAL_1733 = _EVAL_1287 & _EVAL_1638;
  assign _EVAL_1438 = _EVAL_1882 & _EVAL_1638;
  assign _EVAL_691 = _EVAL_1488 & _EVAL_1638;
  assign _EVAL_2206 = _EVAL_1983 & _EVAL_250;
  assign _EVAL_891 = _EVAL_1431 & _EVAL_477;
  assign _EVAL_954 = _EVAL_974 & _EVAL_250;
  assign _EVAL_1515 = _EVAL_2124 & _EVAL_1002;
  assign _EVAL_509 = _EVAL_917 & _EVAL_477;
  assign _EVAL_2175 = _EVAL_1165 & _EVAL_592;
  assign _EVAL_1955 = _EVAL_1272 & _EVAL_592;
  assign _EVAL_1159 = _EVAL_973 & _EVAL_526;
  assign _EVAL_1674 = _EVAL_414 & _EVAL_841;
  assign _EVAL_1300 = _EVAL_549 & _EVAL_592;
  assign _EVAL_1730 = _EVAL_1566 & _EVAL_250;
  assign _EVAL_1883 = _EVAL_1369 & _EVAL_1387;
  assign _EVAL_677 = _EVAL_379 & _EVAL_588;
  assign _EVAL_1910 = _EVAL_2124 & _EVAL_640;
  assign _EVAL_1258 = _EVAL_1661 & _EVAL_832;
  assign _EVAL_520 = _EVAL_755 & _EVAL_179;
  assign _EVAL_1455 = _EVAL_1288 & _EVAL_758;
  assign _EVAL_1801 = _EVAL_1099 & _EVAL_526;
  assign _EVAL_215 = _EVAL_585 & _EVAL_592;
  assign _EVAL_1343 = _EVAL_807 & _EVAL_526;
  assign _EVAL_476 = _EVAL_2213 & _EVAL_758;
  assign _EVAL_1544 = _EVAL_1983 & _EVAL_592;
  assign _EVAL_1408 = _EVAL_982 & _EVAL_477;
  assign _EVAL_1122 = _EVAL_615 & _EVAL_526;
  assign _EVAL_720 = _EVAL_294 & _EVAL_1638;
  assign _EVAL_2128 = _EVAL_602 & _EVAL_526;
  assign _EVAL_76 = _EVAL_1444 & _EVAL_250;
  assign TLMonitor__EVAL_3 = _EVAL_867[2];
  assign TLMonitor_1__EVAL_3 = _EVAL_30;
  assign TLMonitor_1__EVAL_2 = _EVAL_12;
  assign TLMonitor_1__EVAL_9 = _EVAL_28;
  assign TLMonitor_1__EVAL_5 = {{2'd0}, _EVAL_644};
  assign TLMonitor__EVAL_14 = _EVAL_30;
  assign TLMonitor__EVAL_5 = _EVAL_41;
  assign TLMonitor__EVAL = _EVAL;
  assign TLMonitor_1__EVAL_8 = _EVAL_3;
  assign TLMonitor__EVAL_2 = _EVAL_9;
  assign TLMonitor__EVAL_7 = _EVAL_21;
  assign TLMonitor__EVAL_11 = _EVAL_32;
  assign TLMonitor__EVAL_1 = _EVAL_13;
  assign TLMonitor_1__EVAL_6 = _EVAL_14;
  assign TLMonitor_1__EVAL = _EVAL_2;
  assign TLMonitor__EVAL_13 = _EVAL_18;
  assign TLMonitor__EVAL_8 = _EVAL_13;
  assign TLMonitor_1__EVAL_14 = _EVAL_51;
  assign TLMonitor_1__EVAL_11 = _EVAL_28;
  assign TLMonitor_1__EVAL_7 = _EVAL_156[1:0];
  assign TLMonitor_1__EVAL_13 = _EVAL;
  assign TLMonitor__EVAL_12 = _EVAL_867[1:0];
  assign TLMonitor__EVAL_9 = _EVAL_1;
  assign TLMonitor__EVAL_4 = _EVAL_18;
  assign TLMonitor__EVAL_6 = _EVAL_4;
  assign TLMonitor__EVAL_0 = {{2'd0}, _EVAL_681};
  assign TLMonitor_1__EVAL_0 = _EVAL_156[13:2];
  assign TLMonitor_1__EVAL_1 = _EVAL_23;
  assign TLMonitor_1__EVAL_12 = _EVAL_48;
  assign TLMonitor_1__EVAL_4 = _EVAL_48;
  assign TLMonitor_1__EVAL_10 = _EVAL_15;
  assign TLMonitor__EVAL_10 = _EVAL_6;
  always @(posedge _EVAL) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_994 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afbcb674)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b2488ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1408 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da2b7c67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_828 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddc576f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1237 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2a8f275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(875339d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1945 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61a2047d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e52daec3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3884b68e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1371 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cffce76b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_922 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f372e1fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(332cf967)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1938 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adad719)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f41ca93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_685 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(280e83a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47c9782c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1674 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1522 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62567084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1061 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c2be98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_784 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68247ca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2145 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1445798e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2206 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4c224e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df1ee39d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1847 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32c8639f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1033 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1955 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb77c48c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1badca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59797c2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_535 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8636afda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2221 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e3e9631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec400c4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ab9e53c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1733 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51558c1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_912 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ad8fa4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2221 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b0fe02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1457 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b5c941e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_784 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(510110ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1039 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d50265a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1831 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(343f545e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1620 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6ab8b30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1217 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f312a386)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1674 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_537 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cfa6eee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1680 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(951edb50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_947 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(772cd7a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1425 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f642fdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_986 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(583dc9c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1481 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db96ecab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(784f47b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1063 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4f3b590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1568 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43b87d05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1868 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b0596e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1713 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2792a9fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(788dc511)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_872 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe872c8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2142 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c5fbc8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_851 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3363ec83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_958 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53036056)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1670 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7307a2e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_875 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e2517fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1191 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dc28de9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1977 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a90ef3fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_986 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd2d7aa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_520 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be33a8f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2063 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87fbc5a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1395 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e0be11d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_408 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(786938f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_852 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84702663)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1786 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e9287f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_875 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58dbf47c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6536724a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1848 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfd76dad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_707 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7218102b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1643 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0691f39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1242 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b026df32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_484 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f72c7c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1712 & _EVAL_1759) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1235 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bfc2e83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1885 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc568154)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_426 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3ae957b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b66e9de4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_706 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e602329)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1999 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82032f1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1382 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71b4f3f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92100dc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1365 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(770f3e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(117faf0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2100 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82fdf9f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1897 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c7e2695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1954bd2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1831 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92eae93e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3f3dc27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_863 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19929e67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1224 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1526af6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3837c554)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99b5635f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2223 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9152f138)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3dc2294)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1822 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b0062c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_567 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(607db1fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(925bdb7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1115 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de6be9b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_524 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1480 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cba32d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_611 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf269c1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_852 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81b99e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1144 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ce6c531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2227 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc2e612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1654 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51211888)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1092 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8abec17d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_567 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebaeebef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2099 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14cf3316)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_432 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74218146)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2176 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de75c848)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_378 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40afa2b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1321 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef528a86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1557 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10321da3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2134 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e866c1ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1365 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7abb9d42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1804 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84e28c0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bddb1a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_733 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1493bf6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_551 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aed9f6de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1973 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(514b50ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1598 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f11661d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f81f790a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1158 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f56d5da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1124 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9b85f6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2089 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4b8b2ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11813a2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8795072c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1660 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d489e5f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_910 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3dbb554)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2085 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9baa926)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d112686e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1423 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a99515)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba658d7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f74a5ac6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_996 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(979fd321)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_793 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22af5224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1130 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10d42220)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2145 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f6d7bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46d89f5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff53ce56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_922 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49e3bf50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(671132a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dc5751b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1949 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2b32742)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_444 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c144fdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beb7c08c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1399 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a1662a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1dc8a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2144 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb259917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1681 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88acb758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_969 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c88b1a7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1775 & _EVAL_2140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1821 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5919a47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcc70297)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5226be4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_677 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(570ac975)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1018 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e33a752)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45c7f988)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1430 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(716b0d8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1150 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5bbf7f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46cecc3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1490 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(595c882e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfb00dca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1351 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5fc7d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1684 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d951cba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_850 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(327d265a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1910 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17f1fdaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1144 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe9787a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_421 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46dc80fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1764 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ec8b304)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_394 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61e0cf2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2043 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1788 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5c4745a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1433 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29aea2b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fed2579)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1586 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e30869fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1889 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80f1704)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1133 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bca48d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_956 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15a48c28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecb344e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1959 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bced8ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1804 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f05060c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2008 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45fdbce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1585 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f01a75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_543 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7c78d1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1317 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39a51205)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a03dba82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2028 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b95588b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c494fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1732 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ef4ae27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_951 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c013ceb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1801 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(714762e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_546 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b068485)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1522 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e817ac09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1622 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb691e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1337 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(960e9d8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1568 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac9c37e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b84f44f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2152 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f2e849e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4b52ea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_993 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9964e493)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1901 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42053e6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0b07c51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_400 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cea54f07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1465 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be819131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_919 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd524ed4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_825 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0eb4103)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1552 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7507d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1918 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e48d04c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2088 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(307dcbae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(447a19ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1043 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e661a89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de73d389)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1126 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226ec3e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_686 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(738cbdee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1437 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d067509e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1614 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a810697c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1103 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(368a8f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5f81d8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_503 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1381573)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2009 & _EVAL_1759) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1133 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb98e02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80142b00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_611 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1459a6a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_378 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348e4346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_992 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(667e2d47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23c5c29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2002 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(658a0f97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1388 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffb6b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_981 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db7fa00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_998 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f18169f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1717 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(967fa95b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfb6153)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2078 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72ba1dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1428 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bef5bbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1868 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90d29647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1839 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f70be8ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1767 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d0e1d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1711 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d1eab14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1111 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daaf0409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5be9a72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1634 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(656de136)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1788 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82699dcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1158 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(989c0d28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_798 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f97f3d8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39bea28c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_524 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1712 & _EVAL_1759) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f79caa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2183 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3387a395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d38da17f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_849 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3140fbd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0af1b40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1118 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71fd8ce5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1558 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bb928de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2173 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e36f004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb7b9d51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1371 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a81b195a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51f6989f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_902 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1abe936e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2109 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d1505e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1821 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(207f1d09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2142 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efb79413)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1922 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a98b8f80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1939 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6e08341)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2168 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5614aba5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a808b0be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1063 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eddbafc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2023 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1336ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_474 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(434a8b5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_622 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc992525)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1871 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c7b6b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_788 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f902b2b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29cdfee6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1222 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c3c942)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2091 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc9f4a5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_598 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a9e6ec8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cde31753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2237 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80b13a7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1222 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8462532)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1423 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15be84d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1889 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef217589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d356c629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1910 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edd953d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_912 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e7daeb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1949 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7550a0df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1612 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f02a8b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1460 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acab52c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_535 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40c6d76d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1333 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39b3f92e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(948726d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_857 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d303f451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1883 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(350a4c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1847 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f84c73de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_669 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f683acf9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12ac2fea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1218 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdd5b783)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1435 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(524b29e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2102 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97b8701d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_946 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6aa8bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_720 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e34e456b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2105 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3faeb113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1890 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a437670d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eda915ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4b35b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4178821f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_723 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad9b78a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_863 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32ced350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1171 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a752dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2119 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77380214)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1093 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb0c045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1103 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b04170da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1290 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc83ec77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1490 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ce4223)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_791 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e696d127)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d289f4e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_582 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85cb3760)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_759 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59b3224d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1124 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31f9b2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2072 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41097242)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_805 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c70c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96dce335)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_951 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65f1dee6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1101 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1c1ea15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_878 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(103b105f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2191 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(730ea2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_960 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea74d6aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_828 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(408daebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1945 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aea59e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_762 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25896e60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_590 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c246c89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1714 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6301b0ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2074 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c141ae6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_720 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8b9db92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1258 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5483e9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1614 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38f366d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1766 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9bd7439)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f79aa840)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1513 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a09f0a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97425778)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1465 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e47d8a52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1623 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1408 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47df8ca5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1321 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d40bbcfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1126 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c82b323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ca876eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b45c6b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7022a466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1353 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cf996d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1224 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b16e02f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_992 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f75bbf9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_677 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(794ddb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a22023be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1080 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6df33d21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1544 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69e996d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbafa1f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1600 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12035996)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2063 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(411384b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1823 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a39378c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2192 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eba9bbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1570 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(389f3503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1061 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e17fe4a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_821 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce9e3dc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(690f6d14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_641 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50875fba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1752 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ec47160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_762 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c00575d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_426 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd1ee684)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2198 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7a67075)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_418 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37abb8c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2790a5e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1164 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1fa8919)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1708 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d1fcb91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6ea9b37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_734 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e316d29a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6243fa22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_998 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d3d5fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76b8b28a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_590 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54ec08c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_957 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(324d5d1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2151 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c67a548b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a81b704f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1847ebaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1673 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_891 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a65e5946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36717e80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2098 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5af354fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e9b2561)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1181 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db7919f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_981 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b613da4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82ab43f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1999 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5998baf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1343 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(315cb5fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_670 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678d211e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2068 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29b93f2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1598 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0c42408)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1457 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff6f7bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_605 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a020246)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1934 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(661aa006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2055 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7df7eef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40c25a0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_953 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc55ee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_933 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88ba5c4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d166cabd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1468 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a9d778)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ac58bf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74a53028)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1532 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b6d5bbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_833 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e34f636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_816 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9dae05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1163 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce88fbed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_712 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b748df1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_993 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(318c7fb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1111 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3b2c3dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1231 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb46f068)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_991 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fed2d463)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1047 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e5656b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1558 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42507971)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_966 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f64f3cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1797 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6564ad0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1956 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fb8b2e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1310 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a702221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_797 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f619bb43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cfd7a23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2003 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(353fc88c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1080 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92a8060c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6db545bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2068 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4a45b61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1623 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6300907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1477 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5402a6ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_718 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c891085f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d7fa5a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1355 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9662105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1231 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afd3d040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21df74f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d203bb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2034 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc443b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1128 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e6dbb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2176 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a13d1e48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(977ad6d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b34d96d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79ae1a8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1317 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(641688f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1507 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f1fc2ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11b4a89e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1024 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14e03e8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2196 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95786627)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c853e40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1692 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0ead47f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1613 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2cb4c1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2173 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a197b46f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1816 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30cc1948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2040 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87b416ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1192 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7990606)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb2f60e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0e20ba5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1171 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aef1ad50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1181 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cea13cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_730 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90ca53c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_503 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3c9e06c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1330 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc0ebe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_833 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5877002b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1035 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b99a20dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2168 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c518324b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_805 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(401f7c05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2149 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc20e2fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2034 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adcf23a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1622 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b4817cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1390 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ca24a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_728 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77b03add)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2020 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38ee472d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_902 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(902e3bf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_708 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9484efa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1876 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5db246ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e19ded)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1197 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9663e757)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_999 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cba8f9e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f1cc11d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1248 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1430 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb6f924a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd07f669)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1428 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ec81371)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1286 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5d36eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1703 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3801ce8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1300 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eb1c04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1727 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76785199)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1735 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c388cdeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af88b7a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37b02f09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1955 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d6df0d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_728 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe9549a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f28a77da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_866 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d316468)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8406fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2020 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d03569d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be9fdf00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_435 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e822c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_840 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ae693c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1039 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c1a17a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af574e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_870 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86380d14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2014 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3c18393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1823 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a815c48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1592 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c14d6ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1163 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97fc8f8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1950 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea4bf187)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1654 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54081c34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1822 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1881656e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1828 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8566df5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97f18f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2119 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59b7b5b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1711 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6888ab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_402 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b8211a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2105 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d04b51dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1699 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fda3d541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1773 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8ca2bdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1a5d60f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d739ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2237 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fc2d85b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1586 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f730dcbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_878 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a672ed01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a4b94b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1150 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe3e4f13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2141 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a33c2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf3157f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_472 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bdcc3bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1717 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb050cf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(207978d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a68209d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1258 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88bff7ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_622 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(959a3537)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2102 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0e7bce8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1592 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31b0ccba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2222 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(541a2bfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1043 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f5bfc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1838 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8d872d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1071 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4633ae29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecfb6c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728b0b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1934 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e02212)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8217d239)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ed2189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9d5053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1186 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5840dec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2014 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bfef95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1575 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e0e2f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_418 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b961d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9602f7d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64fdbdef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_598 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83177838)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a68b748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1692 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29000d88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_723 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71e138fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7923eecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_994 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cbc69b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfd3ad47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_825 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be0ec3de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b709b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1230 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da4e357f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2171 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f793f03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1884 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b859635)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1950 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49fefbd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1355 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(967efae4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1300 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2513613f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_551 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a3d8a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_670 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a57ee1cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1600 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbcf5829)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1551 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2874dd04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2120 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(188739a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1024 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e566ae9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_678 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(176eb041)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1435 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(925008f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85d6ffa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1101 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d15b5d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_476 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30575a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_797 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3acc10a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1848 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e9bab62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_537 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d125d6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1587 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4876bb0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a2ab8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1437 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(692c32ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2100 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8de4d81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ed16f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_851 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9621589e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_963 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a50b85b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d62b7e72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_946 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf787aaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2151 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7360e54a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_815 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37591bdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_626 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb84dca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1399 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(363bc216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1515 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53552487)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eae2af43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_730 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dad9f40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_444 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b1269bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_511 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e51611b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd3f1165)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2227 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57bb52f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1058 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b54a7dd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1552 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c44dc3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1684 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(686a9db0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1783 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34a227bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1816 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f628d3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1918 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17edf64d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67b787ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_449 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccc4294d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_866 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e0755c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1357 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6773f142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1679 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8340d630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_953 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(425f9592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d597bfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b530aba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8c5f474)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1460 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ee5661)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a87a8ea5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2218 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebfff9ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_509 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cb8834)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1a11e38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_669 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee494bd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2053 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51c100b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_706 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dc99acc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95a412a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_435 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bd77e76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_679 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a99423b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_830 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc1743d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2010 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(642885db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2122 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e15ba3a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_429 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfe3836e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f75808e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1316 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fbf4b17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_812 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ad1a01e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1330 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f31a743a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c3d3c10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a839647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1793119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1542 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2706957)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_785 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc51e25a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1271 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(345bb806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1871 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25010da1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1973 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8700e832)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_571 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55e44097)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2074 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d245369a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7910bba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1025 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bec86bf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1766 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4562ba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(691ee621)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49f3b08b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1382 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aff9bb60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2050 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be90603f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f3fa15c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1725334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20d6e109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9421bb2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b14a9413)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1956 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1331fbf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1891 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(757083eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1587 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42d40531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_887 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4555a1c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1389 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa7ae3fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1699 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caecff8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1122 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(453d3764)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1385 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e26161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1730 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a20905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f63a1b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1217 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a43d093a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1328 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(704ed72d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1963 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd6a55bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_678 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3789d6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_421 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db997be5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b11188bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_812 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34895ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_402 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c433428c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d72c37e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65e46f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1047 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c538885c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_466 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf568f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eca07965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1746 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e715fa89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1438 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7bbe7b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f2de234)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab44cc4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1673 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a748ea83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2192 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef2684fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2040 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1643 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74c4ae38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b521961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1733 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48986081)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_830 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b74caf1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1708 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ac9adef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1311 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb014f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6eecc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_542 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaf1bb96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1197 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24279f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48e4bbd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2055 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a5d954d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4cca179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b401da8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1541 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf7f032a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_497 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5b5b428)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1357 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec5f372)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1890 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11228f27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f02ce1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(861fd461)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2120 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43777c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1211 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac39254)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2170 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c22b656)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_686 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41479e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_448 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0eeea16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2191 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e792b6a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1145 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3c61b61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b92b0f2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2062 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18ef846c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1342 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c871f5d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ee15dd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1498 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc21cc65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e6eb404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_783 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ee383ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1895 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60b1df97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_472 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99d744c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_559 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a27260e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2268afd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1884 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7d34823)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1192 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2287ff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_759 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e6f83e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_607 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53232f19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1703 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(228f0421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1445 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d211b231)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7f49ca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc67ef8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1922 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdb6f50d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_815 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(977c57a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_509 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17eaf751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_712 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55a48e00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_931 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54f1aa2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2091 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f9ff4a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2088 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9e78afc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1186 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0a1ff4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c128c987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d9b851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_910 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(450dd5a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_671 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8992f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99080da4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1938 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4ab571c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1347 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcdb22aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1613 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e95fc01b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(954c4813)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_517 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6c00c48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1035 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d22c1c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1608 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10ff573a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1364 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88a63cfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_954 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d5a3615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec6d5fd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_449 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c5a9917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_999 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f75c810)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_521 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ac2e2a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1390 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeea6cdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1550 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a729998)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(230fcf7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb43c28c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ad576d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2043 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1003 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7389c2a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1316 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(337d1bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2128 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79755d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1406 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6796601)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33ab5f7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14b32962)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_582 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb4ee271)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1891 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2e6bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_996 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f30add8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1682 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(302f1b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1611 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5f876cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41047a75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1347 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(328a492c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8098650b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_546 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a849fbe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a0e4de8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1514 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb14e67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2007 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b60eb202)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1998 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f525e34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1018 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1305588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1342 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90a6b6e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1071 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40f13c52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1611 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(842435d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2122 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b704c7dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_733 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b1831d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1608 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bca6a309)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1145 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db2ff25f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2089 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(676c1a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1873 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f3b58f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1752 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3068cc48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf7dba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1570 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4e5140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1786 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc2b775b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1976 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7affe962)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_432 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e5e0b33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1237 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d457f5fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d410a5cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2072 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0fca167)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1846 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57b6e0a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_857 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15989ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2207 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ef677b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_870 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfff9620)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(705a85d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_521 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d66c8cbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1513 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6b7dbdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1897 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f9434a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_679 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8db6d4e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2170 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee5d28ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_919 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5da0753f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b918f42a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d49b28cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1115 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e15c6d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1506 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b17b55d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_850 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5108dab6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_497 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e01a263e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1242 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b609ae6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f0c6bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1767 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2c2065d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0939c06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_559 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42c3f376)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1164 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db2eac4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ea282dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_791 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a40cc82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6d6d2cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bd7e0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e0efcd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1481 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1059e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1620 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53258ff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_876 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59823acd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aa246b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1455 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a66e5672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aee865dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1130 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf8cd7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1455 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94991961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1326 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9729ad98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2050 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f99ff700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5c37edc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_543 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a10862b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_963 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c116064f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_931 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_419 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa5ed165)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ae2ad88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678a591f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1727 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f02ecde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17498397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b735ec4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_484 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54393079)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9387880)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2002 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c017713d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2108 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f63dba3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1585 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f646eb53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1660 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a8e84a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3ad6e01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_735 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b29615c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_903 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb92402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_954 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab4f1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2098 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ce5a61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1627 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9230b250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f36cebc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2028 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611767dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2128 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d85a0d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_929 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3020434)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1873 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6051eb1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_408 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45836507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_412 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f051420)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_956 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9264e63a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7358898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1433 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(620cd6ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e396a034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c5422b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2139 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a30b388b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_362 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(421fc1b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1959 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e20e410b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93f6c50f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1876 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47f12b6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e30ae4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e840c12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_957 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf68eaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea643774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cea587f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f03f5e31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1681 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a9ebac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc138d1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(510fd908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(113cdc9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2222 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c179fa51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2134 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6164e4e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_872 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(232cd5ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_783 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e964d292)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1153 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7b85ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2194 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64f2a2d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1627 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2c45eeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1506 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d120221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1290 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(247b0686)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1159 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9af2e69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1445 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18194855)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2078 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60ae9886)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1311 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9939acc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2131 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e45b7469)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1575 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19949640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1906fe29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_816 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8c2ec65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1343 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcf41a7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1388 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84a7e3a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1688 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(867f6846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1901 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(826c51ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1936 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fc19ea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_466 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd4da928)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1337 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6955f34f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2206 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47bd22f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1827543f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d9e5970)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1248 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2010 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58d23f53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_474 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfef3a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2175 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89f67f7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2008 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1a8e659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cfbbf28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_969 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11966ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_777 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa06e6cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1797 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a73b6e59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1670 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76bb2a32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_534 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb2bb83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d911820)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2175 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8564eb74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46a4b440)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1507 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efdaaa40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a454b2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1542 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc4f2c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1895 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3d63844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1058 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a053770)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_777 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(872e6941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1838 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeacd948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_923 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf85c95d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_511 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff8d7f46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da8372ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1117 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3af7c52a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_891 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9cc9eaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1230 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21f07a45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd1d8b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1425 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb17af42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1738 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(789cb7e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1735 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d916207)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_685 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(387c8394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1738 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e576fc44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1773 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e18a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_607 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c55f4186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_517 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(302fb5de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1159 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9232c151)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1977 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6358d3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2195 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26179e41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1764 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85d68c5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d27f4226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_708 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92110e0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1477 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d08fbf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1328 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c9668f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_923 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(700f0414)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfd8012)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1438 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3121ee99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2084 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d34c486)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1846 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7d9be6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_793 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44257f79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2099 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_933 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3057e6b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47c5c7e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8b6c568)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1310 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d828906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df65e857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_394 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7afdfce8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1093 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e85528fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2108 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27c2cef0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_785 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d521ee34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ad41a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(176718c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1680 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0370516)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2171 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5051236)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(792a3d73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_966 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5eb994f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b65831b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aabac4c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1211 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f778f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1967 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63bd97cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1998 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb93978c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1480 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63cd225)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_840 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(261c689f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_400 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(570face6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_413 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef6cd9d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2053 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7415612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2149 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ce06717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1033 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f29c306e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_887 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(709bbb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2194 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90d374f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1348 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41ddd4ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd699e37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9af4808)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8b1f398)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1732 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c06d5846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_641 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2587e0f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e203e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f5fd489)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1385 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2571e60e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b87faf7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1003 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a357fd64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2557d826)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb798f2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_960 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3a72ecb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2196 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a88f8fd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2085 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e68a20ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1450 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a46b3e9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71eab08c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1557 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29514663)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1122 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a394e323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1153 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a2e06ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc4f2bb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_487 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b44c445a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2195 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2850b9c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1544 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6e3684b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2062 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c5802d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2144 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c68d7411)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1963 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97c2bd13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_362 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77b2f06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_821 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff13888)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1333 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79e157b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1450 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9e684df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1677 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c6edeb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1532 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36f76864)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1286 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba2fa0d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d36bb4e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1326 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eee82cc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79c2bcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_958 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df650447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1936 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3cabf57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb3e73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_671 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d984a73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1550 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22784906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_735 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd0dc902)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_476 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91b3629d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1271 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30723a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2198 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51f9b1bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1801 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c610332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1746 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53aa8b0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_419 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab255887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_798 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b37d8cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1389 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0d4ab2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1118 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7eeeef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1514 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da42d939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_429 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(336b4a28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3245d0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2023 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c6b8d7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1025 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f12ab7ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_876 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c3cbaed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_487 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e98cfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1828 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b2b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_626 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7681c635)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1839 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22d7cfe1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ebfaa4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_676 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5706d0a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1883 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90227924)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a483bddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1730 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8241ebff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1117 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce19d850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd11de1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2109 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b3e640d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1348 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(454ddc31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1541 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3977bcc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_991 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f95fbc6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_788 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edfb710c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2007 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb08e55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2218 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59c0d689)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1468 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a19bb91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2048 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a32ba1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1967 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82899b81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_707 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98a21e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1688 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ada88f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1679 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2759e76f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1976 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(300302f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1885 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecdd05a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1677 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2363c1e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e0a4d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1235 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(870fc097)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_571 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c3ba4f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1b1d8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2183 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdf8e175)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2009 & _EVAL_1759) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55993371)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d14a9ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1714 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42f1dd87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1501 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea186d13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2048 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ca366c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1498 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de90d450)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(598e781f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_903 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3307e30f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8c46f02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1364 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5779da8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1395 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d92c96ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_849 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eac1c292)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(248c93fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1775 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee384ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(305c62af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1501 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb33f4b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1218 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9102a09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_676 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2834e2e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2131 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96046064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1092 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc46ced2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_947 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d0e7cda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1406 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b240d77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a957fcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1095 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7f3628a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0bfb779)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1353 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f17d6f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1095 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeb63f9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1612 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a0833bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee561b8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13125892)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1682 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28f83ed7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1939 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52de1743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2152 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf34ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17704757)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c939c6e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1713 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4533b28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ebfb03a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1551 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc0f049)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d922ad8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1515 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(694f8f16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1191 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7323174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2141 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39c012f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2003 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1bcb541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_929 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41dd9219)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b86e8b53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2139 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(760d02e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_718 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a07a137)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1128 & _EVAL_2140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7342da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
