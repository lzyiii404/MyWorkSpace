//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_0_assert(
  input  [3:0]  _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [7:0]  _EVAL_20,
  input  [3:0]  _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  input  [31:0] _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input  [3:0]  _EVAL_30,
  input  [2:0]  _EVAL_31,
  input         _EVAL_32
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_50;
  reg [31:0] _RAND_0;
  reg [3:0] _EVAL_77;
  reg [31:0] _RAND_1;
  reg [31:0] _EVAL_82;
  reg [31:0] _RAND_2;
  reg [3:0] _EVAL_105;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_113;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_161;
  reg [31:0] _RAND_5;
  reg [4:0] _EVAL_175;
  reg [31:0] _RAND_6;
  reg [3:0] _EVAL_181;
  reg [31:0] _RAND_7;
  reg [4:0] _EVAL_189;
  reg [31:0] _RAND_8;
  reg  _EVAL_224;
  reg [31:0] _RAND_9;
  reg [2:0] _EVAL_239;
  reg [31:0] _RAND_10;
  reg  _EVAL_243;
  reg [31:0] _RAND_11;
  reg [4:0] _EVAL_257;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_296;
  reg [31:0] _RAND_13;
  reg [4:0] _EVAL_348;
  reg [31:0] _RAND_14;
  reg [4:0] _EVAL_389;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_401;
  reg [31:0] _RAND_16;
  reg [3:0] _EVAL_427;
  reg [31:0] _RAND_17;
  reg [8:0] _EVAL_497;
  reg [31:0] _RAND_18;
  reg [2:0] _EVAL_501;
  reg [31:0] _RAND_19;
  reg [4:0] _EVAL_549;
  reg [31:0] _RAND_20;
  reg [2:0] _EVAL_563;
  reg [31:0] _RAND_21;
  reg [3:0] _EVAL_568;
  reg [31:0] _RAND_22;
  reg [31:0] _EVAL_574;
  reg [31:0] _RAND_23;
  reg [1:0] _EVAL_576;
  reg [31:0] _RAND_24;
  reg [31:0] _EVAL_635;
  reg [31:0] _RAND_25;
  reg [4:0] _EVAL_655;
  reg [31:0] _RAND_26;
  reg [31:0] _EVAL_670;
  reg [31:0] _RAND_27;
  wire  _EVAL_156;
  wire [31:0] _EVAL_98;
  wire [32:0] _EVAL_343;
  wire [32:0] _EVAL_381;
  wire [32:0] _EVAL_315;
  wire  _EVAL_85;
  wire [31:0] _EVAL_496;
  wire [32:0] _EVAL_588;
  wire [32:0] _EVAL_594;
  wire [32:0] _EVAL_96;
  wire  _EVAL_35;
  wire  _EVAL_318;
  wire [31:0] _EVAL_433;
  wire [32:0] _EVAL_69;
  wire [32:0] _EVAL_631;
  wire [32:0] _EVAL_210;
  wire  _EVAL_654;
  wire  _EVAL_595;
  wire [31:0] _EVAL_144;
  wire [32:0] _EVAL_180;
  wire [32:0] _EVAL_547;
  wire [32:0] _EVAL_419;
  wire  _EVAL_38;
  wire  _EVAL_406;
  wire [32:0] _EVAL_119;
  wire [32:0] _EVAL_176;
  wire [32:0] _EVAL_130;
  wire  _EVAL_380;
  wire  _EVAL_93;
  wire [31:0] _EVAL_379;
  wire [32:0] _EVAL_120;
  wire [32:0] _EVAL_170;
  wire [32:0] _EVAL_430;
  wire  _EVAL_204;
  wire  _EVAL_581;
  wire [31:0] _EVAL_618;
  wire [32:0] _EVAL_182;
  wire [32:0] _EVAL_515;
  wire [32:0] _EVAL_273;
  wire  _EVAL_443;
  wire  _EVAL_251;
  wire [31:0] _EVAL_519;
  wire [32:0] _EVAL_480;
  wire [32:0] _EVAL_41;
  wire [32:0] _EVAL_612;
  wire  _EVAL_538;
  wire  _EVAL_274;
  wire  _EVAL_267;
  wire  _EVAL_647;
  wire [31:0] _EVAL_132;
  wire [32:0] _EVAL_81;
  wire [32:0] _EVAL_290;
  wire [32:0] _EVAL_534;
  wire  _EVAL_300;
  wire  _EVAL_171;
  wire  _EVAL_339;
  wire  _EVAL_403;
  wire  _EVAL_457;
  wire  _EVAL_55;
  wire  _EVAL_48;
  wire [31:0] _EVAL_366;
  wire [32:0] _EVAL_167;
  wire [32:0] _EVAL_394;
  wire [32:0] _EVAL_439;
  wire  _EVAL_260;
  wire [31:0] _EVAL_184;
  wire [32:0] _EVAL_136;
  wire [32:0] _EVAL_90;
  wire [32:0] _EVAL_369;
  wire  _EVAL_388;
  wire  _EVAL_463;
  wire [31:0] _EVAL_342;
  wire [32:0] _EVAL_118;
  wire [32:0] _EVAL_162;
  wire [32:0] _EVAL_244;
  wire  _EVAL_102;
  wire  _EVAL_138;
  wire  _EVAL_145;
  wire  _EVAL_639;
  wire  _EVAL_355;
  wire  _EVAL_404;
  wire [1:0] _EVAL_199;
  wire [3:0] _EVAL_637;
  wire [2:0] _EVAL_368;
  wire [2:0] _EVAL_503;
  wire  _EVAL_671;
  wire  _EVAL_334;
  wire  _EVAL_426;
  wire  _EVAL_177;
  wire  _EVAL_335;
  wire  _EVAL_560;
  wire  _EVAL_438;
  wire  _EVAL_656;
  wire  _EVAL_164;
  wire  _EVAL_626;
  wire  _EVAL_61;
  wire  _EVAL_40;
  wire  _EVAL_510;
  wire  _EVAL_579;
  wire  _EVAL_146;
  wire  _EVAL_346;
  wire  _EVAL_456;
  wire  _EVAL_349;
  wire  _EVAL_326;
  wire  _EVAL_71;
  wire  _EVAL_67;
  wire  _EVAL_277;
  wire  _EVAL_319;
  wire  _EVAL_491;
  wire  _EVAL_331;
  wire  _EVAL_341;
  wire  _EVAL_424;
  wire  _EVAL_325;
  wire  _EVAL_248;
  wire  _EVAL_522;
  wire  _EVAL_537;
  wire  _EVAL_311;
  wire  _EVAL_569;
  wire  _EVAL_247;
  wire  _EVAL_464;
  wire  _EVAL_345;
  wire  _EVAL_414;
  wire  _EVAL_398;
  wire  _EVAL_540;
  wire  _EVAL_265;
  wire  _EVAL_66;
  wire  _EVAL_337;
  wire  _EVAL_43;
  wire  _EVAL_270;
  wire  _EVAL_488;
  wire  _EVAL_141;
  wire  _EVAL_532;
  wire  _EVAL_223;
  wire  _EVAL_303;
  wire [7:0] _EVAL_317;
  wire  _EVAL_110;
  wire  _EVAL_190;
  wire  _EVAL_485;
  wire  _EVAL_214;
  wire [4:0] _EVAL_151;
  wire  _EVAL_467;
  wire  _EVAL_95;
  wire  _EVAL_52;
  wire  _EVAL_364;
  wire  _EVAL_529;
  wire  _EVAL_383;
  wire  _EVAL_445;
  wire  _EVAL_661;
  wire [31:0] _EVAL_321;
  wire [32:0] _EVAL_76;
  wire [32:0] _EVAL_653;
  wire [32:0] _EVAL_564;
  wire  _EVAL_49;
  wire [31:0] _EVAL_598;
  wire [32:0] _EVAL_362;
  wire [32:0] _EVAL_518;
  wire [32:0] _EVAL_159;
  wire  _EVAL_523;
  wire  _EVAL_313;
  wire [31:0] _EVAL_64;
  wire [32:0] _EVAL_481;
  wire [32:0] _EVAL_134;
  wire [32:0] _EVAL_121;
  wire  _EVAL_259;
  wire  _EVAL_468;
  wire [31:0] _EVAL_408;
  wire [32:0] _EVAL_622;
  wire [32:0] _EVAL_561;
  wire [32:0] _EVAL_150;
  wire  _EVAL_440;
  wire  _EVAL_310;
  wire [31:0] _EVAL_663;
  wire [32:0] _EVAL_527;
  wire [32:0] _EVAL_193;
  wire [32:0] _EVAL_395;
  wire  _EVAL_123;
  wire  _EVAL_91;
  wire  _EVAL_613;
  wire  _EVAL_469;
  wire  _EVAL_295;
  wire  _EVAL_191;
  wire  _EVAL_396;
  wire [31:0] _EVAL_451;
  wire [31:0] _EVAL_425;
  wire [32:0] _EVAL_502;
  wire [32:0] _EVAL_648;
  wire [32:0] _EVAL_333;
  wire  _EVAL_353;
  wire  _EVAL_328;
  wire  _EVAL_256;
  wire  _EVAL_108;
  wire  _EVAL_201;
  wire  _EVAL_39;
  wire  _EVAL_299;
  wire [2:0] _EVAL_53;
  wire  _EVAL_533;
  wire  _EVAL_359;
  wire  _EVAL_59;
  wire [22:0] _EVAL_494;
  wire [7:0] _EVAL_550;
  wire  _EVAL_573;
  wire  _EVAL_253;
  wire  _EVAL_233;
  wire  _EVAL_72;
  wire  _EVAL_495;
  wire  _EVAL_36;
  wire  _EVAL_628;
  wire [31:0] _EVAL_640;
  wire  _EVAL_111;
  wire  _EVAL_285;
  wire [31:0] _EVAL_174;
  wire  _EVAL_34;
  wire  _EVAL_615;
  wire  _EVAL_268;
  wire  _EVAL_492;
  wire  _EVAL_506;
  wire [2:0] _EVAL_155;
  wire  _EVAL_435;
  wire  _EVAL_557;
  wire  _EVAL_302;
  wire  _EVAL_207;
  wire  _EVAL_499;
  wire  _EVAL_585;
  wire  _EVAL_106;
  wire  _EVAL_413;
  wire  _EVAL_498;
  wire  _EVAL_60;
  wire [22:0] _EVAL_112;
  wire [7:0] _EVAL_340;
  wire [7:0] _EVAL_143;
  wire [4:0] _EVAL_196;
  wire [4:0] _EVAL_434;
  wire [7:0] _EVAL_514;
  wire [31:0] _EVAL_99;
  wire [31:0] _EVAL_278;
  wire [8:0] _EVAL_291;
  wire  _EVAL_301;
  wire [7:0] _EVAL_188;
  wire [7:0] _EVAL_232;
  wire  _EVAL_530;
  wire  _EVAL_109;
  wire [31:0] _EVAL_596;
  wire [32:0] _EVAL_652;
  wire [32:0] _EVAL_65;
  wire [32:0] _EVAL_258;
  wire  _EVAL_314;
  wire  _EVAL_352;
  wire [32:0] _EVAL_641;
  wire [32:0] _EVAL_242;
  wire [32:0] _EVAL_306;
  wire  _EVAL_475;
  wire  _EVAL_393;
  wire [32:0] _EVAL_390;
  wire [32:0] _EVAL_562;
  wire [32:0] _EVAL_79;
  wire  _EVAL_577;
  wire  _EVAL_166;
  wire  _EVAL_255;
  wire  _EVAL_261;
  wire [32:0] _EVAL_587;
  wire [32:0] _EVAL_541;
  wire [32:0] _EVAL_241;
  wire  _EVAL_474;
  wire  _EVAL_344;
  wire  _EVAL_602;
  wire [22:0] _EVAL_371;
  wire [7:0] _EVAL_410;
  wire [7:0] _EVAL_511;
  wire [4:0] _EVAL_86;
  wire [4:0] _EVAL_546;
  wire  _EVAL_363;
  wire  _EVAL_600;
  wire  _EVAL_78;
  wire  _EVAL_283;
  wire  _EVAL_421;
  wire  _EVAL_73;
  wire  _EVAL_54;
  wire  _EVAL_322;
  wire  _EVAL_660;
  wire [4:0] _EVAL_472;
  wire [4:0] _EVAL_114;
  wire [31:0] _EVAL_565;
  wire [32:0] _EVAL_376;
  wire [32:0] _EVAL_249;
  wire [1:0] _EVAL_160;
  wire  _EVAL_447;
  wire  _EVAL_304;
  wire  _EVAL_583;
  wire  _EVAL_218;
  wire  _EVAL_140;
  wire  _EVAL_221;
  wire  _EVAL_633;
  wire  _EVAL_528;
  wire  _EVAL_575;
  wire  _EVAL_361;
  wire  _EVAL_642;
  wire  _EVAL_493;
  wire  _EVAL_347;
  wire [15:0] _EVAL_659;
  wire [15:0] _EVAL_208;
  wire [8:0] _EVAL_553;
  wire [8:0] _EVAL_482;
  wire [8:0] _EVAL_115;
  wire  _EVAL_211;
  wire  _EVAL_70;
  wire  _EVAL_558;
  wire  _EVAL_617;
  wire  _EVAL_280;
  wire  _EVAL_606;
  wire  _EVAL_370;
  wire  _EVAL_154;
  wire  _EVAL_179;
  wire  _EVAL_89;
  wire  _EVAL_272;
  wire  _EVAL_448;
  wire  _EVAL_486;
  wire [2:0] _EVAL_629;
  wire  _EVAL_169;
  wire  _EVAL_599;
  wire  _EVAL_198;
  wire  _EVAL_63;
  wire [15:0] _EVAL_535;
  wire [15:0] _EVAL_357;
  wire [8:0] _EVAL_542;
  wire [4:0] _EVAL_578;
  wire  _EVAL_56;
  wire  _EVAL_416;
  wire  _EVAL_172;
  wire [31:0] _EVAL_286;
  wire [32:0] _EVAL_630;
  wire [32:0] _EVAL_441;
  wire [32:0] _EVAL_178;
  wire  _EVAL_386;
  wire  _EVAL_526;
  wire  _EVAL_350;
  wire  _EVAL_658;
  wire  _EVAL_590;
  wire  _EVAL_229;
  wire  _EVAL_476;
  wire  _EVAL_544;
  wire  _EVAL_407;
  wire  _EVAL_665;
  wire  _EVAL_552;
  wire  _EVAL_524;
  wire  _EVAL_92;
  wire  _EVAL_152;
  wire  _EVAL_94;
  wire  _EVAL_504;
  wire  _EVAL_418;
  wire [31:0] _EVAL_397;
  wire [32:0] _EVAL_478;
  wire [32:0] _EVAL_539;
  wire [1:0] _EVAL_360;
  wire [1:0] _EVAL_264;
  wire [1:0] _EVAL_591;
  wire [1:0] _EVAL_284;
  wire [1:0] _EVAL_436;
  wire [1:0] _EVAL_484;
  wire [1:0] _EVAL_586;
  wire  _EVAL_227;
  wire  _EVAL_609;
  wire  _EVAL_142;
  wire [4:0] _EVAL_126;
  wire  _EVAL_293;
  wire  _EVAL_543;
  wire [7:0] _EVAL_87;
  wire  _EVAL_104;
  wire  _EVAL_668;
  wire  _EVAL_230;
  wire  _EVAL_252;
  wire  _EVAL_327;
  wire  _EVAL_638;
  wire  _EVAL_516;
  wire  _EVAL_601;
  wire [31:0] _EVAL_298;
  wire  _EVAL_597;
  wire  _EVAL_316;
  wire  _EVAL_33;
  wire  _EVAL_399;
  wire  _EVAL_669;
  wire  _EVAL_466;
  wire  _EVAL_559;
  wire  _EVAL_666;
  wire  _EVAL_57;
  wire  _EVAL_548;
  wire  _EVAL_269;
  wire  _EVAL_236;
  wire  _EVAL_446;
  wire  _EVAL_228;
  wire [31:0] _EVAL_101;
  wire  _EVAL_254;
  wire  _EVAL_507;
  wire [32:0] _EVAL_567;
  wire [32:0] _EVAL_610;
  wire [32:0] _EVAL_217;
  wire  _EVAL_329;
  wire  _EVAL_75;
  wire  _EVAL_288;
  wire  _EVAL_509;
  wire [31:0] _EVAL_42;
  wire [32:0] _EVAL_135;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_411;
  wire  _EVAL_125;
  wire  _EVAL_649;
  wire [31:0] _EVAL_100;
  wire [32:0] _EVAL_45;
  wire [32:0] _EVAL_400;
  wire [32:0] _EVAL_644;
  wire  _EVAL_551;
  wire  _EVAL_202;
  wire [31:0] _EVAL_187;
  wire [32:0] _EVAL_461;
  wire [32:0] _EVAL_168;
  wire [32:0] _EVAL_209;
  wire  _EVAL_566;
  wire  _EVAL_545;
  wire  _EVAL_431;
  wire  _EVAL_97;
  wire  _EVAL_250;
  wire  _EVAL_634;
  wire  _EVAL_616;
  wire  _EVAL_367;
  wire  _EVAL_505;
  wire [4:0] _EVAL_46;
  wire  _EVAL_453;
  wire  _EVAL_623;
  wire  _EVAL_365;
  wire  _EVAL_372;
  wire  _EVAL_619;
  wire  _EVAL_213;
  wire  _EVAL_620;
  wire  _EVAL_465;
  wire  _EVAL_603;
  wire  _EVAL_657;
  wire  _EVAL_74;
  wire  _EVAL_173;
  wire  _EVAL_471;
  wire  _EVAL_377;
  wire  _EVAL_525;
  wire  _EVAL_225;
  wire  _EVAL_235;
  wire  _EVAL_332;
  wire  _EVAL_382;
  wire  _EVAL_262;
  wire  _EVAL_216;
  wire  _EVAL_489;
  wire  _EVAL_593;
  wire [31:0] _EVAL_555;
  wire  _EVAL_197;
  wire  _EVAL_632;
  wire  _EVAL_462;
  wire [32:0] _EVAL_51;
  wire  _EVAL_592;
  wire [32:0] _EVAL_643;
  wire  _EVAL_323;
  wire  _EVAL_195;
  wire  _EVAL_282;
  wire  _EVAL_205;
  wire  _EVAL_139;
  wire  _EVAL_417;
  wire  _EVAL_336;
  wire  _EVAL_607;
  wire  _EVAL_483;
  wire  _EVAL_536;
  wire  _EVAL_351;
  wire  _EVAL_200;
  wire  _EVAL_384;
  wire  _EVAL_124;
  wire  _EVAL_608;
  wire  _EVAL_220;
  wire  _EVAL_238;
  wire  _EVAL_129;
  wire  _EVAL_68;
  wire  _EVAL_305;
  wire  _EVAL_281;
  wire  _EVAL_373;
  wire  _EVAL_183;
  wire  _EVAL_117;
  wire  _EVAL_240;
  wire  _EVAL_276;
  wire  _EVAL_287;
  wire  _EVAL_387;
  wire  _EVAL_222;
  wire  _EVAL_47;
  wire  _EVAL_58;
  wire  _EVAL_531;
  wire  _EVAL_490;
  wire  _EVAL_589;
  wire  _EVAL_62;
  wire [1:0] _EVAL_604;
  wire [1:0] _EVAL_428;
  wire  _EVAL_194;
  wire  _EVAL_186;
  wire  _EVAL_458;
  wire  _EVAL_107;
  wire  _EVAL_128;
  wire  _EVAL_450;
  wire  _EVAL_614;
  wire  _EVAL_500;
  wire  _EVAL_460;
  wire  _EVAL_354;
  wire  _EVAL_479;
  wire  _EVAL_487;
  wire  _EVAL_237;
  wire  _EVAL_226;
  wire  _EVAL_234;
  wire  _EVAL_378;
  wire  _EVAL_517;
  wire  _EVAL_149;
  wire  _EVAL_294;
  wire  _EVAL_356;
  wire  _EVAL_203;
  wire  _EVAL_625;
  wire  _EVAL_402;
  wire  _EVAL_88;
  wire  _EVAL_147;
  wire  _EVAL_572;
  wire  _EVAL_415;
  wire  _EVAL_158;
  wire  _EVAL_621;
  wire  _EVAL_582;
  wire  _EVAL_405;
  wire  _EVAL_605;
  wire  _EVAL_37;
  wire  _EVAL_650;
  wire  _EVAL_212;
  wire  _EVAL_624;
  wire  _EVAL_165;
  wire  _EVAL_580;
  wire  _EVAL_122;
  wire  _EVAL_385;
  wire [8:0] _EVAL_477;
  wire  _EVAL_330;
  wire  _EVAL_309;
  wire  _EVAL_611;
  wire  _EVAL_83;
  wire  _EVAL_185;
  wire  _EVAL_279;
  wire  _EVAL_432;
  wire  _EVAL_271;
  wire  _EVAL_627;
  wire  _EVAL_206;
  wire  _EVAL_263;
  wire  _EVAL_103;
  wire  _EVAL_571;
  wire  _EVAL_292;
  wire  _EVAL_153;
  wire  _EVAL_308;
  wire  _EVAL_423;
  wire  _EVAL_452;
  wire  _EVAL_192;
  wire  _EVAL_470;
  wire  _EVAL_338;
  wire  _EVAL_312;
  wire  _EVAL_473;
  wire  _EVAL_131;
  wire  _EVAL_664;
  wire  _EVAL_44;
  wire  _EVAL_646;
  wire  _EVAL_422;
  wire  _EVAL_429;
  wire  _EVAL_289;
  wire  _EVAL_520;
  wire [8:0] _EVAL_412;
  wire [8:0] _EVAL_246;
  wire  _EVAL_420;
  wire  _EVAL_444;
  wire  _EVAL_437;
  wire  _EVAL_391;
  wire  _EVAL_297;
  wire  _EVAL_442;
  wire  _EVAL_84;
  wire  _EVAL_636;
  wire  _EVAL_127;
  wire  _EVAL_667;
  wire  _EVAL_374;
  wire  _EVAL_570;
  wire  _EVAL_245;
  wire  _EVAL_584;
  wire  _EVAL_662;
  wire  _EVAL_409;
  wire  _EVAL_455;
  wire  _EVAL_215;
  wire  _EVAL_116;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_156 = _EVAL_30 <= 4'h6;
  assign _EVAL_98 = _EVAL_0 ^ 32'h40000000;
  assign _EVAL_343 = {1'b0,$signed(_EVAL_98)};
  assign _EVAL_381 = $signed(_EVAL_343) & $signed(-33'sh2000);
  assign _EVAL_315 = $signed(_EVAL_381);
  assign _EVAL_85 = $signed(_EVAL_315) == $signed(33'sh0);
  assign _EVAL_496 = _EVAL_0 ^ 32'h80000000;
  assign _EVAL_588 = {1'b0,$signed(_EVAL_496)};
  assign _EVAL_594 = $signed(_EVAL_588) & $signed(-33'sh20000);
  assign _EVAL_96 = $signed(_EVAL_594);
  assign _EVAL_35 = $signed(_EVAL_96) == $signed(33'sh0);
  assign _EVAL_318 = _EVAL_85 | _EVAL_35;
  assign _EVAL_433 = _EVAL_0 ^ 32'hc000000;
  assign _EVAL_69 = {1'b0,$signed(_EVAL_433)};
  assign _EVAL_631 = $signed(_EVAL_69) & $signed(-33'sh4000000);
  assign _EVAL_210 = $signed(_EVAL_631);
  assign _EVAL_654 = $signed(_EVAL_210) == $signed(33'sh0);
  assign _EVAL_595 = _EVAL_318 | _EVAL_654;
  assign _EVAL_144 = _EVAL_0 ^ 32'h2000000;
  assign _EVAL_180 = {1'b0,$signed(_EVAL_144)};
  assign _EVAL_547 = $signed(_EVAL_180) & $signed(-33'sh10000);
  assign _EVAL_419 = $signed(_EVAL_547);
  assign _EVAL_38 = $signed(_EVAL_419) == $signed(33'sh0);
  assign _EVAL_406 = _EVAL_595 | _EVAL_38;
  assign _EVAL_119 = {1'b0,$signed(_EVAL_0)};
  assign _EVAL_176 = $signed(_EVAL_119) & $signed(-33'sh5000);
  assign _EVAL_130 = $signed(_EVAL_176);
  assign _EVAL_380 = $signed(_EVAL_130) == $signed(33'sh0);
  assign _EVAL_93 = _EVAL_406 | _EVAL_380;
  assign _EVAL_379 = _EVAL_0 ^ 32'h1800000;
  assign _EVAL_120 = {1'b0,$signed(_EVAL_379)};
  assign _EVAL_170 = $signed(_EVAL_120) & $signed(-33'sh8000);
  assign _EVAL_430 = $signed(_EVAL_170);
  assign _EVAL_204 = $signed(_EVAL_430) == $signed(33'sh0);
  assign _EVAL_581 = _EVAL_93 | _EVAL_204;
  assign _EVAL_618 = _EVAL_0 ^ 32'h1900000;
  assign _EVAL_182 = {1'b0,$signed(_EVAL_618)};
  assign _EVAL_515 = $signed(_EVAL_182) & $signed(-33'sh2000);
  assign _EVAL_273 = $signed(_EVAL_515);
  assign _EVAL_443 = $signed(_EVAL_273) == $signed(33'sh0);
  assign _EVAL_251 = _EVAL_581 | _EVAL_443;
  assign _EVAL_519 = _EVAL_0 ^ 32'h20000000;
  assign _EVAL_480 = {1'b0,$signed(_EVAL_519)};
  assign _EVAL_41 = $signed(_EVAL_480) & $signed(-33'sh2000);
  assign _EVAL_612 = $signed(_EVAL_41);
  assign _EVAL_538 = $signed(_EVAL_612) == $signed(33'sh0);
  assign _EVAL_274 = _EVAL_251 | _EVAL_538;
  assign _EVAL_267 = _EVAL_156 & _EVAL_274;
  assign _EVAL_647 = _EVAL_30 <= 4'h8;
  assign _EVAL_132 = _EVAL_0 ^ 32'h3000;
  assign _EVAL_81 = {1'b0,$signed(_EVAL_132)};
  assign _EVAL_290 = $signed(_EVAL_81) & $signed(-33'sh1000);
  assign _EVAL_534 = $signed(_EVAL_290);
  assign _EVAL_300 = $signed(_EVAL_534) == $signed(33'sh0);
  assign _EVAL_171 = _EVAL_647 & _EVAL_300;
  assign _EVAL_339 = _EVAL_267 | _EVAL_171;
  assign _EVAL_403 = _EVAL_339 | _EVAL_28;
  assign _EVAL_457 = _EVAL_403 == 1'h0;
  assign _EVAL_55 = _EVAL_22 == 3'h5;
  assign _EVAL_48 = _EVAL_9 & _EVAL_55;
  assign _EVAL_366 = _EVAL_24 ^ 32'h40000000;
  assign _EVAL_167 = {1'b0,$signed(_EVAL_366)};
  assign _EVAL_394 = $signed(_EVAL_167) & $signed(-33'sh2000);
  assign _EVAL_439 = $signed(_EVAL_394);
  assign _EVAL_260 = $signed(_EVAL_439) == $signed(33'sh0);
  assign _EVAL_184 = _EVAL_24 ^ 32'h80000000;
  assign _EVAL_136 = {1'b0,$signed(_EVAL_184)};
  assign _EVAL_90 = $signed(_EVAL_136) & $signed(-33'sh20000);
  assign _EVAL_369 = $signed(_EVAL_90);
  assign _EVAL_388 = $signed(_EVAL_369) == $signed(33'sh0);
  assign _EVAL_463 = _EVAL_260 | _EVAL_388;
  assign _EVAL_342 = _EVAL_24 ^ 32'h3000;
  assign _EVAL_118 = {1'b0,$signed(_EVAL_342)};
  assign _EVAL_162 = $signed(_EVAL_118) & $signed(-33'sh1000);
  assign _EVAL_244 = $signed(_EVAL_162);
  assign _EVAL_102 = $signed(_EVAL_244) == $signed(33'sh0);
  assign _EVAL_138 = _EVAL_463 | _EVAL_102;
  assign _EVAL_145 = _EVAL_12 <= 2'h2;
  assign _EVAL_639 = _EVAL_145 | _EVAL_28;
  assign _EVAL_355 = _EVAL_639 == 1'h0;
  assign _EVAL_404 = _EVAL_30 >= 4'h3;
  assign _EVAL_199 = _EVAL_30[1:0];
  assign _EVAL_637 = 4'h1 << _EVAL_199;
  assign _EVAL_368 = _EVAL_637[2:0];
  assign _EVAL_503 = _EVAL_368 | 3'h1;
  assign _EVAL_671 = _EVAL_503[2];
  assign _EVAL_334 = _EVAL_0[2];
  assign _EVAL_426 = _EVAL_671 & _EVAL_334;
  assign _EVAL_177 = _EVAL_404 | _EVAL_426;
  assign _EVAL_335 = _EVAL_503[1];
  assign _EVAL_560 = _EVAL_0[1];
  assign _EVAL_438 = _EVAL_334 & _EVAL_560;
  assign _EVAL_656 = _EVAL_335 & _EVAL_438;
  assign _EVAL_164 = _EVAL_177 | _EVAL_656;
  assign _EVAL_626 = _EVAL_503[0];
  assign _EVAL_61 = _EVAL_0[0];
  assign _EVAL_40 = _EVAL_438 & _EVAL_61;
  assign _EVAL_510 = _EVAL_626 & _EVAL_40;
  assign _EVAL_579 = _EVAL_164 | _EVAL_510;
  assign _EVAL_146 = _EVAL_61 == 1'h0;
  assign _EVAL_346 = _EVAL_438 & _EVAL_146;
  assign _EVAL_456 = _EVAL_626 & _EVAL_346;
  assign _EVAL_349 = _EVAL_164 | _EVAL_456;
  assign _EVAL_326 = _EVAL_560 == 1'h0;
  assign _EVAL_71 = _EVAL_334 & _EVAL_326;
  assign _EVAL_67 = _EVAL_335 & _EVAL_71;
  assign _EVAL_277 = _EVAL_177 | _EVAL_67;
  assign _EVAL_319 = _EVAL_71 & _EVAL_61;
  assign _EVAL_491 = _EVAL_626 & _EVAL_319;
  assign _EVAL_331 = _EVAL_277 | _EVAL_491;
  assign _EVAL_341 = _EVAL_71 & _EVAL_146;
  assign _EVAL_424 = _EVAL_626 & _EVAL_341;
  assign _EVAL_325 = _EVAL_277 | _EVAL_424;
  assign _EVAL_248 = _EVAL_334 == 1'h0;
  assign _EVAL_522 = _EVAL_671 & _EVAL_248;
  assign _EVAL_537 = _EVAL_404 | _EVAL_522;
  assign _EVAL_311 = _EVAL_248 & _EVAL_560;
  assign _EVAL_569 = _EVAL_335 & _EVAL_311;
  assign _EVAL_247 = _EVAL_537 | _EVAL_569;
  assign _EVAL_464 = _EVAL_311 & _EVAL_61;
  assign _EVAL_345 = _EVAL_626 & _EVAL_464;
  assign _EVAL_414 = _EVAL_247 | _EVAL_345;
  assign _EVAL_398 = _EVAL_311 & _EVAL_146;
  assign _EVAL_540 = _EVAL_626 & _EVAL_398;
  assign _EVAL_265 = _EVAL_247 | _EVAL_540;
  assign _EVAL_66 = _EVAL_248 & _EVAL_326;
  assign _EVAL_337 = _EVAL_335 & _EVAL_66;
  assign _EVAL_43 = _EVAL_537 | _EVAL_337;
  assign _EVAL_270 = _EVAL_66 & _EVAL_61;
  assign _EVAL_488 = _EVAL_626 & _EVAL_270;
  assign _EVAL_141 = _EVAL_43 | _EVAL_488;
  assign _EVAL_532 = _EVAL_66 & _EVAL_146;
  assign _EVAL_223 = _EVAL_626 & _EVAL_532;
  assign _EVAL_303 = _EVAL_43 | _EVAL_223;
  assign _EVAL_317 = {_EVAL_579,_EVAL_349,_EVAL_331,_EVAL_325,_EVAL_414,_EVAL_265,_EVAL_141,_EVAL_303};
  assign _EVAL_110 = _EVAL_20 == _EVAL_317;
  assign _EVAL_190 = _EVAL_110 | _EVAL_28;
  assign _EVAL_485 = _EVAL_6 & _EVAL_13;
  assign _EVAL_214 = _EVAL_189 == 5'h0;
  assign _EVAL_151 = _EVAL_189 - 5'h1;
  assign _EVAL_467 = _EVAL_5 == 1'h0;
  assign _EVAL_95 = _EVAL_467 | _EVAL_28;
  assign _EVAL_52 = _EVAL_11 == 3'h2;
  assign _EVAL_364 = _EVAL_23 & _EVAL_9;
  assign _EVAL_529 = _EVAL_257 == 5'h0;
  assign _EVAL_383 = _EVAL_364 & _EVAL_529;
  assign _EVAL_445 = _EVAL_11 == 3'h5;
  assign _EVAL_661 = _EVAL_16 & _EVAL_445;
  assign _EVAL_321 = _EVAL_8 ^ 32'h40000000;
  assign _EVAL_76 = {1'b0,$signed(_EVAL_321)};
  assign _EVAL_653 = $signed(_EVAL_76) & $signed(-33'sh2000);
  assign _EVAL_564 = $signed(_EVAL_653);
  assign _EVAL_49 = $signed(_EVAL_564) == $signed(33'sh0);
  assign _EVAL_598 = _EVAL_8 ^ 32'h80000000;
  assign _EVAL_362 = {1'b0,$signed(_EVAL_598)};
  assign _EVAL_518 = $signed(_EVAL_362) & $signed(-33'sh20000);
  assign _EVAL_159 = $signed(_EVAL_518);
  assign _EVAL_523 = $signed(_EVAL_159) == $signed(33'sh0);
  assign _EVAL_313 = _EVAL_49 | _EVAL_523;
  assign _EVAL_64 = _EVAL_8 ^ 32'h3000;
  assign _EVAL_481 = {1'b0,$signed(_EVAL_64)};
  assign _EVAL_134 = $signed(_EVAL_481) & $signed(-33'sh1000);
  assign _EVAL_121 = $signed(_EVAL_134);
  assign _EVAL_259 = $signed(_EVAL_121) == $signed(33'sh0);
  assign _EVAL_468 = _EVAL_313 | _EVAL_259;
  assign _EVAL_408 = _EVAL_8 ^ 32'hc000000;
  assign _EVAL_622 = {1'b0,$signed(_EVAL_408)};
  assign _EVAL_561 = $signed(_EVAL_622) & $signed(-33'sh4000000);
  assign _EVAL_150 = $signed(_EVAL_561);
  assign _EVAL_440 = $signed(_EVAL_150) == $signed(33'sh0);
  assign _EVAL_310 = _EVAL_468 | _EVAL_440;
  assign _EVAL_663 = _EVAL_8 ^ 32'h2000000;
  assign _EVAL_527 = {1'b0,$signed(_EVAL_663)};
  assign _EVAL_193 = $signed(_EVAL_527) & $signed(-33'sh10000);
  assign _EVAL_395 = $signed(_EVAL_193);
  assign _EVAL_123 = $signed(_EVAL_395) == $signed(33'sh0);
  assign _EVAL_91 = _EVAL_310 | _EVAL_123;
  assign _EVAL_613 = _EVAL_10 == 4'h8;
  assign _EVAL_469 = _EVAL_10 == 4'h0;
  assign _EVAL_295 = _EVAL_613 | _EVAL_469;
  assign _EVAL_191 = _EVAL_11 == 3'h6;
  assign _EVAL_396 = _EVAL_16 & _EVAL_191;
  assign _EVAL_451 = _EVAL_24 ^ 32'hc000000;
  assign _EVAL_425 = _EVAL_24 ^ 32'h1800000;
  assign _EVAL_502 = {1'b0,$signed(_EVAL_425)};
  assign _EVAL_648 = $signed(_EVAL_502) & $signed(-33'sh8000);
  assign _EVAL_333 = $signed(_EVAL_648);
  assign _EVAL_353 = _EVAL_300 | _EVAL_654;
  assign _EVAL_328 = _EVAL_353 | _EVAL_38;
  assign _EVAL_256 = _EVAL_4 == 4'h8;
  assign _EVAL_108 = _EVAL_4 == 4'h0;
  assign _EVAL_201 = _EVAL_256 | _EVAL_108;
  assign _EVAL_39 = _EVAL_4[3:3];
  assign _EVAL_299 = _EVAL_39 == 1'h0;
  assign _EVAL_53 = _EVAL_4[2:0];
  assign _EVAL_533 = 3'h1 <= _EVAL_53;
  assign _EVAL_359 = _EVAL_299 & _EVAL_533;
  assign _EVAL_59 = _EVAL_201 | _EVAL_359;
  assign _EVAL_494 = 23'hff << _EVAL_21;
  assign _EVAL_550 = _EVAL_494[7:0];
  assign _EVAL_573 = _EVAL_22[2];
  assign _EVAL_253 = _EVAL_22[1];
  assign _EVAL_233 = _EVAL_253 == 1'h0;
  assign _EVAL_72 = _EVAL_573 & _EVAL_233;
  assign _EVAL_495 = _EVAL_17 != 3'h0;
  assign _EVAL_36 = _EVAL_17 <= 3'h2;
  assign _EVAL_628 = _EVAL_36 | _EVAL_28;
  assign _EVAL_640 = _EVAL_670 + 32'h1;
  assign _EVAL_111 = _EVAL_655 == 5'h0;
  assign _EVAL_285 = _EVAL_111 == 1'h0;
  assign _EVAL_174 = _EVAL_24 ^ 32'h2000000;
  assign _EVAL_34 = _EVAL_8 == _EVAL_82;
  assign _EVAL_615 = _EVAL_34 | _EVAL_28;
  assign _EVAL_268 = _EVAL_615 == 1'h0;
  assign _EVAL_492 = _EVAL_10[3:3];
  assign _EVAL_506 = _EVAL_492 == 1'h0;
  assign _EVAL_155 = _EVAL_10[2:0];
  assign _EVAL_435 = 3'h1 <= _EVAL_155;
  assign _EVAL_557 = _EVAL_506 & _EVAL_435;
  assign _EVAL_302 = _EVAL_295 | _EVAL_557;
  assign _EVAL_207 = _EVAL_302 | _EVAL_28;
  assign _EVAL_499 = _EVAL_175 == 5'h0;
  assign _EVAL_585 = _EVAL_499 == 1'h0;
  assign _EVAL_106 = _EVAL_2 & _EVAL_585;
  assign _EVAL_413 = _EVAL_549 == 5'h0;
  assign _EVAL_498 = _EVAL_11[2];
  assign _EVAL_60 = _EVAL_498 == 1'h0;
  assign _EVAL_112 = 23'hff << _EVAL_30;
  assign _EVAL_340 = _EVAL_112[7:0];
  assign _EVAL_143 = ~ _EVAL_340;
  assign _EVAL_196 = _EVAL_143[7:3];
  assign _EVAL_434 = _EVAL_549 - 5'h1;
  assign _EVAL_514 = ~ _EVAL_550;
  assign _EVAL_99 = {{24'd0}, _EVAL_514};
  assign _EVAL_278 = _EVAL_8 & _EVAL_99;
  assign _EVAL_291 = _EVAL_497 >> _EVAL_4;
  assign _EVAL_301 = _EVAL_291[0];
  assign _EVAL_188 = ~ _EVAL_317;
  assign _EVAL_232 = _EVAL_20 & _EVAL_188;
  assign _EVAL_530 = _EVAL_232 == 8'h0;
  assign _EVAL_109 = _EVAL_530 | _EVAL_28;
  assign _EVAL_596 = _EVAL_24 ^ 32'h1900000;
  assign _EVAL_652 = {1'b0,$signed(_EVAL_451)};
  assign _EVAL_65 = $signed(_EVAL_652) & $signed(-33'sh4000000);
  assign _EVAL_258 = $signed(_EVAL_65);
  assign _EVAL_314 = $signed(_EVAL_258) == $signed(33'sh0);
  assign _EVAL_352 = _EVAL_138 | _EVAL_314;
  assign _EVAL_641 = {1'b0,$signed(_EVAL_174)};
  assign _EVAL_242 = $signed(_EVAL_641) & $signed(-33'sh10000);
  assign _EVAL_306 = $signed(_EVAL_242);
  assign _EVAL_475 = $signed(_EVAL_306) == $signed(33'sh0);
  assign _EVAL_393 = _EVAL_352 | _EVAL_475;
  assign _EVAL_390 = {1'b0,$signed(_EVAL_24)};
  assign _EVAL_562 = $signed(_EVAL_390) & $signed(-33'sh1000);
  assign _EVAL_79 = $signed(_EVAL_562);
  assign _EVAL_577 = $signed(_EVAL_79) == $signed(33'sh0);
  assign _EVAL_166 = _EVAL_393 | _EVAL_577;
  assign _EVAL_255 = $signed(_EVAL_333) == $signed(33'sh0);
  assign _EVAL_261 = _EVAL_166 | _EVAL_255;
  assign _EVAL_587 = {1'b0,$signed(_EVAL_596)};
  assign _EVAL_541 = $signed(_EVAL_587) & $signed(-33'sh2000);
  assign _EVAL_241 = $signed(_EVAL_541);
  assign _EVAL_474 = $signed(_EVAL_241) == $signed(33'sh0);
  assign _EVAL_344 = _EVAL_261 | _EVAL_474;
  assign _EVAL_602 = _EVAL_22[0];
  assign _EVAL_371 = 23'hff << _EVAL;
  assign _EVAL_410 = _EVAL_371[7:0];
  assign _EVAL_511 = ~ _EVAL_410;
  assign _EVAL_86 = _EVAL_511[7:3];
  assign _EVAL_546 = _EVAL_257 - 5'h1;
  assign _EVAL_363 = _EVAL_17 == _EVAL_239;
  assign _EVAL_600 = _EVAL_363 | _EVAL_28;
  assign _EVAL_78 = _EVAL_600 == 1'h0;
  assign _EVAL_283 = _EVAL_15 == 4'h0;
  assign _EVAL_421 = _EVAL_17 <= 3'h3;
  assign _EVAL_73 = _EVAL_421 | _EVAL_28;
  assign _EVAL_54 = _EVAL_73 == 1'h0;
  assign _EVAL_322 = _EVAL_32 & _EVAL_2;
  assign _EVAL_660 = _EVAL_7[0];
  assign _EVAL_472 = _EVAL_514[7:3];
  assign _EVAL_114 = _EVAL_175 - 5'h1;
  assign _EVAL_565 = _EVAL_24 ^ 32'h20000000;
  assign _EVAL_376 = {1'b0,$signed(_EVAL_565)};
  assign _EVAL_249 = $signed(_EVAL_376) & $signed(-33'sh2000);
  assign _EVAL_160 = _EVAL_296 >> _EVAL_3;
  assign _EVAL_447 = _EVAL_160[0];
  assign _EVAL_304 = _EVAL_447 == 1'h0;
  assign _EVAL_583 = _EVAL_348 == 5'h0;
  assign _EVAL_218 = _EVAL_583 == 1'h0;
  assign _EVAL_140 = _EVAL_16 & _EVAL_218;
  assign _EVAL_221 = _EVAL_389 == 5'h0;
  assign _EVAL_633 = _EVAL_364 & _EVAL_221;
  assign _EVAL_528 = _EVAL_633 & _EVAL_72;
  assign _EVAL_575 = _EVAL_278 == 32'h0;
  assign _EVAL_361 = _EVAL_575 | _EVAL_28;
  assign _EVAL_642 = _EVAL_361 == 1'h0;
  assign _EVAL_493 = _EVAL_25 & _EVAL_16;
  assign _EVAL_347 = _EVAL_493 & _EVAL_413;
  assign _EVAL_659 = 16'h1 << _EVAL_4;
  assign _EVAL_208 = _EVAL_347 ? _EVAL_659 : 16'h0;
  assign _EVAL_553 = _EVAL_208[8:0];
  assign _EVAL_482 = _EVAL_553 | _EVAL_497;
  assign _EVAL_115 = _EVAL_482 >> _EVAL_10;
  assign _EVAL_211 = _EVAL_115[0];
  assign _EVAL_70 = _EVAL_211 | _EVAL_28;
  assign _EVAL_558 = _EVAL_22 <= 3'h6;
  assign _EVAL_617 = _EVAL_558 | _EVAL_28;
  assign _EVAL_280 = _EVAL_156 & _EVAL_35;
  assign _EVAL_606 = _EVAL_280 | _EVAL_28;
  assign _EVAL_370 = _EVAL_606 == 1'h0;
  assign _EVAL_154 = _EVAL_31 == _EVAL_563;
  assign _EVAL_179 = _EVAL_154 | _EVAL_28;
  assign _EVAL_89 = _EVAL_5 == _EVAL_243;
  assign _EVAL_272 = _EVAL_89 | _EVAL_28;
  assign _EVAL_448 = _EVAL_485 & _EVAL_214;
  assign _EVAL_486 = _EVAL >= 4'h3;
  assign _EVAL_629 = _EVAL_15[2:0];
  assign _EVAL_169 = 3'h1 <= _EVAL_629;
  assign _EVAL_599 = _EVAL_22 == 3'h6;
  assign _EVAL_198 = _EVAL_599 == 1'h0;
  assign _EVAL_63 = _EVAL_383 & _EVAL_198;
  assign _EVAL_535 = 16'h1 << _EVAL_10;
  assign _EVAL_357 = _EVAL_63 ? _EVAL_535 : 16'h0;
  assign _EVAL_542 = _EVAL_357[8:0];
  assign _EVAL_578 = _EVAL_655 - 5'h1;
  assign _EVAL_56 = _EVAL_31 == 3'h0;
  assign _EVAL_416 = _EVAL_56 | _EVAL_28;
  assign _EVAL_172 = _EVAL_416 == 1'h0;
  assign _EVAL_286 = _EVAL_8 ^ 32'h1800000;
  assign _EVAL_630 = {1'b0,$signed(_EVAL_286)};
  assign _EVAL_441 = $signed(_EVAL_630) & $signed(-33'sh8000);
  assign _EVAL_178 = $signed(_EVAL_441);
  assign _EVAL_386 = _EVAL_322 & _EVAL_499;
  assign _EVAL_526 = _EVAL_22 == _EVAL_501;
  assign _EVAL_350 = _EVAL_526 | _EVAL_28;
  assign _EVAL_658 = _EVAL_14 == _EVAL_113;
  assign _EVAL_590 = _EVAL_658 | _EVAL_28;
  assign _EVAL_229 = _EVAL_590 == 1'h0;
  assign _EVAL_476 = _EVAL_11 == 3'h4;
  assign _EVAL_544 = _EVAL_16 & _EVAL_476;
  assign _EVAL_407 = _EVAL_22 == 3'h2;
  assign _EVAL_665 = _EVAL_30 <= 4'h2;
  assign _EVAL_552 = _EVAL_328 | _EVAL_380;
  assign _EVAL_524 = _EVAL_552 | _EVAL_204;
  assign _EVAL_92 = _EVAL_524 | _EVAL_443;
  assign _EVAL_152 = _EVAL_92 | _EVAL_538;
  assign _EVAL_94 = _EVAL_665 & _EVAL_152;
  assign _EVAL_504 = _EVAL_94 | _EVAL_28;
  assign _EVAL_418 = _EVAL_504 == 1'h0;
  assign _EVAL_397 = _EVAL_24 ^ 32'h4000;
  assign _EVAL_478 = {1'b0,$signed(_EVAL_397)};
  assign _EVAL_539 = $signed(_EVAL_478) & $signed(-33'sh1000);
  assign _EVAL_360 = 2'h1 << _EVAL_3;
  assign _EVAL_264 = _EVAL_528 ? _EVAL_360 : 2'h0;
  assign _EVAL_591 = _EVAL_296 | _EVAL_264;
  assign _EVAL_284 = 2'h1 << _EVAL_19;
  assign _EVAL_436 = _EVAL_1 ? _EVAL_284 : 2'h0;
  assign _EVAL_484 = ~ _EVAL_436;
  assign _EVAL_586 = _EVAL_591 & _EVAL_484;
  assign _EVAL_227 = _EVAL_14 <= 2'h2;
  assign _EVAL_609 = _EVAL_227 | _EVAL_28;
  assign _EVAL_142 = _EVAL_609 == 1'h0;
  assign _EVAL_126 = _EVAL_348 - 5'h1;
  assign _EVAL_293 = _EVAL_14 != 2'h2;
  assign _EVAL_543 = _EVAL_293 | _EVAL_28;
  assign _EVAL_87 = ~ _EVAL_20;
  assign _EVAL_104 = _EVAL_87 == 8'h0;
  assign _EVAL_668 = _EVAL_104 | _EVAL_28;
  assign _EVAL_230 = _EVAL_31 <= 3'h2;
  assign _EVAL_252 = _EVAL_230 | _EVAL_28;
  assign _EVAL_327 = _EVAL_3 == _EVAL_224;
  assign _EVAL_638 = _EVAL_17 <= 3'h4;
  assign _EVAL_516 = _EVAL_638 | _EVAL_28;
  assign _EVAL_601 = _EVAL_214 == 1'h0;
  assign _EVAL_298 = _EVAL_24 & 32'h3f;
  assign _EVAL_597 = _EVAL_298 == 32'h0;
  assign _EVAL_316 = _EVAL_597 | _EVAL_28;
  assign _EVAL_33 = _EVAL_14 == 2'h0;
  assign _EVAL_399 = _EVAL_33 | _EVAL_28;
  assign _EVAL_669 = _EVAL_399 == 1'h0;
  assign _EVAL_466 = _EVAL_15 == 4'h8;
  assign _EVAL_559 = _EVAL_466 | _EVAL_283;
  assign _EVAL_666 = _EVAL_15[3:3];
  assign _EVAL_57 = _EVAL_666 == 1'h0;
  assign _EVAL_548 = _EVAL_57 & _EVAL_169;
  assign _EVAL_269 = _EVAL_559 | _EVAL_548;
  assign _EVAL_236 = _EVAL_269 | _EVAL_28;
  assign _EVAL_446 = _EVAL_236 == 1'h0;
  assign _EVAL_228 = _EVAL_7 == 3'h0;
  assign _EVAL_101 = {{24'd0}, _EVAL_143};
  assign _EVAL_254 = _EVAL_95 == 1'h0;
  assign _EVAL_507 = _EVAL_13 & _EVAL_601;
  assign _EVAL_567 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_610 = $signed(_EVAL_567) & $signed(-33'sh1000);
  assign _EVAL_217 = $signed(_EVAL_610);
  assign _EVAL_329 = $signed(_EVAL_217) == $signed(33'sh0);
  assign _EVAL_75 = _EVAL_91 | _EVAL_329;
  assign _EVAL_288 = $signed(_EVAL_178) == $signed(33'sh0);
  assign _EVAL_509 = _EVAL_75 | _EVAL_288;
  assign _EVAL_42 = _EVAL_8 ^ 32'h1900000;
  assign _EVAL_135 = {1'b0,$signed(_EVAL_42)};
  assign _EVAL_163 = $signed(_EVAL_135) & $signed(-33'sh2000);
  assign _EVAL_411 = $signed(_EVAL_163);
  assign _EVAL_125 = $signed(_EVAL_411) == $signed(33'sh0);
  assign _EVAL_649 = _EVAL_509 | _EVAL_125;
  assign _EVAL_100 = _EVAL_8 ^ 32'h4000;
  assign _EVAL_45 = {1'b0,$signed(_EVAL_100)};
  assign _EVAL_400 = $signed(_EVAL_45) & $signed(-33'sh1000);
  assign _EVAL_644 = $signed(_EVAL_400);
  assign _EVAL_551 = $signed(_EVAL_644) == $signed(33'sh0);
  assign _EVAL_202 = _EVAL_649 | _EVAL_551;
  assign _EVAL_187 = _EVAL_8 ^ 32'h20000000;
  assign _EVAL_461 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_168 = $signed(_EVAL_461) & $signed(-33'sh2000);
  assign _EVAL_209 = $signed(_EVAL_168);
  assign _EVAL_566 = $signed(_EVAL_209) == $signed(33'sh0);
  assign _EVAL_545 = _EVAL_202 | _EVAL_566;
  assign _EVAL_431 = _EVAL_545 | _EVAL_28;
  assign _EVAL_97 = _EVAL_7 == 3'h7;
  assign _EVAL_250 = 4'h6 == _EVAL_30;
  assign _EVAL_634 = _EVAL_108 ? _EVAL_250 : 1'h0;
  assign _EVAL_616 = _EVAL_634 | _EVAL_28;
  assign _EVAL_367 = _EVAL_7 == 3'h5;
  assign _EVAL_505 = _EVAL_2 & _EVAL_367;
  assign _EVAL_46 = _EVAL_389 - 5'h1;
  assign _EVAL_453 = _EVAL_30 == _EVAL_77;
  assign _EVAL_623 = _EVAL_453 | _EVAL_28;
  assign _EVAL_365 = _EVAL_190 == 1'h0;
  assign _EVAL_372 = _EVAL_670 < plusarg_reader_out;
  assign _EVAL_619 = _EVAL_301 == 1'h0;
  assign _EVAL_213 = _EVAL_619 | _EVAL_28;
  assign _EVAL_620 = _EVAL_213 == 1'h0;
  assign _EVAL_465 = _EVAL_11 == 3'h1;
  assign _EVAL_603 = _EVAL_31 <= 3'h5;
  assign _EVAL_657 = _EVAL_603 | _EVAL_28;
  assign _EVAL_74 = _EVAL_657 == 1'h0;
  assign _EVAL_173 = _EVAL_2 & _EVAL_228;
  assign _EVAL_471 = _EVAL_17 == 3'h0;
  assign _EVAL_377 = _EVAL_471 | _EVAL_28;
  assign _EVAL_525 = _EVAL_543 == 1'h0;
  assign _EVAL_225 = _EVAL_22 == 3'h0;
  assign _EVAL_235 = _EVAL_9 & _EVAL_225;
  assign _EVAL_332 = _EVAL_327 | _EVAL_28;
  assign _EVAL_382 = _EVAL_332 == 1'h0;
  assign _EVAL_262 = _EVAL_21 == _EVAL_427;
  assign _EVAL_216 = _EVAL_21 <= 4'h6;
  assign _EVAL_489 = _EVAL_216 & _EVAL_523;
  assign _EVAL_593 = _EVAL_489 | _EVAL_28;
  assign _EVAL_555 = _EVAL_0 & _EVAL_101;
  assign _EVAL_197 = _EVAL_555 == 32'h0;
  assign _EVAL_632 = _EVAL_197 | _EVAL_28;
  assign _EVAL_462 = _EVAL_632 == 1'h0;
  assign _EVAL_51 = $signed(_EVAL_249);
  assign _EVAL_592 = $signed(_EVAL_51) == $signed(33'sh0);
  assign _EVAL_643 = $signed(_EVAL_539);
  assign _EVAL_323 = $signed(_EVAL_643) == $signed(33'sh0);
  assign _EVAL_195 = _EVAL_11 == 3'h3;
  assign _EVAL_282 = _EVAL_16 & _EVAL_195;
  assign _EVAL_205 = _EVAL_344 | _EVAL_323;
  assign _EVAL_139 = _EVAL_9 & _EVAL_599;
  assign _EVAL_417 = _EVAL_26 == 1'h0;
  assign _EVAL_336 = _EVAL_417 | _EVAL_28;
  assign _EVAL_607 = _EVAL_29 == 1'h0;
  assign _EVAL_483 = _EVAL_15 == _EVAL_181;
  assign _EVAL_536 = _EVAL_483 | _EVAL_28;
  assign _EVAL_351 = _EVAL_536 == 1'h0;
  assign _EVAL_200 = _EVAL == _EVAL_105;
  assign _EVAL_384 = _EVAL_200 | _EVAL_28;
  assign _EVAL_124 = _EVAL_7 == 3'h1;
  assign _EVAL_608 = _EVAL_2 & _EVAL_124;
  assign _EVAL_220 = _EVAL_22 == 3'h4;
  assign _EVAL_238 = _EVAL_486 | _EVAL_28;
  assign _EVAL_129 = _EVAL_607 | _EVAL_28;
  assign _EVAL_68 = plusarg_reader_out == 32'h0;
  assign _EVAL_305 = _EVAL_205 | _EVAL_592;
  assign _EVAL_281 = _EVAL_305 | _EVAL_28;
  assign _EVAL_373 = _EVAL_10 == _EVAL_401;
  assign _EVAL_183 = _EVAL_373 | _EVAL_28;
  assign _EVAL_117 = _EVAL_27 == 1'h0;
  assign _EVAL_240 = _EVAL_493 | _EVAL_364;
  assign _EVAL_276 = _EVAL_183 == 1'h0;
  assign _EVAL_287 = _EVAL_238 == 1'h0;
  assign _EVAL_387 = _EVAL_553 != 9'h0;
  assign _EVAL_222 = _EVAL_387 == 1'h0;
  assign _EVAL_47 = _EVAL_11 == _EVAL_161;
  assign _EVAL_58 = _EVAL_47 | _EVAL_28;
  assign _EVAL_531 = _EVAL_21 >= 4'h3;
  assign _EVAL_490 = _EVAL_531 | _EVAL_28;
  assign _EVAL_589 = _EVAL_490 == 1'h0;
  assign _EVAL_62 = _EVAL_7 == 3'h2;
  assign _EVAL_604 = _EVAL_264 | _EVAL_296;
  assign _EVAL_428 = _EVAL_604 >> _EVAL_19;
  assign _EVAL_194 = _EVAL_428[0];
  assign _EVAL_186 = _EVAL_194 | _EVAL_28;
  assign _EVAL_458 = _EVAL_186 == 1'h0;
  assign _EVAL_107 = _EVAL_553 != _EVAL_542;
  assign _EVAL_128 = _EVAL_107 | _EVAL_222;
  assign _EVAL_450 = _EVAL_128 | _EVAL_28;
  assign _EVAL_614 = _EVAL_450 == 1'h0;
  assign _EVAL_500 = _EVAL_350 == 1'h0;
  assign _EVAL_460 = _EVAL_0 == _EVAL_635;
  assign _EVAL_354 = _EVAL_460 | _EVAL_28;
  assign _EVAL_479 = _EVAL_354 == 1'h0;
  assign _EVAL_487 = _EVAL_252 == 1'h0;
  assign _EVAL_237 = _EVAL_59 | _EVAL_28;
  assign _EVAL_226 = _EVAL_467 | _EVAL_29;
  assign _EVAL_234 = _EVAL_226 | _EVAL_28;
  assign _EVAL_378 = _EVAL_234 == 1'h0;
  assign _EVAL_517 = _EVAL_516 == 1'h0;
  assign _EVAL_149 = _EVAL_7 == 3'h6;
  assign _EVAL_294 = _EVAL_2 & _EVAL_149;
  assign _EVAL_356 = _EVAL_2 & _EVAL_62;
  assign _EVAL_203 = _EVAL_668 == 1'h0;
  assign _EVAL_625 = _EVAL_58 == 1'h0;
  assign _EVAL_402 = _EVAL_497 != 9'h0;
  assign _EVAL_88 = _EVAL_402 == 1'h0;
  assign _EVAL_147 = _EVAL_88 | _EVAL_68;
  assign _EVAL_572 = _EVAL_147 | _EVAL_372;
  assign _EVAL_415 = _EVAL_572 | _EVAL_28;
  assign _EVAL_158 = _EVAL_415 == 1'h0;
  assign _EVAL_621 = _EVAL_70 == 1'h0;
  assign _EVAL_582 = _EVAL_593 == 1'h0;
  assign _EVAL_405 = _EVAL_179 == 1'h0;
  assign _EVAL_605 = _EVAL_628 == 1'h0;
  assign _EVAL_37 = _EVAL_495 | _EVAL_28;
  assign _EVAL_650 = _EVAL_16 & _EVAL_465;
  assign _EVAL_212 = _EVAL_22 == 3'h1;
  assign _EVAL_624 = _EVAL_11 == 3'h0;
  assign _EVAL_165 = _EVAL_262 | _EVAL_28;
  assign _EVAL_580 = _EVAL_171 | _EVAL_28;
  assign _EVAL_122 = _EVAL_580 == 1'h0;
  assign _EVAL_385 = _EVAL_237 == 1'h0;
  assign _EVAL_477 = _EVAL_497 | _EVAL_553;
  assign _EVAL_330 = _EVAL_11 == 3'h7;
  assign _EVAL_309 = _EVAL_16 & _EVAL_330;
  assign _EVAL_611 = _EVAL_117 | _EVAL_28;
  assign _EVAL_83 = _EVAL_12 == _EVAL_576;
  assign _EVAL_185 = _EVAL_83 | _EVAL_28;
  assign _EVAL_279 = 4'h6 == _EVAL_21;
  assign _EVAL_432 = _EVAL_283 ? _EVAL_279 : 1'h0;
  assign _EVAL_271 = _EVAL_432 | _EVAL_28;
  assign _EVAL_627 = _EVAL_271 == 1'h0;
  assign _EVAL_206 = _EVAL_617 == 1'h0;
  assign _EVAL_263 = _EVAL_109 == 1'h0;
  assign _EVAL_103 = _EVAL_9 & _EVAL_220;
  assign _EVAL_571 = _EVAL_24 == _EVAL_574;
  assign _EVAL_292 = _EVAL_571 | _EVAL_28;
  assign _EVAL_153 = _EVAL_292 == 1'h0;
  assign _EVAL_308 = _EVAL_404 | _EVAL_28;
  assign _EVAL_423 = _EVAL_308 == 1'h0;
  assign _EVAL_452 = _EVAL_2 & _EVAL_97;
  assign _EVAL_192 = _EVAL_304 | _EVAL_28;
  assign _EVAL_470 = _EVAL_7 == 3'h4;
  assign _EVAL_338 = _EVAL_9 & _EVAL_285;
  assign _EVAL_312 = _EVAL_384 == 1'h0;
  assign _EVAL_473 = _EVAL_7 == _EVAL_50;
  assign _EVAL_131 = _EVAL_4 == _EVAL_568;
  assign _EVAL_664 = _EVAL_431 == 1'h0;
  assign _EVAL_44 = _EVAL_16 & _EVAL_624;
  assign _EVAL_646 = _EVAL_9 & _EVAL_212;
  assign _EVAL_422 = _EVAL_185 == 1'h0;
  assign _EVAL_429 = _EVAL_493 & _EVAL_583;
  assign _EVAL_289 = _EVAL_207 == 1'h0;
  assign _EVAL_520 = _EVAL_616 == 1'h0;
  assign _EVAL_412 = ~ _EVAL_542;
  assign _EVAL_246 = _EVAL_477 & _EVAL_412;
  assign _EVAL_420 = _EVAL_473 | _EVAL_28;
  assign _EVAL_444 = _EVAL_37 == 1'h0;
  assign _EVAL_437 = _EVAL_192 == 1'h0;
  assign _EVAL_391 = _EVAL_364 & _EVAL_111;
  assign _EVAL_297 = _EVAL_420 == 1'h0;
  assign _EVAL_442 = _EVAL_623 == 1'h0;
  assign _EVAL_84 = _EVAL_16 & _EVAL_52;
  assign _EVAL_636 = _EVAL_272 == 1'h0;
  assign _EVAL_127 = _EVAL_165 == 1'h0;
  assign _EVAL_667 = _EVAL_377 == 1'h0;
  assign _EVAL_374 = _EVAL_9 & _EVAL_407;
  assign _EVAL_570 = _EVAL_2 & _EVAL_470;
  assign _EVAL_245 = _EVAL_316 == 1'h0;
  assign _EVAL_584 = _EVAL_336 == 1'h0;
  assign _EVAL_662 = _EVAL_611 == 1'h0;
  assign _EVAL_409 = _EVAL_131 | _EVAL_28;
  assign _EVAL_455 = _EVAL_409 == 1'h0;
  assign _EVAL_215 = _EVAL_129 == 1'h0;
  assign _EVAL_116 = _EVAL_281 == 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_50 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_77 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_82 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_105 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_113 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_161 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_175 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_181 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_189 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_224 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_239 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_243 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_257 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_296 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_348 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_389 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_401 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_427 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_497 = _RAND_18[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_501 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_549 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_563 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_568 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_574 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_576 = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_635 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_655 = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_670 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_18) begin
    if (_EVAL_386) begin
      _EVAL_50 <= _EVAL_7;
    end
    if (_EVAL_429) begin
      _EVAL_77 <= _EVAL_30;
    end
    if (_EVAL_386) begin
      _EVAL_82 <= _EVAL_8;
    end
    if (_EVAL_391) begin
      _EVAL_105 <= _EVAL;
    end
    if (_EVAL_391) begin
      _EVAL_113 <= _EVAL_14;
    end
    if (_EVAL_429) begin
      _EVAL_161 <= _EVAL_11;
    end
    if (_EVAL_28) begin
      _EVAL_175 <= 5'h0;
    end else begin
      if (_EVAL_322) begin
        if (_EVAL_499) begin
          if (_EVAL_660) begin
            _EVAL_175 <= _EVAL_472;
          end else begin
            _EVAL_175 <= 5'h0;
          end
        end else begin
          _EVAL_175 <= _EVAL_114;
        end
      end
    end
    if (_EVAL_386) begin
      _EVAL_181 <= _EVAL_15;
    end
    if (_EVAL_28) begin
      _EVAL_189 <= 5'h0;
    end else begin
      if (_EVAL_485) begin
        if (_EVAL_214) begin
          _EVAL_189 <= 5'h0;
        end else begin
          _EVAL_189 <= _EVAL_151;
        end
      end
    end
    if (_EVAL_391) begin
      _EVAL_224 <= _EVAL_3;
    end
    if (_EVAL_429) begin
      _EVAL_239 <= _EVAL_17;
    end
    if (_EVAL_391) begin
      _EVAL_243 <= _EVAL_5;
    end
    if (_EVAL_28) begin
      _EVAL_257 <= 5'h0;
    end else begin
      if (_EVAL_364) begin
        if (_EVAL_529) begin
          if (_EVAL_602) begin
            _EVAL_257 <= _EVAL_86;
          end else begin
            _EVAL_257 <= 5'h0;
          end
        end else begin
          _EVAL_257 <= _EVAL_546;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_296 <= 2'h0;
    end else begin
      _EVAL_296 <= _EVAL_586;
    end
    if (_EVAL_28) begin
      _EVAL_348 <= 5'h0;
    end else begin
      if (_EVAL_493) begin
        if (_EVAL_583) begin
          if (_EVAL_60) begin
            _EVAL_348 <= _EVAL_196;
          end else begin
            _EVAL_348 <= 5'h0;
          end
        end else begin
          _EVAL_348 <= _EVAL_126;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_389 <= 5'h0;
    end else begin
      if (_EVAL_364) begin
        if (_EVAL_221) begin
          if (_EVAL_602) begin
            _EVAL_389 <= _EVAL_86;
          end else begin
            _EVAL_389 <= 5'h0;
          end
        end else begin
          _EVAL_389 <= _EVAL_46;
        end
      end
    end
    if (_EVAL_391) begin
      _EVAL_401 <= _EVAL_10;
    end
    if (_EVAL_386) begin
      _EVAL_427 <= _EVAL_21;
    end
    if (_EVAL_28) begin
      _EVAL_497 <= 9'h0;
    end else begin
      _EVAL_497 <= _EVAL_246;
    end
    if (_EVAL_391) begin
      _EVAL_501 <= _EVAL_22;
    end
    if (_EVAL_28) begin
      _EVAL_549 <= 5'h0;
    end else begin
      if (_EVAL_493) begin
        if (_EVAL_413) begin
          if (_EVAL_60) begin
            _EVAL_549 <= _EVAL_196;
          end else begin
            _EVAL_549 <= 5'h0;
          end
        end else begin
          _EVAL_549 <= _EVAL_434;
        end
      end
    end
    if (_EVAL_386) begin
      _EVAL_563 <= _EVAL_31;
    end
    if (_EVAL_429) begin
      _EVAL_568 <= _EVAL_4;
    end
    if (_EVAL_448) begin
      _EVAL_574 <= _EVAL_24;
    end
    if (_EVAL_448) begin
      _EVAL_576 <= _EVAL_12;
    end
    if (_EVAL_429) begin
      _EVAL_635 <= _EVAL_0;
    end
    if (_EVAL_28) begin
      _EVAL_655 <= 5'h0;
    end else begin
      if (_EVAL_364) begin
        if (_EVAL_111) begin
          if (_EVAL_602) begin
            _EVAL_655 <= _EVAL_86;
          end else begin
            _EVAL_655 <= 5'h0;
          end
        end else begin
          _EVAL_655 <= _EVAL_578;
        end
      end
    end
    if (_EVAL_28) begin
      _EVAL_670 <= 32'h0;
    end else begin
      if (_EVAL_240) begin
        _EVAL_670 <= 32'h0;
      end else begin
        _EVAL_670 <= _EVAL_640;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_418) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_664) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52382c22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918c4d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_664) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(272e4fad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_507 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96fa9775)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_351) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2015e7dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_669) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77982d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e2d132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f7fbce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_605) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72242a7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_370) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24ecac41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_662) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba42c796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_507 & _EVAL_422) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97903ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e09b719)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_662) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4f3c454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_669) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_669) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_664) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1d5d305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_423) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_627) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42a579d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b34659e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_405) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c02c2e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcb4cdbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_669) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5c2c5f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa4af3da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_584) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ef55c03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_669) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e18d151)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23223b66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e1e2286)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_423) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efaded7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_584) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d183075)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(515dc8d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2ceee07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdec5e31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad4ae52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53526990)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_382) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_621) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b143c629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a8809d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_662) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611411a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_479) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c46fa700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f696ef6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_662) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b2536ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_664) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_455) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76d8675d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_582) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d968cc38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e1e419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_584) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_662) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc779b5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(897c83e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_605) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_520) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b680c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f243ece4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a930e63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_669) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd9f3b0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_584) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_520) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_423) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(339ae757)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4db2120d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_444) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_625) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ada23f2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b49e3ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c847707)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62638d12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2396e2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad580a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_418) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c73b2fdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_620) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(360c5011)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f9073c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_442) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_418) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_669) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_667) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_664) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8f9ed6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_500) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8207de3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_517) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83131c73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0059c0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_667) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caf8c29d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_418) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e86a431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_423) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b81d323d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_664) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_455) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(820ca019)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(483e5190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_442) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74a44400)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e162987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(302b5cc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_625) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2d1f1a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_605) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe75bc99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aba5625)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec0ea252)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_458) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_520) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1802e06d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a9b4e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98817fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db2f6ca7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_664) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_621) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_525) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7f72517)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_370) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3389808b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_614) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f171119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_584) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2999ef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84350161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e157559)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_528 & _EVAL_437) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3fbfc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_662) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_667) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74bfbc26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d0f91e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_517) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a57ddb47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_370) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38a0a437)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_636) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfd30c4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_627) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(176e8137)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8012f30d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_374 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c8896a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29c475bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72649d15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_444) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d03235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_479) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d6671d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e64e5922)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_378) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5b73aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71c5a702)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_667) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_582) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ef66ba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_627) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8fa056f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c4015b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea40977f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_487) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93984adb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_662) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(482456c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb134dd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80ff6e85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(499edfb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_584) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dce5c16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_370) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_462) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a53e40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_457) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d09899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_457) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc7be6d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a099cc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_525) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed249b1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_385) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd4781f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_667) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d3ac770)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_458) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf1f42eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_487) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdeb136)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_664) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b131741)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_520) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_405) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe73c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_662) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_446) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f1435d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_589) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380059e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_642) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a309ef4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_582) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caa3789b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_664) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa4a97d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_664) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_669) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(340dd7a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_584) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a616b07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d8bc61c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_667) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f233117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_351) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a7c9dc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a109775)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_382) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4694c43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_528 & _EVAL_437) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_642) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db895fb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_507 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_584) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db1d514d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_507 & _EVAL_422) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_636) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_385) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_582) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_605) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad8d5f5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b9e8859)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11ff4447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_620) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_627) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_500) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
